-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NrFIuk+mxcwQ2XFvNDV0QPHqHQDjbhs99XtNZCgA/22RpZHHdX5Oj6L5bQOv5/9edCPcidepFCrN
o0hpxZjr353qjGx9v854Btths1F8fm5bjEUWCyRO18VnUn9tTt8QNk6nUHmpU5gfyl8KDa4h1WbF
u0JqOLC4yvRn5p4zWZVdhrr5CYgRC8DVPIU3ew0UPSk04/1Ziz9+sGJDsheMUQsGy9snmOq7jcBq
I3I5DnwuYUJuNq0hvvEF6HNo81GskugDVcI7j/PFbkQ3/pZfxleMb0sZ9bBY+UkdBI8dpoUlD2ve
YdcaGSWBn24gU13TuDhpGwg+IClvex5pNS9DcA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1040)
`protect data_block
wvouTT0rXiXQxZzsZt3G0pGAG3TkVkNuHdeVZnPmexX8SWRoiWwkFFtyd790pBjmRDasDHbkK/cu
eJq49e0O7fyM77GX9WXRDSBCKrFaLLac7Y1i98w3kmFR/qfzAaevt2w4WuZKxGbP8reBqteC81Z1
tqXuBcS9Ufw485JCzoMUhOATmLSLN1tGYjTbAbHMLr1vLKbwNNIlZ5n/zPOLbFtaQ+0CEpTjOa6t
nafQUbp/JWKR0yEW1PdyY/oVSKREiGjp3M5ZNCGIo5+e5uQ0EHF5qICHoICFPtUwppz9i9ReMvty
ve2Nblgmjr9UJ2zzvSuCu3gw0VmfDQSslCE2l1RzUYC2Ek0IloGMQ5M7iue+S/S3FQwDfR4SqsuW
i6b2c6LXQUOvLYloRGxCG+5eaRcYastwxYnF+1dOGQJ6QwR+nML3ni3WLZeeYXJF0pcUpDkUpWM2
Mv5IqQAtM+soxVRerSQS/gRIXr91pRd6rDkMe24eWl0z6xeKzoD9VmtQDWoG7fYLQOYdAxpp2bDt
rKtM1soEv0n20XgWUOEtFhX4vzHZwbdPfI5ZjB650ih0JnK04fAJDeUXAOXlEqOnciEqIaI6I5bu
ENTGXqz3Eo/demzmCITPw7rSoL6fMyuRM5vmuHoIDm63irpUG7fOkYT7nnyaphBUjZmyav3P9rRo
F7aOq8b1JzmdVG342cwHlkCy9Dg3bq2bJPwZBYYFRLKY5pqznpxGBqG+CJN5NAstmO5yWg/uhJ/C
q3d46WxDEI/xwmzPn2cemq9Vj/WLYOq1gmVtm+gSo3q6iu9/bcrrqyJ/E51OvDQVZeTvQU306Bfw
6ZmOIKKhGRoKed5MjNvi0seljnLYLz3RAiOisbm1SwuhnoIMs0tVhFrVzZMIbu0iEuPqbK2H5lsj
n6Ckuv5HPgF3zxzGLiVeYMInd73boKb9yVf0ec/rdTw1ttsMzbfhhP3TjdwZyR98uu9s9PorxQLL
DAKizKY0uKHz2tUKJ/NfyBUh1XMquB8LXMbk1XuW/z2drMEc12gzAlMg25ZfRcA4BKUfgNHrvuxC
EyTxWFY0xb1sALn4Ea8zElqXuOJVZawWLyBFm0GJqnHGkZcGTYol7UBap+wHHNU4IRWCudorSidj
8MrIb6exw5cHdIv+2rXYRLmKCXUYwuKFFZsqI+tPGKeBaxcnGjTpeIZOerrqV6ObXT208kFs+uFG
Ykq0S2bvH6UBLhtxOjXbG/fZwj9+k58UQcQLWkQrJDXFz3UL7H7Cohcm4rn05nMj0TVOfoXLqXVm
uCPGXxjSeKCq8XbMBOwPaBt3bzaQYmnKg6hCJ0e2XAGrGAoPy1FUgVk2uTd2kNnx612jCbR2wc0V
P2NG3FPolqjA1OCQ6RI=
`protect end_protected
