-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SC069JAEj/jbhfmDEwXQt6/TptvnEFUtZj8tYNoqx3x/OVoZlxLjLdO9nSHpu5adkBSNHeVOaA+G
LAL6Acv+HvT5aYUxGNZfCArXkWDbW7rj/94LJV+3WzfGu71RoRRMLds1I6L1MnvGc50+LSEjSR4T
/vWhkbvkLC8+KuP156FSEX7wyU/tQ3y3IEVTr5h2fdBbgiocsuVWLcBTrwILyk+2vo6UR+n8SseG
fMDp2m10F9sI675WAzCxJ+0y5YAFnoi3RGLe29as4stzIW6G3bzP1OD145mRIPxtIUglgjhU+sZl
ASLcDWvJhFSpdw8ghciLptqoYHGl4RW2TntTOg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11552)
`protect data_block
n1Sh0JcUwHb4XB4mMOTdArkuWcckcUzf/zrq0cosOGz7nZwX/3APBbXa5YgHxNCQuOqXpQeGcShw
0pX8iST5F0skZ5dG7IMURI8c1wB3v4J+n8ltMWxVbg07lHXkRYM/8/9ZlmVxwh6p+7sTEGxcIela
m8muQaunDWvgQ1N7c8cBbJ0IZeBGSZsntElVZpyzUfeIfbCHJwh5tOQfR8Cn7VUvTA3kL6zyOHMR
CqTxtPeXUAu/FX+ID0ZHlL98BtEnVIi/HE9DOhsBwqWti5zm/00VRqmnNGOM6GOqdyxgskFGSe1W
8yYur5NAXA6j22pse/xZGcE04Y41t4IHSZogq4aWswny+LWny2sw3ncxhcqHcOCl0EE5PF51YdVB
yCC5TwmCnr5yq7zLsaAaNzN12uvGjtulgS+oxE9YwYcz8C6N94LgTAYGjdgB9XB3BZscI/YzZwD6
7K1ykUyXtGYzEy8aFyHibaXKhD57HAdMnTpGaZEuyAmSBlmnb2X4ehS96STuG6Nob9pVdu5/GkpF
B+8O92InH90z9GB00zGbsdrS+NjQh8O0IOLThDqNxm1iYS2z3GLHi35ZUyswZV3lVRxJn3fgV4D7
OCJr2q1qpjzI4UYlahU6pGeYXUm4W8dvTiWd5Dv2zoyM5Cth07K7UI1x7cBGB9H1/mqaFu03r8IE
eiUVE+sQv67hN5bMrq0BGGbH/Lw1kPYR/0rzk0xr1zMiklZewDWP7S/7OOJMoEBHIVf/I+MPrBPR
B3csE0CfMtZphmA3C7GP95pazTiWHQ3WXWzhCUJ+8LL7FLcbdiuWAYfA3FosZGM+TiVHNwjghZly
Trij+D6P1oTxeBHV2+e51VQxOuWtQ/CJkRyOrubgqltwsfBCNPvx6zP1qi5WmMNHVpDw5Z3OqRcR
2z6QNTj9WHf2iW/zuUblZU6d5zU4Pqj9IZgDg4/6Vhd1dBUxpDtl59NMGOQ/UJPomyVNVl1PYYL1
mgRroSGpkso6PF9yfax6Rv9KaG6uyhEwP1UveJs/wUTmwfvSkApmykP410X0mX/g5PLoMIvIbn6P
0WN/1rc0u5ZX1P5pEKUA/7BZAD+SPSrbokhVytTsGkpo+zN8uOTlapRiBQ4xU1Tab7QoVfU0bXkV
nEQoqCqx9hPnOusbwyjsWUJAqGNIaPaf3mvHAu5H0ULC2eFH5xDekopaV/CXWa/W+BNdbnCwhAUu
9bq6wqRj/gQguH448D9ncPcM3V9zwVjHif9pYxHWZpCKmQfZCBbBNl8heJQyqQ0p4vjXroqbKZ9F
lJR3HHAmwRGrzwsblbTD64E0d/prWFdSjxwwTcXaVsHiTbF9mm9KHx4nts0UNDLM5C1o/luQheO6
OHWe9SQHLJv432Y6/js63M0xnegGC0PanSSgWGdwQ0RS5oGXYrF8gSVHrajXrzyvfBoIl56uo2jz
SLgd51/KYTGr3MUFp81zhhBVmmctKvgXqqm1XRr59Lgw8xIrvtenqo0cRnp6QUGILpVeaZI+y/yO
BQd1CeZDRS0XbMpug7xyASm9LCbF2sMVw0bQFENI10HhJRBE+ROfxGjthyl2OqgSrzvqG/gRmHdo
YASw7a2Q2v/ODl6yqKW1eSa9wtVZ3JttEzZtTvcbUiRn17mzFZY6mTqH1+f7S6Yi26At4MfsDTOS
c95UA7AO/2bOziObxjsJjd03iZ+AMPV9FSeLR8DYPs9pXUCl64CUWEOF+JextnkBd27t5WDrr6YI
Inl9WsyUfWvTOWfWL4vKs0IJHxxtSIxmNrJHBUjcPhwKh5PSi+DejWxb/WRnHqsgq29F/aNH3I25
gPK8fo5qom/zx5gFnEQUWHGn92YelEkHp7XbSCS3RAkNofs9YBW5aPQyATBFYV77rBhsV4CqbwJK
wjL9qYxLAsSZOQyi+hvhMjCBW+8w50YCIYWxDbB2jzmLgIbQjaitg3WyZ0WEz9hIp/Rx7bMydybX
f+clmWuqCYGaD3CxyXPHev5xykYo7rx3MiE7myFZRD0hUSF8ph+4Qv0HXap5kIi8RwJ25a8AKi9X
tdhrIcbqbA176ET//oxb7Ob1YJVWfwLqtgqwl8C5JfJo6W5uGq+z80p8WD5Bx4T18j0+VOAvSA2M
SIoMWunwViUDblsOEg95+4G8MIngPp7OnL9qYIW7ZGeYGRh9U6Z1MHFnge7B6Qp3dhM48KefqqFY
BCJhJLs9kycATJqI/CiWCR6rjgPxnTwZZBYCR8yTOBKdrchbBCEca6liueA0gCxMv8R5t2Cojtvf
v83XBohVp4Jei6l1b8ZtHoUpCOkvDm0cwp44w0mH4quMUjy2Sjn4vYSdLo8w8OxO/YrSbKyXvhTG
IvfT9jS2hFDITQHZ/pHEEmqaREf6zAPWx1/MD9+NYrnbKwMG88whrQoE6m2YbskV31G/Qm39D8P8
tK6lllf1SPbB7lFo+S1BYJ87e8dobybG8aaynV364VjBQnqBbAty6gdge9MDE7STp4fD432slzu4
eoP3qaHKGfV2fAGbjc8dchMFKAJPKYOzQdDq7UvGNRy2Eo01RywzN0imios50DIjTwyyv/WIJ/o3
e51dqJZlzOJe0Jf7xO9/y38CZCh/MfJQlhp4hr5gvFXnbBORXVtZ1smcdUlb82LADMU0VLKnOH0b
suQEYLDW0HF9K5KUYQ2gZF1BYaITbPvmx7qXmigkgp2oIGCxueefL3vwP3gGiYIf9Gt/Y1VjWfxp
LntAMLgsX4L8uoMUc5UOppYDUA4CBexrBfhXVSainByee1RcH38pu6RjMGf8uv4ZKWrzw7T5dN/W
VQLEq57omREcm/HM2Nq/pD6bRF78moee8NXikNj82lxYKr0rcyBtZQ882XOooDp6wFeL4zduORRT
pQ8RNCF3CTpq1QNm5K8BD1xUMUE8uUEZ8H7n4QQ4cXdrssBhjeu/yFl+VomynZ4nBT1FFOKR9jtm
zkcrcm3KfmBpMp2LpKAojKdSSZee+fO1pkOcGuOu4yfas5b4DK/8y5+PpvhqsUL9o92GIe8YGtP9
ffSreeefOfm7cHk3t9bWg3xBvyTn8LrCyY8I+q8C5PCfUSva8rpr4o+MGqSvbRrZJYj/r2ETTXZ9
XOM5bkQLFek0Cc0cvEF09hQ6xyhReQ4jYwRYJqlkeA9sURvt2CiNEr8aWmpfe1d9QIhqjKTeGViI
C12t7WNkGOQ4qUIBUoCg10GhWPzFqpd0LRlUysKDbee3aGJ8lIFs6jA+Fiekv4MVPjQciyslIaim
g6Gbu1cs628Tj6/XEf5uewasJcsphmD6alCP+0Wbq4tf78nRdAgqE6LiEjmC26ZeFGjzGOtKo6PG
c6KD2d+uu5xW4RVtGETFv2i9HYKcSjFGh40rKGfx3lP6e7fXqXX5VvCrFzJWVZXSM3QE3FCH0XUT
JG0Fpr2GZZAVXcLPz8le4CbXiFXvtmqJwn/7Zt0AgSlpe77Kw81iU6U1OLrtN+Xw/E26ozmYriew
r7KhiErG3y86Vde26l3IIMnA8svO5N7rBn2yE0AqxDcqqO6pftxWIIO2dRwfb1qeR0VuRv/hY6dD
jcK1NdFUVgoWSVRWndkb+JOTIUa08em8HMw05O+ir7j0pm5RAJssuxSyslj3wotV6CvcB657yqh2
xaUIhVnlXt4+Ck8MZkkcVjGmLlh3WRGmLEaJlmaSPZgifp4Ac2mNa6hpOAtYj30wqm2k6Dcoh8Ca
Gh1GBd0ThmmyLG87CD8h+yIgXubuPEDSp27CaHmOKQsv360msCk82jLeK9eGlYBa+2s9hfG5YoIR
qoknMMB1ZgbiHMJP2zbIPUrc1g6cFNM4POfR48H7KWJtq6IHLtjZkfwC2zVowZay+pwULPhXm9P9
0l9pk6AO/B3yvyztWnetnayNhGu6g4vRTxwWYMirjQuwSZNl4nsCn9DNJzCbM0ty7f1LI8qCecNz
DqTA4LC/E3CZzdUS0BuhGpIOpZV0GGcdBbwAOaWNKjQ97VZdiM59US9Zwr+iRiMarl8XywXnS2mT
PSIGnk9fzGbr1krOcjo8+wFEg/qtlCHb9LNRteax13Pqlz6ePRdOp5uGXKWBHNaTwjUcEgfk/kNc
LOHDxwzaYtUY5gXnjQTUCQRoLYk9K0HRUOUg2LX7/K05Fnl8Y6+3ivFgVptUPTew5Er1a/R2Vcs/
HU04+VKuLEf+6UKbkEVpd91WQK5v/Si1XLXbmHRD0loe4yzHJ8WSfTLFCcOwrXBujN7BD5EYpIyy
0gMKMLsgIusgy/FH2j7yPhKwzLWcGoognkN2YBGXaW7VewU9oYu2CiTYFX+g7yfMS1e1Tb17nA21
CxoOOxa0T4N29XroegXpSnllT5L1tQh2YriUviYvRz5I6mROeTTEdY9dJuam5KZTTDF9hTYd7t4F
LlI/WUDHXQSWgLlV7aa5CIlVaTD1KcbRaI1KAlKLViiPQD99PvKf8xbLpRjBCu6u1UgjU69KMr6P
JiY8hZfAY5l1y8B5QlBTo+UmUHURmYLDoORE9Sme4j4qdnBWZhi8tC4P1/ot72p04T5Aism7sRFe
JA96bHVgL9PZCTPcwHfpHvMuDYAz7G7g5yYbMFo6Dkb35qaL+wIAEuGojQ1gKaoSX9gGJ13pqD55
M4Pyr4ppc1TAIIiBPZtkUoKbW5tbLbbLjZOccGHZHJdaSU8Ol/KU3xT/Pb5Qb265Roab4uKN6B3+
hY/hHCVI9drgs+2Tl79zEbp/Vi+7G34+SBXWsI05nA4bYwXrI/WlB9xJ0bsNQcEWy7E+F65sfsu3
5JHa9kwHDmzroTiRjothh4ua/il9fIJIwCazDDDGpz6UphJhx+6DADyz9oCOykEgYhaVxyM/LCxz
Mx95cHYnN/XSmTbKZqAFQcrF77pttxYtQyNr6vU6Nl4HqnBDszSp9lR/T+dHjDf6nfgv1bTmSX0N
CKlJUk19dAnRsOGNTz9hIiA8RPnMYd05Rh3ULFVWL2VhIRCf2nbqM0nPE9tcZRPLIU7TYvYReiI+
uyZwcHZ2MvxDk/asQduV2CC766/DqJvMkgc4H3t4scHL6lO/HEIVZJ5SSmntqXeG4po36ctRgz72
kLXg9+EFxZMAcDvAp6okCR18QkTMGXr7uUyxtohbYuJgyAnyFEdV1zxs1jq3kw2A3LF9ia9mr3G3
dBs54zqKmOuXAFOAbyB5Bs85x7MudEbQVpkvK6K6dxIfW2FpLYJfDpepvfeSUI4jLXRIWx8AkgY/
nOaH0mUbqTZlvueUEICRZ4m0dVAbpXaJeAMbDR8jNW4sCxk0UWBDZVU4BM9XcOrnpl8MNLYTHdOk
YSKKO0OB0YyGABBtTZRFLNv51viVMIDqKd+IQiaBV4Nq4tBmDtCCfYJtCGPNfB89kWznIoevOMP/
aZ1a2AGeO64QI8xKRZ0rb9QW9zpIOmQBlPbuaw+Q9JqmFjyiJ1PV5K9FJm4T7Ivzi6pn4yfPfj+4
dVS/GhsJGUMwHpJKVtfmz/lzauWbdSBCkjeZFdSL3CfT1VBt+x+iUS8t/4yZ5SS9rAY8E72K+xJk
ImhSw1AtdO92yLWjapL4Vfc6lSJpB7ABQ8DHisZxrmAvVVbUypM4VQzMt6JSL9pqisb6vyeFbLNb
CDLKl6xJ3w3aXOl3QHoCx2acJ3yCUw22Vd4Itiot4H4D7k6kTlCy04szIqKt1+abNpCbE7snY/xo
AFz+32JywA4IMDm5dRHOCf1FFVBAeYMdORjLqbTZvkPy2kN4hPYE5ogdoanSn36WEZdCTRpdyj3w
TtBOkRSjZid61t7zEBUdVPxtHa+SaVaxrQBRsdktfjn/JGATqVIB9FR6aPW3KYTB14/iCz1V0j9/
OFpQ6zitG3FI5pKmcPn3rb8m7ni/hhdtWIjLFjfAQOeM3wZcgV/Obp5pYJJv2tjQLSGTLASzrCl0
cNvCdxAMbwYGcCkLh/fyvUN0BwIXlH+RMg3lp3RsbaVS88ord+HnkLrMCTeXaP0IFPgsT5vAoDqp
O1FjcsmRYKhnyeJLCtN+7x76/maBwPG5DfyS36VZAty3acBOLkZNCxB8OgBK/CiaS3PJw19NWECx
irZS8L3QsMBvJ16ExE0r7H0Iskk4wujya7PudHj9dbIUckKvqtWErOIxBkRAdaKqLi0GEWwZN6yO
g+S8214QwTbWFbZuVNSfz0+NX+l3GA/XbDYiXEr3S098MhkCyRa5v7sGj5qNr5HTL0Zm6QQEB736
krsiLJA3zOLiE3DBSzUtlRU2GKfuJlh+yX1tz0uHVM9JEcIlfVl440XBYZNQE/x1Y/H8b98n9R7K
CLuxh8eSoQTCLAKWRBJUpCKCng0ijMEL4oiEMDBjPUwIsYL5dNi6gFK8ENAz+ECxJDEOZgEiA32o
xY0NIWPxQ6wEhvTl41dCPQeSnOgr9TYS5I4yIPOSjVGbCcZKZSdxpRK6IJuXlnZ5kg77bbTwnumA
rnnubNG/ezvyjwHdekBR7M/mP/MSCI4daeSxS1jQBI4WT/iw9NkpsXrkABvS1XptxwZYezsVy5fD
ppHDK+C9Fat0nLWgo6fkvjLUNRb45HREtxPm53LakPi0u4ijCvvBeu3KKWYXtDHArZCqMjNsivnl
A0FkzMiVZlnj7K2TxnFzZqWe5Dj5L8VnHUrVmupVBZepTISe/YvXpV6K+wpSLqyU56mgeHEfoBeZ
hD4lj+BQTeYk6ZKKydcLzW0Eu0v9UOuS9a5F3ebQ/0tDIMZ7YIwx9M9dPXFrVnuD9/BmFR8YzHsv
6lzv2Rn5S43P0IzBJmAfBJgATFxGiBVO1yKAomDUiRh5Bx+EHdVgZGR6btX8R6zE0HQHRWNXpmXv
ujPxc0q3sPl+GX87gEM2PzZSyqVyvNoFBdNdTAk3zva+DVm5lUNaV5YvqNj1qbEZbw0bKhDNuPVb
zvJAonfa+EA7d2WdcBGPyDwSl+0F9oy6xa9NIlQjv3mJNMSuqEcb8O0to7/K/GQvRnYPzYcw/qMf
89k42aBgKxFYip7f8PNaT9Kqg/G+oBdoEebr1nU03KnoDnWZYg4S69OHeOuFLktXlY5BasvBxMJL
PHkC8uy6NLybmVvf1ZmYkEEm0eggPGntlA1Gxfx/GajN8C8ZiGs6zlzB4tKvyjCLTBjDOgMPRfo5
F8iBaKU6B3QHYdlcYGbdZu5EyForwjvGBRa/vXmJR9qo4qHpXfNJ6eseEr1QjPU6WKX1FYJY0F4i
OS4WfD2xdpG8RBH435UUvwqoHfvc3gCB5A+a7J3v9Z/asrL5g6s4/VorchQRRe4VsmLiXM6Cqi/a
srDQGXsYLCUdSBtPIkGvijEXJAw4uQnPjbo657rKkzmDWtPBgV0MM1Ql5M/LLO4JVHAYk4ECZv0y
Fwpn3elRlY/7e7G/eddh+hcSPf9iOCGU35YsAKthd0QGccCiRl8tO8YaC+QtUrgKS0ERal5oftPH
4bF7gnDjfRXM5ABomg6pcCY4kO30Qkn+JLjBbUXUpfTSvsv1ZC+apglQz4suu7pybRMUoMcIJhjf
0kG3Pkj78XK09N3r3MCfbFCQbTiYDu8MCVUfDiMQ1xNfCKmDB5VZCv8YzjYZjBeWsT7ppi4jUuyk
b4V+wncZR2wKerhrUdY99w79cMKl5PcZYbr6zNB/bGmi77K32s1q5ACTucanqhSfsl6QADBYzIBP
Awe91xOzggE1n1QopUXQS4lUTHZC+CcoIhO46uI6DJ710NFNVJ+ZTtFhCHpPE5YxIthKExiH4R5L
GSAHmxd+pnD2Kq01tdr1V+ySBcNWMXW/hCn3ZXnrcKx4IZ7widPLirnl5JvMI2xqzHcS8T+4u7x4
A0Xy0M9+2fZ/vFEoU+MLSbLBQH2OODuwZt3ZCIp9EiE2WXFgMyF/CvpVCIFhRrxdy4G55ObiVMiS
hb8vxi1Ux5EgQRfE9FV5AsiCnLPb82hUBnwPN2hmZH+UgRPd/01JblYcgjdWVd41cD0lMshgeB4Q
h7+flAzwGboY2/FKnTOvp5Qv6hiZGgtn2BvIxrIUBqi+y4QcfYz/A6stCGhZqQonD0j+kzaMLFz9
91890e7UjgJbNZkD05ZIQR91DxY/a/RPSmfawN3zAXiMl+poaG45YcNj+BCwQ+nd+YrqxGxRC2do
VnkVfCcfYzQpIywP+RuKHbh3PKwI+D2KuLuu4cAR7xnVU7QkriSY+L1BhlxNK+xithZGagWF6lxa
HEqxIVZwmDyfelwvbyUfLEzQBx5fY1k0yncVt6d9bJxUKzjRl69mI9Qb28XCIP6Obz1rVa9vq4cv
fntB4LPpBV02EhQVzOHTqBBlqyLDbJG+d8k9UQEEviCtmI0Y9QXKP7q55WHllLgV4htGbAovQgTP
zaN7UGzIb44GEGDF3K6i3VB857THqpMWQ0YmF8rHc/EEBvuhw3VoPnAyqoprDUtq3H13g9Q8pmAB
StB38US1cwSd8rgAl6Fo6MYoxepmBuV5sKLk467d9xukoNoKvzCyFxZ25b6RRijKQBKptXwsGuNf
EaVhL1nXSfwQv4s1qtV1eam42t+kfiZtLo6lJSzEh1bvY9K1slV+GdOPPoaKccYZu8WvEl2ILaLM
lkzAsz534cv3UoMWLwsXO/rzCa4eOefDTFLV8XQbJBYxaXM161FN3WsK9HIE3/rxDRB3nHWkQwoa
dB/kGy6qq5hnHRThWWOmQasqkZOcnzdCMDN+6T25T5K0jyR5Ze0Rm7BpUJJwLG3E15GeeGDS4z1a
k22TBtEsAJm+k1xicT9olJhPGMzSyPAeItVmrEzH60VUzbRo5iesKHaV4D3NF1cjO8v8CdXyRmi/
cj1/y3y9XtG6S1w4oDvmCXU2x0eauRSWQ8JeUpQGelVxxn0433E/7wlpKLRpYZMrbssBCnoLgiAm
YRmymh9f5+JUrkDy8n0jHDnzSAw13dCIy/T03a8897okyaAlOwiMqh5aHZ9RBnnPQr211cDM0A3l
f+N2FQTKxY93bW885pSBsImiSfFpxiYD+pszPYCz8ySDoxkO+WU1TegAJRWSTp9Uou6knnxbzvar
XbpZlD7RhJTL1QUSdK/Cbp5lfxiB6jfus5PPY8dNF7PoB1KAKXNvYtFfZlwMHiP1SY/f11lSyM58
ViOztpAsbsvMyR6KpDW0NHi7DQNNqxVE0I6DIu6heL3g3/TOyJR1QnS8/jT/K/3RAZtfSNI7j6Ed
g9BM8bEw2TDEa7214Q8hOJIVvqnTZsNIuL5SNnU7/WPKNaw3fL7w9enSEKUDD6UmXKqcUWHgJkRG
1wGqk3mdyUSwKlG4QlIssVSPzaGq90pnRZC6ixu5Gvex9eRfi615BXkdbem+2tft9h7/eaOO2P1l
uzJxYqzd408jtHFPryVPq8kUe6SMlSeKpOfvMRSEa53wDTDQ7iEBJgyFTLmo1kVv+W0kCDyihMeq
u+XTWL45ZkmuQIm6B7PB1C5D1SIDP8/B1JSxRq+6G9Tixq7+iloYSEk6N1RERVR8iOHrQEdcMsmV
3cZuq+GOcq85gAyxkWRjzt0aRKwserpH2NLk9HVE9Sozhbg13abVsoRXvO19xq0cHyGzLlNdTpcw
If1L5Pvty3HLlfx+oZP76Ka3YRCcmfA+bDRd47qt4KcPQ/QCCaGlUEA7d3Jbjs1VKPapwUnJ3nMv
gCJkvqLfIBce5KgFeLFLazCBgLGnukd0722i+N3C5j4JSIKOz7eqy3yf/kQfV+AGEd21jX+xqeH+
cKkI+RBD9VuO/llYAO84FItHMTde8GaKazlxm/uFWJlgk7Kc1mD58mZ/tlEoYW41MCl28QUB+5Z2
6Hq/vf/h4D85v9GUXgo3n/sWpnFzo+sxMG+hr2cLPp5k8sICD2f142od95EovWvR5OxCyoIFxUm3
wVenOxNNrweecJDbB7A/BugFCW0j30gfaTzS04zBXO3VVgHw1/ZsiSzEPfCraqgvcEPpjy92kZqr
wKV+YRiDAod7l4Hp0QdqXPZaucQpGFKvl+hDFjalhzE3gjX9F1ltgXwW9lcDhT9gK9XhJpqS5mYB
lveAhQllh/KWy1W5K/VvlpiMwS9Oiq+otwrMjqqPlkDtYcVtHAPYjoLyVZoebC0w+HIGQ4jXBi5o
ly/yQhIzffehkL80WxhR4eTAH5HIr7hgbOCDLWjgcTQu4oUEmR9AcZKOia1y11YF2crKTj0YndgQ
vkkWkWMVTh8F1BtZAigE+BeWLjueBiQZAI+iEzvXLkl6O+PmZ/bF0aep9oirxHKbKotCJWpl+apk
YUHdxu+GTgdAE2RjQRSs2MtWk1jLzauiVoJPjzBIwOgfruI7f4bVI9+NjqFJt0muhoilFlNSwgeg
0o84lodN8BNLjmLJrQzCYdE8ketG+99k/mqzk9TOMtYSYuwynsGg0ByJ22GjAstKoo9rEuCP4eG4
/8NV2uT1ESDz4cF2L0V1O6B+GrceEo1JVGSDnpCPq6A+9fqCwq1QUhVKC4VFB6wW5DjVzg43YlZQ
1gz1vM5tc+AHiVnjihKcBfwDIc2DzATijPzUSt75dW/ggHqy7YNkhY40VKnI+YbS1B55vI3Fu+Ha
UNcv+xcGKaF6mHwMtHf1O+w2bpG0HDYMZuERzZC9JSuwx5Pf217+0rcYjImHY7hl46Xduw/11EjT
+ktybDqWjuagx2+idpn76Sm/ISniGuuekeBcocdvAIydTbTu4mdJGF8ZiUDTuQ6TYNd7Bm8Rq8pa
u6v4Ccsscrl18lyiWeN4ck0fUOWtPse2xH+CdQuCWwB+yxwMQi5wcqwiOMEcd/QLnYVaFAiAV6r+
hvl2KQO4VGIOJDFq0u5oUj5IiF7gOdwJW5PG1gTVcn1wvSK7MfwI1egf/YUa66omtWV54NmPCXjl
fmxefCTFnqc9imkasXWUGy3WaIwM7BTOM4lXc/Ao3ehCrPNgCONJXYPEXR0/Xe5AN/Zq9aqEyGnl
yw0ohmJWeFWUyUMChL9aYiGeA8ouF3JaUGBkek48unWjmhViFFJO11/z5Fg2ax5x95UH3LKyg9dA
bFwoGZJ8JmOzVhyyFYx81vmc/fidvqZlk/yZy2YmJbSXEYzTveQkNbNKK8dgwiaSkIe9ZHRBGk4n
EaOVlUmaTV0233dgFH+aCMRQzRrcsixhAEvdFszVulk0xb4giKMS1aQivUeccfKZQ5CY3sSfbsxp
u7CUI/Lw8hjtp5VNGX9WPJY5RgztxolnD6eGjwwRQFas+eTud3zpqUOYx+3tVSG9Hg056exVf2gM
P/Z+Vgc9PDTxn9eWmweYubP2fSyPA9sSoPeLVRskTEKYxkv5TSYRTNwOp4XOSWpAJ5E6JzkdAqQ9
dKkUVCeAONyeez1mHaxWEwTfB7Fmed65IdKb1rl9ePTq1wpkDxVUQ3lLPy2I27CD2wf0EjkkUo1u
Zy35t2TgxXtq+vW9vrHpxWmnlrMYs1PcrAV7Gj9ypfmXbDO6KPutfW6ocsxhE7mKQa9sD/YkfFjP
7+fr8qMC4HwughalZfqtfM4pT0XdXOGsTf8UmzdmuUoUar4D0lR+D4EUZVNkcSDL1g2YU1Kgg437
zkxTYzAptSayVFB/Dm7NS+/mLkaYnGMHrkGw47G/0Aw0pkgCoWXcawsmRzCevRcK6BbHinVPX+T9
aBKT749Fvr2l6scme5pTJTdgRWLH3LOzeXSZTSmxH5jhLOU4Mxu1X7/S6a3X+X6++hVtR2ViYy2S
4THgMtPQtxrzf1otLLh7hcHAK6DRkkDgHjn0u9qPRMS/MkytIBgS5TWSqt6v+tdDrHng0b9kfsUj
zVkvKFka3nsl7XDtbDxAjJqiXuJE38yxsWydJ9l2cD97GqJsfQy//UL2VHv3ErE6ZJGvNxIM0QGs
gB6dm1TnFCVpxfYGdzPMlvxSdtMZjnM5QqdKsG78hvREN4jTbOVc9IXnAEfoX7NAm4dyTGCGfGKG
1sWdB3ecJ5P3znDPIxgz3T1U+RX7l5UO3dM2UccCCMSZQ5SlhYnMNmqIFlb960LKORTBxgK/Mfpe
p1Nz/bYult9EHu4RcMsCbkDLswik7tLGpj2X11g3J4KwhALDRPt5nH7d9ge3QIQwGTlqkh3r28kH
iimRWMGBgQlUBJhBBBnjNC6jB+jdwcalquS6D1x+snatDgzN+xfDc7yaIouNF0kZnGrhOTz0gNBD
gzyL2BrXQNVaba+RQVU672yOItj8fFZOu6FSoRFIm8nsNZkw6ReZG29jfDalkUHCPKEeE5StadaH
3MUOYz6wvVI4iu10SCl5kVezWOlVXvSOy3oHp0lXx7B/xC651mMjv8FSIr2Smn2hy/GN1S0XnpEz
Wk7iXptaJyHn123f3LIOpYKmMFIX+Lqa1/BPQFEzGCS3RX+shuEybWLOSND59mryS8Gv29CVzhlz
nhODZlzWBvPnWsqlkkFmV6/vo3dOiltQZIkHy58ZTnCAqtUDKMBC3oJwsSB3S3A0dtNUwHYiZWVp
aTUkaC8fldfcMUA/Z7sNS2U0O3vAEBk9/JiuXy2buOueUnHcz6jo6woV07Fi6BUIUly9J3D6wTWS
L4wI6HxQMQPcCKvO9pNpOMuLdPVk3U4/tF5wAsR4v5VI1+Vop8DJ5VXaubA14j2Ggore0JF6c+Gi
uSIi4LX+giRMikA10XfI6+tUWNffyauiWVkdOUWXijR23FNkfFLBLW/pVM4YGumRs1+Dpb0wY4j6
JPNqQE9199sCJWNc1kEPB7asl2CplK4s+C1S/YQp/8G9KTjCPtcbWxbPmYMwswNHEDs23SvLgNsC
yO0nrsg0VKiSXjEfsJUA6ljqyq9oapkuJqc7FkoZvn/x3Uw5pa58wWJTm9ZK6GHG0gFXmfC0gjaL
IwBhaaMLKFFfA8po4uCKwogmoBD5MY0Db7xOGUWiBqkWJ2dIT5GKMD5CCkN1aFDXHbW7p6xLw+rS
DDl+P9Si5ZgevCejUAIa9JXPH2rgMGSPdVxg34q+haJsBf/+hu2Oec5sk4pPGRDdA8QpeAsmJ63C
IWNMJdr+1X6qmKAAj9/zDm1GaUJbGJ72afEtN11fkmddSE2WC6rK0EB/Y6k/Z9Wb/owgkqBVJYgq
uehwcg4+Rn3/W8wpnBXdnSpI5KZdQxGbfVuyl55EthN5bwd5RXVfSlxK2iEi5yXVmghjcaAvjI9s
l/sWzfbOdQGeYV3Bi/8SZnLA5MvImQHW4kYGtzPGFarPzm5Gno+bswijBqw+RA0v8vR3zBOsSe7T
4KZ9QNLvxgDdOXreKKVg9z471jtjuK9uCDzlW8u2gP2jop74gASfdGkqhaFzKIsZVLqP3HmhQHU6
U5eGFBWyys1B0seCuoTRW6mqj5uI6vY5ibpIYhZPWoVEPFH6sV+M23knUnt/C1Nh41LUmu9iWj5K
8V0CQmXwp+f1XyLJ+v1i9D1a/F0J7ub+jBgzSnBuX0Q9VvsoeTj1/9ua1rOgubGofUzPpgdx+nd6
Oo+eXTtuFTabeNWyX5yX4WBSq6+EytSWTLkHpkakIPHoxNRTwOSWwkncF72eL52G9e5yHomY0U0r
zTYgPBHKQQuDyVdtYrxlpIT+ThvhK/7B484zwym8nRKGOW5HKz307gT8pvp98IHCwdbB/BV1vfJ1
0d/tUOyZEIvlPSsqXHuITOlIqXgSWo4aL4P+ZcDHICwu53DfJka8LPMp0TjmxCBDgg9w8+e6gm57
4NixqIDPh7k1fliHJ2xgz614mLZ1d23u7IVRxAVUOzJ1IDROHNI2Jax14p7lE8EQ5GuByE5RW0ZY
Vdj6dFlz8G1uCR9Zvvk4LWVdnSQMdMxYAqPCxJpZB90OAfTnb9izmljh7joZdgeGl21LS3VDFGPc
+Bde5mzsuHMOywHg20Ng/7U5RNYtjVRoCsz/1DNlSkWAAOfK/cm0xOxx8+w6eOQU+3jgWM5JJXmw
/I/oIuGZm+qX/r+dzN1hlrN7LgLH3e8ppxEoXB5kWuTUGBJBPF+8sFaHHiLUuoukov0q1C7HfI+/
q/f3oyGB+CMgyNsuxoJYgwoxXw2L0w3FMLMkp3yDVtT7nxPEHwpSZVlKntlIRaKOy0ukg5EavMS9
d+KlflC9cSlHNJ1R9kaRODcb7JYYljMFQ2zcyRfBR4uA8e9bZOYyb/2m/JGkbLThupGnCnNqs02f
5UGquQ0HYtAvqmbhSAU3kqUd/2lmMFRuvDv+8pzPASRv3haG3/4hzXffHFN46zPjAkZPGYGEAyH1
JIEpDHCBcVtGQzMZok5cb/IVkrssorggbaZrpo31sm9xSSuPe7yAZHRYzYz2Jg94L80wo3UE5gVX
3HnfOCalNvhq3n7LFPbnmRjSVIRrE5+/VjcX3DBIBLbj1l/XTotoKS/Sn7cEDhFeHmtYLFdLDmK8
cMYi2i8RQFp+P0ryllNXDs2khpNoP8VZiX9vNL9pWj9SygKs0kCH8/J2VAnN4AIV8zX3u79D7R6x
JICtT74GCXy8m0IMX6yHZhLeU4KAymepI37EEcVlXJvjKWaWLYtuCzcRyNIq7HRrMJLvQJuKEjQa
/ijfEPKeMmbtcnfBcC5RlmRA6vHLbD+juasn/UPCBY+Na7Gv4cnL+LP/4hqyvAcOPzXBD3rTAVrq
TULdWRdt9gB6A9G+xLgsxNttRObJpRA2+HES6951gN4t2kRV/UEoOUAgssAde4L1ZOSBk31giLN7
zByAbgGJK2KpN1us9XY/6rr5fd4cieKEJIjzzL714fDoq14cSvDk8xTe+UMzLm4QOgo35fDGgxVj
KiJIbnaCpLJ+c62UDpL2TUj5/GUfvJwEs58+0ZMtPV8tfIKw3hBKX85yupB3FIrU3eQSF7qw1kTh
tiTk3vVlhdW/KCSxDq/irMBhKXYPG5S968HoyxM6vYI5hKbDMomdlUPzYvFccCR3Q9uUh+05DliM
gM2MpFhgBRn/EEqatDtzchgnzJYgQ8uB8YqJZVD5F0gdz8cI1Vyg388Sx/g2h4njjIdF2sSpHwOE
sBvFTI+0xVWB2pYn7PptPfu8BCj/HrrNPo+5udi4kCt6ydthH58+pucH8teRGXEo+IWPeX2kba3z
umOALEaPQ1jhdj+52nQofSgxONi1Hq9Gwgo+32SWRrb6n4rpCDpkNPNjPwoQVaqGywyEqtEnqOSE
pQR/j+HQnojsLsH7ZdTiXsG/gY3SnPQTSuO9taLKqENF3xfiyXaWsekiFX3UD1LB2SwvLBh+x/OV
uAmZ5g5qDoOZJpaxmQUgOEiRd7qKZn3ga6+WV1+iHX58pr7y2mjT4bt8Q0JXul96fJK/Srz/SL0h
Osoj2AlQoHUW4gdC9KfrZp8LDwrMrYFLWIVoe1lVpUUEi4JD/NXCUJ6/0oQCES10L8hMHUp11d8g
yfXMxQOiLDRLMvePNi1FegctxgTY0oh4Q/yamVzaumNt1ktI5KI=
`protect end_protected
