��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki��Ы�T�����Ǐu������D���u4��`u��Z�(g�Ü�q3~�1�f6y~�!X��-�f\>��s�;��Y[d� �FXi�kD���jz�$?��>�����%�O�>���q8�͎��n>z�0=z*�g�4!��CaW�ͧ�d]���pb܎�DqY����D
_���m��h�I#��iI��+��q*�DN��5�&�f�TZW\z��6��O9��Ϡ��|/1s�*5!�\G�����9���1�I<�k�q����d�LV����τQZWm��IZ��tSYmdm�Z7�&:�p�A�TQ�U��k���l�Fb��N^��P��t�D�ÞU�d�M���	���#���5�,#A���y���2��I�1�4/�,M�U�~���<K���I���u�
�a:�u���|X�*VP
x}\F��Lw]X������Wˋ]�PTA������a?*�L�NB|- U�?�6��&�<�U^�0��10�t7x��b�(D�OWjs�L�]K��*Q��-ߛ���ᰉ�9�k�N8-�mv��ko��H�@ ϳ�C��Wm
�sq�K�>�u!�L����2�*(��<�Y��VH�9��<p� m&����$�b�u'��X�l��B��$�/�_2�)�"��ظ5s.X��ʮ܎O���4_�Rg���]+U�a�������j1�r�uԲ�y����~��Y䓲�н����U?q��;���/�\�+2\�����4跳�y���!�*Ѡjp��,�\*��i~+0����qtj�Δ �2&�Z�^~�������Ŏ��2�د��9y�4�ї���&���Ț���6���V�fY�U�����I諓G�w.��͔'��@$�$;?��v���1M�*A��j-ܩ�l��$d���^�P�Qs�� �p���.y?���uI��W&5i�!�>�y�
8;�&b+bކC�v o{b���9�Xw���Zg���$���z���k����?��6�a��s�l;�Qȃ�t`��t#�v�d�XP�
Ա�L��h(�M�5��3(����5~ung���ѕ�S8tU�o\��R�i�x�b�D��]���,RkMZ��&�W%��hn�3�.���5� ر����\QOժ�s���d�K��N���o�q?^�(,M&w����b��B0�[���ԫBb'�K�6�XD�&-���x���)�6����rNyY	���2J�U�.҅헁��` d����}�\�I�{���4�C.�H���ц�����98r�`H����Z�p��%G������j���MO$�
a���*����.�0�s�b�0�DF�0;L�2+�P5	mw��+�ȩ1�L`��f�d��ؒ��~���6r��x3/l1��#e���FZ�)�Ի�gQ������_��1t.u��� �\F,x­�.G:;������W@�H�<�[D�"���w�;F��6y#q�I�~�E�I�������4ҷ�-��oIj�y��r!fFB X��I���M��Ƈ��C����TD���:6��E.�n7�nLz�M?��Ⱦ?v��a���8��|����"g�׏L�c����<X,�)^�x���n���
�}c$�d�*8��ld/� [ �v�E!�MAy��Z�5��,��O��Z
��-=�>��L��Sի��)�/Z���>]��7�U�ŀ|'	�-�#�m���C�hP,�*�X������c���da5�[��,b�Ct\p���цI��If���c���|�g=�s_���m
}��Ű�I��vW��s<��7�U~B=��جB���������V;�)�!7yT�iₑ��޾Ev��R�[�3	��%�FO3aap/�}S�,�r�g���m��=N2{�[,�i��Cɓ��'u���3�K��M�q�J9����	��ԥ��P)�)y���Tn#��='��[�Rp4I��L��.�E�fP[���~Pe��p�e��2?}��0E��MC��lY���&=?���T�Xc\Հޞ�Q�'�1��BH	���Pt �~������6�6�m2���BR�94�C�Mؠ+�d��<1�m��R�ƺ�F.�x�Z2mK�� X�v]*��:+ � 6<������	��"�B2)Zf��77�נ��������	s�)�In���F�5����hF�� O�Js/�A\�0e�QܤG�Ԣ��"TP�~�D2n��W�G�d.�hƟ��܎X�����\%�B��O^�Qc\8b�5��Fzȏ��,��0�[.1�ϼ��#�9�W�~�]A'rǑ��"���V+-dٴ�qA�E첐a�ϫ���ZI^חI��S(�.GV@~�"A��U�z��cٽ!��1��R����kآ�ViO`=�Q��<���;�l��4�_��"$�#5~u�-u�  �:h�{���H�2�4$��h1{�� �=u�RVZ}ʅ<w���o9� ;�j�1�a{���I�PF���B(��n���Q^L�����O̸�a�#��WqO^��փ	�Q6-'7Ŝʹi�X�%��v=`�����!��:����-ﲹ�u%$��/��4��V2턥�H���+�aF�3Zr~���(�,{�y�L���̾x*9�֨�����b��&�����9��֖��'�%pۃ�><So�@�������~�_����Hn�k�O��lR��o�EӴ��#���`k3�i��.���:���e�Sх��Ub�VzԚf$7�;XVH<���1,/��ע��������y��/r|�P�D.c
��p�cW���3j��QľM�'��x���E��K�k�dk�`۠b����g�����2$(��h;tg�
+؈�_-���2,!�X$d�>s�<f!�IA̫���ǵX�6���31��IAz�p�������	�KC������S�'(�"K���p���Lҋ5߆n6�K-�:�ee� ����e�����q��1��^8�n�%���;94�fΉ^��j|p�#�AR�����f��6��1d30�r���K`b�H��,
��	=\�.�J��t��̋�?N����p{��K��@�'u����8�<ɛ��A08���gt)�����K����{�zW{p�}J�}�y	�΄#�ɕtS����P}@����0O��y�Y�`�
��Û5���	�`U���exC:��c�
D��VPcÚw?��+�L>���hR

.���h�ڦz��J���tE�u�G�����aR�㏘lK�@Y几�o����R�G�A��N�t>�d1J=���&�k�h����Mm�>Ժ��n=G�����fNnv����t[ϣ#li�0���F7��pv�o��P�[~�ӧ�C)y�7�e�����$3�>��b����R\�Co��d�H��1 �XWQ�6)D.I�����ax�7���U�m WO߅n:>�LTf/�G�U��5ڼ��1��d)Rc~6\t 3��ZI昆�>)x���kئ��� �]�������������XREP��d����2NA���B-�Q�����pL�l�����	H��0�����y��c�V�u�R�I��ٷy����.V�����4��C�TxЮ�E)��(����F�7+�q�<����/X;n��DZ_�YNuHF(2�ʥë�S��uH�Ԛ6�������t%���8t�X.�˚b�ݕ�����y��?�����m��54�e$��>���-k?��^}N
Ev��&��Է�,n!Ԣ���ε�����0���֌�G��QƱUG/��m��)��In�p/M�29im�_
o�ͷ�-�[B��\��sRi"J*����VM��]=^�2MR�:0�Ll����\2�����Pp�!@,�^iw®��+S������b7t�2�a9'1���ME���"<�����c
�7�H
n�0��*E+��\Fr]�k�!��^��n5�&b����o´�Mc���M����y�������˺}-���l`��7�����0=�L����S�����2t7{[9�3#�j�.V�a�8���s�{�l�U�}�+u*��[����\��b$z���1��x����8�ZU�����	<5���JV�O�d��9&u1RR���@�F�����Q����;�:@��p�[�R��%��QF��G#�`i��j�3b%�*Q ���S�+�1��q�C-�:_���-����ty���R���$[S�`�[D� .M�h�<VD
+T(��im�o�W�Q����)�;�)�Q�zc
��+��RJ͖XH��#�희�.Y��� �,�<-N,�È�oRQmƹ����v8f7���=�[C���K�p}w��[�Ϫ���<K���Y4ƓQp6O��2�?����t��$�%y�㱖�-����f��r�5gG/')����ѯ6�;`������i�"}����[�_dcq��{�p��TTZ��;��+�G{�۩ow����{gG@�����+�6���]Qז��p:��
f>5�ٲD���H�_�E����h��Ξz�]t���iX��L��ٙ���� ��|�&3��n�K��T��"e�層��� �o�1m�ve�^؍ s:м)�e;�C�%"����dL�[ R�/JŬ�`���4b���G�ӏ�un1'���]#jD�x�B�u-U�Rq�v�V� H�oŇ�G ����y�~̵�8'3{�
M�1iP]���,p� ڣ5�^�LկƙM�� �9y���Ll��
`�E�YMYH!���9N,������ <`��}EjC3��9߷m�ⵁ�fbx�.���i)����ӏ�G�M���b@ejZ*-�](|#Hb��ݰF�^�4=%EJř�zD�+�������	K��|F�]IZ��֦�L�j�!�X���a�^� R �wD}.�`�h�L�vn��N �P�#���[b�����j"}����Q���1(�{~F��3�6�3'B�ҡ��]��9*�{w�U\,�X����q~�`x��%��-:����n�<&_?Mt��ٯ��3��$>՟r����&����5Oc̣�^�g�pp�b`(I�kMƌ���Z��C4��9L!�|���^cs ���"tcA������,-
������q�j���t��q���Z9HC�ü*�K4V���q$�Ҝ7�b	g��1��0�d�ͭf<��5�S�Z�T	�b��2kxE���U>�&m�KJ���l"�B�U��@���f8wr�����Mm�羧�/�sߙ��r=?9�v��djX��`�XЦ�m��-� �����&R�L�����>����N�LUq3x��Ts�㹃�0�(��V�����E�x�C�Cz�����!g[pZ<
���&�d�>����Obj��b/��{�J1H��&|�o�]��݉'�J��Z>�3|Q�A�6�迒���.=�S�pF"/�yЎ޼5*ţ^�=X�:;�K��u�����e�x�<G�t�&[��iM��z'l�\��ʅ�M��o���&o���͛��n������8Rb�e2G�����7Ֆ�^�>��j�[:���p n�<�e��4qD�L��`0�\�߬T
c��Q��d��&�B��|of�嘛���"�n��V���Puc�4f�)��R`�n^o�
P&#u��6�K8���9g���Akta����B^�H�0nδ�]��Oj����K��G�፳ ���B��6$ȶ�cDǫҐ�4�ŘmI��/���R��\d�Eۓ�8$���pa4��}dr�bb��(��Ƅײ	B?��+���.`*��j�F�b��ꃿA��g�5e.$���z��+[<x�1\�̭M����4�d��D�U� ��l�a���+Z"M"�:QNw�d�f�fYy6Nu,@��ME�@Y��w��W�+�p�����y�V� :|���q��jg2q��U���$�U�7!���9+4W��1${��=�B�9�R�`�ڃ�u�&���,m�/+Wٵ#�N�G��1+�D~K���8L땎��u�G�Ǆ.�S>�.N)�d��ќ2���E�m5W�N�]�
vh���
$�3��"V���+|��I1>I��ͣ.���Vތ7���4z7H;�����#���L^�?�'��*.��	_T����]�^|C��zs����
�i�Fb�v�j^�6������0��aR���v�b@���v0�%P�5�K���`�Wn�S��%�Z�\���{}i��Խ��@�.A�K��IҐ��=Π3G�t��|���3���9c����'�%ĿW)9���u=��/��kS�M��II9k�!�e�JL' :)��@�O���P2@��x;V���2�kN��3n�Q��
W�F�F�/ز������~j�\g�k�%���Ӓk��$��&��'��}Ф�V��`T��6n��,�W����1�A��A?�r������gR#|��%���r��8e��\��+?w>���w}}�<�ܪeaݽ̏��yYк�5qg[�?�vP���{�}�ʔZNt�V���u��5�ZM�C$������|����0;�+G����]yT��l��)��<u�6�Z���[�hSY���Ƭ��k�#����e�2���n��!�ໜ��_t��E������uFOsν�b���U��d�,�p�.9��O:���&��?�fS��t<�n� :P��t�1{��B	���V�*3/tׄ	(���'l���CK�OQR ���X��R�����OQ�d�N&K�ּ��O!��f$��f �~
�����L&\�$P��k9hP�/1Z�L�Ͻ~��Q��G% uz���Җ�A:Ma���2o�х�'{{t@����rr�5U�68�a'�kkO��dz�x2w�y�$J��'�9 .0����eh��2iO��:�T������$��n-`\s��
�E�?�٬,'ˠ�䬠�r�ۭ���i@+U� t���i ��my��c�y����x�q_7F4h����o2��'nc�ks ���X���U�h�YA��'�<49���e��e���+xc���n`�{c������x���q[q�o�
G���z	A�_�
ER�ǳR*�Þ���Z�5`ɏ��J���n��Wm�Fl17�8��ވb��7�c� �������/��s�\�\ �8!���O]�1�̥�k�T�r�8�q���Z��|�u�[.��o,�xg��7��&v�|��$?e�-�������>��;�>9��D��9���;7���D���.!��	I��B��b�y��|�b�^*�l��\i��S6O3V�<~�Ю�.�bA,��?�YIT�^��?���7:gI nz�-�	��[i��Rd޹?�V,Y�	��N<�!f��v?	��A���t�M�ҝ����pU�^�` �>�<�G�nfr�Ҫ�],-a��f>�R�K��kHO�����m��gA��kE]�X��
͐w��m��_L�V��#��Uy	��1�0���A՗�,�����(���Kc`i�k��I��L�2O��KQ+[K�*Z�c:��d�6 {n�uK��@>7yq���Qž��%�@5@�3e(Aa��R35I�,y�k�!<I���$=��| *?u�����)�L�T�g�Z�Bf�T���,�*$��X�;q>ua��~%��/��!ڟ�lӻO���952�q���l�`4ߙ���֢k�`�׻̾���sC~pXO�D6�؟#�1��O�Nkqs�K�c�Dوeԇ��0���3��Z���mH��dv��Q������W��;uU.�b�j�T9)��X@�C2�&jbi�}�� 섨�����M�U��S����1��}��!v����GPɵn�M��=��Ex�?\)���?��F �U�������T���1QpOf�����s�B�O�f�[;PL��6}
��AnF�ZZpM�f+���	alf��Byt��A���9�@gq)��j����C��v�{�x^Dp�9�S��'�X���v��}�?ʙ?eo97p2f�N3r���sDDi�0�<}NP��߰�0��,��c�wk���x?9����;Xl���+T��^�x?�k1n.�a|z�a��YbW���x��Dglv�:�հ̺Y�d�2�9ks��n] 	�4��9"�y�������o�tKs��^�~ʬ�AY���	+tD3@��Z'�Z���J�~)dYڨ�2Xjom4C��Cлw�n��B�7�a�ٺ��j:��/D�3���PA��N��xu��.>)�<��I���aOTZ��]� 7����	���a �ﮏ��W��C��&h%SQ��A22z�XG�g���<�
�".�;�oaGL�E��M�k��.����p�!p������j���5�_w�xL�c����Q������1ɗ�r⅏��+��$�x���bҢ&��s�l�^����|����l_o�u}ePbP��s�7̕���*�t�L	�I���|��NX͐���,{�� +$.��h&�w��;������e�ǜ� ��|\�9��h��B>�p�U�/�,�0���(A���\�w���
�R��oj�l<�({��I|C����F𔩪E�;��^����nJ㣊3΍$�ɼ ��/Ӄp��+�w���20�*���Ƨ�]V
����#y\�)��N8]���-+"����A@:`j�2���&�	�1@����%w�2wֶ�gT�Ȳ:�-�+��`�����@[tg��,�Aߓ^_f�Ok�,oJ֍�W�R!����<{S����::*ft���bHH����ȉ#&��)�����'Uy�S�/�&x�hN�(b����
���p+u
�XZ����_'S�B4Hzc�D{ ��7!�h���}�;Z�]
\����Wlnn	`�v��cϲ��5�2��ƽ"�ИZ�X^umH���5�����	���:V-��
��f|��34C3\Oz/��27��I�A_�O����M��ʃ#^3���K�!2<�7�Tm+'1��e2�,�L�κBnÁ�;=O��
-��ï��g�J7�`fR�U�ׄ�o�.[ zJu���N�\2}ЗMЫ�$)�܊��8q�[��߿u�Qq�y�<�{0��pl���y���Hps˿���7����������r L]/�n�*�"9��L������ǷNT}O<+��߼_5��CW������&��6r�?���q=@���[�f��;��u����_����n�NH����[�A��Lܰ~*~��v�rB��$o(�4B3J�3�� ��qE�!���r�������g��V��������IBy��m�L{�'�[����g��Sw�����Ԕ�Q?�_���EHΉ�)ϣ��oI�F��`+ʑԯ����t��ZѸ�47����'��8{�`#+wj�z̬����T�o��8������a<�7l�>�6�@�嬘E�9䂉@�ef����06$���
{��(C 5&���m�*�
)�)����Z痴W����z��>��R��Zf�ۭˊ���Ɛ�!�E���3e�vڨ�d?K�P�Om�4�w'��8�F������@�L����wW�d��|�����<�~���FEC�9;5�0!O���GЏ��#�G�h�q�lc�x�cm�Ŭ����mLZ�|2�5L���������$���f0{��X��)PS���q<Ϸ���˄[9�#�86��K�����E�6?�	�'�x��/J9�����ۖ>���+��fhPf��Y���F��Qh+K��%�v SfT�b����M��V�w��Z��7���}N�H��e�#��\�m�zcH~3nC�%PjH�1�n-�O�z��-Iq��[m�jCc�R�����קӲ���©���5��l��=�l��F� o�d�F,�f��G��Wǈ�"=�c����/[I�bs�BX�����#=%@��.�_f��S6�o���e�Z~�+ #�az�a�2
D��N��'Lt�����e��&U��m\.=�9\3k�K�);.��L���M���zQ#F<�<�Q�{sK��NL�!����!1�+�Axq�J��=��q���2��*!��qn]�gr�>���u?裑��[�_���}W�'�����,i��ݨԺ�d����&��Y)W�J�LB��e�gBםhŞ�'�>qW�>�k������?�����ʙ�:�z\n	ZWZ�J¬X����)�q2Y�qS"�����jTJ���$��F��`�)x�����8�/X�R���i�+�s�֧5��y7��E��<�>p����y�y�Rwnz���D�WI0t���\�W�Ԏ;5�>��DoS � �s,| �;Ư������h����!�5�{V��s磯GB�����Nc;�^j���tC��xo�&{�w=�q�83��*6^ ��|,CC5��{^�S!�!��;u�����{��X��#'�(�c2�yx.-�^)�Kɫ1.�i⊒���l|�� {�B̡��OMQ{/yb*#�:#فZu=��w��n\�޺���Ae�J�!��GwW�^>,VeeZҷ��/<o��S�V�K����� XGJp�˚�9�k~72�O@�ӑ�Z�BI"��	�#�CY�8���{�$O��a	���Sze��l�Y˶P������f
�����^�K\�Br6���N���V��Hw��if�́V�[:ߙ�,٣Qb5r�ke�ߡ���u����s�&���q��&�F5sO���r��8�\����)���Oߧ	в��	�O^j�
�0�s�
�M�V�Nuh/�O�^�d��� u˄5|�z~��PС���f���>����1td�� ����H�%n��ך�T��Ȁ����{k�nZ�����Uj���[��� :�� G��,V�H��U��Ą���X��ڌ��4�A�a列.PT���R=NY��������@���l�/����
]���u���6t���	4�C�y=��l��{��f�zXs�ڴ�р����������Qx�fcD�����>���[�X��"�����Z��	���<h��Ig���]G�
���J�QS�*�!<���g��Iw? `�#W�	�ɉe5��QtJ�ۯu͠"��A�ށ���Tb�Oi���cKy�%P�~�u_b&y�G���%��$�[/�����8�'v�� �7��q�r ��6W �����fqM�#�����ӯ��G(����W�d~��ВJ�����}�{5���0(+�#�p�3GQ��!��W�{�)�H�o��r.�S���%�xϷf�ʺ�r�ZeA�'Y�[j�����'j��*���+_kp�1���j�R+��cɪd5yȒ����x�Y��2IGY���v!���Hj~D6Hx��4t�IcL��<��w�xR�x#�M8 �51}H��ir�L�Ջ��7e�U܆��j��~	�|��j L�B5+�����dd�jJ;J[�5�[��9G�=/"���͊���e��-kM�k�z67SQ<���'xU��WB���H`������3R-W��<=���REI̷�S�'nǐWZ�����(ǰ����&�u~�������CF�"�md�T�8;��YK��C��Ю���D�E�����o;`��(ɱB��{�����z5�l�Gh�ˎ'T�cޗ���P��E���tY��6#�>�IH]!�o���ڽ�S����v|x%'~���^�LA���J�VT��-U�	�G9G��h�`��g�,��/�6�����!�
5�Ccxi�I�0L���I���A�ЩڞF��F�+Gq��'����I�;�$�.
HC�ʱY���Ju�脌W�[A����iS~��)���5��BZ�j���,GkN��r�Sa�<���L��U�>6�?�'�0(�>��hJ'��%�1�d��|J�v�\��3���=}nGc!9'm���_���[�o�.�����Q}_JF+�e�5�U�f��rY|��R�d���3%��b�a�o%�b~T�����	W����@h_+������I��qA.u'RMa፡HN�Dʣ���l29%k��WI���Ҟ����e�d�!��oX��9�xK(�+�Q�y,6��N����+J��k:��V.~���ɪj���{�|m��r��d\����џ�̒�c�sC1=k����ѽ;�C!�3�7�UʳWm�O�e }�ڔ�4�YC�i����E��Z�FP��E�lu�j�_60�V����ݑ�ۨ1�����nNKc��6���*�b�<��Bb����<^r��H��5�s�zM�Q^�Rf�焖�V���9X�BUwFKM�
L�k���:�������螭S�M��~�?I�LI�tM"-"�]��I�j+�ҏτ��{e��"�����&aB�~��x�T�|��b�~���ڻ�x���X�Hڝ�A�"��*\ʤ8��.�M0���~�6褦?-Ŕ�5p��RDl�DZ�i�I�|Z��&�|�'7��K��sb��eռܒ���c��q��҃\���F�.�U�|'�w��pf����g��򰵣����#K�l�n���Q��]�&�2U�I�!��<�x���~���5!�|�Sǩb CP˧x�(&��dy�������K�_�#mQ�{`���0����G��e�|X�}$�>�r����*��p�Jq�`{����9�֪��oa��������9����$
�E4�\��s [�ͽ�c9?)���p�_{tLWFt�E׼�>�J�o��d�	d�l��*���j>�t"K���#D�](0w����m��5`Sݺ�$��w9�{�l��كk����J&����!b��̙V�i��M�J�T,Jֆy��CZ!5�fb?m�8�AF7L߈̶U.s����=�]���$�*C
�gE[�h7�:G��Ђ/T�.�j&�seU`�j�e�*ߛNt����5s�nqYT\��M�22��;f(�X��N=_<+Z#�ЎD�d�aW^��b�Xd>��i;��[��5�4T��(G'r���H�de��$%D�3�?��������q	�Ѯy沨	�"�ԱMe���e�a��K1x9Z�6~Cr��,��J���3yz�T�F�w��=���?��%%0Â_K!��Aq�q�[4j�v#T��\^�e�ʔ�D���+�}���ax��1��	���y��^�/"��
���=��ag�_f`%No�����ݣ�~Ð6��#꧖�}<�ʦ�wN!�߶isYŏYJB���F-�&03��%z��(/s	���\�O�Ze�wB��t�:�ղ
4�xX!m9X��k��[�Ԋ��?cN��*��dN���g�P�>!(�n�/�����L-3����l��W�L��5�`11�R��x���X�ƥ�źQΎ!M:܈�{�/��Sꮌ��dL	���Z��q�&^��g�$j�P�03;���MM�
3�ͧ�
�������w�w��𫲳ϛ����7{�#84�[MMٙ�_�>
��x�N���r�щ'��'��"��$ˬ碸6��< Ąs@��TJ�!E�Γ5#�õ{T�N3��Q�.�6�>���K^p9X�j��9$9�
R�7(Ϳ�ŉ�����H0��JP(�4�����'�lv�E���H�I���ɡ�ͼQ=p/�-y�;0�b�D8fƉ5�N���J6�:�lȒ�?f;�3��Y�zRl@��%�dU�s���?�廴6�n��b�ݖ��V�y��#,.g�8�5��g�����"a�>��������ni�4>*�ē�\�*W�O�9��L�^Ԏ���ʙ��4PrC�s�~y��`�������r� ӠJ�L2S�/��-=H6&;�Qa���P��t��$�:��4,Ҵ퇎2m�5�������P��I�Ϯ�Jƾ��"�щ�wa���R�59�4՟>������?9{,>E�>%�o>����WN��f�y����!D[9q�3-��N��9�{`��b�l�k�]�waM��k��Z!��Ԁ��a������c��U��'{���:h;�t���Y��?�*ņ�HhV�Cmw���~� j)��&��p�᠂�L��N���:vÇ������$���M�V� .��K�X=�(������6u��_��&㜝=ES�s��g���F��$�l���ٟ�)�EqU*	���z�Z]0xG��;s\�;�Z7��X&����Ӎd�
x;��0�b�u�a[j#��R:�Y}o>C�).���1}��w7��0�B���6J&���O�ˊ�C�c�N�샺��Z	�[.��-�Hۡ���/�dڡ�e=_?X�	H��}8�G�tUBNѯ�Nbq��=�R�|�q�<udˢ�%q����E[UYyWG4dr��Gqi�MU�M��;{�Х�4�M?�k �`�->�-�E�����T������9E�H s����;�pT�y �����ᢐ��T�䫢-������S���gh-&w�=pG��2&��5�-���wJ���.v���'ۄ��c��xz�O�{��{J��� 8��j�
v"s��O)�u�������Sa~���"'m��t���̨��j�U��|�5.��6��'Je�U�����｟�i��kX�
۳�y\3p�����9"ȍ֋�G���w�Cޠpg;G��MǶ��0|����������MΡ�� ׀d����;���lY��]���I�/1���~o�M^K���W�j(6����}���r/~��1�)����DO�	7+2����zv�`�s�{ʤ��C&�	����{γ����?B�l]n���;XG����5CM���4�tC�=�/xv�0�p�~_J���@�G�9ʅd6R�:[�@�71�s,BrC^��o���k%$�^�/˪A6d!w[:�|v�S�?8����D�"��p�@1�#K����������_w����s�!r�1z ��pq����Ja�h�� �����R6Ŀ�[��]�4p�.>�1)8R�TY�ݻ-�yU�b�qjMk.!D�OĹ��1uB�4�������P;|d��RM��1�Ք�K�~҄j� "O8����������
�j���P�
�F����V7��h�	�3�q��ף�Bj�ŷ�{�qgcS�T�G����@�(4�t�Ή�:C�Y,p;�̚��l_��B� ��6�p�>���J}j�.��c8$7�@c
,����Pe���0,b�D�m���ؘ��iʢX9>��ĉ˴M��z��:�K�)�`���\tu��o���4�����T��!.1��/���{������|!�f�:"W	��u߬��'�օW���.Q&��GtmDl*��*�CJz����b��R�r���m|W0_�b-�2R���Y\�ۖ
[(���G��J :�y'��q �(k�#��8��&Fo�0�<�yKO����iNL�Er�(�p����
Cp/0��������2�
Ⱥn׏��m����%�� ����ZX��e5�����^饬�3Ŧ�BW��3X♫������Z��=��mnܫ{D�DC�$mR�0U�����J�x�o�a135N�����U�2����-����� �V��`��:��(��#�7U;t1@��X�L����
A.�>g��Qd.���Ùf��Rc� I_���$����oH<7�JJF��EjъG��<��j�@(_��ə�p�})CiW����ݝ,��ư�۠�S$��m�|*~FFc������!�*� J�D�X_����75}~Q���~t���_��^���߽��g
C�ƽ����MV��I�c(=m,��������Y�+�x�B�Mc�lؓ,��/k|m�OL~�+�O��)��,Hs�	�h� ��BF���.�`&#Z̙zgι�����9<�	��{���a�g&P��߁�X�ЮC�0���/�́���<�Cn�6"J�(5,���:�b�:ٯ�
%d�P`:?�!��?��i��[����ҙor����
���H�(T��7`�J�QB�Pwq(�7�q��q<����������ٍ�������+|6Y;��&QX���~��
$ڶ_��A�ыnhH���lv��w�'NoRWi0�z���w9+Z��q�Mf���r�䊟�<�d� �ʹ���?t�Fϣc�˩�=���b���P~��%�L���`t�G�H���]O<�W�Z�Wm9�&hM;C��P�Yi��N����%�Eh�LcQ7Ob��#�'�R�.m�,Y�2�}Ԋ�  ��������_�l��@�� Fɱ�ػ�:r��j�22V|9 /$���9�m�*Fܩ>�)���PB�+��c�5�BGd���Gő��1���?����?ldЯ�˅��PE�ñ��10����a<p
��T��>���N�`����T�^�S�P��0�]�;j���/r�m2������������y>M"�[�;�}������|����Z�KE�;~T�|>��b�a�\S�xY�o:���i�hdȨ���@���c��{t;۬n�u���naҫ�<������p�w�Sɫ�8�d^t8��#�#�`�<)^V!��m�L>�Z�J0�B� 1���:��ؠ��ǘ%�������HBۄA�i!P_����`;"���}Q.̤�S(�~/]��~2Q�|%Q�ۂޜ�����f._X`並�Ԇ��L��M���/Y}6�NԨ���U��fu��ڰ �	-"5di�yu2��� cMvc�\xC�f�c/�� �`>{�D�x���z@LA�L���%L�� CJ8�j����ې��댋'm��ƙ�v�z������\ 0|�f5�p��Υ+�1�Hp$���t�����X��6��@�K-��ҟ������_��v�g>�Kj�v��r�P�#�PF�����)8�k����g�
B���ʾ���x{�<
�8)����v�1�Yz�V�;SMw�x��LUTpg��ژ
/�sy���X��4H!�7Yn$���4�Ѫ�~>bA���ǰ"� �2�P=g�3���/uf�*��M�����p��Y�$}O���(�̅��3�s%��aw�{�˙���EH��
U�}z���nkb�闲0�i�E�P_-�s��'�\���'J�
�v�8��.F�R~�z۞o���>x�p�L78�?��;���Q��*5�)4K��X��&7t�5s�k2
� ���QJ�J2$�|�M%�L|��=#���6��7�Y�9����Ub�0���ڃ�hjai�n�$U�M�W⋐	Y0���=|#� ���w�0Y%l��M���>6x5+�;5[iI~]���� D)WwA}S�qM���:���u��$C�
��5Ex�W�1����.[��/�Jw�m�͔[��/�>H^�@������ʂ0T~�x���wh�\�i��w�����2X�!j�e�&���e!.�#�u]��Œ$�ZW��r�b���Y��&j�7�SX��7�g���Ô��Q5�W�un��6[�������� �H�j=��S�,æ��(zD᰼]�	����%��K�Sn����ګa2r�P�l��w�ŧ��ٝPB؟ ����4��r�2U/S��y\V�՞u�0�۲Z-~B#��W@僣�p�2��{�B(�ˎ8���F�H(ZJ��SQ��*�S�~�Ec�UR[ų�M�����7%=����Y��[E�[��{��(���ϼ�W��Wg��2[�qp�H���s����J|y�Q��:����|�n 5���7.� �f���q�S<�<�$I��<BZ&4�����vdP�k��S䘜��H�ʲ������;qp��|3�#�Ke�&�[�;��J輴y����m8���q��u���a�,M�>k�[�^�#�U.`%4m�F�8�j� ��C��2����ƛ�2{ƕ�V1B���K��I�,��	��6�9��L 9c��@ڜĪ��h�Ӣ�x�f��q���1D��H���*/�_�_��,K�	+��*=շ_t���a��t]hrGZ�57z�.�D�>0*���=�2�v����=�%*q�J�k�!|,��~pRZ�	�M9�F�\�K4�)4���K"�����R7����H���fA�ҳ����T��I��vp��Ph^�r5Z!k�^^T�+"̭fz.;�;��k�\yY-���n��h�c�8͝�J�ەh�D�ភ��=1�Z��ӆ�8�g{~>�!8���d�:�d���Z�_E���s�hq�}�Kb��l}]���o���?HZ/������(a�v��H�ъ��4\��+�#:X��B���~O	8�?�F��0d��9���	��^�� �W�&�'�G+47��?�6�mԁ�u���/���v}�x����|�^��m�酟�1�ī��.]'Zα+����9�Mu<'1��S���L�
?�g��=�9�IkfA�n�/���Az�kA�h/��AF�H��O��e3<z�����{�c�sq�#z����S���ӄ*�����42?��2*�y�6^_3���Z��Wm��2�`�=a�Co-�������/��*+$��J�,�����u���M�^��P3�٥�H�j��MT���Ȇ�Vg���	Ղ ��8�L�I�O��
�2��mA����g@�o�Sү�|}�yD���b�����14���F�&�h��M�=ۋ@�\ ���q�b���k���Ge?�� Ƒ1ػ�; ϡگMj ��m�0�wOc��e��xU�(#�^l#��'�~���%"]@��! �#�=�-v�����_�~턝��`��8�k������]%�\I��(��LEo�nP�5�I쀉�m̬����u��Qj�=�Y+Kٶe�V���>5����H7���-�g�����q��=㬨h�
]]��>C�����5w���!K���r|m�����I ��-�_��o/���ߍD�+�#��W]�@�őf��9�>ǁ`�Bt[�5Ql=Tw��4�r��5g\�z���lJ��љ˗��3p���`���k� ì9c/��	NE�|��	-��P ��v�i���0|�8���<ϝ��q��`{�Qܟ1$j�9��}:����V��-t�`J�N%m�$�5�6���j�8�q�a����EWL�Fy׮����v��+�H�O��Q��a�3"�g��WD�z�\�\�~(-v�,r�DeݩK].����T{��\�����	��F�9�/d�����Z�m���n���M����-r[H�[C�Q���z�t��^5����.zў�uj�W���W��)��A�.��g�\D-�O�7���R�,;�-���M�󸂛���exb�Ŝ	΀>���i��c�`~!�x4����!�Ɣ+`l&�J�O�-���e��K��m�-XO����~��<���gI�t֍9\׺�J����=?z5�'_��@���Hr��?�_`�]\��$��X#W�ʘ| �����-dV���f���z۟wW-� s�e�A��$��W:>Q���8ȃ���t�gYo�k�u�������q���4����θ������2 ��-��$*<Ќ�N2d���(S����"n���*������0g8X��D������j>ٕ���
��ۢn�k�}4P��T|�A��ۻ�8͵`\�T�>1�&�\#����}G��'��)O�}�Q.w*�r���X����w	����~4$C��L�9~�!# ��Rd"��E4n���%�Jz��8��6Z��X��
��f��)���2��񧽮�����lQ}��&ɫ^=�<���^�Rm��u�QHFx��Pë���[���!_�3�T��6��?���Kj�F��3�<M��ۢ0.�0D�F���GK��B�?%\h�|v�<S�gE�h�6�V{p��R���2Oԥ��s����e6@�6@�a���(\W����
�j�Ǡ�@>��w����M���!���y 1��]��G��}����X�@'���,ݽ}} ��V���}�z���'�7���y��kJr�.|ˤ�7�Vjw%=ẽS"�mz���� |�ޡ�:�dS�z_sx����3)��xx[ /	{�B��^�ѓ���D+��;
�\о�NԻq�Sሷ�[���=cby�ț3:�A�U�P�o&蔜�J��x���2sp���W}�֟��������%�|,8����g�:+�.O�js�.��e�_Q/�,x�T;���{ �Fp���x��~�?H�d����%�d��Y��h��"� �Ex��J��.�� ����_�٢���#r�%�w���Y��z	�	EH������аm=aGae�ygF�Hכ��"��� ��E��/'I�jE��,�;������ ��[�J�=��zet�[ƐA#o
��f֢�~��iC6��@�G�:a�~��i�,��	��q����1_'ߍ�i�<ѳ(��"�hN���ϐ׭â��Kx$�ʈ�恌J�ц/疟�6Y��E���*�8x�E �=L�y�ea�y����9�X��Sl
+w ����
ސ5hR6G�Q��T{k�:�/'NT����-!�P�<��r�:oo3�l7�T �>�F�&�7��	�&06_e݈Z9j��
Ճf��Q��:��y����f�>E;�ąC���a�#�|�Ot)�
�{�\�H��̆�k����t���Z{��G��#j,"ޯ�K�IT;ڶ��N�~F`n�����]�B���'�~����,E6��5���η'�������;�-�{���)���G
a�X˖	���n3����ꆘ�>1��|	�x3�����^a�8rL¾L�� ���a�m0��P�"D�M vԒ��w�n�I��(����A$�1�6��Rڟ������� s��s�!{F�x�:@��a��78��P8��X>�����j���Tb���Y���@x^ "^G��g'4+��鰹�^��ۊ��s*ư��&,��t�V��1H��e
�L3�e���E�1��+�I���QGc(�!����K<[W����a���=ݐ��X��~y�ۈ`eBS��� �A�P��IF���l�lB޼d��dz�I2i�qk��ӵ�Ҕ�&��r�o��c+���h����G{@a�	n�W��v�j�	Ӧ�W���4�!}�ιY!1�چ�ĉMƽ�Y�PEX}�i,�p���	C��7y]�A9cj���+/�0�O�,@|��'��0��,Ͷ�S&U#;|:9i����6bmrpv^�+�Fߪ<#F���� ��yW����+Ikl�-�4��Q՟_ñ��8d�!�D�X(�7�@x3�`� E��\m��k�ځ%��X�PŴ�ᘼM4~}�z��"gO&�������+�*<�Ϸks�(���\�>�f��(��x�h�
�[���!f�?�>Z��;V��O$�eЌ���>�H���T�`0z��v��F?!ot/�ݾ�F'���9q�ɷBO�����,���o�Z��l8zH���z���rF����2Q�f���$�I>40�]g
� 2���ceHwZwXyN���2�fD�f�|E��4���@B�t�xS9�5@A?����vA��: �"Z7�_��Q�_�0���u�G�,@{��}#�IJ�M�����p�M,
�FQ����>$�/�8%z��l�2%���.�G����)0��J���	����j����Z_FZp(_k�N�>�45�|�p�b��}0����lXI���~�{��$[8+Ŗ��O���4XH��M_�7��K�FG�Qz�x5b9�s,?`~ps_�����VN��9v[��"1_n���ؔ}�e���bOt�b��3�&4cѦ������9uM�	��m���1�06���S�n�?|oy�g �~R�lHTq���+I��wG�\y��l�R�K�i��_�����#l�s� 1	q�՗��0�G?EW��=��0�j�9��ج�HR�M���Д3��m�O!�v��PP]U��M��|S)ёl�w�,7D���m!���t�% ����S�Ѝ���6��\:N缸�9	�L�y�E�I�^�ǯ���L8�Jr�<��=��q����[��OF�Bb�W��5S#�H?��2<tۥ�$���kõE2]3+��|R�����/�II:��:tG��P%Зs��&żļ����a7Ť�I�^ҖM�Fv;��P�ۤcߘq��;�J��KyqMѮ�_���O�u6��		4ז3"z@�4xx�c�@�����(����܊�;�(�絡͖T�9�.6����Ⓧ¸���̻. �/�7J�
�ڋ�"J�'����2چ�Y�F��Ȕ]��Pt�mU��dy�?��2	i�)�Ą�p�	�9Q�(���j�h-�y�&��Μ�OV��^��9y*Mչ�/)Y�@��ӜPڳ���t�_ߒ�S��2*��Q�C��!]��PhRȑ%�T�|�Z�՚�a�D$�Bc�:��!�87�kz������*�|�ڇ�H����f�m�FIŻ�^BAT|mB�����hq�Ҹ�i �e?`>V��+b�]������-g�K%!������.2��^��v��7)�����Fo�����<�8U�ã�2�J��W��Cq� �(�g����42����: �K��Ò�y;t8剬Bg�ƨ���BĄ��Bq�_���;��²��{ƀ�S�:�yʢ�4	�gPߑA]#zn��*ם=�0���S+�D�C?�@74�rx�S�8-�;�hp
��5��ѿߢ�CΎ�5ִp$������r���86y�#y>���6"�����5zg3�iJ��^e}���_�(��4wLh�a�#�X��B�*" ���t5ՃX'�?����{5*�}������Fy<fl�znzhqi ���%��p����a�g���ڗ<�]�N�T73��L�&�ۡ���7;�
j
����u����+{Y(�Д�Ke���݋��	S�b�������%�֞��VA���=��dV�%K�S��x� *�Ԕb���$ϰJ���
��|L�X�e}��&XW���[�)�����:����P]r�)$\��{1v �ؘ�|���䓁҇y��_�����9�q{�9m[�&kτ
��A����
9q�.�\Ul�Ԣ��u,�Xcɝ����WXP�� �.������l�m����m?բ�7�[�m�LP������w|���u��E��[�@. gX�ʲ��	L}�cY27�i��H�|��*s��o/��`���`QZ�3���>�HV�
��=#������:�yhvN��%�w|�N{Eӌ�6i�(�6���z;�7���
=�OT�qQ
�s�E����WI�V� �B<_�������c�vh�����A�$�F�#�F�T���-���\���@�̺�Nh'{��,rtx��pFœ�+��×E�����0�0<n���J����LX�n��!Hơr�qo�ر���� ��e����0��R4�rש��Ihk{��4����>��������*��M��%)�_�2�딗ֺ"��J�u�
��ɭ@Q�a¤��~˳ym���s��d�J�U��s\��{׵+�P��IMl�l�g�s��������r9)��z_R	���DmJD3��?�n����s
$bix����Ε�:��-�Q.s���'_�Z�}E'��c�M�YA�ђTP��1�S��.�����R�g��r%D�r>'ف���񔴦�\��B�1��?l����o��3mY�`/�}�$j
�V,��6�gR	��m�c���ϵ��]�[��r��/X��轲�>�����i���ɭ��-E��S�f ��U	z73>��z�G����^�Dy����0���I�"J���L�pޅ�}��f��Ί{y?ˤ���f��jt��*Q�S��6]��F���J@�ʾP��||�ݷ���7&۰�C+��O�U2޷�Z��߄�^���a���O|�7���.H��f-�����^uL�&�F�Q��������x�פ*D�*LwN��xXq� ��ܘ��&�����r�ƃ+�]�򨭷���@����yNt�z����rGU�_ `m��<��>�Ŏ���#5X�΅8r L�)�3gWO�YO�v]tCJsW����z<'�� E���5�b%�q.�Ɲ�v�ꙃ.����Ă�Gɫn�MΖ��EcF8���#o�ݖy��!��J������zJO6
�y�J��6�&���#f�ȶ��4ĐSÜ�kr'��y�š �6U3@��#j9�r[��@�&`���؜����On����ܴIU8$ʤ���Is�V�%�����`e��������e���ۂ�y{;4i_���cm�Sd��Q�1e�-6��h�G͐����a�Y��G�6,�X%�ꭥ?�y��$�6�}������EG�B��#;��޳{���Z���h5�>1�4��.F�ҜD�ޭQ~jV���j�f�%�nO��U�Y���bZ�b����Nx5Ϛ�D��#30�o{4���_���ֶzk_��r�V׬ͧ;��y`憒��uDo�Ҫ�W�/�Nh0H�#�5@Ӄ��ɟ���]RGA�l%�X�� �-A�f�h�C�����M�\O����1�['��}�
D�]6��D��<þt��,H۷�'���6������\�6��e��%�n��[~]�s���}��?J�`��0io�k0��u��h�����oț��մ"c>�g�x� �Q�ݩ�m(r�����S
��<�j)ӗa��_�Ƃ:�R�p�zU0�V�t�|t `��@vaB��QdV7��dHn;��j��t��!Y�y7��L�oI�m�J,_%T4,$ڱc~��v-v�|��@�˜�:%#M��y'��^e��y��y�Z���	׸6ہ�=u4�f�D�V�gkM[�cr9���S���˓�-y �sL!+>|�U�(P�X��6Z�|%�C�m輻ʃyqk�3 ��#�pB��@E�L����APW1��E��H�����sn\�{�-Ά2�r���b����P31J=��*�s��u��-�ur���gЫ\S���Ƀ���u���tI����Vs�:v��/���Ja��Jy��db@�l��X��p�H�`�j��$�XBY���� 蓑X�dj�SLȗ��ؐl�a??��u��>l�%��<��X.H�Jw �R�;%O��Ċ�����M�*���G8PE��,V��!�x���Ǭ���Y��pt�C��Ђ�	��o6����F�;�:;�9�3B[V�.31G+��P�d�W��*k1ǯ���vGʠ����t:��܃�����z��D8�s�Z�Td��=�Ǥ\I@ �w8��X���ɮ�m9���c�����Q
j�Fw�8����}e�?<��7�v},]�J0  ?�^DI%31߭V]	i,|�(���"��_A�	�[��N�sV0+$�V������ɒeMrD������e��I�B�e��v�� H�7w8}-�r���fF;+��=��%����o����'#sn�,i�T�Bsі��/���D��yw0����M�¼ߙ_Tj���pyC���m��_Ƅ#��:�+�~\)��n ڠc���L]�3��&g�ʊ��A�N�u��;�6�n�V#�uرs��k�_�+�~�j���_l�4���I���wm!1߆?��,�5}�X�P�Y���,�f:����t�uSZ��Z���	ݸ��k2sdA�EB�V
�� �N��V���ĞU�,d����ᢺ��R��6���B��Rͺ��˿�����{{?�̟0Vz4EbC+i���Z@Ly�F.:0��#x��Ɗ�����nW����ޘ�؁�5*���&�����[|���FtE4Q�%~�,�V� ��Y7J��QJ5�碛y��<�W`w4�p!�bއ�dj�o�,��F;q������aGΤaYаՒ+���N�FfN����e��A᫽&���`���<K8� �W��']"�,��T�������8wk�uTy�:,��$}���b;ǲ��_��`{;����C�P�Z�zޕɀ��E*�ٗ'�-ӊ�P+�7f�y�E׳���m1ԡ�^X?y �H�msC�����ߕ���fB���0O�?��"x&��=�����r k?k��aR����kA�Bt�U������vj�Y�	��DLe@�r������.#�.�&��kd͆X��
�	�md����Ƀ"��u���"~<�?=�V
(I'��<��C����)�:V	�x�a���(�s.F��~��B:�\>���Z�7��:S� b5��5�0�\��niUA�%AnWڴF�p�� ��fe�+��Y1�|�"���p��w$Y�1��l�l���.���