-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rkgurBehUiZ5vSrOMPhEwIvzyzr6+IyuG71WoEW467qJuqRdO8apMCjEPgfX+xA2bDNaTNOD5w3E
F9kdDf6oZGQl7cltUjQM+wkqxMNgxuAoF8yx5r6DWKYGsthtgkl8qBD1g1yXSDYZeHte8OfhWh92
+5iO3kEyw0MB0imQOV6lRK5iHhnIm6KUNsX/R9kUruf5iOg3s5JWt6AaLbEIuOTakA5r5seXmSVO
B3UEuXRHGlFlL/hKVMbogsXK8Bjfq/OsBbyvuBOaO5Y2oiEHJrQRuz2VGKNGHtVRKn5LR3BDGbUn
Vs5c+owSgWwh6Mqn3df2jzvqkboezaPjlGeMpg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 111872)
`protect data_block
QGP6reFRpf7KpEEQe1tBpqUof0+OcWkIFqNcHi1ht98Zs0cHmIFRFgvSZouXvUN0k04Mk9g2wPoq
BQvz37DOaqEQ5lFUjzSGbCwxpO9WPLH49eNWdkOO4P4GWPO50Hw+vo1aPzNmw5VU0n3DTtNOYYSk
figC2Wz2mFWmqOBQ0fphplSdJBPQfPRt03IZvA1ba0GzOE9FXBc0iRBTt6mCD7GaqaBz0HxWnezj
8CB4IbWUUrewYrzrW9ypvz/D8yLgDoHbqRDsGExDgaxL2WW27j1OPJ3/CbuipMC6jQdgkcuz54OX
KmG+04pES1TNwTPOwwuV5AFLiQE4CiH4f17SuhdUPOAq9FWOEqWIeBxWnYD6ntDucOw113spzfGf
c6Ry07NVoK20XNRb0OtWBdP6si1d5MTWxV/mMdAOmjvYy0TNgN/7gZFzjJOGrK+2MDKxDLnm7aXD
65gJP3djnujotTtDIHL/IazSId0+seyyv5b0cniXZaWr+Hlcrn0oIF9qtG8XwIahLJYVEJj0UMSP
zizLWHzNgx2iU0A3OfSZ9qqlS2nvdZdyo17q037MgwAgany1GuiaERBNMfO6EMbpJhnQ0xwsdf3Z
7uV6kQ0E4TMDFH2zd1rFSmNyUguNvzvyDsrC7+uPvGZflmJ14nmM6zImHr+QvrAUyy5DGtlf04/m
O21kXD1LRNjdBmX0sdMCpKg6g3qGMrmfVLuhJ/ruorsNkvVO/0qoBGzxcrC5ya0IK2tMF89FHSHj
4X6XYpeEf+iN1OE8WRkRHHx6LGhL8jufa8Jz0oI0p3CcGVbapA1q4XttIICr894X5EKivk66+TQB
GldHw8I+6uRrktSiCIDqY8x0UJhHm6/UTPSAsjGXi4G2GdCRZ7g7GSkpCEyn8avsoDtARdSIQDO+
Zhj8m/ng8LDj4sRjyyOgJPa2R3qV29xyqtoBMYQqLQhg94XhWm414zITg7mN025hM5rlh4kFXunA
bBSc0gMzsLl24k1mn9vwVcWAo/SztDcF/3+8TLjuStkh+Tvckv2JhioadZ2bJjwhsl2ghujKXNBx
AAGcnd0JG4I8bO5TrlH7IUou74rxy7OQ+3NGj8d8yesDlEOODqpiwjTyOuqIPFL/LzHYxzqDMI3q
uzM7PpnXjyifck40EJptOUDBedEf6008KsTIAhbCYssgM9gnbIBu4P+ktH+tzMK/2hwqVOY5b9k9
DRcNqfitPNilajdGjjqxpSnjsLiA2WXQdVONVH0b6+G9agSvHf09dEm8GmEuYR2a9RHmAzV8Ji0H
ErfIlT1lp9swrAOxrj76WLdN2DHGBgFnXtuxZXQwFvD2eTYO/bXP/CyTewq7WBnkxH3/zHtgHXZ+
uc7jsxNSfYfY1ewUTA9X4Ng8k5QDHrX+nqGFkLU9Wl07TAc+PWvF1LNIvFaBOcWwPww/ePSseSP+
IkM4AuaFwTB+CSEjhykxJUZwGDS1J1qFcRB52Z+FumgMFA3EaYh6mYgBlT2xy7D5iQ01prhRrVoy
33T6nBta2vkaAaieJGT4Xv2mtEbvXlRaps/N72InLaS8UdcYImHrCqzp2XqWyBNtGevBmYboCyOO
Z2ZfAZxa/E3iRjI/OEPi6vy1dOQcO+SR2IT3EYwv8ZtiolLElbpFk1qKM7Kl0OA1kVMYBNet6Bfu
W0yvQHWiobJd+O35W2VN4lGWHKjiX8EKum7Ry/2gOV377KIAOOMmwrDNmxUPh3K/ChmExNIn5tuR
d6KwmjEQg3wcqNp4SZU0dXEREVlc73VXcsxBvevCCjcjXMtUaCUQPkNVLcbo1ahxc7SINdE6S1yV
KPWVEXlWHITBm3CWAZgqwOznVlMTP1M/C0NlY+xMM2RIlfqJ6PZEUmli8DYxqtAppviPyK1TRCme
E4O801Vu7lKFjM1nlob7bMgSrIa9mCvlkH5patSLEy4G8ar20N6vXQ/T0C4aKte6BWRqf2rODmX+
28Ced1DclMTmvuRVp8m8sQJYwWHYSBBagGWb8u6sAk6zp1ncj+uSm8dqH3Jo1o7wrBFJllz3/6RT
u5DhbVDuo0xjM/+5oAgCc3sHCtsooDGb55BVnMXi3RVCOchEdh00zwP4O4UenBv7ayUBfEn5tvuK
KG6Uw5NFeuaUUD79hjA3DFyDx2eGBMafKktY1E3w0dVbF9Cvjl0Mcuv4HQohiiMw+GQ6XS92R8BV
spc2wcXiSqSxgZp2yMzlT/9WQ4JHzdeVxRpNO9Wqc2PIX1ZP/MtyKfI/Xjc1xScO1xPvm03vyuO6
Dtjf+twF5ZYGOdLgf6A6MCjGcqq885z7K0qDJFCapJbho0Eh0QDJiwGnpm7J3SZiofvMqySutcs5
4lJV9ZN7yiPnYCRjt5cbf21HiEE6FE6qhD796Nmyefx+pZDZXw9vxwK36UdWjYXJ8ZbNhGXOvyjK
UwgA5InFMbh5Tl9f53AqIhfblbhsWnQUOOe54iokXwb24iTMMLijGKC5QlrvwrZ/rEW83JA657Zl
K7m+NYduEM1TE+62nwe1SdfCF4PxnQDOJ4jGQpjOW96ZKIkAMcO5qzsfyEjKbLxkB+nU2rK6lZ7F
5SYYsOloorM0qhP4N61so8PN6wdThy1zlWpVfrgE6gEb6X8RdxFE6QEQbGtU+4b2b8q3OBB3sW22
4GeYT0lNbaPaObCyPCzbghhNhNvI8FDbE1Vx9WX6PDFahBDm4lHt3QIRMAM59WzTj5ptt40Yi/yT
TElEgTvZtpH1apm/PO231aHcWU6Us4cwJeq+JDj7gb7Z+BZvtuZdzXGOKnVqTT91XoGMRnWtAvni
8OunVRFOaJKDb53H4sp+SALX0AH+E++fy4IuE7EWMslh/rVruo5L4PYQFmfcXb5uYBLOw4t9/F79
v2smEHNYxwXLccmUMqLnFHljfD8A2KeswJ8IDbtrb7/mPdKtgLYMnNPNA7YhqgkFxwsR51DH58yK
dQiR+e5syfBaYeM487jcRafo9UdMACLRkcSXELUNDV8lB7AciSlAgS5ZOKdZf+m9BNs8wLnonnw9
wYbmlAh49GYgY+53ESEUkNt/si7kdk44ko/0J/Zh5RnFXMsNM/x3B+UU5YVKltpsu+yt/qGo+Tiv
boEy6JLpJcwZkzdrxAq8LCtjpIN+/zw4O/XlxrykUxbu6+OyzPkVeQhvwRiOH2ErJv56P6XLKOh9
j5m7qQTKyd2USIUeZm5drX25zKkAr8EKDCCnO7BMPkIKa5QP+0K4DsmduE0hKVsfAjbTlKs39LQ+
etVGhNTegow/LvdMbR3JNxhdmCxXfCnH8rBxgpt2oUcnbrKSb49us/6v51fc22CvPiURrb5ab9EJ
XkDp7brM845OSs0JcjqG64R7YCyXYbYejyBFU9IPol/Vyl845KhG4vIz0Dt2WNCLxTFwVMIIw8o8
QpAL/435TwoLTpOXMUBP/RtGDQi+8MzPrbD9mcAFGP2eJI5FhzlExasREZ01FXMGDBrMztZJJPzM
g5l0cHipFWp635H+ab47zYcpO4FAFG11m5k5LzoAguXwSH4lh81J7kF7lmfvyc5lpIiO+GskKdQ1
wQDtptMPv5YJYxkzB6j6k4FBGDfPtm+3m9LbUAKov8qXaxdefdCfY8RRix6y3P0THj7vc0pbjUXg
bsr4YJ0zuGmG48x16hp1O+nf0Dkv8oZcmcwr7/XO1ML5hg5y55yqihkva+74+ugqshTUUpXIxACN
iASB/2piMUaR+184vKioS8lMUiINUiOr/w1cNDLa7PRz7VhhYz1BDmDrJ/9fwQQ30DBag3YHv4S8
2QL6pc3pfaSnsffvkL8r3ozIxVQ1dfgb/bJoM2k40ZRjtwM0DJqy1yUTj+hMlkYq1+Tuf20yAIuZ
KnFEGMakpZsAb1DCWBBt5w4EAX90gvuJojNByc6+FhHzK7C19UaFHso37ebV3Mcte/s8+AQmu3aO
GsrJZ7qK4c3ivJ1ZA9qBDzpOGts6VfWmPAfpZUKTzSIBxVAf7w5PVSyYW5ZH8CAWgK5ZJMLiu8OE
/he/XbQNKzUtgrcM+GAX6m7JGtpUNy8a71MNzzOX3m0pZzoAt8MyQVynGrktLjYBrjLnCCCTlqPw
YR8WUnOZAXFgF9V0vcPS6Q8y9eG//iJQBOVDV29SUho2occvcDq5FP3FZV57Q+Je2LEWps/L7Rxf
j8e/6p5m20DLNRBASPLdRDfY6rE8vUkBTqB6zrpr7lEEdhZBJ1tFNY3Dt+GbgcgqTsIfTep91x2r
2f5jOnnuX2SLzwsCCKzpQezw5yUWbtRw5Vts74Sx+NIm6kYpiGgBFhB+br3SYpSC9Xh0jcjlaMbF
DILLbN/5thsI5f/jd6wyZlBv3Z2LH9/yNH9koQVhhGZVD+T0pDizLzIX6E7FELhIExCE0HuCkKx2
nWWt0r82iIlDXKSMHKdcS2xyJuAqKOFMKaHgEc9SShErG4KA4hQgeqQ26VVAyIHorejzQaINL4DU
UCrTpNCPgvm3frfL9uX/e10c+xIJtwV37tpi8uwELB4ueMDuDi9DxBEpKOB6x1ha3PFI+imQoD4A
f+iYrpzG3T3ZCbD+VfP+2NeypaPT+19QQT+vFy6nCBLlY5YAwPonMQWAVeH6NrUqDewIoplWoPOh
s/FFMdLVUx86R1f9GmOSekiP98knAWnbslyQTblGOejJ8A7SLcOKaHMlEMo9EF28Uwrcxs5XtzA+
CvmFVO/+7dkhaXN1psthImM8snM/i+81/8yRLf65VI5586G0G9ujW/B0RpwBc+eytM+qMSkYK/Nx
tEdLqDnnukfin/DSav7369ZPP3XQ0unH/Gn1lbwLZ1CaPx6QAaE8o7stvWt3mQnJMkWwQuohmeMf
cYfDjYumiNdeiBdRvo8fNUVtFKCzuUmq/lyoOcU/o6Drv5+M0wGvLzwvsArWN7jWzHqM9IcMeaTj
5YV7dMzaTN8ywQPu35s7b/n6rZPLZtvAQydQOCMLsEi5welQmNf1jfJv5eTq/pHkaouJAuqY7gx5
XgOryUM3pbxPfevjHsjs6H+HcTTRTtZUnxKgO3MW7vnvfWVpZeIi4uI1QOdI2B3M4TUEslr4y88c
u1phZcKMbwu+L++Xi87ShTPdLSUyGpqSXglNqGuW4UAPj49V89AtVoZZTnIMs3EQiv10NdOasEYL
j9JYoWEk6GCSiO0c5UzaL1NOj6TmI3zMDw9XGowRXxfrd0dtdSyLeLqkgZ7UaaveXlj7ihvSDL4z
855h9Om+NDvBZ7pGhWFy9M10anG82NPizK9wfJAxs3X4c+1LqOmjzzeEBI4EskxQHpHtDa+3xxrh
T91etFOd3ibultO43f8n3/FNBBm6zjQzJcWm4cNleXhqtJIrzJlza9c0dGfEORQptso9xtK4zKZK
bEW7+kDHbBPtlaLcPZbJxz3zyLRdIq+UqYVdEeoaSLc/Eaxazzl1DTxPehZsaFV+KekSmUnudnCY
bWyr2ckGVkh+zjrf99staLuWj+NdpKiOyZrD63aQw2bBWgozKn4kWNKM5CNVezJj+MAYHG9q2jSE
7oDobpRA2tehJYrJSV4szcUTDyR7rvI2bUUquBhK1+2M6R3UMp1dW24+/+JQVSHJnJXNnPbZa+3g
IQFMdunA/NWQhPoYLJFxazHAy33oe0uhvKLFDsFrDqIjH+xBgSIxqp7W3Sniz4l3ZL24RrIUVd29
uGieG+doxnLdI58O8uxDtK7+E+5K+Qx45NVQgaRlNiIXp1rMnQ3I6DqwaMpJMFa9KO/qBCZZQcw1
8yh4gN40apEiFALR6NSyWUAbgrUw42EIPP2yXPVaAX88xqxwT6AWGSvgTkLpSVmRvfUDVXoA6t/2
JB5khhYjnVh2C58YS1jpG66ZwatIXkgjtZJkRbY3a63Adh2SbZ/+64nydbbjMI0UFKAv6Kv9XcRO
Wz/X85SbIgQbrmUc+rP0WwRJ0Lrw8vXnai0MIoxkCkZAIGYoPHpiYJtkZ5nlrfB17vDpO6RWnlSE
NrqHanP8vdol/eMhASvVamLGGBAz56+ymHouImZ6NfAHDfstzJdOue/NDW9VPc2TBWoKO4pVh//3
DUoWuokvh4c6vfN21Y1Qv5AFlud405SOKy6ubrtzxLii38zHkrdaXVFHGeAT1rmxxHjgfaUP+1qj
6ynB6iqZMwWRSJbGA2PIY+v1rym+IX/MZk4+Nvte7eYwxA64xBFYAtPgmpFiIi9x8muRnyWHF7wW
rP7yAPkU7+30vcgYIW+U50GSxiYVosO87sgtTXmvfg4XOi13lIgAYSB4DyJUR0Z7jgrtvegEsgKp
ksX3+b58DDjrucNtZ4/TutYeStTUVerggl+9fHzPdkHv2OENgLOaFFx6IBCuOnhdRusqxRLIy44N
W0kILspggvW0rKTNPuIlaXOJH7fIE8Y52oSxFPEQpr/NNkTHcQA5RYtGTKFZhcK40Eqh4E6kdBPu
gjaZr3nYKDbcLDaW05r3zvra6O5/3bfOKnBIa6IphT+qv4bySvqrG65ljjYdm2sPso16/4YrYzVS
nvR4OceD7z2vHzxhurDcLMgUlnTLb5JFdRyXygceOAgvHv6pGJ9c0LFbn1lYNFb2E3B2p3n7/V4T
OEC/7KGB+hkTFUqgsOJfeSxoluD/zu/6/gK2vRLvEdRK1iKhu0cFpVal0Ani09v7jPAPt89GHtax
Vv/MREoGkb3rzZ37igHPUwOS+3S8oadEkQftnXXVDKhR0b+0Nm/IMXAV+mZLmB72QZ8CtNALJUqS
jS4OQBM5Fuia9d10xCvVfLcMwY6msxwRIGafN3BQFGRKGW2SD9S7RM7LRXhbbvHQhZGXzuAfUhwc
yRjcgk+47M4wSiede14+YKT4XNQ4Pi4VhYRZatSCMegr0suIvHmin7U2sPmOvkARx1UQWGIY62MO
6wr59umeH9wHL4AIrDKHRPErHSmABKNUjYFx+XaSyFcbO9hwNsZkSkNL2/TPxKA09iv+TZzEKS0z
feTEp6hPkyAv6GuzaYq1wXfLPlc66zmEb3mFmLrjVP2HtgMfTQmpsV2PoJ0wOS96irNEzEoTD1As
jJKC12ppEIUxpiPGIqixWY+Me62gptnpbn1yVuzv+AhR0+gK1QbixvTb+CEdF0bZdXFw15/hZ+NG
r+qbOazDuBgkUlsqYWIZ60J+bUs83fkDz8z8/S0lylVkxYzwB+QK8S7Vf1dc7Z5yjPdw1FFrb0ai
GNT3BnJ1JTBNZTBB0NRiGA0bPWRWo0PiXmaesVNp/5JVmemf3mlINqdUOOSZBa99w/c08eVIov5k
ZWTJHcrLzBKLXgxIlbU+trJDP7Fs8xlzdoz2LJykGSaqt0/rHH7pj1aTcCA2HyLphoh8KFO1OO08
8WPcF8zPzMFHFaPGIEcVJ5Up2eknf34HrSu2YXC9LSu7u/vJYRxA74NAlnrzOjomAFYCKWhpTayG
DyheOah8zuQu/Ohjw01ql1ZjNCBmh5xy+JStfvHjApHtOZs3UYJppu0JFb/DhHIvB7V2n2C9m2XC
CnNSHSdW6fMcvH4I5bTzvLYs3IYmHS2Ghrf3ghTUslznQSVLetSp84DTWIQCdJB5lW9GijMZ7GVu
pPi4QPynh59CLeTHO8wDe33A9GuEWrHpW+6PyE2P/gRdtS1yMvB8BGs1Ce7gnK8OChXOY2y2tVTY
HbEUNnoc+OLCVwi0eigs9hePV1JtYj1XiIdMNjHIL7jb9c6Lpi74P2MvAjC6Ix0v6ihkLX+TPwAX
jbWghBsxOVzeehTtAJPvJL1Vx4rG1UMmOL6af6yS9+P1eC8pvZVRLQL5O2JIedImO+PXZZf9nsFD
M8ea8NkZ6VlM26uU7odbasNV7xCMuICZwJe2exJ8bLd68Ki3szs26TbsTRMHU6BwwolZTOJ3s+Ia
tP+UesmlV0+tjUxpLTCsClc45DD0towKxzb66aTjFz/x5pWaPdunlEDVR7k2Am7yQWkwfkX2icNf
f+ygvp1IdyUX9z7QJZAbDM3yHkKXFjaQyZbB0vmkH+Iek4n4ligQqZnu5HK1nezsTcKMBlG9qLRo
8NVEZ/wzBzgC/KHEbJSS1/QEMP6Z/XaRvS7aKsONfFd/KWnqBfJu54eFNmtl6ckulOWi2LX6irOq
xcRm0NHr13+Ny5SeFPwonGNJwuqSDTInM/MlmoSknqIZmHcxleKes5DIQvHCP8HsWNrkqHxSmyXn
f1VsXlNR6kkCmtQ41qF4G3idQXsJ3lhnG0CZPI2G8ymqxqdWLBEn8uYeOeFmeFcnCnXWZSxWddBW
cXtSfzWJ4gY3HGiiOMe6AbUfgz12g9r0t88ptNRtxnKUpJ0KtIEJtQrBvWk5xn5+mXq/34EPET5B
kquL3v2AzHSUKyh8yMklPgEAr/GU6qM4YCccXIJsXIvbsCJduL6aNgYvxtF2ntEUZPQokzsatCKa
spSoscjd5iaRuzeroDOAKPbMplbsLYlAi2aJoI1ss6meqMYM6pU2G0EUFhnvWUxXMEnGK1aY5+df
ENT4ILUGh/tDd5+QQhQ4JRV5TeOkMbysDKfnV3gVR0Vv8VW60PSsinwVKLszc3AyCu73JLuJCP0A
zx6DnVvFLR8sj74CVkxQ62thHY+IdhsN77lC7eqFhXegjP3uNBC30aS8U6qwG8geSq+8AO6LU7W5
b7iTUl6RwRUERqgNXtsTpMtK5gJbmjwNgfnHEKf/TuH83Q+dh3c/J6pb8pTkbBihQmfv75srxBss
8IvPrQfK4OgD6ASw/+Kbrp47DEFPDzX5i9EN5L6fNHBwqmF32Q8+aBEgwY8G9gYUcWwK8jXDlDBW
PUBztdB+hdXPi68r79J6h4t534v0BXyTJrA/niVZr1aFrzymF4wnafXZiqEAdpmT4Kf/TZQziIXE
WfpOiBXwqSvptUx3jVlQPF14qk+d7Qp70lXJl86dZ1ZrKpzv0/c+QQ0fbRmZdtNCnEVtmeHejmwO
qbSufzQx2hAkj7sFuzLL68ZnrXFFbVrHGDAKVxUeLI7KswcGHurOYKQxFpAjjrExbZS6AastRPEz
c85FaWcGtgEdUxtCoKB1Lp86xAlhoQCWh/+1wCXw4FZUq0AjDV5fQuGVAfRBiLQhgmu2vF7IuLp6
Uqz1qzwh4dEe6RG2LruI9RADTp4eRfRnOdeiKTQycsgnGkZR48wvLH6AVgwxJ+znBnjiJd1toZne
jx+jLiAeS/+c+gWy6KJqdoak93zTRMzehgLN8uzabFK4Lcje/X2anJVWGlqP5F38a05EJ3TWsMNO
lds2w4DzWq07tmq53fV6CN9afefj10kp7mJmv8bTuJwSYHhNN3401bkjmmMEjfVK/hZfau1bjqoc
XVNaa5Bofnq7M51FNbxzOk0rqfq1tL9+SbDBIuca41jzz4rKL74Uw75WIQ18kptsilmndx5mB/YF
M2tvdLXg5EuPMVH2tDOzrwHUldnzCrd41k/zUkyR9xm6iqCFqmRGFBc3+mdJKuahZR29XdSr9N/D
4JuhqGcpnKi+DXPApNbt6EnoG1BLlNzvJ+gOXq9okbRJlRPFvRKrPNFNpiVvH2lM7ILohEwIdx2V
Te199WbD/P8McMtRj9Qa/rCN5WoK9bcoJ1X6PUM1fm2cL5xabUfDfRdKVFw2cLooznFhf9gkgFdD
2XvblWVOXtjejHJZCs6JRDvFnQufVFRLRYe31fCfNKGhdPkIGzvDdD73/94ud6vUJa8IoKEkI1Lg
WeJ2R+TZ0HA2xZ4kCQMfsfWWaAs0e/xA+3gG//sLCHF2abLTU9ikaw0jKpPkUb38bpePOcuZO8ub
odpQFHlZHd3OXTxCs+YDMZ9P4WCNEhf207WD/3FCrSC5A6IknxH6khMTulnNTJR2h5XO7nrKYuB4
mA6y0dOM/edGTrjEL/43E/X1tuagg/eve5N0higZCEIfK17HEK2UwM1wrsmqaEh9gPxhi9HtHwVe
8h4ga0rLFKyMPSU88YYTYWzeSqyRBlAMlo1XUDPNbvWkwUcKQQ68FJRin06NUVFhC1n/+MRIlaku
OCpvo4tDIzV1XZU0Sy80gJnYl6pshtZDiKB2CpyAIg7b1yaRrvaaH9ZkevFVI7eioGFWgzfQ1b0D
wBanRlfh2YIeZ/kx62isHHgmW8v1Ht6N78bQuzu8F1WpxtVq7x/R6GeMB8QjkA4nmW1r8lFctIgP
cVKQUuVR9kCsxjoHZKcb6XwUtbYf84lbLkNXFAaXRqI9lbx0z25fazCY0BoWDJIpkEYgfjD0t9vT
QoW9rbee/g5fa8SNRgUA9XZKa7A0ZyHjWu3JTCWbbsJlZ0We+QvHndq8skun/0XepC9e/I15OM7j
I7vCPFOXzwyCFA6G8m36ekIPU1SPNTeYxKcxpzK8bf8zVhnRLxmp/os0R5HvZ/i20nVglQRNeTJT
NT58ZpsoBSsl2kU0S84kbqHGAsbRWW/zjzAgp+ONdbp8rywldr+sz35y5L7rmyB4Iv2NwxJz2pK+
A6hUn5hCUfWxANx0svLaDvPTmaMxll/R8UVILTwyhhm9LtBA7HpGv6QvV3UKQpX+vpLrUfr2T6AN
cHa/9yBIwY2SGLZUukdMOuyMXxPgKZv3xGTxIZ0G55UhX5lO/eHVV9mHRR9gJZujwnlLKDYWGvXf
jUkIpsU22pg9DRTNxmayX+lAv6MNfuXFxTlh7uvPTttjVOtP4FzUj8bXIrbYRzHd8PjdWSnJbSXy
lgDQ9NdgjL/LnSXmrtX0CflE7UuEtt7VhVJEF2TUuoznlTyfJi3pOJ50dWowGl7k+iAc2tWqSt7a
9plRApQMYxFicsVINX14o4M/rzdjapTyOHW+AndcjWBbrmFQv9Q5ta/BPeF5bSWwM+saJQdMrrpo
aLVJKbzfG5Fz6S+26XFCOPftwMjOid/IHPesH3SF0dm8a7oS1lwTMfEKPa6xdbNbVGpva8I8XoU5
0Yz37cm62KF4HuDnbbAVLsktOMVltLH6KgMCdzavsfNYZhh69eg/4Yjo/O0/H0ygko7DCpjFRs4w
d4n9+E7rsK1F1uPtRc1OOIi3srsW1iKYITyVkuOcEvSiONS8Kk9W9f9FeycQ3Y3KwjrNWW4YYGgS
s7LRN3lVxE7R1v0Inx18ZsYTBjEzvsuLOwxLrYeydFN/e2SJQ3FfzCKdWim3KLEDVV36Xl6LXKwm
9+mmr5eKYqcIsKKcUWXkd5W/CkvxYmZE5HtaUljJ1/Jh5w05mUTVGN0wXDzXv3OgmeXoEvot6p74
YbD072FhIrSpsR4YM2eJKUKdVl4+uz9PwHmxx7mIB6filrZsoT6/ETMyePoNSo3qJryCsQOGGmej
muXqDCm4Zley13fmNwqCV7ORX6C7X4To1ZBp1z+umGBrltNCyrKK9c0rMjMnCUqB0UNkWsqviBxh
y4KeAK3doYIxrmR8XagDS1WR9zDjMaq6zfo3lpjwuFWm/NXDykbDlJg5kl/Z4hpvu3HClpdYJp+z
AzvZTnlIl5eotOQb1n75S6PkRd0oqKg4KZNh6jhTu63G1xHUXZN89yCNpL+Xq5spMJ6a/YBu8Lqh
6au22zcInx0LKRlXSj1oyKo02out//Ca/6WJ9UkjoQFQNbrXa5R4u29OVFM2c2Dnnh2rdH/gL/lf
TFIFs/7Sh8lKaQIFbjnGKhkqZ2DpMInOKPgheMelOyZQxenVKsM5aJDzyibafDcGKwhXdEDgK5dc
LnXSsy0xHlx6EsXvGgTxgol4sIEtf8czGxHBWymJaV3GU7C2YdtGmk2GLq30o4GECXu0sPB9vsmC
zoXXzb9O8tCO+jPMQipUtPG3sPmglSZDQj8LfausJyVrEMe0cB2khkS0cDb5mlpMI8lq5a5JzO3O
XgeYQ+LAxLhInVDvczWiFsOuL8DGFGqJnXI8j6DguwDvCtd4rg/ngW3uor7Lz4wcn60LyJ0NYB2j
BDELD3L8d1Roai3nIyNdWnHU1HYDsC4PdToxRBhWddtYycYvG/e7jmmmald1Y8uvnzg/QuYmo4X7
eAIRoXYO8Jo4NzwjpLHO1dbXGZfOnFTXvH5HrjRVH2msJlCRxXMhC7TrwAbAQjwD8svpoF3DjPG9
W9uEXaIXW+SnP3EI7EEzA0o6e6rdybDjtWkYQ3zFn4YEhrd5yIu3dArZDzSPRf2kRcGCn1Knb3qc
DqTnUzwiBBGbINsg4eHYZhokN4k+6W3YHMdS8JndL31N90zVsos9AO9EeD3Fk80PTYUFAn3zpDUk
/3rZHCzkmJ0+fuvk7hDWwTFxBWYBCbljRasrLektDWOybCOIBt2fRkakHTiYVVfNLpGzfZs7zkQl
Z8q6xKO9CvAL1qLDiwzwobGy3ealoGIvh4sMqqrxLo7nr6i5DAot1GG1Bhl+D9LyIAeXlMQxXEUc
9gFeQ4yngP3cY+UM4DJ8aW2ik6Kg6dnN+bP90NwFP0gmoVZa9SaWlKe2luFXfuFY/0VKpeDWp3NX
800KgU3XOc4xs2/JjmviafbthBCnqmqG93B1S21IYBrll3h8BtlK1TuAU+xReMomuJj5t7qcnEzs
tYYNIx19Z4MEusJAG53wKsFEBKRHPgFEFKs3Gw6c1HI3y26yMPK0RiHItFa4fACu6TY253Ab3A05
bfrTOxauv9+hrUEYTjijNesg5srUhW5uiZ2Xc92cvVoMxdZMZrXDR2T5mFp9E1Hw+DrGU7QHmyci
0kFSMSEHMT2CdRrx7ZNDrI1lMAwKqpzZEP3mSe0oP7ZursXQcGi6RBo4l0AoDEe/4ErhiP/uHF+A
/KUred3r8a2ytb6b7M2skVYKifs9CAhyYBlNAzgRJWCpG+OcBSQYmZeIuLOre35pHH1ieIxX7uN0
TATyw66vfG402sEPmqkW+zij9t/Mq4nR2kmXhCWrO6dunmc/9WgqwD9eWmfpD9s48y9/lNecP+H5
ZRJu4NbGGld02pFLh0iYX36XUklZgwmmjoNmzyI/IG7Si3jXguY3nqKWogNNtXe05NbZgyAfCJe7
bdUSqRDyXO1XZ7ARL3fzZ99jnS1eSnjlZVKNm/xs6KPDJ1btlLVRoXxQ+lS5l2bqax+wXXZO2SBu
R1KDMUeC9CfPB7v/BPdavOxHgzeeDxZgu+yX9YTZB92ZVnXJ0IFYhujkBIdsM36FaWv36sZ5wvVo
KcZJsufSY+V4gE876R5hXGVpjatjXFGqpF5ucNbMwUE8Bj5fIJNU/laJx1oMDbjprTPao0oVqG6x
11/OdkPHKmI0wFiE5zNqCDLZqXUAsEPESNvAP0fIheAIY+rQ8G3kKVo4u8q9edoPOL3c1Fb9Frbn
MnMF7d5anVaXp2Ri2gj8jRWyNuKEG06+dNpw10JVYAPaDYvdT8sr2mfVOwNLuF8MPzaC8FCtOn9C
7DmvQKiP9Qlpw1aSthIvnQ1JaIcmf6iv3NsfHJAZJvRHUuc5/kkrND8wUytEsfZzbJh41Ipvde+q
+9+SW9npqMGl4uMxdxjlgJBii2EfwLuHIp+XIQzDJvwRJajBPH+Ou4IGfUiVXD95RnWf7+wMpDHw
VB/INVKIl29iCH7X/6gY9vvL/nfMfGZlpDnP9rUeUUtZYh+r3uYenUuKceRVlSrl/vTRyzRGSfnz
SEf0DjKAKwqqsCsvGGrr+sochu2ttz/+LW9kXYLKeJFI3uQwhVWg/GlifdidDAT3uRV/5QkOoz5L
aVNSphDE4uRqPqyHPHCsY36PxaElJNf72N5J0YnYk5gQbQRBTacWASSnTtZWo8rrFxP5RF/kLgFK
Yxf7rh4sedjTeeKpO2+Cle3vm+rIXPZOW2BZIVVyct0FivBcjLfs4mJC4MZrEWZ5yFgmiwYmh0yV
7GxT7muBbWdiOxg4KmL5Fk2xOv5BHQr4MD6R9guMLoujgsAKFdunNvIvUpd+3tIij1vBKuWjPjjP
Uh//DE4jYFNzojUNGefIlgOQP4Vezl4l+EMmKCWwiaSQTPFjx5DSscFioGkDDWzhRbxEbe3aLVFs
wnBw5ZBHyg7/PzCveW1qF8tJxr62KUhv7pYthWMda8vBhSn9Tl7FuSAMgeLNc7P5h+6Disdmqx4G
pJ9smp90mQ9rUc4nBp2p1DeogfVfJGznuTxE8LR44DMFD5BtW2n6YtjJs4iYYkKSx3k1Cghmui++
rz+3tjrIwS5n5QdzLcMcdCqjGbjO5jeyFSlWJDAsiBiWVeinb5qB3oB4lg2A4iD76yf6U+gjInJz
5Mo3oUbNKkX1v0VGCgcgUvYdS/Z72qwugC0HKG2mZlU6LO4HNhck5nqOzt0Vvynwa+D5FM+R4+BR
WCnFmprZ3Zvybq3RrFM/xtH353Eu9aWxSypPm0HVjOhkLsS/Vc3rO+cvVN4KuMVFoaxGgQtp6hFv
ToWrHqRy3qcp+EhQqRcjqXW5gg5cLADV2rQwpd9E5un96dAbwnfu6j99XZRR90kNf4+kREIbT4To
eycONYDjEDzSSpTU9NGCyamWeBbJbRIErN4T9CplFbV/KnjLZGPJ41T8ezgYjvNqpclXMFBJLbv+
Ee2a7euKL7pMhBWTUnjg9MFqYT2pKMKAuy/EK4QfMrHiTMtaGTXBmfQUmDMHUXIGUboCvL3oCewP
NC9V5ZI8Imx7Rs4LIwCtSqlrdzF6qiIuvJWSkAROt3GdFKYjOdTD38UhyfBmG07dMVYnwkM9sLBD
SV2Xkyo/77rnGsodaGNJIqD2S1KhaDxZ19du+2Z234X+ySLMRPLs8wmtMo6mR9efQ/k0k2NTNgib
mQU5t9bqkg9h8F+RRnJZeDntMi0x74YsUpkNdWgCs53Oqcel/WsSGzZj3Ym76F7Z1+/yupJbCbXo
Z27BhIccKk/GFacOu99SH1tR/+dhZyfCgSWlpFUL/j4/hbXbAkfMgEeDIgINmUAXYI+pxOH73FtY
ucu0WzUMAOgjXZpqMviY/vlqBa2HxUeQiY3SZ8GiNX/5w3rEwdnZRv+R0c/u3Sm//55k8ctsFEZQ
7CHpPwHcQ8b23kRZBpH6qTc3f1OLF3qb+ViqDtXygo3Fxc8sK02Ucnq0GRBN6qKoPLOBmDn38dfi
mN3ods8veBhIvJaLbq/66OATJDAJ7rTV0bu2nKG67Gp0o2hLmAkIU+rNrhy6A9XRMX68TFa13fNf
/CKmoaAFKR0d37QTRKsotrNkrfaY+Bp66/P1eul1jLbZ4uqSDFpo29NrDlLB+rZ75bZAisNyp1QX
DABFTnZcVSgwwEa9IQqsw29RThJ+wq1rbHg9c/DbQImag1AHqwLFOKvi6oPu/J9jwvOw+6JPkMW7
MMnj7xM4Oe//DUiemFk3joKz0PhadwnIWUHc/YZzTJaIvD86eGcb09VtDqA8FbeQkJJI4FlmO+/t
OVjEA//BwDsgfkqvlh0XQId1rtgtp5dM9xKaBDD7fTt5mK8EdzwF3xgj8p4HJm3tUN6NA/60t1xA
m06EAg9hDUXKKvsAJzAL01h+TN6L9v6+GEtaEeMTc6UH2KDFHnbpqNBBg+X5HyRMpF2Hvhxy9HP/
7takO0gHZLpfskhBGvauvXa26mW2IvT2sqqdvxcMKosMDWQInMmfEX51jt4KS8EGblMPYZ7VxMO4
UD3JY6daUftr7ZwFGWZgMX5A2jyIlJHReoQyJOjubFXovQOXs/K6SwVW8v1Ed0XblpnDS6GwWxcC
Szz2G8iClQnsL5NUwxY1JCR+OWl0uPMTdsWdDAnBgGe4du78+GlcG2HaDbGRkjhSXAdQMBlUEOB3
cJp2La//gBjDct6PAucAONdoe3kz3JkIMK2fdfsU46cSnTrTXkpW/PwyPyr/8C1HTbAZFJvmFiZ+
y55e8Zn4pjJPPGYWsLLM+owdprqYslTmazG3gPoLmamnSQZXgnyQZnSYv7T8LTvlyfGWPJTyddcg
PDH4wdCraMqf2HpdEUz/yTADMJBVWEIRW78THQZiCFIHgEALNOMPiIQCS2JAHJXDLDUvFv1oN/Ew
Klqtdd5PF9gFlkKQp6qXYJ1qFgn6/ZtP9qW2yPiCJGm3GXRf2Cgn/7Cctczp29ApItFjKfwgBRw6
5fmdQoKx0gXp4UgxDuVaTf39Gj+SBY3Qlu+Wj3y3J8PqrcNUlPWHcUqNj96Trhi6IgJITH1iCv+O
fZ3fso+FIM5DiN7r7KylBLDwSRnEUKsrC4Mxwh8P2090PN4zQzlX6lxF0jP3zBeqXOgUYeCiFh6n
Su1puUFAdWWrrzHBBN7sdNkSWZgj0L+s2gEws373sh5aO87YmyzpQH2n64iEY97L5PCX2e1bQ2FJ
7l+duXHO0AHtXHppj9yOuOchgQNR1q97/Wy5N0GkYV+eSdjpshutWcAfb/snmlG0WJ9vBnNEsCQD
XQLeh0eKzPYNo4tF8UxRPZxy4YTo5/ytCD/dhFYaC59CEdJv75dQOt2AKM6JHYeo3xhOiC+nC3b7
cRtWw/whthFVxkTwJNV6YnjTLxpcfrL6QCkHDyc4wD8P4wy0ksFpYWGC7eHMcRG4P/uicunfLYT/
0yGzpJKFQLR395G1wKhnJ4ytZ7IR+jWZLG/bb1CPFDaJ3EVcjPr99+wktP81VhcU2NAmqfyDxDir
K7D5bgYmEOpgVU2ISB3agvAiJiRCL7cxJo1W9w/7so/ALwwm13HjBV91LcG+RBgAYOlF3G4n2Pyd
hNFYsPalUV++bdGhgkw7as8GSdIlQlnyqjw9228QftfhPWYCvwi73oqktOjIIKFTuXwrtQGRGS/d
smp9k4NWXleX7UVG+nFD2yrW+sCrUf6wjDGX0kHKGUNuS4HpSBfrqRLIWcoBisO0FJlE4s91oWSe
XQK2TJLchZynUNL21UajvgzuLwSj8mWR2/AUUEsbQjaDuOVX0MswDMp3pZp7eqndCZSHHD+b9bur
5pi9jWK0+tOwORDQN2bmm6hIoA8NMXQ1YNWXbEfN78YymoJQWuCLJ+PZJJ9oh/1BcuAl5E3DOilo
8F+35uuQwocfCctYSnw/bFnS2yuFqYeKOJ6YoLjVpXNXOy/Qcmd/G246UCUdBjl5IXTymLRK/niO
Fp9wb46ZE4hL/vdZJV8pb/lFVC6QqkXlwMHhtnUZNpJSvVpEThoxHlaONeMon+f7cx09hOHY/zCg
aElDqrpkA8ycqaqKYW/6A7KnWNvY3ix/axXDT0fSYzidEGvZEfUGdthjp2JUh4eHPwCvnXm7oNDp
ozK1qAnfD+ah/fSKLhpMldElxbtNcpUJbgTmxjx2XoPvmJPvQK+j36PXV0i8b8hrho/uaQEJAtzD
uTQRIQQX9IYHp4xohAtjPXswTa6sm3SlwlXM/j69mHREVSmw5x/33R9utw9q0BOoEhQdLr5+BB0a
HReMhp8/L78Goynw64UTQcCeSPRhxAoIaJNt2E64VBqaY8Wo3eS5bnvDTx5nkYt5aNqC+wT8KS0k
E/e6FnLvjBUQYZoSCntu3mfq3bf5X+djmiEpJ4swAkaBny4WorABbqoqKbOAqy3MOz1EVzUd4LSB
yOx6UV6sjLXa21qS+vHiMDWEdWRJzJT5YNPCYNhmvxPoQFBnNQPLRnU6El50UL2mORbVMU6aOS1m
7qIp7P0H7GUQY/fRdXtUG+qPh/0aRQqDSGt2zNk+OVn2Kj0MOPkhkF/WXN7PAJydj2gUHyTTM7r4
8yu1n0Jrzoe2mF0w1SktvIC1N5NOv93LpbXGJ7fy6Dksg3HfLmxYa3eL7PSVw1I0f7thGNqRVqz2
FnslDlzTaapvpbPk3QlXesD7mY0587E5Ny9VO6TNQM5hwExgcs3n4p5L6/Q8n8PYyJNzOLeuxKiy
Ios/u+rlWsxEzPC7Re6VE1HXVIhv4FkfXBBDtZ4eVMh5eDEnQqNOIT2n4h9jsnIxOFd8Tm9Q/1GP
gWts6F8gmRlCK0PBhqiZCDKn6zd96Ymzc3lYDvISr2wOyCkKz8bBwMl6yu/AhMMRCthmRgZ0Tzk+
vNGOtdYTBTMchtjweZJl2l+WKiFRtE5KiB8T01Fyl7DbQ+IZ432bKpWLNb9LOoaMrsER2hW9/seU
HVS8qRzmNNEGYbe02uvH5ss2ePvWTr7mCaX2e2eOGulOBWjz/aFZo5vXfU7aJ+gdNNOV7Bo/Cyou
EYFUi4aw3XVrKpOJOobueb0rVmD3vnv0b4hyNGFTWihuz+kNhofJwaCtuzGQRo286pOJpvfuOeac
OpC9kMaF+hvD/T5w/Eko5e7TiAO+0Gdpdzj/kv1kyz2lwTAb1Vem7lL+JXt3qhy7NbnOROjKgCes
y62znFjLHEOfwTXDRX1iJx282M4xUB5KGI6o1eR+rIPshighG0v7Vh+UNEi4/1kpGonr8jjTvZbv
NfKamrgjjd7Cw87VcrgoKb9D/AKueg4JReOQLuLI74KENT9J/UUp9SAgYwSNd2slcKO/EskeeWWP
xwnk3jNsqkhYsMjNO+677RwePQxgrJFL8HsyEJBqKQ/gxcB/j02yo0/msX2kev9cXeUjw5WR1tmy
4yqFK0/fbJDLRam0EjmXFleyPqQXTWplV3zxTcLBOJitsTVMFlz4drUVAh5ltt/Skbu8U9ziY5Lr
+EI9gql9j/P5gQs+squnxDtgb1DlJetqHLMQxNLb1Hiw29N9x+1dr8m5Ugfj4K1P5qUgW7ScVFB5
MuyXDCyX5VuBBy6RIHl2EVwXVMFS5fRR5j72T9jxJBrGCrl1V48LPOqPJzYTP8bwP+r67amK4Ax0
+IytoEcnpJmuC6r/z8AiYFHHgAnh/q6sMYyV+mwXGgvfOpxOPC+SIO4FbeG15ILsJxuPZEppLm97
uSKvBJilXF7qfc+CJSDmrPSbCq7Rdv/vU2WviJXOljrBNSt7SZQMf3Dh5lbX+2HCkCg4jnf1M0dh
1z99mpnJ3h3zpgwuxVsTFNouPR9J/jBH8LtBUyOUuerkJYBWIytHAEyyWYmrJukWKJmRoIUKzYvg
7c0mxrga3kvqwuzrGZ4Y6B+uU5E6klCSOAanS/wYE28Ig2ckX9r+bjQraAwaNz5KBusJxecKLF32
Bf/yfB3l4svS8FDhXqJyqxI7OpRnvTRLZGAvWsD286m16JmJxECvrYAS96jbIMGxb0pKagXJP9CI
yln61FgXJqqx1aEcj9pDd+6uNuwTgE2uJdThojOH8WxDuTygLVYa3xOb4PMiytSrij1UsentLeS8
NOeUKkQN/cnpYHVca7gMBkeND345BqF7Mh9QdvSDiIicUwHss0DewZI1023TEOn8q1nvIrBJOQZd
0ej65nzOS160RfTy1GfvnJRBpmrEa9c6/IynNWJtZm+FWsstTvFTPqIaYQrTE+r53EtkJUsk2NX8
9H66MRGLfGCaaIaDUCsIzbU0y6C7pFIB/QmLFuRbr6C2/XdlIklY7UCW3A5qqUPkuRXv7KWcEsti
BsvwsIWttXS1Pr3z/AG8VbScGN+9plhaAqHRKgiXrCQqj5eVNXiuFEm2Ba6SRwszBH1kEdymHnG1
yMQazOTGCnInWhBP4GiHoNeCKFgxg6ja5aLB44duXNJX/OxnCbCzyOKBtJLUI9XQm/7QYFPCU0El
3Q2Rli6vYf05/uGe/Lim3+APoTUn2Gm20vtRI7HiEfu+Y6vf+HQasHwRzUTXoTQSVfl3N3IgBCAT
YPLJa8QkueJfV9kxK1Q3jtql1BSI0qvRGA/wt0d8jxSsoDLZJzTfByc8qN2h6q+7MVByg9pV3At1
xfOdjpQoo8Fno3qpfWylMqzN4bgCi72n6FCEEO/dWAgmSf7tNAdlL7iP/8ljzC/3NC8KA7vyWTiZ
WimI0TNvRetXg5CLzo6vNo4KQ26YQ6V3pJ3luM/LLL2zTHtq6H2QvIUSvffRS4VLGrTnclBDu4Vt
XpQnv/cyW6+4Qbp9TOYkn2TvgP2HvIf2KEvGekqWNxcZA8BGJwrfCklpglXBmC3wM5NlnnawdQAx
cw3Mv7eDczYcIeu4kPNrYrrDuzQObEkYMfTq2WpEMT9N9xE+88zFVQdpFOATU3mzK32cWDPdICOa
T3Oa8CzSwbXx4Wv2X25jXANMaR74Zrt4ZJ8Ag/hBMacoKC3sUUPhi4qiv2a/hVEFPUXCP8uEBvxU
5AQgV4YtTPOhkrq/qmgjPk8fT8400eL9/9M8EDyfIq34Wy1Mys+NnkrQ9etZEEOSUB/qMWx9re1V
4cMFjJyraDAVBv2SIYs+w+9E+govfjVmtZOrzmZiY8SaHp6vM6Kjy4p9XNAVd+0ml0H9wqnedkla
Y0IEcZStEMmgAHZJ7Xfgi1YzSOi+E+SLQ9hOuxK73UMJfFLMztT/HKn9LH5oOThZuiYm09+87jWF
/CiL9JAbj30sTkij2/6gaebELAUeipXn7Cy1b53GtaPxrlQNjjhIveQC4aD9cPBR5BvIyzK3YKC/
PIDzTIxtpvSD13ZxeCRGi89pjyioBZJMOrSYD1uACQAEIvYvTCyclBPTQlQDZB2jWj4A9VAYf3jo
rii2eLmlFpgjDsbvDteqZWvBarXEFDfddVg2cOah6rzsRybUBwwE42ONkcktluPdocStecu80WgO
L/B8GMHw/scJHGJfs0wtGsTWg0r16Jh9lN3L0Kj1rgtQ8EqgQJUPG0h6vVf1vIoCdRNDXX1dJq1F
tw/wjWvenBV9JID2S3GZ7QoZTB200bmxdkRik5khSW0LrkfO5rcIg+K635uWY3fJcNPt+fpZsqBk
9NZmKWJ1zxR+xDaczltXG/R//8EuXF2vXhPZFt/q6r37/9PCbBMFdaqFi5+PzD2L4btitOp8R6Mb
5FqmJMDntpGnCpf24oPboLG9MQIIVuj65i5/vqmoXIooQErcLnVacgOfZakKAwMziNG8a8ibA7m+
4IqCIDP9c9T9bODNRw1HiQ8EYICOt5R0GaTCfpDWzErjNIzR+r3o6NIMKwcX1izI7+IABHb26aV8
a0DvOrzNFxJR+UyVK+Q1KpJvLcTedYpTz1r8RJ0aEs7+l897MJpZ9YFUA1tTqAOQKAa9ln/BVzvW
GkNZCKUtJXLXcyx+XJe/bZdL4Bu6vYEM7PkXgwlqt8dlfWZfdvVAx4KY5lDlRT1hxHVRhc/5zj4y
DA8V3LntyvnwRQdFlDc3vMzI1L7qTnKhEk6kdCek1nmvkLA8jCSi8rOHxkXQvf0CoPuOKL+8ssc9
ucnRVsvDxAZBAWjlb2m9UCMitIh8i+q+piIYCeilk05vzMsT1AGrt1PZOGje0Z3gbocla5x41c79
Mg0aAWBb9KNei9wFTI5Ym12AIWojzGZxm+0qXiYy523FKiaPs93/9uWzQ3UFM5YPVgSd1xtuThK4
QRz+PbU3Xdnj+kd7p2VzbikTikky1iglIdm5KfTXWzUFHu7O+wSXJ2OtCkF4hNMGamstzKtW/Kj6
0ZYWG5RUi/OgEW+jdsGxwhyVA1p3+K6M+P8C442tBPRXbIBPqnq2lo4fqhrGijAvPCnOcFUrWVt/
BrDK6gjo9nYmjwuGa6sa8qtuPzfVXLIlOQyYEnxVvRE43glscxTkCbuKAz5ntWM1agHg8JN7qbm/
J9WtpgyHpgCbgMVMIPKILj9AssoP6DdZV1ywrMvPQDn+Wd4x5glTr1On8Q8qNBLUUnqpy/ZcFeFD
IqdO3Op4jjOhUTFDBdo0hkzS7ILJHUojlsWNOqEO6TEvvkcCXoXxT89JIQeqRWc8FoNYsoZ6TPLR
yon6uj+0Upi02NnctT083bnitAVDzgGJb4ffk0yPHxwa91uvB9GiU+t8jueYRCel8IkBx3QshtqT
pVwJIPK7FCGHbH4lu5a/I3gXw5GBs8mEjtjQGqMiLKuXxdTEe3HMDnnVzCNcT6jIh7bfvAmn1L33
4GYKNB5w1cSzng/MFBfHgdiZnbq5W9VkfVS3AQgfE4dXTziDmufyFmScXRy+B9jsEmM2odH6y/NS
oJ4Xd7ziQsByX1FVfauBaYHB83ueDkwxF5lkGaJOnDrOAFCuKPBVkDtiRQIPuXfm+G0WQ+seh4eW
x53NnvUK+HY7JqSvn3uYBOKu24s8KktTRTiTAnidyuDkjOZdNTAMKacWsCkIM9nJNV6L6QuHoAlD
BINbN8QeqUoGv+BsnvpRXW/OzRUAiXOH3T9B5/9poYtcGQJEFByopCu2Ut4wY/7qbQ7FLWWjWvqR
MizCGza7Mj2NLPvAZcMm1hNUVOx1NWJM3QDZR0nwMsYGMv6nyTTR09eYFQNOJz7xcRiLZLpMVjEP
3aCsN656DDdYj5pajkxyYBZuxBl5Chf85BcjHyRmrYFTcxhBzZ5Jfxw+AcM9HuecRIo4mv4VcWdV
zcvAcNx7IMxoEs4rBdRCIeSTYM2wvQbLI94eGX718k1EqIOwRjRTyb4NceXpWW01ERK8FkSfgZSm
5sLvnMscG2ZyzKEIkurztWHi916E/EL/a/jffEGeC75O34SWlwH/N0qR0TKVS1K+Kqf/b7aWvc4V
8BG2qYYfGHbUBgqRa04vDPohSwYt21ah1fYlA/a2oMveJwpDgVEKq3RpwjYgwDTdkZ6ifJ+JQkBo
3ZgFD8TUXPSQW4hV+aecbPmxk//1UeIjuD6X44D4Or7Pu1BiTjkgTyd7oxdSmnS8YHMh8Ng22d6C
BOQgWzFzw+UPf/QFZ/QN9OgICtjap8GWsIPxVgfTlmdmxAq4g8nl9ueziNGz5USSmDxCSwcUGRNK
trHwVldEaiS2jF/VXVIUJ8yiqo6i3d3myQdSXk+8tOrNA0SOBsA7Jmq6kXIYfz0bGDUxAo7pDtD9
O5InLxLznYY3lTozV2Ie9R5bihpEcogS52ryWuvDeBfpPyQ815sR3t0dN8R+yHY4tUJ64b4Gir6o
xivNYGxd61T6rQJ4tMufpJRrkHWVj1Q+8BMnoLWILjrRYqr5zW+pE6PbCwyJeVsVWkgHnG25RV8W
K7p2djTQlHoEuzLz0w62Fzp3szTQO3B835+zubDEnFuvTPhfPhfz3qn80udTS9jWl/q8AjA7MMeX
wOrWHc2NQ6SY4qOm8QMtqpXt9BAoGIGwJacuiNhsrf785rEeT7MhCOxViTC1iqYn4zh5GQkGiEf6
4GHPd7OkreSXNhRLPjac3uP61zv3gj6GLi3G2bxIrZEr/zYFXGgzqRIEbMcnTogA77Ok0Vt4eshd
MsyOnm6+1SThWrehX6yrmP9a9slu0MTr8X/go7otYXdnysF9TmpNlwiYRV1+3l8sniXnys8KO8ew
g2EwrJL6X348YPbCIQbtM2yEXgwrYakLh1MlVBFyovP8XxibcMz9SmLjn2QnHGLYWPgtumZFU6dv
kq63wo3zw2I3KOQ55wCDwEeEj2/igk+bgLv0DlmQ376WxEeZKH+1qf5du0XHAq3eLTrNgrICaOEs
H2Q85sqe07r5zbcF2d9avsB/fG+nXqKjOWd5o+4KQN4rUAJXmi1b/opdA4O70W+SUwqrGadTpung
VCJcZ5lpmyLvFvKAy20c3r0BXabdL1zY9weKG9N5hd1Zp3tl9djO3EBZ7uJEB41u0mn2NKbZY+r/
z8uWLPn5su4/8ozHAItrjT+NO5DjfceUseBoSkG1AZMkq6vre7HkklSpfjm+fs032T5JxyK31dc0
ndACMu83lNxy/4mqK1hFXpUV43qHGq2jrQMIehtQ/oLgbEihaSXRsHvQrnDIER0+XrxOvdSbxG8t
BfkRSbbBJAS+9/y7fKXFTafsHTJrIlfU8Gyvrm3ZHXaehqww1EsEJNdfEUYPYancuiLA0zAg/t9K
kICwYMc0mm/exu2ugLeEVOfFIPYeRd28ssJENIBYLCqpttz6OSmtQt8U4hrxBuLUfNwUtec0jnxS
9RL2b1TNczi9P9N4pKNHyKvcghKxM09HemcHbu4bAlz4lwfLvWeBbtlbqzwjbmNzXDT3kgVpl5ap
tRBzuo7+jEEB6Ki6BxkljuWgMgSVStk0NyXqR6UY6pzjZM/+D/Zhtq5jRdRd41sxXTMmNkBa7l6T
koAbZvQgfXRwDAHQT8AGPTd9YeBbPnklVhob8493pYxJamdfKljjkn06outrqYyP+EIq+9pUMFoH
zDke1W7U8YizAqrMYtm4x/NiYGh9ds9JT9xIs02l/7zPndIJuGxMqjmMYZiPQ/Dll/M3/G1actum
40aKs+MWhTSSJSkqvkKThV4IFV1VtsTVRE8n8FHe7mGc8612n4GfzdeIJGzfnGYgH2ZMQcAE5WuK
AdvUL5uX5AqrganI+qaeiamgtWmQz6FpRWDU5RrtovxY9rvr7xYLMO3ucfqJbTcoPjEzJlQTiigK
A+pbo3G0IM+QPt9VIL3MY/4ArV2HGEtYnr0mFZJBQPj2RRJ2jIem5aKWy3tnbeKEkBlrYkzUsgBt
hyMzT9GtmBgf20MI4ENlJBNMmZcJcskNqS3y76fxQMtUQ9uStNgXZ44dkVcKsN4mQ/hKm6deSvRo
+rj143nhlx7bMIzGg2l0Ff4NCzzYke4WaW3h1/MLY2yJhPb4wK1m6nn6WF7G+8M8Susv0pHOkHWn
APMgtdqaDLH4VGL74LUd7JnuV6+MHg/r8MMb/LeFWoMJZcQ9jDacMO0ZNntUBZZJn68s5NjK2Ocd
U4K48c2ZyNzuAQT9fzT6lRe5nakKLhdbDe6jhCWtaFx6RdY1Dyc5mJWNSucYO4ur2BQgi+p9Xv3V
F7X6qiQlQCU+OIXtcbxzSWiRHyUd1wL9ATT0Q0DzkMttgJGKOOi1JStUX4ae8pKDATV3drIWwAlA
2h65j6rjR/nuDFjnLIFe1PKQ6qKxR8LWqcNP88cA3LLEWgDskw/HtbvKu/FMDFnF/AIqQ5SATPA3
FuTxlZ5hf7B4x/+khp8zwDPnreBIZWJSyS+00Ru6VeoijsCdsQLnBS+e1vIehCwlsmUlqhTXkGPm
eFUMGlLF+VgTdrqAZfzKc7etJfBG127hdaWaBvE9dX9Q5/lKZgHB5d7pZjQUzxZNkhk5Gwce7tbC
pVEDjdL1wBfUhgHXYvagjVa8OE0SNbNSkbMkmu288Zu+p6JaCfA/mwylERF3fRbLETwyi09jo2F7
oaEZ0VlbGrLBVSdpdwOwpYIq+BHVVceHVVgluNXB8wa0LEkckeXK4AxiF0tsF2Ff1QcVSfuyhEuK
qN696ljwJ3oFmQnhKsMiclEoYLRc3nubJYyxYbace/mcE4WfujLhELb36Uahih2b6kf6vXll0buu
H5Qnv03KQNpcnTTjP7MgN6zMLeuVqR9ztNQ/EWVtTXB+2rmHgjQjhT4rNUBYKlp6C7YwuHDGNAYU
yZmtRZ29CW7EFnbERx/ejrUdjOjuiJjfM2rF13bT6N7mini+Qlf93lAskExGwgbSAPavNecPJDKF
AW6SUJthmJkWEdEzb1CGrgtemoP5mbZg0BL2DZSTnJsdv9a+bLDBqcMH8nmYAt26ll14a3H0mXlq
rHCPsHQlPSuPd8LzRdhwai1RLZ6MmB/gwB4rdkXG+jrLPAWsLMQtkjIuCqd63uXu4UHqA6UTuu75
EvnKTiOW2PJPjDHr94w2AJRZpkFFVyqDhewN1j3W78WrDf7ULfPAuTJBbhZLJp0WdJYLCqtQxfjz
4f90CP/GQdMY1LJJCj/XmReFEoFxc8re4KPsD8e6cmI7NotZSDrJ4yGFCYaQgyW/OB3uisnACu7+
3KoSxWvYRAyzUKgykuQIUvVg3EQuQyn7x+oCAc9SxQOXDoFe7c7bDuvXt/HkBshaQ3l4E3VLMbFG
XdYDVWwXjpL6e1AzDiMm0aVHdaPhAoKOCTr4KXbfDkU/WL69Yjt6UllYrEm/73dwcBGG+iPhzV+K
I4fze+MsmTSAXAPGpK2xNqtMLuPpYEmcdnLHw09B7ha0hMzaFByK9NpoxcdJlU3SMWKLmFReYtcA
MEMx9xlTrmzbJyfs+0EZ+nVNb6iWzsjqhc9JjP4hm+ecnVvqUB8zVpSNXAbs3WyDNuBaQMdcatdj
m8p9IMWmXBbDp7mDhGHGGx8mkvmqKSHj8ncHdh2mBWvm1CIcwl2mjDIcVQmxQxUk4A56jdLNTMLX
8pghTaUisttTIXhRKqlzI3wCDHg3uBMihr4Yo5g3I7KdGWY6N0KXtJpazZNhf7d4CPT0Wy8GzM3d
47sB0d99F+Q6ExAHQOFzlWDDnpyX7TDqBD9QqWaqp1fb2thEEIexBROXMmlxxgzYtH/T89sM6YtB
C12WXezk4VlybRrGnk0oyTwqztytmMEmWSia7QHIZlf8hdJsSF25U9VjLC8GKn2dzvGgn2JzM1lh
k7pvgg1dD1WYMZVYd0/jEMSQPxHcA9Y5/ty9TVjsNRcq5pNABs7TLwUa2JBOd4JzQn+2QxMLgfco
JC+7YewTWtju+8mdn+DUSh2IGxAlL15AePlTTffiNGr+bHq7ERfRjVJBEp8rFvb9frtByzr3H6PG
KXyAAh5Lsu/cRmCp/jaoWn7eXFKc4+zpGINGJFvMbLbU1O1d7pgbEyPtCVrUvA0FuwUvPrafRJTL
QgLjjSIho0HZmj2W1OwxccqmVpHLI0yOzfijh3GNagI25i5t3D2wjE6JkmjnbvrHbUxOOk8qfVT9
ekBzvq1TAKRJ0YCZxP6xGwXYCBCBkB1zGUbP2fNbUojA/n5eU3XeoXh46VSlFqbfpIu0trD8ISTN
6KHcG/tdplqvpY++tyDzO53fKqJJzGaxjEVfjLdeoHAZzEIWsOxrkB8ug+N0/fbPLFCvq9zjDJm4
NN8DB38gZ8iFrMGPYK2ujDswUQoQ57K+b4vmSB6QCe2iTOcWXXzygY0q4LacFvqpqJ8wLrYiJbPg
QQKsX/JdiDe+xyXYmS5NKGq1uwGv5xmN6xOJvnIwu5RaBnH0EEh1UNdhOST2eD+KnrnaEmAveP3K
GcjUwRKmB0F6mDV4W9OfJGQC65GiJJ3u1Zq17Oa8rA0QpKGP+2hL4MrEu4oAyL/fu10uInUwo4Pb
E3gRQsmduUO0BKvztT53jXPixw96EcwSeBKVyqG2v+BLICU7jKx3onVbWSZ256Ty0Hv73w2f7A6v
tA4jRQ14JfioUJXVgoow5SuOe7yJ7yQimBMoq84C/qKReuu2zHqaDIRfz5RMXV+jvLaABPJziqrd
hHWWwmsZYKd0F10DqngWUKjrnapcEj5NOS57I+A+wayOSu89Nb2l1QrLnfJqVsH0CsF9zpfgc4pd
jQ1s7WXNBANCR9zxkNugS3cRDu+izPLxO3uQkiwtJZE4QrM+VXmFr+bFHX/TcL/lv9EZdBj21cDN
BR/DpHc8KCoHvQCOa3cV6TKIR7sXcnAfEFt0On99mBJ9sIZZFg064LEgEOEyc3Nh/VcULgxDnWjT
AOluAiJHzVsPFYZmGvoOb9ZrUzVBQD8cGDgysnTeVtBTx3pZ2wERTcFNC23jntGR4NyyNWYE4mKt
8oIE3AoriF2DM3uK1jP7s0go4ti25J5rTwB+LKhWiK5WTJoyambRk54/Hg2OufZXn3VlQ4kflxCe
x92+wqZnaZjbudWdmD/orFj2krD4ovIKztzcIwDBD8TeSRA5dCSjzn1cZs9opYvlFRGxWWtu9sX3
aGmO/NJEKKM0qSJoOOEoENEhaAkUf3MLZOcG1J/0ChFhXc2g24fFcODrp6MjPunV3+KwBYedKJhA
cwJhQ0Rcbd6oPZ84p4mkJ6IUeKDn6K0LkKknqtYjf15PIJZuQLJGYogIr1jLcAsFR3/zBCCvLVpM
xMNwAgo0y6KaRXC/1uxx2Vg8R6LqTQ7HeSeoWeogVkSPSe8qIOP3G9kLzkjlebRgcFjBtpybcllf
UaZbCc8rbZTaqHb2z8W/iANG74NXGFPMeKtjUfkuiiBAXYZYiKVD8TfADWug+zUcgPnMABVh2eKk
3ETUJ9B+z0rE4/EqxZC9Ry5SS+yQnnpmAdqynNah6/abH8vk3eQgbCKcNhgntNBW4ouI7dJrwejd
VaLHbG/11TqYJ6DkLuECrZG/MwZB97Pf6pi8Pes7YxL3CjMy1Ib6PFPzUQe2TYS7Bidcwq3unUBc
yWZW18I2XM29kRHxk3XCr5Wsa6KGex9TU9n/ypFowIAkuJpwqRl71RKV9pd7vOE6vm8fwj/QkQgl
YJijM/kUZTq6BA6OkE3issg9FZzM2sSus6EnqTgW1SFR5VwGJOy1YL2EYP+nuNVjN3Hl5VIaAWLC
5EfMBB/2+8i+T3oNN3gNeSx/mrtqFet2UBpBEUMuHwlNdo2gFFxVIRjRGsfcaJOv0N7fFOdDIt6M
tyRYdQmOFWN3lrs8Oe9K/PEvqi9ak51heXyI7f8gv3vdakMYKywIlmaLiWd1pkMrEvnf5VweoAEh
/dT52fIRHcQ+p8x7MNcPWyXM8do570SfGL0j6PU3jWy4ojfGvd1cIjdJTkV6mahGshFyma3Eyk6A
FXA3wPRXYPOYjMYWhzwYRPvqNTFB3s0sRvlI1uWggoG4nHH8nQxTG7i7Wjh27ceeH+fPyFwwMdDt
P0m7eIWXqmtV8+cSCjnFJXPBi76dnGKGNQbppSrBDGlrDieNjcUt/jCD7vCeuN6dAEf11KZY2X13
Zz3OaLUTxev+W01a7UZJ7uYI2hzz8WGgRp3HQXOJw7rk/Ob/dbOFfRCcpueS8WXZH0FtTL1loEh5
tlAinEVpqxqqWztMIt9SRxN+WcnFkTyyPo/mQnNyCTSisOUFqkuOYiN3moeXJ8e4cRz+OgQQpCqJ
Yh1+E3qfZre/Y9nIokTOwaKAG7FcUCHOePmqogLhIgkH15JqihxoAGZWgKks/ApUl/JkroXmVVJ3
739TAShdo54uAzjJY5TDXysEfUmA2E8wAl1yh6epry6M0Q+qK703PTv6c32HMIFhI2So58mTr9XD
ghChNPOoKySEvDB4zJSybAmjRpZIn9bcSZkY6QYD5PUKLInC192wnOTc7h4cwxfyZ2G5y3zbEdyA
ImpkC2Qcj7LblU0rCObKkDJteo8d5LIR3f+K67ieN25CKRmvGu4Nlc6lfEYqTDWl1RqGZTUG2cMN
4MDtPor9g4iitcz7MWCDGlQqkRSmjKSs6l3lFDExali57cXJrMcB80uszYoRuZgsnJ07UhmRsmQ4
xsjc01KSUr609oTHCuCpEOeVJLDDSsEC3tU2cFPYm4wpLFadcYDlXCoikPb3+12AldIMD8aXajM1
dpcfg9hCz2iE9GO135Ny7mfOoqYEGKaQC8nkZa1AEJU3yGCfYPCCF241tqO7UPX5/GYT2vwcyNsw
hPGopvfDSKdt20j4BPqHIw5uPMOl5w9LfZV1s57p5jK6amzwzvpayj0YYSDkxh5IGPAwE89j9ybi
0S65YbFFdpZCC/XIVTeUUSkEspoRJvbPK/pn1DrJaTg+9NCbraVfSIeY/FvyUstmqWIKTnTX1opB
KzPwugl4O0A+CZGHy9lMZyTdtl5S4U7mI4lfsdr4tBkKHDqCQLXZFC+/s0jEFYyB895LGkqZO1Kd
leCgzCc4Xp6FvXAWSYQjCiWpM8J+mBHYh1Kemd3IHWJ4CtoFUOmORiXx2hXMupyr9VA3CMIClKSD
3ek5jDZ3sADxw98FkL7Gkrjcx4uO+o6Ck2nk1DM1Bt2xzNNxA6gVWAYHHmAvVJcxUT8b/4IqkVEo
5HYhh5yfKiboCv05t9PHeKy8ubeBJOB4jzP3zu0DcgsTzIwCaFzC8sUxtRIL6BZcFlXDXOp54VJO
HRY/yxoTUagKJDdmWPJtNZovLtyDC/TKXujkuyzOLwczxbZ8LosDqsYnO5MI4TqgPPPQc1VlLaEq
GcYkiBDr4Zf4yMjCDpJ5eg2H4Tb6pfW28hBqqIPfKtjYWWMsX4OU5qh1KCZ9m/V7DId83468kBNM
4caMtvb1fwPmoZJfVOZCA8Ki2Oi+NY/vZjT+B0NkYxLsxnf+cKB92YiDWC4D1LFuG4HxBzu6477U
tZS8jx8kqo9i9Tth2g5UNOMLvUcNsqOEAqh3ZW0oCDwiNZPpvHKw3015ZDFciKn/BVAEgCv2Zx4G
2khT0qgUlzcYWztXtsVJn+b1JHGxAASyRgYpbi/HGKPknvrUJ/WO53n4NLHCT5a8UBgkAYmC1g9e
W0JxiBTpxsHldjOQyHS3hGqab7Xbu2IEweBJblYTbQ/8w5BVElRPUMHMejlS+PIHkl6SmDj7r+W3
Uc7xg7s1LbsCtNn4my/HXGPAjAM1LfJX7IkFinEkAhmZ2/dHj6hjVZ3aQIw1/taVf+z6mw7xyzZO
ngyH8FmJMdq/pJ9TPNfomSvldk1JO4ksfldfz5tyOeJguLT9U2QK0cgjWRgabQKTE3edarowl7Ik
X5dzg7pLvqDUG7HoMg4fFRffgohemtZRcroAwLjiYENueYS6sx/Ce0zMg+wfQveNA9IKjdl/uX/9
lplprGM1pMkuoeH3yd3C0w9syv28CiqCTGSjNjUizjxAIrNtcBiOc3dea0a/GCkcpFJZL14ht+Td
pCZDEscf5JxaWVCV7VBEhPf1ABF72JKs670IdOz+fMgXXAiWEvjlt4HodSJeE/eXzB/AOuC+4ayT
sZiwHD+s1Rvg5nlDALsCdKyVhmbvSJgHbDp1eQdGsK8J0tc1krHUIv57NzBn5IdhVLMnT3ycJxr6
uwWDlQ04yn1dNZAhReva5E8Ux5Fu5I/4bqk42e2KrPspqeuEZECKhXBiglV5LWYTXpmWbpsqGOgJ
xVLTuZBRzG9W8Bngcx0PMmNud0WVKvfRS/Z837D/fdTpAJOChtaWGp3kz/ve7g6F84/z8CffsMjc
WMu2oFDMABttAIfcMWoy/yckvOEoVaFYE3pwGFux6AYgVFldhzO8la+U6oEzxp0yISuhoyCIpp++
6RFv1n9h/39kKbBlUajv6t+sH8+3l96mwh4z4m+ip/0TFFdNMHoWRAqgdXgty8fHVgm/kWb+bwI7
PIBhLRmDsrZZdjamas5Tj/Kw0Hk/xb2vgquWHs9NKgik1HVt8vXQSV7rkNzLXwDfeiKMa1BX0zX/
97L18gJVO9/HW0s86g21QPf7hijwvhMGwh44o2woUKTF05oTDnZ+GkwA0GWT8E691r02P/W8KqJJ
FiUecOnJ89m+YvIvbRCR4uHYBYleRal1HODlcWFAd0yxWlT9nQH4ZawmqrtMJoNbp7oJSLscTUxd
EnppQVI6zjT/4+k9ilSHvmrmcTrHQ4LCvDLXDFKydVdU+qutZTVlO8JoW6XEY0OdHDcTW+XSnZiC
YO4Q0osEANmt7tBtBUm/LAgpDx5vck12OdsvTOaY3583u3lmqEVBZoz1GywLQEA4uwtILfToSTbW
+BL4BxCd/gIZjYdxrrWFHlaKXh0NDwdGZIW9a5mM/fG01GSNxu6meqj6o9L9CNW/BIOWs2ckkYEY
2tLBVvz5PJ58O5+DOgMqRawiY95TDCpJc38yMGob1X/K/lLRoNjsRU+eavwOtbXezIzwvrCr6ZRr
hBADZgkn6jBpjDcMGC5NPlp+jsIyaANYyv7MNXQNEDznGtx6UjHL2usH8yCGRolPgs34w8scb489
aweaY2adXlUeFGB+1bd2Kamw7yNmUFfhy4vma5UN/2utXv2ecBZ3ht9cCE8epkb1MTJQ9xKl0IQn
gg5a9Z/aySK4jwUBhARw3jyDpelOqKIhSoULxDwx6hvHZqrnPumqER0zrTwDzaRsMHx8AmLnlEpQ
Yux3hJXawjXpN7Dw+xLIT6bJypAsfw0wXXE48EWT4JlQSu7IAOVFVd7d1bAX89XteQUmBJNyGoG5
dJ8LkMoFWbrGdvI7bT+oGsoszSc6DORGQp3lDtRWqRamwqwg2d5CQt2eNqyHGE0/IbY/s1sAck2V
nyroG09xFSIrZdzFXEI2jY71sZAfy0qLEnG1tBnbZd7coNFH7rVGX45rdET8x4KctkNByPkdiba3
iXAOaS1F9ndDnnccwfAOXEzt1vsybwS+bJRUdXW9weZqgiXOQ5GqBPhuGONNvyT9r+8bFkOgT9ae
TefpynkkQEvWGfLn5vjLYAsZX40SO1JesE3N1RetOus+j24za6YH8ephlCTEPUzk0dSYBwJVIMPh
Nqx1lIO/BnHFx/c78EH5y26Yxp/KRgw0evy4V4UfkGxW2PMwTdaQ6RPbSK6X6IWf9yR422CAgOFu
netPKJ66Lo+VsJM+WWc3cT1J5YeyT/qOfrJdj3PVboJRY7HcJmV28NPIYkxNmtM5uPVcqINE+hN9
Vz4Tfjie+LFtdVMFc/m66cacVZJV2L+edArmfxKN8/CIPpc4eV4IR3cRrHhn8xIcwkRpyn4w0f8y
n62t0CQdtmYsCnNNEpfrG1AFmUebXSK+LvGPQ/28VDvFIiGmEiAOcFPDFjRKeS8FLs1ODoCCE9ua
vmriZCGec6sCO1tIcd9qL0gmXk/eEYM35InFqCX+grsZDDn7NwcBRpvSm0zIoAOv6enOUBPdR5l8
8fX7KD2T+SR7vj0jl3gAMPj6zX5/NzaVN30ZG4IvhJhanRO88ZKL2g7ovOTsdqFEYIRxNpJBasA3
Ndn1eOzBjgItAw+CE79OYTMJZdyE++nbdkdXGFrd/AwRUMkMKPPDqmxsTHeDuPkU7zpcNGe7KREY
/ak9IZN3w5UJexAR5Hlf2yUVPPXbKy3RJtDXT9nQqZkOoyNvWhbeHbUOkdn0+mvruaSagQIBlxYS
Goq7iTUEVazlqXU2bqDPHQIqrRjnVwXi6pKeOMjiKMvaJNFVYxzoqUrj9il8i/gXkjZ0ZZsOjhfr
SPrTj5jK9t0TGFgST2ymDURuX5pbKuwfFi1PrDXnR8obVRFBpkgVmhktF6D9ebt1fQCEeg+owlaw
hd4NYyo7wfm04Xz0J0py7iv41gjixonqP9rsi/O9aaKnlrd33NbpKQq9eRu1Qyy2jgtdICInF0HJ
V6qbQKmvxhryHSJV0hYTcDhoahikkwJlXttf+B5nDDttksQNrLmJ7BXsLASqnpB7R+TQGlqQAT2m
bsOe2S54n8kmmpkaJJnkfCeaYnFop8V3bWuqYVvyRmvlesQGFpX+hICZpWj9rQhk4ezl24ehP6Sx
NvniV1zKGtnXq6ezDJHiUeGV5+duDMtrESrVDPloSU6DGjMAtPxyHXOZemDnid5/YXaG7jG+Bq3+
YpM8d3l8/5rtuldXdo76h6moKfLd3s+6KsBRll0FX7iqwD8KYjbE/VAeoPW68rBtgLGlRvyndhIN
qJ/F6zQbEUKsTGd99+JgLjxhp+Q1TCqN083tnrabBS+dthbA0dm2dsBsSzcVKdJT8uGu9HGqxWL1
rzNWaYax4luBrGSMUk+/KNyIbsZX/FmB4nKA2d6g3FqZT4E4N3qZUwXXeoZ3J3qQu/44iBzLru+r
sMYXmtMVP/JAs00s/iIWPL5bjPRt11gdAwNpr+uDNLxk8XYsCmGZ75cyTuZSgl9IMVOZcaYym2Bb
WOeuJ3H6oYQusCYs+G2RAqELNk0j82fdwSQ7u8qGiCyR3XYw1T8N3ZbBCg6oQF3EK1O7ASFwH7ZU
01Rh0EGpY8DrS6XPfFRbkW0Jo75xhP1HlpkBO0nLaOzkJkKYMPElREwPS1/pWjl0yPkTbeQzw2I5
fTnegdm46rYO7mtF6aCfN8j8XEOIaXQqDhUBHMpjZm4JUDSCitCJiSN3QN1d2NPDXjQKKw8VPGHd
UIL6b/PtQQI4hKLGjNJcDW5dlGHmWm9JE79chWNZ3hJGU4U90ZGwDkYIP2F0cMUzPJSehSF0bL9v
DyyaH/tQ0b3RyHKWcmI7AoELQai/ASjjUv6SJDNdtaV1vEBjyXxpsuaF517vWMx/JhiMiIYClvca
Ugk7ErPXWZftxtB4xqVBTbNA+cwqrCpEDSbOIAnua54BFIMkUdp5slkYXyhu37clZ7RnQxNM2UpC
xcfSWUlkfPH9PzeDL5DbyEqPG7Nbu30zo8YbA7ihNwzgEB4KdsBScCenYOlVeZHgS57tBbTXaLaa
ivzInd5gjzjtC3+ZL7vUEzGoJhktHZM4P3J7A9aGpWYHbZJEh9DWepp7YixFnjTMFh1VISJ68Gae
EG2WitSoiAF0k6L1wUMEaSiQn8Z2whEH7d18IVblxPb+wlBUHIkRBYLeU93nrJZK08uMgkoYn0t4
Lw5HwIEMEWPdbfw3q/lo/g5ljRbOM8heioxMw/gW+c+tNuW7I3TDeZ/9VUEFDKQyE4bVJZm0fZvE
3kh0g6BnZBn0U/jiw2JMDMoRxvdf25K/bMTocVfB4eyDGvR2gJxfsa92N3oW8+i+YTneNLdH70UJ
tNbfPvyWcWFaYKQYZhdQfyzT/p7H46qS1IdJin4QuTQY6+8kEf6jIFPTM6cvIKWrjDdYbToOVPr+
fo1NM/Qwc7rHdpgPnKmD+nJ3B1fn5FWLI/uERkvMw4t+PiaeerEs8yQ8Nj+gGsW70oU4G7MRraV/
DQjx66gYD91EZwLOIHZHZWp4QtB44bnoU9cxk/qawaf65HoFrYJuSVdtmcq7xZMBBCZB/HlhJ5yL
l7IRHAXOeCNI3vKMK1UhkRVmWPhCACOm2wGKKtQFpzNRl3l1wLhy7CfFD8naLskt2S4SUEtVWc3X
Q5ew3cS8gj5r5ufS9MsM5FJ+XdQJn/spFeRSRJcZzMbdCwnfsGOK3VwJP+9dxpOTilQki3TmKJV0
sMRE8orY36EeyhICF5K1iAhxwgYHSfJ0NJTh/jHxdne/Kcuuy2Q7D7t0cAT3YEuZcO7CJnGO+UeB
iNb9N+mlDbl3Cj4p7/VxCcDYG40PIXFRvtLtgtn6Rbvli3Tgq82tkLfGtLDIeYJL1PuE/AQNr0I0
Prmda0mX3/S+LsV/UQZX8pQ/giqImauZ389nY1HhZq0BDryEQKJfDEJcDEY86LZQD5Q3LnbXfzj8
b+q1IAS/VPEHrs4998Hcmx1ixpKWG6fnvO0FO/SheaHqG2CQPlMMTiEV3VB+xxTTo2LbQfeOHWf4
Yvh59rKHO7msfd8cHyuKA/OSe5ilyY2LE5m6kfk3JdGaDj2wmqekTHreJ/2lc4Hw7Aw0x8U810WE
jfJpm2BzZOvuWQxhYGq3lQGaimaYCdOW1dG45P9dv2koUVMvcaQ9mK6wGiZzNVn/g0oeAPeLCv55
tgVSwnOb23kWl0fUXnHLxi6KHKyvnlVt/8uOn4C1m2870JsqaZEvovEf+SomjLX9M0jzPSJ9k/9w
HZylhgvn8Xbvny7TlTtuyCqlOOZRTgA3XVrW6YT8fP5JKYv1uHwfnkm+cv0R8hV1k3XiOxq9Om8A
7XWk4bm4xTbPdmSNtDZS6fS+ZVR6XF6d5fMv0i9aluXLGMwnpPFroysoW6amkdLI/dWDr6aoLaiI
Iqru/+ElNleD2g4BXB9z1Dt/tBASd+TpMEdiRhluT4VUQ8UghV0YPkerWq4pppFi4OUwz9qS3ZKC
OXp/8ZkF9eJH0Dympi7DbSBGlAuDd+2KJMzYGKjmIloa3AnSP3ZS/bs83ooJUcVLohNiiae7s+G4
ks+iFptsYkoVQ6upFFW8j0vwgMu1pcUIKgSmy169Mem2iD6qj3VeN+aVEZy+AVfwWzTKVaUvy/A7
78ut53OWikfSKKla69ZSsqUbJeRI7wCoJd6kRMRxiKMHM1poVUSGjAg3F5JMj4HeqJYTh3tEP3RA
NcLwDVrH2vnL2iV+KgeVBEjd4lKLMr14CBn+hLS9a5d/MpjLOjlXAzYPS+tNukLBbw18phVETbkL
x9d4jUsbrvK1/Tvpo57viHUzj2oELvJVSvN+mOE4KNnGTgZzcmPIO5jxMFz7UxdRhq/VGvgdSxXk
zSD0fXyTQfXmKGtVQjL2jeiod3tyxNkJertYIkTiukP+Oc0RHVX7VqUuObSO4HCC54TyvVBYxb7H
+hTQPS9uLKo4/JJTCFbD4IxOT2xmhEMEqfzQW0CBSeqiE+BloGzkGoLsI/aqjgI5kUu1C6U/aZpC
D42+MxygaqEDo6x+8ODd9wKQyE008SoE6KqgBjZm/QjDvqodQI61Fa+8fzy/HMUnh6DkUcwa1llu
pGmr216K+QPvpcABvUPzY6Z7tSjfqVPPcUavUM3QMDjp64OKLSCTfl82jQlFl8817V6bk0MDB9cP
fgydHqeNFiJ/WyDPjvLz33KQ7nuaTRD2eJh6zzYyjTqzTKzT8x+iK7UJ8KRqf5RjNwq2t1Sj6Yiv
BVEa/eJ8o4roTQYY63zAR6KuuMW9KO7BxCyxrN2EcV0JwgD5DBzeq6GdgxWa7MiNFqG12X1Ahug5
a5x8qNpMH6yG1Ob6/RDNp+mF/VnXH1mqOyiz4A17Y6UvI8Qq+rYpTgc89Bb2T2/pVPOl2h9FUL4U
Wf5f4XFfT3tBRPevpC5AGSBquuDqwc0GSkjBLkcWRGtW/m/W+fxLE6bFHw4LznSE07m3q/FcMqsq
KW4n+z9VhQG9hFnZulfNU+p8Dc5o+FBYg0NFEs08WH0u0Qx/6FaMnlaDCaT9L7a9sr3GuaUrva39
Z9t/0T5Gwy51xceoFuD3BdoVUtyiC8KOZVno539A7ZMJBojIBF0E0Tg/H5lrNfghrEKRZxcEa/o4
1DWQ7pq2zxRbRL0dY8PuJ2Q8XF7M+57eg1wJSCoI4rigzT3vdRwZG4KbWj1GXhcvCXC5fN3wC7j9
PlS1H4BYlcU8GNssrzNuaLmk/K/gz20frzvjsg78HRXtzJJPUjxrs2xIOl3rwUkSPK/9Uqgi/8Gs
/4jDNxOvi/M0R5z4abzAftk47hJj1tUquXtC5FtnAzghosTYP6NFe9hWqMz8G0Qz+GsOQBTjodeP
B9EKv65NxditSLAEhn7/R4WCHl7kb8RLgDIRaai9v+wNgKzPHH124OlIvthAwYxQxdXKt8wj3O4t
BCy96FV8tQHx0zR4N7LE0r1VfibpR2KsKGk9rSbqAuNa5V1vzB8lWgce68VkhGe01fkaCn0owZgj
ihGHHYQoJ9LnIJzJvjvzsAKqdi8D+UMLO4ywQ8FhlXjHocp+xGP9FHb8g5ra1o91vh1I2cPnIpxH
rTGsJyCUqj/QfdqjND9gq77z2VfNQ/KHtm76IGBRahBT5menMV5gkb/k848A9H3QUyFAgk3YvG0L
qlcRUpFlgVbgF/KtmH6dOXFkojVdYZeIcAALhBIKHmPgRReTEqvLgOxxxkU+STTo+krPPBUcPeOi
Vh90MeJ5f3lubPR+ybyMWs7xwq3bXSsfHe8SvvotLEEnM6XdFjDF6nXJD6sHUPN/zc8jzzxo/yU4
Qd2+k/fEV18k3L+XKeS8AgcBHj3/xgbQRFuyCoOZ764b1+h545ImT1Pi5lqML3HCfRum7+ao1JLZ
8zmOQ27htMT2vl3pJY1W1mJ5sHjFgj77vCpUMlF5jOks8sha4N/gfyk0CZjPrVWhKe1pkX6tB3P0
xgCrQZS9hV+ckCAr/4+NRA9QIXMQdWeY6G7h85VDizut6LL9kBjf2CBYdOasm9OBOs9s1zgSGEkp
uIpKPqNhcvEJEdvpzjJpi4Ib+2vPNzwf6SbtjDuqB3OlLUrEoPlsiEdIFcTc1XGQ35AWYkvDeNtn
v+mcfx1K4eupVyWAHOugFfy3GAg6fFU9CcxK4c/p5IDVPuQ28yhHgmDO0VcgcSm9DHhJ1ZRMhAvs
SM3U2aVGQtOskzwX4pMt75lLq+ZZyYglx+Xh4Fmd0e4Xjk2XjnVYzFApkSlW0AOjpCf7tQNwvRQb
ZPsDlQ6nhBRGnb1n0HuvCcec7x5NP3cSQRNKcM7WPUxCMoQfM4zHK4ZDn5KEpCZJP2ZBqoAyJlUw
1UwyJewNnlm+RzaceCujrKu6hYIaQ3yZVJry+I3nJCW4XIPiCKX8KPhp9YjZRAiv3EXFz/X8YZb/
i0xGuFQwyvMH3IBLGrRTBAhsUfTrNLZH0WMrzAgtqyiXCTAwrb8Azvaqdm/ejJVJM5m9l/7PVna4
V8akFG+P33Qrnis2E1TyePE9Bq8jw8Dze6Z3DVRfOLCKB88nxHFs10RtWQGee5P0VsYR14P1aOPv
496L45GFhOy+Kgz6hQ6wf2YDzJOzyHGPrn7LAFiUf2BqjtgxDrD+alhRj++pYDeKKaQpRHarLgZf
CrXKOI64pJrEnVwbbhL5kB+Hlds+q42uWGcFdBpms6l6JnvV96qOy6nx7PCjE+pFDC5bk9wLcQu0
GDL9YI+2ahoeDlW3strJbl7kK1zTuDjlbtBIfwdxEBgJmzGY7lASvitqhVWCDNGjEReyeOc7PN7i
+9kiKfe7Z5s/2my7LCGqGRG2Mf2vTYLHZ1EBJifc6H9OERWbYd2lOgSxuoTOALOa0iYD7OHZhwtl
4Is6gMYKZXNLl8eQ+4GaYsywxu2PXzo29swL8bggn0HW2acsXA9oLz38Iiq9MGgYIkhK7xtJ5RJp
taZckSZgMMJ2SfMXn+R0os52az2VAl2PvA7r9g3I15zSr+KQZKFZYgsmJRhxCNiIh4sf+vgQESTW
ydK2vjyvRZqGOioJFN0KgfV5RVa4254Xmxi1hYr5QvqSQg0ZiEVK/fHmdGS5hGutJaIDP5E3P7nk
fqFTWmLjzYkpTUmRCSGSEwqVemDAqL7imtPnj+AOdEwXCHjvsX/rndO1/FdVZIUjckXaldkep2An
mabj2I7rNVaAnRQpxAFmycwQQkvGBI2ZR9EepJDwUk30aaMipJFymMSQChocZDDWoN9eXTCX4NmN
qSXBG3rJ1LNRzwvBjuZ+1xBvAMfpf/7/sqcc9crob+DrXzE8uCWmy403yUhHSkllsTrYqx3oPZu3
02LGLY5ap78/1KBI931Dhn52P1l1IPNwwv6pTrmYlI4hS0Qs9dGqiS5T5yjoweRh7PLZ6joZ2N5C
7/Lh4VX2/wShYyWeLkvCAS/ECWUhST0bj+eIDeq2lYZWmu9y6oEYvP6hR9J3R04eM/mu5o63bhoD
6KhiIVDEKolbgyXuW/ptaKxpd4+KgLMqe7rFKRdBW9WpnA/EduCK8lImQ1lbfpuR8rJABBNSnmeo
tFEOv8MPU9iCkeca4ey1Zz+3S6Hjrp0g5nm9Enrq0myYaFy+0Suza2b3LESfMgpxOlFUOXWQqFM0
FPSctjsWVkKn/vLNy34bYqB9Tx6U3QoxlXOyBr8ePXsT+s3mrlLXyiMih5P8aMNODVQARC0P2GRJ
A8DgBmZ1Yz/vcRr4BEmEtomVJD+RCO/lkgsqyVK+zJVFNn7XZMOwt9MNw10StHucXrfX55T0GS5T
H2aZSzMGRx5ucmVO/wOzKp8TgYrlArYmOkCO85FfUVTHapDU8qPsiO+eMFE7Jo1uZXAQabZr75q8
9WmCcE2D0IHSMUzu04rXCTH2t0/FCOW9qql+3d8TzA/o8Ye2OfMadcbP+gZLZjP59PwI0X0W9Gvj
JBI+AICVadlgZHbkmt6CpCrziAwGBwl1dBkKfgHX6WmixSA3WkUU/sM1WivSzVONyLpraZGwM2Pt
GiMk6pTMHbJF8XYAeKZO9TL4Ul0GQzqCmfHtmR0rhVVGUorv4flDKB74SH71AKbvNQrOPUmqfryT
dIaiyQcRnuseVOgfBE+ykfVSHoLY0a+1lcnk5FhbZdgs2FdvGCOK7D4GggLXAD8/5gtmMnZDu6nf
REL/G3jrqJmey2M5wxa895LWeISuLzTQU3WKVS1E0CgtEA5+bWehZBb5ZhWmz2N5yT2Qgc+RDB3D
UCiS8yNtGKs8V3kVUSnu1Orc7SeE3ZuOnA94e04J9BK9usSLRE8eI0NBF5H4plCT0QsAGetvzcUe
XV23Whz3giUgYDpomZ49cbR3eSqapIhU4g+QuDwE2IdkPzTBl5ihjNA4CzyaAdB1IrltbnSZb45/
2Aesulqgn9A0sjyHoUDy1Z4VsuqiHQZj3Gkd/zt0gHu5sfAZ9k3e9YcNMekf52eh2OjES7cwOY21
GELvZPmN9NLQ2mJ3z78OvTAUrN9t1anxusyY7YZdkF3Q1S6arUKjKy2NolSUIOb4MYjabxkhE/Ch
Qte7lI/Cv4t6eUUz/SQj/q3xiBfWLzclMQ6ej2/8YdvZVENDVzwvDylywt1+3BPRuZ4xZhg6l2hO
a6BiLyEN2EtIsCeDoBDcYLX5SPIE3sWWIyoH6dwOVuijKCzanBrKdu38AL6ESnrpJuhxJNkw67fc
A3towsmIlboVZTiLm2JgYoLhXXX4QFxYVyqdeU/kyHOk8T8gmQS1V3HssENm9ufZlEvHe5uDiv+R
l2XXYE6IzWl6iAtjnGBywst+yxDZtyppcFXomh/mxAL7QN8HgrGDI73df+RHsmahKyqfNJmfRm/W
5je1MSdtO9v16m8K1UK+KYNojKXnDOOjb0HN1OK8IMxSGrM9qjwTMIUqAMQBgmL1ErOpsnKtoAI8
gvx96yojBivjOB6RLV7V0ZIAX6wJEz5WT544Pdel6TqXEbcnMIAg5MbXnUpuZNjk6m50IN+BsZFT
KXGMhbs4X104Hkttp8J5lhrvKKqY9naQZqmw4OfENAywcZyYKNeRlck05KsTLHW6J77s0scVZ+iC
v9PEdfsnAGuTkiR3LIlvBvLiJeVWFOhdMrom99aOZte5HXK0iazyGIGqzU46YqqdrSbxGZVW7PGe
eqAg9V8PKghIkSfRQWZRNEc/K4HX7kMdq/aiqt2NwA+YgYmiqtuXXMhxienhJc3wdICLgHeSV471
5XY5OD6Z6GhxT5zAlzmqsusgCb1ouWzCUNGgPGRKWpD9IqyWiU6UrxebIQGrZ2cXoUyhPq34Lidm
r3Rw75pP/Epbr8Xeo7ehEQz51lbnEiDavhluT27otVLIcdgVabPxCl9u19+TrNONTmnzcqzoVa6j
N5G6kZ6mcQzfqajGKzKZeH2ZlJ4iE/Nn7tRgmClcSiCP8zEFlWvMSEIlRqloCVlGg3FGJHDiGXy+
4DU2b/IAtPGMTsPU7F7bXi4XxLxnN2ZfUO49WA2nfGVwHMf9VDWDydrZIrxewjRn/S//n6ugaMl1
Sf3x8yGgD3xe3HcpextKn822FJx2n3WB/M+RBzxwor5AMh8wwedQuYSnszqXQ2QbtKyM6nzcTZBB
bnloACUxg8BBEA80BHwWcAtgaAn20lY6gx1YB4XpSLC+o9s+6UuVTFb5TBlgd/kDIBHGGiPLMdcm
jQxVm4cbaEPBmp+Lm+TkCkl8zp3HH/jsJMh3xtPCgmSpnItYDVnhzKZ3Jcwigt4BjwSe6CK90ZtU
VMjIdVEvpA/LSwav4vYgBoLBN26PN3WPfi7B4kz4OZZVa8peTWaTJzRJNKcknGwgBf3RZVg4PM6P
ejdk2mK1XxszAo6t3+EpvYUfEl0pMsooEJp77wct2QSzhEC245iu8QJXxWb/L3l8VjjwhYYBP+RY
ISQk3qJAOxj3rlfAMBMhoOBJiVnCwFOg9C1Rx2ukarJ+A/kDJQlKXR7u1l92M06VaukyzwY4zi91
ZKhHIBhmpwYYNoEdZ7OjWLGg2jqUU0TE2dQcazFT/G7LXC+r9yVt/UkevOmTtUyoh2IjhHlkKwR8
CWnYzx0FTMPv5qIqkWpfPcfAjt2SYJf5jKthH/K40oI3wbjGpYHQHg3YG1lVmjKwIHKKsZBZAk5A
A/AiL/VRTgCSi9y5KkJP4pHOkUZaeYeFZUT90krTm9KxRdshCCLg21EKSGiEuGvYZr1GJoQE3K/f
M8Uv440qL9XIZAg60KFSDyTDusc48XVHIbxz1ya13bxU+gSgkb4vVjS23lPiCzY4e/5nq3JeY6kU
HF7gUVhyufjhGkxCvl79Zc9AeDqkQl03EsnZ6bLoKNIZpNJ93TStIFuYGZuQd541748HVpcS3WgP
kke3jd/3fjcZ6k2EksXnLYt2/GY1aGtsjAQzAtopMPPApjnpxbWuQPnLYP65Reo9ZxLX4cAziE/s
sxZwPCs5xq2aHvmN6vkbxBHSFkj7zTLJmiPFuW5k5els8AHAxlc/T8CBdfgMbkVzhTKWhbbgNKBA
mbwkKqnAhNUWFvIdYGeEmWNNq+5OW0lJcpxtlYrDqN/M9BPVNHYAmqxLDostVCDC372shSZjqg+r
Wwcayj73AfQy11rSNYKirohpsWUwZ3auUTJSUbhb7kLGkdjqkd1hoS2OlvZwv6YpobC5r/gQr81I
3B9HTp5ixHVxB2OQncokx1yxAXL7InuNJU219ljtWCBbmm2F4FtG1WXu+dqJeRgBOhJlNGSeu2MR
bcd6nilHgXihqZACHzm1+EnM4yW3zfbJtoii8t1dv7Va3/jaXOWmmFW5Dn/g4zCh7JL3YfK4EbRl
HxSHbl7Ubdg3tXZnyb8T7F3g8DeKAEYy92b5l4eNoWr6NWWwZbVaHDlYN5c5LrMYSGyeT9Slwbqb
r2UktMtFJjzcnvwyG4jqbUa2TG1Svy15vtDd5ViWhLBqP7dsiduBNJhNoeJUy9q/lfVcpy2lTUwh
4U49/wr9rQe+9qpHLRpoXwWtMlVgxFgdp43AKr3rSGYTuYHeHLfuRT16vuh5pLS7dRQcDIjDEe1q
W4b+vd9Mnan8maIslIuQ16k3T5UJom/+kDxMR0CyJnc9K2Ndolf7uskOas5UuPUAxgvMllheHEz7
BTGRdY4EZGVn0zombvkeNmYCvxo9YZ2u9eb7QV6lNsAWDYfASGR8oOwL9wUO/HpucV7lPjEIt2b5
F3L26oKr2HOzLhGKkw9bxXeqiCm/sCi6MXLjneixFMry3GrlatbovlURwkDTgRVXBXdMJ71vgGZb
v4x95Kj1v8DZu8YVJhK+0KhWvwfmd+ghI2J+r/L3FrMBcn9IQHKtw3+XVf7KVw09SixjdTXxurIe
MVP+WR7M7CuJwWud4HNcucyJkkadY8zvwmrso+FgIB2YJssskAYjP5DRLQVbGkPEKJEj4OgN1Znh
90/h2rui/otqBivzUdcLmUGiKCCSSIV7GR46HFlBkV21Fvgz11AZOMTMVZkRNwF8RJKVDNqDf9N4
LDLXQBarfbMdg3zspxPg9/Rcet5ePlAPSZUwsXMvL9F38S9078Vd/ngJvwuSztlsIXLWyHMXyp4t
xn7YXPp1IdPZDkD0t1eBmY4pW56F/0vyqkib3LfeTGyGivKO5VexDgkqK8zZYViIgmD7ynZdKBe4
4FlSZjL6s41PAtBa9irjt1NGGY+qwCaNHn6PN+ei9wRvk9s+eZNHp24pnCkGu5cwzwj4xBugC1y1
rpv41FpBRcd03jYo7m3SYU6ktJSOc79qdlab6VkvtFTNluUXX1U99JxJKofj9oGnqsJ0s4ufkCcm
BUkkP4B1d4uwAMwrRZPqyz45GWH7XmoPrYAOquQUtBboluYeN/W3MBmDm6FNcyM9Mp19gRv1GmWi
9HnEAdr/WKBR83bYKYcpLzbB96JscyIBFNjRHg6bV+OFH3tLDWbJFx88TOMM9alC9yDsJicMWnHx
Zl5IYoeWuZjN6FbuI+/EU9GBw24lXj2euSr3v9p7stv8CJaXx1Bx1Yc05ieHdLd/Kdhc1SNv9DUu
VlXuQfzJBELFuqFkU9UjCn66Alh97Tb6pP5iv6HJhRBX4913eq2z6dYXY/m6o/HS+2xlDlJczBdI
ILiLBhFYJM+W56vrhjEYhMQKAYDRppMucoASEFsAqFgCq/IqAEDO7Ewxisk1if9Ip/MqYVs0fF9A
BJtM2pQAsMt7dIf2n+y1fgulJXWWozwLEPOzoW/PO3y5xRH12Qnco0c3j3nha+W/OHW4qmUNHgRT
WGOA3vj7BZ8liVpSOa65V8sA/Z0RiWfW+hv6Z0Ehqli/FH3IB3g9PAG4TDLdzOgIGHnWJKu7cVu/
Na32yHO/jgOQnnXt77XPVbT5mybgs36V9emQSM7Jd56PoKfCV0HFtvNzo4Vjz0U9orDWQY7007cP
gfZ7peDLkp+wrTgIoRGIDzVD6BJfRdH7rcdUxfIDuYc9w3jqe1ab919NeIJ3YKpOvqVswwW2+oUk
QrblJxjbGFyOz1Cx4S0mDUsyoh7GtOcNHEzVKrqsJisLBSV3A4d0JNeX08g+RDig57Llm8F6iBKO
rTYMssJNSL17Bwxsh+XqfxxsHScgG3Z/JjorDD6a+pXa+IIFlVSwTDsNjeBepuGcVOKjcEcBUHLv
GeBJCi/lEuLBJU6u7zbm/yhlbgGBzNIr/lAYZ7fVuhritbqT84L5qHWdHqqWbAoSnyA5WwuQOUvR
SX8ggfUiAHWAzSPpntusaxxcVePObGXPhu9ck0cHQHzZsoX90/ScD6DVZrj9cTzhQ3wxnap1PsWy
fMbzJ21BSbk/drDReszIlerNLmmN0Vwo/xHVJllrlVkStcgLjj254ThcARmtrj7YlRshsLqTFuzW
n6dkHd6DTAFwcdopelufBASiqJsyoLHELql2LXbIuvfvhS+OAZDk8l5wB0px7xQQO5X+0OvbqTvH
tmIUhPIo4BuprrZJYwN9zJmQ/z0A1v829qc0b3TdBGx9laAGmNpUdaftlJhh129tBMAYn33K3vgD
wtj7ANBSjJqyst9aXZ0ZPFZPLZjfwYbwKZKsPVk8jkT7JtF0kXL1pkQcrZpZUlUIrcIiD9L3zRSm
y12uAN7BYkLH6jy2Ovm3s99GlVgaeH1baQ/NrOJZzWz7ICmMmglEhmmqqCRgBOEAMAjg41p8eBvL
lgQnCT3vXgI8meh+iwh/WJqUVm0Le8jOrhJ0Xm1NL3JvlwvzR7YT0EcF48QMk/5RwVXy5Y+skc7z
98VqMr+fSUfjX+vU7cOBZ048SdWkqsOWT1L0JZy6pq3ANNMd8pZMd/bijQnZhV3XCViqum97rQgj
Nadd/i5ogB+iPycXo5nUz6gcUuwcZnyhoZqYLi0x58O1I7mEHjtMkcAFcxUFMV7NTpjLM9+AbS1D
hdgVpMfRK/5tiZdst2j2LHCBKdcp49/N5Z1leMi/g40jyr55+siiOmEUVOd1Ca9X/tc6JGekJJcu
MBLOGh28+pLvTMtg5SP/i/SM+OwhiMZ0Dgi/9tXA0hR3nTE1Wh6+IZdsTOEvWOSqhfDlR383IKxU
XQAxCkEeO13JldJ8pGXSSb/3t4bBYPGuevm4S2y7YOf5ZpeWGUFIrxPyHKoQIu0aauIqqp268CMT
4EAr4hnC2mbLZAZDJOxEUc5wKkJIPdDnTFAmIMDB2tUMYgarraWH4gQYI4spRswRBOu4dQoHjiIF
f18ktF6HumKiZLfhOQAGhae9FpDXdSHZFMycuHx75SzC/DuzB9PkAGVR/feKJ2rmjAskALMaWHEu
Chjn0jXjmA+J6EF016z4gTaOmdNg+ZVimRnZLscY0/kc5ikP4uaPmiz9B2GtdMyP3PkPFxBnSUby
iJTuyAHtsgP1Z0n0veLJx3SQva6LmikdHxFMaJDzBLFoDxsyqVLVZwyuEcE0qSTKE7Di778fnt/2
m66B5UDi7R6w4d751f2VnNP/h6PI/CKJSoBt4bN8Bys1pnUHkQV3SJWfJNdTCmzMeItmoOaAMtK5
9eZHt5eHYEOB5qfic0T/CI94MYekp4JibTcOnDppXSPqoua3WFQWtV+Cq8dh5gftYDrSfH3LWWCN
x7gfyO3Q+dJtXH/5s9OT+BTed/EHvU6B/mP2j0pJaNNzlvDDS0nxJZfP+4Icw9fuao/2YdOMUevX
GMVShf8At9sjkyh+gLdeZ9yhN5veAl/iav12JSJHjUGB/JfNizqytZQIbHfJhlERVxYDHGEB0dxy
WsXm5PtPIDQIbNjALbH3DDbak0YarOkpOKoEFY07ZIMMN8wZ6mEyC2P1vafYFTrkEvFMjOAgmyKN
58ayIUZUNsDhMFog1FD+b2MFVDvsgevpbeplH9hp28jDAE2UcvwEBG4wY2gtx2QyqhiJqwfauMWg
xH/Eh0Rt4LI7VBFtiIlgVrAUs0mIHi92aZWgTAfbJIzyxrXgnNff3St5B1eH3SvYDIPQoaXgveW5
C+dJJqCFgD8XYuzohFQebNehBHdq/1AzxJVIIMrA7SbdMKUPCR24GSHR0wEHIoggThTRlOmimXd+
WrUrMH7tVbSeBE4WUIjCVYDgpxixfNPXD7R1akXbmHrFJa1+AXlchvskZCS80HHBw/2e/DXXJNbp
aRFbaYDU1U8JRszDBWQCQzzbNyH4tKcZwiuAb0JQKPJzkggPmKXEtwrE27f0DqzUXFkelBVPxUHy
UifJCTYcIiUjr4gIK+Vs+CvfpKJjR/cupcjclW/YamLWT5UUJ91smA4FlP5FtOVHQw/VVGHgaWmS
e6vvyvWDyQhPeAwCG/wKV91l6hG3whZNioCnde3HK741QcwTVIg77ycHSmNLyUi4zacY9vcWtvDJ
am/doaeJ99A2JPhnRbznx+XicZTWlM4zQvcwx0APKm4EsImfzPPhDIj9S0ipoga3qkCA6sf98yr/
sANsQbqBhv6/nMfT56RoVfIklNBwO9bKysShY2akC44/ObrIY98bKyv2bGWAaRaVX9F/jZwyzsVv
/jv+D3hOHAaEHfmQ5ed8nnkepkk9Ob+CdGsS8kqw/kaSWjscdIA/EDny+GxEsBhqEg+3gLR3rdQD
4iMJJFuSS/eVJCrPh0z+ZsEhLefspU3MuXOEOuw5R2YCoKa1MsjjEEw6dh+BSAWivSuTxF147tAb
69/KOOJEyRwAjtIiLWJikj1AxOlCTdxEloHQ/TBYmtDa0M1cBzgVYzlvL1W4DrR4K8gqeO4EKDdA
bK1sAqxSKjRV9N647i7OYB1JolOOfZwPfNYYEIBLXkqlcDZYbuZQmnSgBjZ1KO76BB1OD+BdRJOy
vfV4psPfw5zUd2NE+4Lqmwkdw3FK2Myw2MTN5jpxBtbcXg8B0DoINZex1JK3Trpd2B4BByE6ts5W
k871bMBUfGpaX2OxJF7W2s8wdL/VFAo2c+Pw9cNzi25SGnG43d8wEaxBrSkRkXcJomi+xnajkK1e
PrKOSOqg0woSFAqwsz5D8QyztMaRpwAWmFC63+4VO+irni/w1FjYRwWlQm1APzIyUUkwtpp+3kb1
qTuQiuuzWU5I2kImvdhZ0KTc6q7Qyr12WYr8DcuIhXrD8YMs5N4RIDdotfmNIszcBWtHz6anTnha
tCFjg8HnR6JHITSlaaq+YZ1kEWEYWv2E/wraRrAe09gI+D4JaaLgVhk+rA+h9AGyJePvS4ECl6J7
BHTquGv6Sk3O5ndIZDnmkPIqj8T8bD63vEg2LMoyozofCi/WvnVBw3UBAIscav8V0/+cyioJEAQO
Rx0rmBeH2WpBSSNMqJtSwv9Uu9lE7PdMlLTyW9GIThyn8YQubz8zD0z4gGNg+vEGGBISOIwoNwrA
D1EsYDbvBY64Pa5fm0LvM1X5RSJ2xaDYEhQuRWFo44WqmM7xTANvXavzg7aWp2379fVdu3dFg5aP
B0Hg7or1xOCC82VofdZIoyNKpq7Loa2NocpSbryjew/zjKYzw59EebcJN/plR09way80+FjF5AxP
g2gVjHIY2w13kEwqwVVZ26uQDEwy+76b2JRZ2mD8fGWT+43dxy19XSgF9ojttFtPxCLZ/nvT2aEU
k3U8w/NpBngDlTO60R5y5Mo/XsXew7JPmSc/IlnM6gWvhOeS+KqUOBC9m+EFIal1LQiowRh9ALwm
gZ+MwamkM3IrAwZfpXRrRF6rE1+hQz1TlHYPC18YcFrKeb8gLxU6udNxbYkWrmshjlvoZbWa8hs9
Jz6kWdhtzTANCzSZSvbAxpfHQSdN/301YTVZY3A1c5yaZe+JfSCcm3yf6Hgd1WsZ8Ogyb6gyyZ+r
2fTL1w49cdOVEOpPMj2jq90BPP0Y6CL+xt5BguKjH5EE88m/99sUrd5FoAgpclAYwU/Sb21+lObx
8OFH2ib4BCiN5vbqpKMvkFZYTtTU1L+M51JEA9Txw5dO9krNkGhsoPIb0Z5rLsf/aMLCBQGqfD4s
7PzcYFUyWdTGaGHA6YICJTVza1/BGsJEJWBK4XFQWlazU0UM7O4CxFp41sLQgt1Al8bDW793nj5W
rMJA7+vg061aO7uNnEEpVjUnvkR/PX5maJFLv5vAghp+vXmjnjVvZggtd+oBAHNT8DBU0/Xjczg9
y0AbeiFtjF9OaSZ2r4pcaQnphi3UMuUdConEZKoFDGhY64eKqZNeKnvZ6IEe3uH0r8ayJi7x7grj
Vy0mkHrttiob/T/lUbpmzaZSe3henxVlK/hSK5HKILqunPycBdF5BiK6IhZvQ7KDlMFteQNEusyI
dvyr1J1MTce9e67Z5SZ2YRBJ00a0xN7c0hUgBltqU5cgRiXCyz9heU4+xSpABmTYD6fmHibwASBd
LgpwItwAqUASxZ/5RjWHd58yZ4yO4iPNbpuSd/KSCnM9Z+eU/GTiU4RPqMDnCi34J7jTe8/cmE0h
x+e5JdUcqXBo+bzqJ/oGB658A4uO0Djk6xQceW2gWN5NiC8Dv7DsA9uMfDratFiEscm7bsiMf2rG
sRfIFUlpXGqaDlGOAgRVNY2YSJ1RS7NkrwWf1w3XQpWm7Ctv5FTcq+11zH8Jo0kzmb+Mh2ofCzot
unSsRdbpF2/7vIG+PZODpmHHjTvOC2nR/+L4LlpostZuGZP6t7eZfmMuUpfAywfXfTgWoIAnGDIj
WyBaKSXzJv00g481z6CSqEFCUooTp6QT+lZFalYFUbOMvA3mlLvJWx2LL1uUG64i5G2WOmk8Mvqp
pmD3ibyyoIMBngp2U5NdGvzWUjP0fz8E7wYwaglVPsIjlcFYSnDMWvm0SezGcaHZ4WhUfxz5IP82
p/vx8G/tWvn8ZOQqWg+z+2CJBnetx8fjb6Dnrx+GgvYA+ko69Wx5zhx9suUdLHgWWncjt+Kc2Cu+
yr8lcg/r9vtSOjUntiHmrETaqUUo19KaJdS9Ih2oi5KGUNc4hDxqDEPtX7/YM6zKcacQWsVJ4LFX
9XOoft/ELfd4fu+UDeK3UZXiEMHFDM8cpOI65VZ22FVloxqt0u04ld8dgKJI6hARWEvM6S1h2BFL
5LNLmqkVGXWJgypQE+mBtKjJO5vltej147JDnYWFnp/6sVcCOhj9zaeOzXhsFE1dyZFQaI+6MY6L
kFEShWt90wbz1DjGr9AVwiaSCTzkgMa9ObsZy3WGLVnHttbJMZeBePDCImuAlcY0B70Llkv25Ure
jPgWaRaSL6q3wS9NcQhw64erea1FibawOFFJBhbCFwnzfUsuggIqPk7ebcvDQax51TTshfWinHta
T6DDjdkjro9ITqDD4hZqayvARXeUqmV3KUwk34Q0bl2vRsBfdVDHO/V2GmoRyrQDg+7TLvga8Go3
a1EcqFOMKbjc7ePF959tlWKCEZYHOipPKdVjrlf98snXCths5NZD6/viteo1ZpwOZlG4QTUK7Cd1
q5GP/GGrh7bkj3/G3P9lFjAxrM2ti6MMoaPahFSeg1FVOzhMYYJ0iSDQ14Ked6XulRTQPBxwdian
ChOnuPn5cb/GFhE5+VV7UetgHLmbAwGNSDiEg8hD2DKnXOuB9PwrYJbyLZj6d5+YOohHEp5yAG7/
TbITK+6lRtCLWNP3+nQbbhmq9llJNUsHK6YF1HLP1nUB5ip6CUmFCJj3CUPqm2CclBSC9WbgoChO
uZtiAp1MHRIFv2DvAF+ao3qTcI4gY5y3yisjkfXiKkW7AveyVgbUFRZQOYRKot16E53oVsGb/pQj
HW2MvDlI827S/JzDQ6LDMO2aUh0wzIvZi8F7EhjhHMxIGu+dGTJk7d560I/iBrbjsPxLn+xCfKHR
hYWLFOArpT/YoSi3GcMieuMQ5ODf7X09bgE8vOhcm0wX/pBcf7xxANzsUvexl6ni6OnqBfixq+jn
DrKym5Z6KIIb2uTNarAsZd9NMkJ8n7pFIL8kehVejsMo+oHlUhlfWZuIlu6O+YvYiwuQCj/rsXGw
g+hnfUulSGwZcN5EDtxz1hAB8567TLYEd1sbgoTb45aTos9e6WHJmKQ1XIq4qJgppV4LLKf1B2qy
Ut9+S+HuHwgB5/K06aZ5QeB49KOuIS18mDq30Y/4bwsZgFlGCiTPsN4D+HeYrmTxRKT4C2UiJ6Lh
gYP46jI+AttHssBAtUH8VCaQh92nw6DiYgRfylYu7VNcl0z+FyXkTMJ3C7r0btOjsEBSLhR9mfTO
sBQlym/eo1GyGDex9ybZ+ZDhctF3YFYSyuW1cAjR1NzusdpdQlwTKZJIolxJKSCzpSBEcEeRqGul
g4B1xfgdJu80p2eJNaduPb2xHBaJ+5veEI0lvYmDTtKGASejO6TuSnyq/ELYLc/UPBvNCGn1qQuU
9/bVqTJqMqiEECTIaefcBK7PJI0ezXW+NUNSXIIpvK2vcEvtvfia+tbX74yHu3KtWQZneguw8u5e
MniG4PRM5KimaG7xP8viy4IBzFtemAHOBdo/+ayfz5a7iaTyLFEPo8+YEvtLZGkzxLuDvJE84+q/
B/4ZJtZ+/zmpBKgm0ehKp4+oKXAwk4o167E+Yg+qdemuytPrXB66V25ULuQhOaUfQpXa8/wlTPaz
SvSyT8sgQZnJZlSTR/GA0QEu8xwBt5ihrNNb7powCEJvJm+fBB/aBauluyAmG4Rr/yudf4YWqAGv
kLkbS49Ypr+OXyu6bE5nEGpDQfkt1Tz49C0W16qD/daTWyx9aeTzz2ojNq1ll8s5LuGtstDim2MZ
vriaqwEQtBiiJHUTbZt8oOwfRCaZL1+DSXDXVkgpR8HpiukMHC4qRcUCuMAVt0SooTL56ywx8eLE
rUZH2JbRnjtqvLNEpBEOwUchEpjhvHi6W9/xT4e+URxoUCB5+k5AYUAXhOl6z9CU0Y0Ry11wHlgK
7O3CyAQyj4HLedcxiPh3Fybxaj1lniWFv5/LeBSru9lepmFY7teCPLlhKR2tMlge+InDZ7vHF2kP
oqSzF7SoWKLVyV2Uc0FY20c5ZHQhCFh8xQv++Vw76DghIiYdcWIU36/6zKWk6QnjxOyiVWuOILjJ
WGmbChoP0BW0AxA8Y8Yh3htRGF8cpWi9O+YaRaE0H9M6VGziUg7kF/lgOQ/nCtuz77tecnPK6qwK
BVncOmdTwr3jDBRbx0rIpjsI9xrhf6DEW+Hn6py1kK4D7lIE5QySVGGBT6TgwLY9sjBG1zruDrM9
IcWZlRzAjaCBmajkU45orgF/xj/D6G9b2vMCnkkDKpV9r90JfqlQt4V9IgTDrW4paGeudTBNeg3C
DDecAI3a4PaVYHRG2XBFUgAzS/3O4Jvpth7FyKJaUVEnSFYW+hG5eVRM7c/2gLWsntuLgqB4uhdL
b5hafmox32IhKQSjVzIh0Cx3WqTqjsAK6a32q06UkRo4m/RKaNmevFBmJg/OsACYkI44hkUofT2A
rBzWv9p/CBVm++v8iuLs3+nZf+QJD/PXquYalAo7zWRsTlQDXLfY6G5DNHgaLJadfyHGDZkiB51d
e/J+1SayOWkbPiGE8JgwySXtCb1esL88RHlZhyma6hrKDc+gmdreTk7+gGbAFb3JKalZRWiJRLvb
0ds9TqSGLOW82GDCUi8NdBGoWP8MCbNx9Pdd34ba8Jf2AlpktgvNf1QndjTYxI8VjfZxLsGN0fnd
BVSOe/uQJY2qFQCSHonWD63ToOcLqHZ8fR0mxxnocpX2Vb8C+5cklut9FEjxr/LrdOVyXeRW+xZI
albC/DuQpkSUV/h/kaHW0ZsHiXYmE2wECIpDebO4gJYUIUeJhc1IvvTloboKpt63FV4wzqLj6g/o
vPgrQMDnUAZ+y4ygOzgzg4KBPOgZ26v8NjDynvX5d+n3Y6WsE67zv8pZSjPn+K37G/dwBzODqnBC
6XMUb22eXty+P70CpEa2Qn3JFGKTSyZT8N+GeYrfmDkl0YI5uCPsCotpwmGppq1c8rKpcPbVAs1W
my0qupDZ8aKXZ84nmHoO0KW610ih6DA48pQxN2Qr/Xx/MaPDr9IEgtcP07eg8FeQ/GAVOTvuvgWq
wehbsfoxTQxkSKMXB4gPmmaXSIrNVsd43/1PUp38bNusdcjgcFQJ2ZjkBDmoR4dBk1WxoOjwoiEa
SiEB1tzSTDow8SMejyaTPJ/JGRejsq/qHbSymtaizRBvfT7r2lp8Y1a2Vz1D6SUdu+h9Q/OpmUWj
87PBoVGvBP9QJ5Gshpdeeezk9hh6TDtpVhT0fWFRQ6G9e0Y391On3kwuSaig+H3751MxLzlTMcJc
VUqV1IQ//zf49fwV7HddG7O+EWF8fzBc5A3KvAjT1M6zMqW6SwHQiQw6oMhehRT97ctibLPyzqVX
7vQI8te0zuP3rQqi0cIUYoljMbfttqHvZ+5zhu2ELpzLW+JerOQMrRKAqr8r4/e29o7RqZYHKaHW
G8HRjKxDwRP+Pit60uepIPFf4cP4KR6mFUnMsDYkwpXHNDRr0F+PadUTrvzu1RKo17holWRxaji/
3i41DcaLIxdyD79P+Bi47eZdzIpnS5rLusy4yNpksQcOQHp6y0xFV5VTwwN0Mj2+tj+khjSKqIcS
+ZeIB4Fa1QChGyVjZ/QySJ1BC/yFU0XuC9pTBzY25gf5OE7qldk/+UR0kpf6nkfVXsx+MWfPUPAa
iPEJKfZOagv8jRebQZJkVaRTTIw2Y+oDwTkhVLmlH5H8PsRjJnl70Z8Zbup+9nyf4SPohbeZWyMG
7Dy8ExhHuUFWs4XMVcKJ6HhN9MS0idrRf2jF5Z6CUhEfNNJv2SSBNV18RXIn7/+lSPCkTQNzU5Kx
iiyOjv6JF5BwdRD7ZlwQBG9SHkkSDTa7+psuNAn7K+PC+jESh7+45stWvDNE2qg6qZmgi43tOlw9
PktKzznHrJWJNHixy76Hp9K5+WTzufIJzX6/iRq3Q3m4C1ZYMcEZuTFDXOmQlQO3EqB+L3EBF3cX
c/ZK5fJM/m1tHkTYYeNu9c8j4Rvgo1J1eP1YmjhYJ3Cr3ZpFhKeta0GKQ6m58TBBjOAQo4J7M90M
Aj50NTOYahnfnEXyW4Lfc2qy7tUeGXKihCgR4Z3l+XGuuyJTczAld5YBdNdV+86e3HwTInATE/oP
WDte1K4th7W57o10RNQn9WOHmr3C7QXS13ZG02o1UcDngUeJijvQEqZr7m991Mq6mMp7ofSFjQfy
K25JKrE9wladEtTeAVAw6otvDldzqqx40pPPwlmlRe7EloaFw9fQIVoKDNVnY//FTSzvQbmlxmtr
IhFoTT4VIk6LYUQxchTSUyternBaI4N/Y+xGNC/IdOPqagV1CTsGZP5eX8FQici1/Yi2SVX8rcEF
YfaroHFmpsMcdxC4o61KXajRUFgPt+17HgDyC0sNlPuq32pfeow1GSWu76t4PXClasr55A/QSvaA
gCKy0Ph08QoVKpKOOb9doF1lEUmk75ey8RS+TQxwDjypDXYAV3KhWW9tMUcT8QMdJPtz4mjJZbNM
gFH7aDjPwY0X+6MsZ+oLELaGawPYXW6KOnZh4OmPuLC20htjYNr4Sl2AOM7ZzUffjiaIv5b9kkGR
fHDCC8/sY2xJXNGQ2WcmboshcWigzzpSN6HmKijyHD4DKkVs48Ab87G8d++ajQnUtb8TYKLoBdyj
c08JcMUmq4uToc5qwjZb101tYP2jvRwTQwguP1Nmv/LHEZoCX66m2oj46LsGBCHyIkKM2mVv2x4J
TDviUSk5nb5C3j7rKTMvBSwXSq1CZvmZ872BhVaoVTcNrL7DM0iE7y5l1kjk3LDB3bCR5dcMZctj
awh82UYTb9SdR2Bf6zNB18RlKu51jK0wg2vmp4QAjaIwoLTvWmP26cmy4QIKfVtVw7/ohQS+dttT
SwpaZOhp+0FE1TtC3TIF5Fo+h60nzVGyYqtcy/1SeQdxe+raf6qHEkGyrEz58jS2DCxRHeQYWq7V
QifOKWtDT8d8AyWv6vjqxGnKxHnDeyRuHCs6/nVXiug87MHkVZzzPrDCq2aMjaGWfqnWVyde0Yxd
8UtJ50eABK4f7fAweCcgm4TBvgDTpHa1bQKLkTagQx6y4ULnn429ciZPP+WHzkX8C5YkS9PihyBz
5F5Zu1jWI41/wkrPJiIO9XlT1Wf3uTFdSFNz9WvU86xL1tU++GROsEF23hYnO3pThd9ArITnTb+q
6wkO9fKmSdNAfWxk66MdIzBNNJdSHXU/pPjzjNTStv4SMLFhkM8rt9S+jhTP4Vu+xpIqbEFMxCPj
kPJhybZOerLYT2IMxAUtzR9YbYTLLI99f+Etzx82VEhi1VRnJaQ8rYq/yEjRa6XzP+j6wLdSucoV
kY2gzkS+t5j6AXWx6zJqxiIDtEHQnmLLa77dSN4Th3Q8CC6xT+ObO3wAdu+CLkNKv1LPCIBfWeNx
jo4RouuBaBVjN04IVtlQga1pu4Zw3Vesb3p25jUh9E2TFqyZ//rSOwNYIHbd3BF+3UM8lgVPtd3W
LAdC6OtyvMoF9kYHZDcLpx99eJvsgq4sZtqJbSccqVsOyublZtMWs0+RDLgHoPxqumwzjqFx8f2x
RWPZBeHZZMcA1hyVsShnx9XBYSQ5EiavM16eTQM2w4OoqPEuYCbUCE9uaaa1lT388WW/LVuPhVw9
eIEN+vDyaU4bWcEP2D/dLDpHpvuq8GWkX1JFlaPb/Plb4WpZ40gfK06G/s8DY7emELS9ILN6qVKv
sy2x45uLA5iyhamCHK8TKHzUpXuMkre3f/vN3dVX/9mgAczWyEoYPo1dsPQCuvKEi1cHT3gN9toF
2+wshibxWrercDvVMXxSqiZwT0//t7VRSzZwlvLGNUXAanU2ES78igb89dKw8CTO+/Vm7xzePoS4
CFaWnY9R8RfmRgblVgoX2ZmxBVyJxir4Ya8YvPqszADeKx5mS1lzJL+5jyeMsgXU4YlHu/HH9U/X
UOX0huBWJ5bYjBGXDMaYtQMV0fDaK02InhvekuuC9A1TFMESy/NMcRFlfH2WOrIaN6nmUQU6vI7J
2v9W2NS/DJp2F5EX36oOf1s+D84c5ry4kdEqV6vkqv8LnL+GPVvSv0cnq/LmI1hkZ3nFLZ6KJ1TJ
ui9sYWnPP+SFuEE6fzg/kNZFIzSsBnIjctbX+P902T4Nmo7UOw5y3m6j6Pfo8gFDlSkx0aWt5uad
DaZ9fj9KlthCPCf/s3TxPjHdaA64ca2bR6VuV2cNzc7fSAS7vYyAyya5DwS1F6o7AiTkDHtPAe0e
OTNEqLbTy+zHqzciZWz8UCnKNvl+NPSMohqEV4wKO/D55vc8I80mDxXXQBJLu7oms/ZSn+AykAAm
onWVBqC1H+Hh8TuYHv1+RpakY7eEPwVd0nlJ1KfXtZc0qs+N4pTsIcHmkVPQJ9CweGG8Uh74X6L+
grfWxTLKEMJa0od7R+mTN3mxkK8rCleMioQebXKX1P9Jz0uO6yHntBQ6sduO0P/F3LeYfda2iJR9
nbSt5DtmGQBZufqgs+88qGcJuBRwCtOMfb0NGwbpCyUSsYzMU96mMi9OmhwIyCqQOPgdtzCB+lfn
3YozXtbNyX6v0EtqO1w09gtaveB0vZUWDm/OcmNhHoT+YybgsJeVOWbwp0xFNDKEEX7VpdiXJtKu
nYCm9h76HEVFNLyAUzMx4wne4ti73s2qz4L4uEb2oJRogCyQy9UzMRcKYleEMkDaQGGKxEteXKWk
TCJiw1NdzEiNxXm4pd5M1DeVeJE3ZGlv74ZPMXM7VHSDoZbZzVpSilPNb9UZZQQkV+7fj7BZIP/j
XUKw3RuSwHIXgyErv5kW2ntcSROr+22G2PmeHwm9pzZfouZ6lcQ7xoPkYz5DSawfnN4//vuDizyl
wMXTuX0SDJoOHxwDt8jR1nyXO4w/leFBtm7PcKq4xWce3CXJ3IwUuZIdpfbqlPLNLYTrOEbe7XeF
R2O3KU8B0tYfnjk7sDzynAL+Znl5jYzk0CW7cGuPueSR6K6PE6T4ZZ5uSEoHSbrqWYzMoNjjJt3X
IlMdABJLjLxvLZGVsqlKMId0ra0T4OxOFe0jjwE0QnRlXa1oTqV+GfPdRkw0ik58s0ChapqoNiPo
ay0gHf90H1PX+08iYxVNBIUb7iZYE+joV6AqdZ0++ALewKlKwW0fUJs/HC59ATbMlrOq95JhNmB/
aemUr7gG1pR6DUCa33y43sbtisf5T0OKGb2PsTVKxmPxkbN8LYhvoEItSkC3b2upBvHzksb1mAGB
+fZJEBgmDn5JqrOIVyT7uazJgYW9+nxGSxgOfCTgiDjI7I+HYFdkXdp6Lq76GkUPXH2DbdjNRCpA
wj9YlacRPoM60Y03wa/m7ReRfIOoPoigUoQbGz5TVXiMtA6/vmfw/agUaCX92T0vFjHju13k0myF
XKe6M83N6GGXyp8neMqsN2M+oWUM4/Tw4T8ny/L5d2l1bm28RNx3dFQHrcbYpcS5EEKDIdbfIE8o
MOXjI2nesL/PL12k6qtxY4dc6W0TXjOzeNSxMhAFTZLD23tT31xPRO2Bb6doGOszmd9BB9awYvWl
ZWV5+t+rYtJ52bciElpvsEzsQKSeW4/UQfoQypn2f5RGIe4ABii5Sb/rqefgPJf2x2iJXi2B6/Yd
REd62SRFAge7/1i7eIyKH5IzQpziVyCfuYPVU/0xP6i2UpHdOIvS7MQvQ7gpABpl/ULhLAojoKoW
wWxSMdxCDzW+e5vh4zp7YyGCD9MS24TLNVRUKm1IQ7K3F0PWoxpns0OVpDtSZ/uPRhCsC8ILxy7B
L/g6Yg3oD1U5Iv9p13lB2O+x7N68cAqDpukwSwAFbPhtG7x8v3arNKVyClqOpGezT9Zb3a9r37IS
Dgs2vbJMw5ce9qlcg1UU/3+QcZCvhUuK+oPBZcb2IMgEyYR9OJMuOC7gR71w8nsOouSqUZfgZbbJ
nVrZbz6UW3Z5BCdC2cmQNDGVKVMTKbkI19dCdSXcyguKuyc3Pjgu1KKKflUk4x2imONoSD8R73St
qTFp44U03mbHxoCsRmwbVACL5G1EBpZnZgo/QbmfqAMyPWIM+JxzUKk2YnD4qcnMCP+GhBLJ5y+s
eFR1qKJToPNH6W/3u18Y/QajRKhC+yqspAQS5d90/6gITxQ8Penw9FrzEiVpBLAcxmX9HlZfdwK3
kUIZqU1ljcwe/CKUdxswiwwXFEJ/ma/rbabSDCU9TNPD3HxlSEZAk1xQT2TDEJf09VsQohUyVPPY
4v+7t0fHEziUP2GmXbKNAoeqzWvex0GG3/Yjn9SkmOxIDwJMERPO8aX23iCoOxhgdxMN2oGOjJO5
HbsMX2AqmcakIst9x4IsRXjOo9mJ9VevC/t18H6hmMlYK57dHqbr7gI1SxV7S7YZBYmdp2q1cU2M
gCKYe+FxW3JvKCfsst/5cTfcpMBINJAAE9Jr99Gpci7azmh26WZGm3qkxTrJA1x9GsSomjWebpQs
EXA6mfgnWTuFMKgqCix6P6EVOrFUx5UPum3lyNIY8+7FGS2L/1Nqkt3sP+xPh1iKcBZEeOH8q5NK
hrOBzh6SbIS/7WSxdKDXRoE30bxFjm39wleQjx9hQKQ4lERmpJ1Ln7GXjjS0iQauu74wF7BlhW1s
UXHkG2QXoMEA/88Uc1xvIraYbdgiktLUCigBFt0yw0AQnK5CudOc6mlNctEFqxK4MtM84+Td7GTq
9Nt3r8kTliq4JCrGdark3fyNGWaGTLhxYGRMj19OrsqNc2YW81OtAc5qkNkEbwUL79+tjh1DArtU
wC4ltKQ5BlDDVaRfqo1M40j/B8CdF28yHdXnGYdNlrP5hoqDxXpCJLRP5OaUgwiAMOD95lIpuGMR
3s38RKiMFk0B1cq2pHW9SpcCMtqotpgPh4ZonZAxs7JPdjBJCrSvG9dW0p6j+XnCXcQYTVKE/cMZ
gvglsHj3juvmTu5y+G3hBbLr3nSttd0tTBOBQIWH02SRpIGodQtnln7qE3NqbkKlW1hxsq5Rc+fo
nh2ipGp1dpsNlpr/M8y7mxGvuc6Gkk3C3h49zAplGXmJOEcokoIbpyBDOVHk7DUNTIsNU71bscoF
xwmzGIb7xp6JQ1wUIO5BouTZYe73E4vVLfs+9Eowww9lbxQSFkZoep/1BPfk6e6OHDwSPULqtnl2
jUXH6styyunbAWNPeDR37a6GG9ETAJt8R2mvT3YDVUgu/qeMnVT8qP+I3qJpFu+NHHrr/e6bTpSp
uLwo1C+zELFXQXTnbp3oeVK70A7xFrQ+GB5X5ufPyA56zRr7tesq7SjC+l+vIBdln1i6PIfwI36c
OqaCe41Es5mZC+5L90y406ylX/6DX+vV63my1dcG4aGJymscy2rYiSl3GfQ4wFZ/MmosWjjqKg7G
AWSziCa3JfvYZ6cl0lONznORb1VsX4HZGDLmAoDSi5btCC3HLruuUqoslsafacvvPGs5H84iFHjI
8sJpz1ZCSkdqxgDUQxDj1363UwmcMszFVugr//FEHvaDrsop2iGwKnsTMggpuNG/M6aO9OXkIsJ1
pxXWCEky22zRThZkGaOfdj/1Wnfn5fVufc1k0R2jRsZfAsZwQXLxH/uZJqOJM1gVy5yFvLZp/0s+
FD8sN5iJ6a3mosrkWtLMVK/t45DlkXylZldWDxvPtOjw2UER+NdTlf3IxIikg+Q3AVqeGQMrVnOg
xDytQwIjXzHb7lQvFw2ZOa28Gf3jRvrqS3pP4/X1SboWM2XVKr1lcHME/0lJuNbNQKiAJ6wC9teD
JwTvJuBbhyV0tlzTw1Tai+o37uMU0cBAMUbP1nbcYKSoDFAC9p0oC8Om/V4XVMmz2h31jh+1LDAE
VgHsOzgYfNTjO3VNKQsivrrDYzS5TCHuI6YvwxqGtJpRGEg/uKeUvHboteMMXzFEIeX/L+CNOeNY
eLdw8s+/exCOIua7/v8NWrEK1/ROkasSV6h3N5K0pxYkJeSXDnsPx5yWmgo6jDw3TUruGnCArYgX
wfqEmEiIevIyfc6S7TGIqj9SqEjJJIN3jqOfX/oXUPjIsol98VbT3UOwfn6bBBPbSTZMoGGoy4Cs
67snP145DS8eTmZ948TD6VH/rPj7YOk6++ZpgCBr52iC7aNUzK14L/CFdHUyLJXYgZQ8ehb6XGSC
evZonlvGFsr3WGNTHuas4knR9p/ROtz/KHu8ERfb4I41vi+6By1nI2C5cvBVKZh94ZFriyRC+Zar
+EMx0vspmHk7ZslGGKDi/dej1wugJFJtQDtJRbFx6Kezxo1QktxEkFZckXaMdhwhB054hPzFVJ03
qRAf/8coGwiuzZHYJrdY/J5nYIWx/z1O+3MWfTqP8EjAf8zfSPlG9O3ajUT53DcfgQ8P9ingwzFP
b+K82hI9v1IksqroZ1D3doOnXqeA10pAdPhCkxutUQqfP7JY8VFIx54lfUry0dWNBKvLCOyU0RGi
uhQgBMqp+uqFZ9+d33cUME2b4RD9QJ2hLCrYnhkS8QeswtX6QmRrTMsE9+LQjFoSWYzcoEbgtfTL
1OKj2urFMXop2YlJp4aFtnDF52E40nRTBXjoSY2uXR27dH+OvDMTC0DMegf5bZfMPJ6NmxJXoW+t
pFhoZG1v1vcVS3fdVnKcTHr/GDjUIKNs8Nn155ZyMhP62SoCif43JuHIeQ2NIe4PPksIuI2JFD5N
kMOKoBLy/vChHGEcMrcUg5fGgN5qlOXeDE1bMVH6AlaAHiwHGHHmUWredBrZvRxgCL0cFWph7AXi
YgWRNSEjucCdi+QlptoBY10DbYb6h+DYWgh32NmQh2NDai0wMlGirPJla6DNrK7UgxWYW4FM690x
bjT4L0xRqZbKzKXGcZqMrPAoW30UMIobV9lH7Dx5E3SjPg6AFBE4O1AgPRylQdB7n2bg4QUijNN9
NT89CMCRfHU3JS5twPVQ1NrkCBj/qj2BsaN5+FDtVHUVX5ao3MvdPbnJM8YRTR28q2VD33kH08Dx
lmsBeXBqEgRn5mnvGb6fURkUSI7tz1ASnWCEbRh/pKz4CaHe877oABo5CS+aFaB96/O3ov4bEFJy
cHPsOKBASLwKyXKENdSQ1D16dUyVhFeAhwhprojHpziilEtXmlv4JmjM6PLvErt7sEGNB60TMX4I
9gHWA1NRck0dkOzc4gns7vy1RQEAH+GOhyu586CHwgH0A+W/OiFidrBv58NgzcIzoXvHmEhGVwQ3
/FC1UluGEOUyxg5S0/Vn7fidBHToUtowwE9d/NWDPWL+I2hYmNRNujIHCVMw0GwuqDwQz+7ZkcHV
qrPtoaKpZFK/b6OvNTA2YXah/BrVxRATslIrD8Kz57GTyfqDsgMuwrXA5ZRc5bzAx1a290jCugeB
2eWhlqilnpZHwXKlPPYNMzE+YYCU0qd12oCl0qqrUXXFWhyUyNvdMlWwhDGtnv5eh6xzbjmKtSPd
1L3g6FlGrQRWQv5oSzGvEeY2ZiUbP3JqVYKO+B2ZLdvfD+fqAMIqSVBa5l2KwzTNzBKtL/gUoZVp
LkUM8xUTkxQxn/O4k9eQehz5bx5S0DtqIZTskP8LR1R/z7Jyx3zn2tlrwx1dlKh+NJcwZ+NzKExG
2Gl65mMRurSy4fTVcdEG9wzTaKJeOoSOyhrdGCbTErvXfk5J6bxekdD0ASBqErgfnRvOS93Ytf0J
eHNAlFXFPKxs/nRTa+HoZQiS3w77qB6poDZf5TaHIrUaJ2erJBbTXaRPEW/0DYP9hvnV57f7WNIN
nVOBP/1RH11XCICTlvDt7CIZ7TvV86Qj80giepP991uQEPdb3xGUOOQcm0uFObVC3K4byB7/fm1w
TPd2BT+Qguh1ea+0376krgDYKQcppS974cZBohMBBD/XuyF4fGVE84QMUsezFR38OQjs31pjlhSA
68jx1kSgT3ut9ThF0TotKyH8sUdoOCx7K3XbLNGz1lPVsH3mysfao7+fDYJUnKk7K/LgFlY3OTe4
W4U/zWyg+pnMBbcyMjb8UMoAmRzxc5NV1QB8/SD/+uwcuuk0Ro0DEsdefeo5jnbC0p+6ZG45mWKp
+EraOC1KwDq6vPDPnZJPgBn6iD3JoCtM8ES70gIyrSqp+FYrzwOAKJ5C4pNp9//CSb0P3L6tETvO
j+ezFnHaKoT0JblH4sCSkmeD+3ZuSQygoMC0/Mul7OifhvPw7L49LWu8aGDn/zM+YMSR6Cap0Q3Q
Rhs303D2kpo5FI1vl8rp7Wmb2N1utntnj3vvT6/pN/MBS0HrsTONBosTyS27gcOOGfNPVjSneuVE
6P4iNGipNDoaGCLs6Deyln31GyWczsgQuywxT0AvplsQVvaMsbMV8GZ8830CIivS2+rdVrJqR8fm
isrZ7Bf8CPc+ufpojJTQ2U56UlvzbV7N8KrEn5CbCQj07Rl2K/qC/zxXBfBduibKrsAz7zDyiXcr
sGwaiM1RZ5P462lrnXTmkuvYlgqxSBu6u9F9ZiTQ4ml7nut9aiexS6FpyZdXAxGz6rM47l6jNQze
FSwfL/vnXinuZyzY9bOX7oAam+hFvPmDgLCVlgOxmnYURljluvqZV5zer93xRjyihxfuFePThrho
gYDaQTt1tos3BjKSYC76i9Y7H7bOgVyvz/wV/YBWsxls+krMQP36Psqb0AgTMqTzhKVLz1SnatwR
fONnQaV12XIRo10z7BCtqseOj0Tfa/JlYs1r5hPX5WTZNKbIHdIeVWKVVS+H9NbINj3+5G1Dr8cl
iljjMZ0acVmIQbUvxaFpMMhgnccq2Pu4+Ds0jefzpiLIkdyKW1O2xHaaieniLXnHAinUF8LOsuax
RKuMPtc+D32jvM5atw/vyjqggHbMRJ6S0udzT0ARtkY6OzIuNYb0ueb8PuKw3epjdj4CDskEpd75
mq1DZxo9Up9imelcRqUPzNYL1z8VgneST6eRiCJAeYWf4kA0KmUoG6OpnJJLiZuiSAatUaT9xQVm
6SL1b4MYv2/2RdEdzGJn3/8siLyohPDaqAEDVBdSqVhs31BO+viMKwBr/IC2fJV5uKDH68X6d8Cx
62TWIT3JmUr4u4Z10I550TgJlI3xQReDISQ9uGIbFpOARgW66fDEZGGr6qEg3t5DSnKojKhC8ugN
QvIgO+O7OgrXsjwrYobzRUMAoU+BLd8lzzaehg6zLOi8GjoApygLHsxaipK7WJ6+4WxrkU/Wwyht
OEVFFx+sUDOhPBIkxe/K5ung0d3z15d7C8cGVdukdILXJtWrdl53fH5zdsnncGRGO2ZpPEYEVdOq
XaTAH6F1OKmd4zzc6RwlZlFiYEBVkUzv651QkyHRiAfMcPS8Mg+aeJOBlfYJLB2Vi7Rk4qunLMt+
3s3zqaWufSAh4qTwN95dJ9E+S67DRGqPNXX35XulopR1NqIUAi0Vv0NZFgw5vw/83RQQZYydJ/E2
rJO51LwrxUWq87euQmLs3G52NVSjMK5NsgcaI3H/QzN7AA3ERvCnszsCpOOcRf2QI1OaOMtYzuSF
xWlAHBA3RWQz+EhJDYrWQQ2YZnVeObfczIqTC4KWja09YAe3a7xkwDQsyLM2JyZOfu98Ir5R68W1
PnTN75HiU2ALa7ox3luzzYk5Bt/xfQpApC2Eg+FuhDy904s2J128KaSISOCR6R3C5UJMN7QEea6P
DBZQpA12SUcUBOuHzhufs5DGdvXWlMuIkCU3A8FPAuDKWHyKme4ebEnYyLyJoEZ1rkAHCY+IrqMW
RVlQp/XSOiUZIWE8LtfZMJHY3XLTQubieNer3EdV1xwbNxfWzOilex/dXADSzXCDt5D+VnQzC6T4
9NePxSpZdQzmJcWE42mu4yj8fqxI8/8d3iE63qvhLExsZ3roxs+8XbGoYRmjHJgODVsRrGc8RDLf
hHQxLMSnhZLJd+95pTGhzclVRmH+8vsjWcw6w2WOqERDmHukmYRpP6epE1uRd6LHCNCqaNO3zDP3
9d+B7k6dElvEwmb0FE0/3W4B7TTs3owNI1b3+euzUefNWxY4QWaScU2L0rzim0At6a0ukxemi7vj
D5L+7EOQS+RjcrNPJS5s4FyAHUXyGWJi7uOtKAe7h8gTJopwvKCAv/tKLFO3M2eMT1ASZrchIKUN
0/P28ndCB0iR1n26vUgTGC78CWQb02RoocAdNgBvctGwfZO4lcC8EpKuFASwQfBJP5vh96YqVVGK
43sYaHYJGJXnzHe0CAepbETbKGNlAmVai9jI045oa1XlE6f5wh7s7bkMdgPUGOm+WDZroNMZbTsB
zzMf4OjN8RD+NfCmA8zTNZX8C7w9DdQyKpmAp/kArPNNHQshZH9XV5Db6OXynbIQQQmbPOPFf2ss
rcF2fxajnqrB2f5GFgh9PjQp4rZS30BJymQPiGzEMMnv3fvmbfBHyQcdrMsfAxm1NrXRoV0bHr4V
oJXJ1Li/uBQvs9sMo+eAgBHIjRCS0DUfyPcD7fACKyUfyJU3TzQtlEgBI+dsxJ/vKqPjKYmsHF5E
FCe+fT2A8RdfbpLpoe7Xom2OBNTb4+qPeo2FI/BJNpiSjhLE6k29lL4Nexkcj5WjvsSsRVnIN1EF
dqx9zAlo7ttJrmqeHi2P5gIa9Q89Dh38xkwiztyg5eQffN8RbiaonY0+Nh0faoBeSv0AGbsmo71y
KaIdrBmsxiJDQ5s8/w1cs9dTW8f0ad/CTQuQcPBhq5xN1bm6npKyycIpb8VdpTeTtbFpEnGJv763
3ZLRaXFm5F6T1RFrndtVFUzF0jIBWMWbUPEeXIfD7ONPncxV2rLYdvOUHXW4/D59YbKbDD1MzEGc
jzNhI6aN0R4Yt/xuPjl3UTVmx+uUFVJ15IIcWEdEt7fyTz4IIUxLycSP6txZ8bm9hNbt+ejbyvPX
9xS4yMd2saiHau0LSmJAiBskbm0j4NHKTzHj2mX4eyMpdf6KnvQWt5t595/bKeVhzfv6ez8mnEyS
S9OTq+AsqBUNRr198xjK6ZVnkIgRomnX4gInv8JcZ9T9BLrtIwmXBTBsEK9L2AolNcuBbnF3LTpU
xkFSI+REtfNixL7llNAeRgYAU03PU5YLYraF2oUgb2XaEizQ5t7KHgIka0d5xczaQF3mRB62KLj4
NKWIgB8QppA1bEjA+/3ZD4ve9WT8P/d0Ll6A/lHK6bDXtUZxiraQsScbsgBJz9zZ3OZzOSaHJ/Dk
DIJVakbAGb5u853rirhQtyqp97NZvdagA8jz+mnPLmEZn6vaXHs8llkRUdouCSw1fsC80IdFxUHX
c6k10juDC/bwZlgCW6zqqpzj0NtaKRBeNSTtE0W5hW+yH3msLuQUd4N+Nz8Io55nwXeECOJd5EyC
UgrKAtyfiyzuNkKRenzT3NVykWW1CZfXlsKsyN7pAPkDtJY75jWDvcfAEb9OVLaDXE4sxIY0tGjj
wj6q7HF5aXQhFgD5uoZ4X6oW88hUN5IkFfA3Hi/mti9A3kEhD2dZ8kv/7zhGku8VRULYV8/eNsMa
a8ytcP4hFxhLbzXEpmOC0JhpfvbXXa2G+KC5BB1mnjFnG4e+ppm6QfOknxDBHpXAURC3IlULoOJ2
FqPXGbfqN1MSQkNZQj7X1l0M6TbzVRumJjKiudCiklkWL6+DRzEeciUXiR9Xgym7g1POre0Q6c+A
fExzOIdwreQrkY3UR+Mtps0gYr8KrMAWZc20NFEs5/4XW1GYjpAgkQ8N2skoiov5gQ0cD4dIoITK
px0tVkScAzu9fIb+E22iWQz83+0mqMTTHJOHO1Vw2PENET2RsFxvtX/jB4jR9dCyLvRI5UTmHq1P
tbDuEe16Fcz3QL7h5wvXWXVpfcEqFGIBAH6z365ggqUqMlEaaSfcBQri0euHPZ48bv08Bw2a9FwL
6rduglgqQtJqmceOxKaXbfZpSiG9Sxh2kEWTGcNGJ/QhYWi3uq6sTgH779M6gN9TaRPcLQknniAs
cyTElLVhhEekbX7GHqIs+C2kKlnojLvlQ04fP/HpYtdjMo2EltjMUvgaB7OrahGGqg3HlOGEC526
/TIpO7Qh6trvo1+ElXw5cCnurdtWz8xyYfiH0mb8bt5A659pPuvUAkQFnKE3s0RlX6CcgeDT/dE5
oCosrr1Ir/YE5AIlc0yb7lk+9ym+9ASVBoB6MSU+DDyJ62WYNafoA6mJ17NJbfPu6pA3lAmuv1CD
FnwKdYEmO7r2Sa2bD4N+1+GbBBmO82KzE3iR7NDf7IDdyA7T3i4u+tYVR6e0ftuZhIpngC15sRQf
PjJj5TBqKQ7tYTAdMc/AoBTcP7GKlHhnTcC5kOP9LPK5PxPQrhHEgZ7mvyJF7bLeVD2rzj7eh6r3
NreUSIIPeiVba1ZIIQ+pBvhZnZKYGcUM4LryBQ5uoEw1KdLO8CHXepCE7DGQf/X71x4HtgoNSboT
SW8DNqD483SYBiwT/y+WVYBgtNJsgFkyPnk0n0/OY3Qal4fmLEh1z1LAhGvV/6qlognT+hi/pe48
TKemUuHf0QegyiGW8EskZBWtMPFY4r9p1epNEywrDNN3TpJTxzO67FBQp7ectSP+iGY/xicT4Un9
LYjpcBoIJkhoHVqqjHyTWd39qnb7xPdJrPNLNcsZudCNjYq353fI6QvXqUow4MmRTiHTb1WVnYyO
QHlm4jrKrKiT4eXPaxoi68z7sPBaeZlf5lwKixL6kp0U/sKlz1DiI8rMNV3keh+rGEwEk58JlTLN
mdGkZln0LT2ygydhnp+Cf2ASk3MtOSnwry8zGdAgMoSmmYLgiEPdf4ZBHhDdQMZyUcQOKhC1ICUU
Wjz0hzfMjsj7TTel5dn8Abg6cPlQYkfyLN7QscTjFzxVxdgwbyx/mJjZotuc19whJMKvm6FFB5Pj
JdRvlxEvC99KPAzdHZLt970Q880Q4kTZb9an+QAeGKBXDqg3+LV8bQfX0uE+MBu+S9h/DrlANeph
ZSCs0WR9Ax6/S4diDwWq9oqXQuJNs3iYMWxJzaG6ttWAYyC2BE4+u6ejZMJhtPkSp9Kn0D1cBKC9
eVOmkmqQ4ClyPIBdYGil2bA1W3+m2ziPylka3Z7P3klZ8+4sXyifiimT6hMv6CQT1yeCzdtyDkUX
CSg5fo8ntO1V3ipmCcRTqnhB0jMJJ3P68Egc8MSaMfIvbYiJ3+roGrNPnrnui2+Jxtyozu+gxfrL
8/9+IR6ipzsKHqc4XdWP+HlMafNVNoUg/8i5DNttpZQzdgkOp5ZetHfQuJHlRueSqae0dtmXBm2c
1PJlgQ7yT0r9hNO8kNUHy7LHD7LdR20WISGOONKCUntRjniP5og4HBGi8au4V2o9NzZsvCS2qh/d
5nWLjocVQslaywU9MxhEjs1s/9wNOtcLd1GhQkR92GfgKVXm6R7air6LPmD3gtZFsyjiOQcXnJIw
a6SxJB/rsfbHLQxOjvGAl0ZiS0OXPXCGtXycvt7vJsdpMQHS8B8p+nb/Keauo9tIX6wKZBtt+BvY
b/hgYme/npZk1B4jBNMda4pR1kWq0gs5KMP2uDPyJVGjPjDFVC5qTXTxQjVkYqvTmPAZOqbVUtut
fkk63Q8XKSnst89Ia6YiqWhgitpUZq0AK5uCRY/xYtoee9qh+jSpClpYNKUxI+dtcb/rjW/EbPxP
7vAj4hszeO5vd4WH58kqJgpiZCZzmpV3v0igtjWTuK4rh5cyC8prdtExmDKkRSKVt3ape3SgkMPY
fWGGFi41/Xs/2bC+UW9b7f6VfhVaZOoNWR6df/BDIg5JGSBu3Fvbcpsj5OJVIvRWCpyha1+9bOBY
UzUjaHLSGm0PTQevrBrDBajpRVpIMA708PGqw7ZBOZwKWbMYlaRTFSuAuYkCTXEm39a91pAnff5e
A5CWikeiaKJ8Tbe1T8IGtF+omubqNG/RkNlSkw9sJljqHIq5UAgbc0UU3sPoTneL/uwk2cKFzfP7
5FFLjn04MoGNsQRBs1bsuq9NcjZ2CglFxuR/h75pPDS4Tfc7+GAcamnadbeVKSJzcSYyksq/hYj8
WwEzBMTzOH/m/q0LmcieToSFyZqGzKUS1o8BCMliUpNAeaLFTE1RBQV5mu8w5iTDqKI2Dbwub+Uc
F8FagWMyQKG7sWsnUQaLNpbwU6XkBFHfGpnNPQ5SX4bAp523IqD9MXhPgHPI8UXe8o3EAqWx3g2w
ODp4EtH1y+z3JOZ4YOSompEEK/n3VYZTjbG4TrBnQv/IlDKq2f2YXA6ocoyiCwEvF4eGZ1iYGbmV
EuJi4/lQuU+/7xDAfXkLKKSn+9uhz4R7B1zBqnjlpfxmL9l8z9HXJ4k3upXLy20CbZ2yZ3FOGh4l
tLnExxNCkfP1+PVMQv34nsxC2PQewlGpIgH0wliQBPp/8BrAtu/CZOXCX1+WSvYZEpZ9cdO6Pv0y
SSiKrhjTGbPH4Iyb4C4TpUKEMpqc8fG+iEOqcgSoF0SLQtbJLk/9sApzSg9yfKcfD7ykViI4bXfm
YN+UysoJ/3Qve2mecfJQvaAF/5C1auNAu1lq5uGIgxiuOKZ5J/MMFabppTFn0eLxS85nLeMjMV2u
Dqii6UV6SDcDRJDJPy9Lyu7NeWRPDhvikqmDcYV29DRGHXnPGCbkiP+JK25TK8sYt6VxlO65Yx6P
Wv3VKyIVJmicsTgFbkef/dexrZ8n4tdcTiFHccfZ7hjJsVvssoijj/L4Eq6P397MKqWQYnfDZ+Ge
v6O7b813wZKHX4m63Fyc6jDBx82ZA70Wvq2rO5srS1S4CN/ImImMTIy+xsWH1IH3PwTia4OvOOqh
2JzkIryiMKukDJvlCLPhbKcAmq1RkYLBh5MknsBnNXeqFzL7FCTlubZ+E/BF6JjZMBAJ/kqVZkLD
TsG5FqsXx22MDAVvk++V2Fw5mb5rrWVeN+MlPp6Z0a6HIwrrP+NMnvBNdavdNKuqvxYnZEzkPcYR
RXEwbx3CD1UF0KyxAItZLSCTjbr7CUfC71m+jAWdB4fGHikaivQAEQkNPVYX3/cFILCV54HDkkFY
X/wqIGv2+yYPh95icm84SyI0NkD9xYTcr+tDYJM/6X9VcY7aJusj192KPaiotaQkUx+Mpiu56e+F
+rZUge16kZBJ4w1jFE8GLm3HwCC1AUe5/46hZEAmuHdZbJTtjxOFLiuUgJyKpeLnBttgeW9Pi1+F
z8HD3EmJWvOoLWtcwNY4lNV0Hc4cpcFeIspL2xfDnJMTBCKvyzJDk6anCZ7twtOjTOlq2XYRBiPa
qrFrbJVYk5OnEpxkPARaeZwIFwWD1KL92dn0gyvB10d9UuONsHfw7oHNVB/0csBrKoU22BAn92h1
hcoCQ1fZjG7ltwZv8kUdeEQh0BruuwW0AcamCrWzdWTDZOhVYOWCBOoT86N8XvwO2h/4tvUmskch
llDtsZzWQd5xVarHCzmNniin17jtfprUoCfgUJ8crwqNtsC3CCorsfG8OsO5JrXGpq5tmFyo0wS8
ju1IwtB2MOeLs6PKbFT8phhmUWrKOzi7BRbvcTK+jMLmV9jIY+rSt9ySbpMLLjBi4NE15EbhqDFz
zFuJN6FoLqCiAVp61pFb8TINcYvpeWmJymRulSEjTuvn+0WMAGjZzkMVVrUuUhWDEq/Qm31m5QXc
at53XWPUoOJzHMlFLaJ2gigODy7ab1NealUa5jsn2VlUW+rTYK6AGQEPyYCJAAMFt0zrL3sOG4Bj
gJPOY6+nvje+EUEdYYad/Fw4t1iG+mLQWd/tWis1zUGLiXwcbqUc/DHzs0x71sDhu6XAwog2C6xX
0PGiFFWmahkWHQE23hc1ahMXfsi82uss2TvQU4i3I+Kjl1prq2VuuHqV+FYXpG9RpayiIkYUooWG
0MLVQVCEeTeydZ7NEEsAh2iiGGZ0DkUZ8u/rk8j4iNTQ886fys43oL51XCDuiakANeTDNNGiIu7X
q4vdQ3Z865ACbs/y6Ns6yN43B1RD1mU2jYnJQ95XSvPPhgXuo1QNRNEDSACps48NjbQYYnDv1deS
Z0gUCuTswXsJLiBBCyDi5CS50r3L9Tvo9+NLTwed1BjrXYjkmnejP2P3IAKX+TONhzY5dB4NVH8p
RM7BMHSPMVSXWfCwWVEcyqzcUrs6KGjk70lROHpclR/ynyGYxlMOSkaO26n8sbXFSibfGHIdh7uI
kMnyoXGdhQQoGCROItCEcDEBlILD4GwjBmhsIb1LK11YMs41/DVQwCoW1hycdGXjCO16Ly0YLJ9L
1itF6USE30pb79eft2wPkp5a5SWHRs8QswNG8j1rWJ5CsXwrut2bTG/OKw0rb/m8ILVR6XM9ZvAb
GPQ2tQ1C2d2Nqp4m31zkkCPSkf70CZdRNpxovg+BSEWx+C8N549Fxtjw7GGgswfwtFqJCUmHm/Lm
seh/IiLaHFacrkJMcMI3E3se9YHWHceoTXNspT1SOlPazlQ9/tkVTfTPVnPDdO4PnaBKvRYdEst3
GeyZEdJdMKiX5cHVA3U0faahrSr++Q/hN09FxT3To4OwD5ffW/HWUlYByAj6iGWGLfRCHI8XQqH2
1E4iEVOGax/6tyRBZdh1RtU3LkykplQB46MEvhq/8JVMplu/U3W0HBDo4wBU8qc/vbYmnYvn9f4a
qiQpLg6EUhsIcp6G1VPunanetbjv9nb9UlD3eYadrnEK24AOsGqDQAb03AamiWQy58Ai6ghiZ+Ia
tmFRGkHbQVBmCQRigwqzJ1zDZJL+0CDvi5AcY/EsvaERRiznbxHRnzXmE8S3HoHRp+O639yYXdjR
yHtw6N5+srbF+BKOy/55LV8GCEGRkfDxllpi03HlNpyKsts2808FpKwtqqk28J3Q6cXw/nq80pnA
o9lyLKp7ImidbSPbWkacR8j2hGRdWKecIr3OcerZPmKBUbPbMXnpQViibCOdapxrWguNYISccFIU
tjgoCO+kkiTAaBS/cVdFTMVrS60Smbsz7EaCZu1OnbT/sFo8y9y8pu7AiZcFMYkArVtysXBpJzcu
yc/oOQ7hhWvyU/uSxNm4Iq+iZP3fOWtGB6go75WVUnI1hUVRivQIgTJEmVEjnhUn9u9Xc4qZ93Bs
qGQ2t6INWXV479joRmYjCW9Ssqc2hEmqJ/ed40OW5uPEuasU5amdOTh5DcXO725IdGZVgyOG0ZUT
/cydCSH8AiO9+S2D+2mZN+6wv5OkSNFbRG5nTljHfBhaBaj0rVp4/VXKOO2HLK7sYk+wwa7PenvH
P407wMiExerrWgIe8DIIyqZcvvEwq8lngduQiT/+5bmkSk4ZeaqzJ6X/q2j/qbRPe5Sxz0zT6JDM
oTMKuf6hxyLmtJMFRJ09zyjW4unRsibwR/M2/udcCdU+9o4B+p+eFfPAoWBblKS4nz/0o6AxgK85
N5y8cm0X4jb+mTtj4HEbNhsrljPUy5qex1Agogdiq8ecSnXPuRgt8CjTLcn1qfJvOZtcjgPy9zm1
g7IDnKJXn1IDGPegnNDLU2jS2jX7GEwaOXG2oSGOTVPYB/ymtn0yujFfUy05lM2FvcP4S56dMggQ
v6UjzeTP8BKG2o2t2VTGFnL0+dOzhu8huoBGOwoFVnmdlNRHlZxS0YJqLncF03ga9dsK9MqcpLD3
hPUFJm5qgq8vhwlpMebT0LXeeHM4JSeotthlbFlzMmtZgEniAGa3CvoXqq3IbQIGjd/z9uNpICqc
MP3HbBJPMM7KMbZeADqRy2IrYbanVwW5XIFiXdo08OlZ5vQX1hG0xZ8LcSuEmd1v9MHghA797ADd
hRPR8vLdObzEtn8z5PgzBh0ojRg/5xDp51HIhqQ3xW0r2u//kF05CiI/0o0JSWUiJkP61I9CMX6i
Cqvlrkxfgz1y+Hk8ls54EPqWlfiaO5o8/OLCdN318RGuCTHj6vtxXbEdgdiV+ShkCiddR9RNHbAB
7O1bv8bVCQy+/dJSw4aCxdhEyx1NUndFmxr3A2zx1qP8rxmwe6Xdh9ecp4M7OSRg1ugZzM6QwHtD
rJ4VFAXIkPVaITuSp4hWt5fuZbuwnh8E2arsXu6HN82rgcDXHcvapLSNPtrBqjWw02/s+cxy6ZnH
DW8I2SBx2YTf0jIhrwsqSOMREUcHoviMLLFOHVo/T4pMZJl29PTlhUqX9PQG9OshCkp+FkN571b+
sVSGC9A659CoqBW0eR1w9VL0oXQ+u+vsjFfCG5gSgPQ1T19H0D46gl8U7YWgGUK4zqGnxZTqzLPS
7gbo056ZsrZK6Sk04/Tkg2xSE+K+IKNtU6NpZ6LQRDjcmiU+bUlqhEdFWrUVYg3+10A/Q+eSFxB+
qlRSxY5sJ85EjZ5UrWK7/iCjb3R8jU/GRj5S+h1rq8w6W493VisQ1z8n1LmWOD39/NhfWgI73JYV
ETjtcO2Xd0x7OIJBaP4r+SY8kqXU7rhWudTReMacd5kiq661lzO7CBsbDJCWUnemHoFnE2oJLD+L
UpuDBNyI3ebMpMzXIMMDpu8fL4ID6ekmH+pw0nGSLCC80+xLgKiRvs1mTB6wLA41XB2jbfUjjT4P
dr22AIlEb/FcJeT/P2WKGNgE/Yny98QcOpZWL5SBdszIb78YzQaQ8juBR0t7huzQaQCmfouBPgck
y97psSh4zeX38++MLU/75XU1gsB6yNuObYXIPCdO6o80I/xCjqtLE2TDz4cKMmC7WUVEDhnrqSmg
uJVNFdc6jIzNacx5pYzahCdcRi7tDuuo931UTjzsO0MeDdAgQJkMu0D7zV44gy2/VaQbyotnV4rb
U3JReDG5SwqTtt1sc65QdiZuvve2JJP0nT1ZRKgv66Keied7XneKzpiJtDiZUKjHA9v+o1/2WOul
agqfvfhEJEuMN6jORHYSzpy5186Q2DwBJL4MQT8AjE6yLD7FEQYVawuEx562z7AYUDLszh4gRwF9
D0hT/tcDF+ClsheAQf5L9k6JOKKxGgwjdVy7t3UvsMEhD6RZgrpr5bB00dyhFw3nkwo2uT/ye3fI
a6QQvKbwIbERl8wHdyGm37/cZng5q4KrmisdRADopXCQEWX6j9yUlb8V1U4yrp1HOERuqUJ1JHvJ
RpihWlgwnKru3k5ss3oLqlAgV/RvAUTuKqgmufYHo3gcXxKQYPMNPHo0yz7B+1X+pwYXJAcJYuUo
cvbBPPV0ftiNoZE9J4cxcMHVN20TFvVEJDzfhBx7Sfrnl3xz3FYDyxHftpMRLc6ybl2yTVos/dV8
L8Bm0K0NDhXxu4jjtXSMIMnXGUVDcL1JbSo/ghlQiXhIAacpqTloJr4fuE1a/avVgiEfryhhJo1S
vJqatJauTHTDvvIAtuhdhPpqMydRXEDMygkRvhuZEJO0cbsaIjha3Z2TOp736glUE9ldhyvg5jlb
CCLdkcQTyf4yhdykHInhb4o6ffgeU1jmieHVO8OBQiFMbpdt6YCWPapj0BGuLfLsY/nVVopTNtPi
kkz3MXCqaGGgMANFFqA5HHv+c30PlPZxNnBJZg8p9BJnV46+iAUXOSb/WyYct+XPg1jxt7k/he0t
Z78nmWR7od80D21kzhxK6ulSgMI0XWWS9bnLDzXbPZwhYI4xOamU5n2ms+U1MtYjhpau4m63G9Dg
OG3sbxjjkPgt/BQeI6eQRctG8LVOES3gllbU1FZEry9H/XzvOlKYMAAfdcav6rUFPz4lOhYDObzL
CDif9xfS5c3eGFYrVc5gOpH91q5jmkxy66pXn1qXarSSh5reAcJa7SWD8us/wp4kLsx7//VHqnDP
p8FAjl/BWnqDSbOtOyn8N30/ZT2PesrPzjPn7zs5KRQ23WM7krZAwHZmnmcrOyTaLDdFqP/oCtTW
ZNvX0ntQSxkswgBWxWxIqNYV9tSqcDLk/wBr0Qaos/NT4S+tcifywDy8LfKsRY1dUWtjeupJwGbe
dMweUn+a1AmF8H2J8VHo+PC2MmiztYxuH9kg8u2mWBaa2XAIleBOD44bmTYLqhzfWbApmcw1pqSH
P3EeKD6TCUfQJXXgdhVBvGVjdnvWMak3JNYKY2PaC2Dxfymsx9/Uopb6TXAX2VhQLiFQfLqCF2Hr
FVTg5CaXYuwrVZ9diswSCkra4HDXruIIHVs/PttWv4/dxtfGmUkPh0Qr3BzqOZ0P191vGGC2oep5
4U9h6CUx6xqbt6DHm1VEM4QayMXmiF3q/oekK12jsiarIT/8BYfeBhZdtF/R3h8doZKpZyZbBQqJ
NxFT4SWAvC182Yrrsnh1P3gdz+lMI22T3u7gFQi3JV/nBaC7m56uMx30MC9TkyBBGJ3pTyP/klTC
Ciinrf6fr+5pGfzA7rZNzoL08+I3Moz9XTelAZAt+LXv5N2puw+s/mPqK8FxNz7el2MLzHP2zPUt
qDV5rcqojzKdulDyIJ4I6FhYLO+PrVOylc9iefBMolAgEsS30vpTKX3x4lXNolntwWAlWqTZKTtb
ohjnaniKfTqd27/BBxju2Vjn2uBbCwBSZYuypjWlTAUYaeIp4nH06RKRPOtqdpp6r7nSuweGXnE+
aq/pj51CTrV2+F71is1zaFMX3QEdnlhBCMOtrXHV78Qp0gCgSpUdbnVbhyl8a9L2k4YXzIzbYYL3
5RashFFJrXN3RzdNedObpUS01GYIM75Iwf5LNBBDeWM8lA/NMUtefUmeiVZCj/rRDHtEE/UTCZ+m
/2M8RHgnpEDt4C38dOsksWX9pGeMrx2pSR68eiqByIACO8QIP8b1o7a7hN2fxqDEOwBLQ+gqgozy
jlSsweH13j1wMO0CYzX+lxGwGF4tUp5vQ8QXiNLjppIeIjFIass1nQ+cYiBkcPwsIv4h+u3MFYgq
NZHqidYT7J3B6QBNaoiqTyLglDHF9vata21+Zil0U3X3mkSFnNxqOdGsJgd+jJjq8/Z/EezIk15z
uvckdj1Ca6DfakqSNuEZyBZvjh60NaQgElkpHCsxeugOBwMtGzjYGVUJxCHN4fl+6sNi9yDWkj2/
T2ZFvIN8/M2Ph4F1ne7UtPQgMxSD04VDBJuGR5dr/HkQ8l8ZjNriWfXTv4lzVdbrNtu80RJxEpZV
1duc5zWDNRfpn8Cn2rzTs0FpnxLQjX4i8zPq4DZiet3VjSJ+RuC7VueibR+4QacMPzK+lcQaOyr5
uRJhb5XeBbs4EUpyGTIV2pVJXIJIhmTx2mMKpw1xKj1BzLBEdJY9wkk3LGptHa1lj+hHoMaDQDh/
nU6pOfs0G1FOwrgmX/HAt5nV0/WsY4hQDDeAdpyk7G13sI0fTNKx3R1sGD9cDhNRHY+P8gD5CG2T
vHjrFaH7esWQSWjCNMTZecjr9gmHa5eLgEP0nPOE6fZH6ANHA6CM9yv2/r1q/X7mcBdHfD3y0anf
oy/f7/gcgZRyGSRVSXN4aY+IzeVaeAD7BQhPw6tJnB50nbw9SW+mgfIyrSedjfRlt9exFHgkjdS5
uQBdclGr7MW1fTmyteAOmgJ/TUZerOiXe7FXx8b5t9V1mdSX2L8Etu89x0lWvIPfjK6IhDnyrYK8
0nEDcBn4gCtBPj7nDNZeEB2eG4ZpOVaR/sPYJB7vgc+BaQcsqKrV8p0zKlEoK8d5Mjyuhycr0Fep
HZAw3eC0OA5InphNnBrZXzTRdElC9AvYAKrS16O1INBhpre//a2ViBggzrl6xexaQC9KmEXeKOC2
c4BkS9dAGZAlNNqirl+dBMrC7WmQ/0yiCH45AzUrcFV6mQnjgGx4icLIHBxCwDaoRPdrY4NXGroI
1L5oTpNMH7ofZSN2uR7LtcdDN7FrwjWxl3EWNVfsoI0IVWC8uYnmIvyyBQIcibXzzBekOcRDa/63
qoK3JX1B52PBEayC4La1sy5LSOQd1zJxba0IQjfTeddzbsmv2KkrFw9Of9mfTUYbkt7XEz55DFaW
09X85/hFTyl+lXM9jGkSnFKLO34UKmeONnCOgi94KTpfbZyaAeP+zlUZk2cp4Ok0MyoPTJEmelkl
V7GsCVPWGKOqvvPQLT3h1H/k9r/z2wznaWIlz3m8fQBGsLRK4LmE/2qx24liQzsFX52gBeZq5Izc
Yk3gogyAqnxA4M0ZqJjBo85tPoTTC+kErJbBFu1uqdQlVL8U5dHNwu2UDv+BBZW/KMBKwLm85EG/
nWpz6u/dtciufpsLPs1oWWm7QQ8HsO7Sx9uWljcKQIzxIYVXsNe6DHY/RebGaQ5s+t98iP89HKo5
CQ38H7SEaa8czE4LOpdlI/JtDqJGARLsNJrSwaRVVEIINzKoIYZXdVJMu3Cnc91bfS/aXwWtYpNu
pAcgEiefUbtXcRnJEq7s71koeAAxAvSx0pie5xyYLyMvzTb3mo+63PS1EzCDrIanHx4ZPFkqxOYE
hghoAceb+F8v1GzfpMteqM5QxSKy3aoMN4S+G3G2ZPrfVfjBAoZWU9hb6fvjsx7AcAP6eM6l9W0q
ntt22VQ6SUcsW9XBbsVEhbuQpV7MGLvF65tfrhTnHC0K/CfRYV861i1sS5Ek1TbBpp5tlJsFtd5S
QdhqjRhZ73Lv5os4lh8XIPAFB65KKaF+GPYaDiuYRRbSMxO0OdwQlaOewJe0NBNdo8spjo/0Exml
c7i87i52a66FkLlP77dTznlyeaYsjTZoxdTsV1UdUgQCXymV9XjHgMMt1xmO63S/qEQXHwneBXSd
Xuy83VQEsVcVNgJvBJKHGhLus6cD7MUbSqR+6vyzQQVNP08IG32Gbz1LDuRW1yxPiVsf0YjosMHI
8TwWvei6HphYb8XM9xP1vpyHkB2WnkY9jv7o5OBC9CuWIiQZSYdROBdJLgcdyVsxmwFMHtdEY9sp
CitVPr6UGy5xUe1Qumjm7Hd7jyFPadVtnuhytXYOtI1qSdkp929TWBwqCRX2X/7k2L0cQVNY1C6o
eLPf4VgcBYisJtOaPdEfUW9xxP0avcOUfxVGuK7Lptic1gAfHYVXdsiyl5SeQe9XrAFBdZB09Jty
kPOU40JWF+L68ddUt9MIctaI3jbQNYPRA0skEDk8XatsAdOxuyroYunC3PQS7ovW+QmgoW3GWVg9
W8e4NFeDTFIztU+tvQz74A8UpHLTmGlpVV9afvs9olYRSo2EXyDrfyaGfHmCZ5yDOhBrEyVJ9ygv
iiSUMcWVi+hiTQW/RmmbTHZdUyJQzd7aco0V33rOS5yFxl2OJmUa52YIXK4kBoJYMbe0+RpyRrDf
0f40cFd5uf91zQKv0Is3KKpvsuEjmst9k6tvbvJlqrq6y5tnU9E9qYous/K+Wm7n13HnA3rkdP6a
mD8MTtqmlCFd9VFf1mI1izzofISxFgHVMv0FKsZxAAVL/SliOcdQk1r59hAH2FtmsR0o0PCE08SO
BZTmp/YdpRzF/Z8FyIhL0OcVzfewDbQ1Uutrw748gJ3S+UP7Xa4cRwOefmW3CF+KzAdxBFyJjYbY
De30oLXTEwsLxx4l2LEd9bjj50z+Inc965nl8Hkw0mXjZ7eUAOzgexzl7yEEWfQT4E5KmmSYislM
FGlrJe7bxxLQ7Js+StaIZ4YshaGfvp9eECobK/vZ2wxLx7LanznlYEMLkpXKfJ+g1+USiVHvRnBA
75jHdp42OC2I3GbnxKoeJ+gTUakIodrEFTRVj8AkObznB68MXccpwg486A7YZQFSqp2PH4ASjw2X
c8lbEmsDOPXBXRdzuMiM0Ghke/gMoDGK4guvkvoYt3wzeT9tBrZUc5jIAacL931jXNAbLHkqVAcB
VAZ28Drnlk5qmgX1Pj50bxmfA3nrF6aL7MAOjsfZVtL3Vu7S9uMOn9JQ8pnEWUylYbypHQjIPYcy
X1dR77YDdInPl4wK/cXgoeV9rlFhs89g8xTdqDUZIFkjCwljfTpvJcurJlD/ZI8mpdiIyX8ZySUA
NU6VEzZNvZi9i7ei/aLYEQEQdpwG0MdtQtz5ydvERMoEatmeynqd6VXX+ZaML4MdXImAoQLH6Lsk
lHpSqbZgHWzb4gl2SLGh6XLHDb78mhKh8tXj3N4I+UemeHQXjux0e0EavV7s1US76PJ8MDN97AsS
QmdCZjY/dRG8B9Lcxjr6J8u6mm0V8VOYRE+f1/sgyf80kYTEXuqwFTCu4UKJvSsVtkNIckG5WW5i
3w7fssW8L1MDPgObC1bUlQXo7rYXsg/OvCf5HYm3lx7u0uG+aPERglmAdZ6Q5vH11cw735r7ydRg
U3Jroxzmi0mxZEFguwMZiZTK97CIKvkkDZJeG9yYAF0uBHWVEKcBUOl3Wan0MyEqfrE8PmASd79Z
ggzqj8YFgIBrufI1GhA5jomljo+KM1gGlo+OllM5hOr3lzp6f/8DZcNfvIWOZPhtckmWxT4UBv/O
qpj2RjjIGQsxKuzSaFNmWWKpqqWrujbFZgEHFZcsIK0vhk99YdBfYi1nbk70XlDCA4A+OMUzCCNi
Ze7UliQdph1/lYV/ysUDSZgPeFI3Ln/Bb66frFg/OtsTanOMRBPHgY7BPnqMBiVxhzTkhWTngHaC
GeGnPYVKP8PVZYLmFmZYe+eWCwign0u1RQOEEdjiVhab9kbbeyQf48OwaWFAoTz9XsdFFgll11+r
nZSlAC5oIp66geO+kiQwPzU5BokSqf+MAcAFKXNd2iuFmTAl+sMWbuQ3ew7Fvuvw3IqTiaxTmjBg
ZZvIEJtHEMSI+1OegY9fgLIliupgXkQx0sT9n65Ro6UewSUPJ87QhNt22mZ7rOR/3LZUPDHC+q7j
o5ZHdHIXcE9s43CWH2E5BBaSI5zF30f5TaemStOSgXDR778NDCLUZL0AUBz5cn4Oan5NWUv+UCg0
hNZMc9a902fvEuF5UzpFBsMt+jA1ZGoSiJ2JHp7SbfYnEsUWdI674OnOqH4PNAPzaaezGgTdJhvM
9nbb1oUaoglGBCEGIuDKBsqMyX+/JMkzlXVG9Mgumc3dxnv2IQhzob+UP+skQdG8hjBjXsdkoqxu
+Jm4OLbGv4DUaAAb+ZTlcpoQYrmAgDvP3OC38Ru1oKV/QE/HveV9DATDHG26JxceSdYJ3GlFMg8q
QBCrKwmOOXwDTFUxoIeTu7+z+Y8a+qLRSl4wIb/xfiYhf5GcAbsbYLMHCLv7MWAUXQd8M/mDRC9+
KeOAMa32Da9nTHlhfB3CsbB1THV29T5dSjyu4OQVqOOBK6mHJ9epPDnFY524P/9fvywzGTPNUy9M
WgD0Gcqi+cs07QgbbjRLix206wb0/wmrl78iaNMSrUbNmA/lrgo7U2fM1PEa20Fy5Y5PhkYGveoX
yXQ6T/djQ8eFCPzUFHuRPuCnLtbtJOkgGMYy+w6uxaFTevOnbgkbjDKFt1Lwa4ct4aLfU0jt9TYd
sFTmBcGmbJxtlR3EAxEV1W+SZ2kAElb3TYiDRT7m+M+jCh2VKO3WEwj91feF1IEUySg0JimNOIvI
PkkKA5GDqx0XPLn9dxVzrEU0YTLVvF/L7t8q8tPXFfjTnMytXR+HV3masdMa0IJpIWieih2Vnip3
7me/yWMgPatHEfrI2RzBlNyYtNVdrUgG3cV66dvtLHM+8Q8yWeROTTLEg77HkI2dMMyxHY9D4Sdf
BXWelBESlAbLHkWE5NcH3bJ5jpg6b2Vz5Ad3rw8YKf/W88ibEDlDWgxEOzm0vE8736aca6mjMd5q
6sSoUCISKWJaxL2n3hmyoch6Isn88N9yTeQFt2Co5Sy9yVTpSmgjZpL1mEdpSBjkgnj3Uv2XKNmH
QezZ8ugmCYlFg3v+7XkOowiizk+mqVR9es9qLYN23cEb9+eHbGruAwYo+WNVLjJK3Jplqxzx4hFD
7WRuF4rfirPmdfHT7YEN9fgvXmKVhVGPRSem0A/cy9Zg5lLh10c2ECVCohSTivGl5kDqP9lABMK8
9gJA/Nw6HFeh1AfmwseY9TKldHnT5HPp61NxGFFT66aT8TW7hOwV8mKzvQXc/xYJ7XSLz5s5egcc
uiWGCgsehE8JkzI+aadpd3c7Qg7UAMOX0UP3sEViVvj9epIXkf/u7PmLiY98EjV6J7PxCXZ6Xn82
0RVEMY8pQvs/XxOzn64OQ7a/bAhutOX1k4qSsML81MB8YDMn4bKn/eWYgVeM9C/j5FuySQecz8pG
hBTegwKWpeOgruK0jWYgcBp7n4syg6P5RQUzTweGLd2PyraSAD2j+JZ9MzboNE36Id9bU0E1SHFW
LzmSMQkVTuFGfa5hB867cIH0OYLhnZKNvF2pghD6C9FlSmSHnuQiWMUGrkyOQvLbAKSraCv8RlHI
cdMWCapi52yinuQCISsafbX7SM9PUn+3JlN3q6AMUmNuayMdq8iaNFcaYB4j7ChRNkoLWcvL5eB+
bANgnLqh7ugya/AndAuQmyhyJsREQ+VJ2gv+D5VHdC+92HZYRzT9WT13FB9lV3aELpHlRpVjpZea
aKInKuYZbpVs/hadDD1ANCaFvRb7nN9jLytVhFvpdvD/S8EiTpnTNcliIzKuMv0sDZMw6UDWrHvH
JqTk3GIOtoPyGKd+OeZVNK9ejl6g7gJ9Ky4lTC/PUubSByK2QjkYd6LfXBLoa7wpSnoIi41zGyW8
HhYR4oqnjNMYM2+PNTry4pW9XafNdq2ov9K0p5bzJzSFoFCMnGwqtpJ4Y9hJv+Rel9ffCBgSoiMd
WHB3xh4qxnhSNhzqeiizeWMw0vJoTJ/+VBhXP1+aSgKiqtZEGI6fgbYZjhxOv6eIcLctEu4Id7H2
+3UcmGnYWC0cyGZl5M4JjascU1YWvS2Fd0aUjad4vMhOIFBbTEz4jz0wOO/q+PvtcxjCvkB31+sI
v4twJCWIAQt1yqMMYj0fDSQ2ixdTyZ6skqYs8DYsVO28VafV+X1YU8M4qdFJuGHUKySm6+NQo+6W
vTulAC8tCn5avmUjnxhU/h42ItnG37wfIRWPMPujr9Bt82x6lqIslPib+X41f9QncxHaBkn5ZASk
Is6oOJpTnZudFQ1syBnaE1zcObqpKgtcUbXZPG/hB6yyKv7ahUwxRrH8QBLRkJs31E/DRNIkeAvL
U/yz5XyBkSA+s6GWoHz+TAOkEjDvqdqxW9Ou9gwjqO37+KDoZdA4BcGF6wb5+JjQXNQ622WKwZHP
0bh2uAyFbsxGgDeMSbzDRUETyoWlHkYIFiDgVVlToB0L4wf/RfD/R/M1sWhL7bCT4XxLq4R+sNHx
6pXXL6c5CxP0zqGKGp0XeIJ6szh4XtFHwjxGfdBkUh+h45WrQQo/yK9/iZ5CZ3bE+Aa9pCXZ8Ngn
LK37gJBSE5DSS9Mk74ETr4792GbpzrO31R4Xufmku2gjMlPsfgx+5dklKVdUsvlaTdiV782nIfPE
lYJNnrT1v4XLNUH7TonETQfAiladLx7AL1YW+nAN7bAHoouDm/wglNL9lReQaZXPEkPQ0tniFfl9
tBg96FnwRi9tg0D9dFD9/Xh4BmGgNHtWBTkCROD9tWA1XJc5cWHMMVsud5i6E+UcBbYSCxKXL9CJ
vyvwyavVX38v81ZLyl2q6Pnq3ebJ+zmWU1CCpetgcLROMYWw4W/lPwAvEJunXQnqgpmck+MDW9eq
EM5qOh47RbwiGxy8lK2PodjJMKyXwLWM5QJVVvlT4nTdy2YWML95CBbt/0OYS+q8co6BhP8cfuS7
U2sF+2qXqpniJr2AAFOBb4TOHPuIEETmZGZvknD/2P2iCHCbSjLjIAfim7+zw0e43M1FI/53wSPz
B3KEkati37pNJBgcJPoHX8TG8t9mbSxBccesH3mvqiuO2w2qooQf9PQkvvVqpoVIoynoe4piuM9q
DY0pThtSR3oe+dtntro4oTCogco4AA6wG/o5bG9QGKWFEj5y2sNt3CDt+aAxfllywjAWyYt+/j/B
BBC8SX/oKw8sJgFcBYIWmL3AHPmzPzGJQ9rRD61GE3MTiTraBJjjx970dpLDZAD3vAF9KtovTotu
gTYdN2VhoyPfVtd64cXmCOnm11D5kSyrOlKXnbhdjfMyrqTGUBe4fN7EXqeA05/b3kXrTmonPdDR
2UhJWrukrSSzMlRC4FJPuwy+VTfSz7Hg9PPABFHmTW8TYTZwi/MRuufYm2EpWetBoBKRjeyoGwNU
JouE8FEsfJuXhDmXzZEsmeMhY0Tc6ehIUFEHk/FxmDr4jvRLO8RjQ4qCLekfvL3HwVdbjGPh7Mp6
KpaVjeOVp9eiVFU4durQZr7XDXKYehMdSnFzP0HmSrGwX+fHw1NHHpKxrmtF6qfVcgIfuvnytW5z
3ZzVMHq5ACDBXVRjZXtaPPzbGes4fnfKkqGsiNPEOnQW3EZ21Y1LI/7rVdGERQM/6owdq2mDKvvj
ajF4FHRsEt7C9uBTONpdgtxPVgz7Gjk92E1wjreEUifUsKUhy6ZApzbQDESiGTeH0F8XrxyN8wVw
f1hN6xGP4vBlIsTSCP+1IroqMECFYADOXibcwkiGwzBWven7ErliZQStM0ru2AoSTshfnHi5vA7O
FEYWuYJuuRaGtFVFkKKC+ZnHpQMjqVydZa9RBi8OCgOgv9ukY1nkoDkufQaVrbwyY9DutMiVtCA8
CChXMY/TIWu+mcM61wOVyaOQKMb/J81Lj7Is4CKof+8jxLO52ziVGCJCucu4lReKFq46rCiddQWP
Lm+0heDx3aRadEM2kUDIwmI6DTzznwZwkcobNFEl1blYtz2BH1wtR/p4J6mUTQaIkBmqoz0lYLKk
7f1bxnhX2QiScUiQLPZHSmvms15jbsV9l8A/oHMkNJt7k9C0oHKciL6yt1HAYPQs3zq66eKbniKt
YIC2PSUOlemVBQHBbhPTvmw8CrE4MSXSsjN/FrLpBtT1U38txdMrmXPyY+CvgCf54EPXMCwNtf0u
8sT/Wfq9bWztW6HYap5k5xqqNihC/w085Odql1iYXaYq642KipiMhb02pr54XKa12g/SCi5eWAmm
RogqktJ6bvHDTHBfOW2/BBy87JPZ2AgoQV4qbxUcLiszwDtEKea1IBR25ppCJZhYgl8vP3tfSlfV
i+cEygTvZQSQdyy0E1ORjfUQk9j8KBZdCVYFd2aqdExBedjURimT0xNdmiNA0rp5/kxBpynXGvLm
tl4SlRDvhEugJwwC9qhzVdscnHSUOmNeol9ECUg1oLoYoH97pMxohsHy/0LLmNXuYqJGcK048EI1
YmY1VG1O/UMM+X8Pk1iLk7f8OuhX5G9+CViFS3Zh8zO86NSI5iKgERtKQ5pBsXbZVs/blzc2Mkdj
CSvz6PjWD4o9cAf2LaYuJR72hRCPLH+71GmQGVEaSQCGFza08/sG2BQv3+ikDl73dWISICru73VI
8+X0ObE6cQTClzyK5tHz5gDuLxlBea7N6EnMXHUri7qNfHYwwGPhryjMj0FM6yolGRQ/cjwS4+s1
hFW1CJwZ+qMp65ySDsEQXpFr1GnOv8CVnzjsRTFqXhfoG/j1rrgbsHnkv6BU7jNS0fdREcYJ0+qO
nNBYR4+/mLbtcNG/ZNU/TYupyiY+zWeSVsletYqmzyhiWB/Kfc2LMi2kehavOiqezOGUrLK0GfBT
Piw34o/Ss9HLwivQ2mtvdxH8Gv/4YFA5y0taADPyogX0bsnYhMcutii0yuZYnRJsWNacSWcuHULW
A+4xX9rgYxNw8XH530GpQoQX8lWlOPofYMmeaGFCbz6shQWJqJHsBsZMAtiMn3sfBxTxxct37Dgg
aQg6Fx/Uh8naqTYaHIBfVrE6+kZCAeYyt+AFLHJj0sEdBG69no6Fu2QRaSUrk4Ztq1dsW7ShQDpP
B0E2gqNhstWWtIw2fRBufGqq9v8Wv6cV4OAHMz7RWq/TpcbljMY5LYbc98zulM3+aGcft4sRz4KA
9/M0Cw2Nhcf5z5bX4/wHMu8VACHEuOOsqMp+FgJDN0Ep8bKxaa+xy8ry9/9+We5tkeiwpz9zEra7
cyXElPjPtOjtSoDb0K37PraivL+tKvgANqiYwOu85k1Es0UvoW2Zs6qqLVNvwZQ+En+EgGe9VsMa
AOLtH5pue6HBc8TOSq2NqR8iGV3GvQUdHDhn1r/bqWdXDbDFhwk7h8XUNAJuNWw/0t2RkL9jhfR2
Y9KW6TGiqztdreKPvAV+/nXIAvNKZZPkqxIL6tghS9NQbWUGJir5lHvC9IQd1rpIkRp1E67wbG7k
uTxZDpkW8tNo/8oo6EtYZGeFhOMah9CGfFOUdQydqMlMK2/+APuayFsnpI06r7apk3TYsyckHslU
wVB5wsGjqLnK7oq9EMC5zCsm2Vci/Dm3J4MSWslyJDf5jCzVOiCBDfo7VnLu0VTipC2XCpqW+9v6
8BKQbAlIjfY2Znnp3jtdNIy0vBNXS505srcyGSKfW1y3DcW0fEk7DTZCioxk2bcFIvA1OTF8fHLR
jYherlUSd34oH6Xb6JQBceQiaXyBwHsLulLRRz591oE3+UkZTkLH0uNljHvvqO+rFrGT5F/mFD2Y
0J0iHz0vZNvdfdgvYxgmE4hOsLL0qLXapocPGNrby/Dd49IkQaST1LLVoj5Nu2fkIy8VaUyrhaun
NSQFslJwODlHW8bj13+sndnkABIozqyjrKCuCXPagdwxWGLur0xlrQgdiNZJ+cOF6bsfOmK5HLbC
XnGutzpGeVnBpAoU7VYzTI6l/xbuHS/Zhd69zEO0XT6fitiH+l/ZeDrCXhZfQ9HDErSXbpPfFywF
fWWB2naQXlmm4HMXXoUJoy4x7J+QCbpnb7YUNbvduGD2PpUihh61bYfa0zYZ0gjnhPX3aFYcomOZ
70yX0CKVJFasnyRb5Je0xKPMXYlG7JxAemJmxQfoUjiXbcEc69AMQLmH4yWvucbgbhRxaxWOAs93
3FYPLR1VsewdFi507Ft6jsgurlGV9Pclf8B85u+4KOar73I9xhbEDnJuh5ATwkCZzh3pcpD5Fs2i
KdDiwo7Ka2pmR9HZmxv9DfeWMH/f/pWZP80xcKXROfp+Xov70dkrevLWuQEH/um59faYcBgZp/jV
NadEIYP+oOcIVGbSjERPkhHAiT7+AeN82B0J6PzIu1kIO/URsQ/JyhnRXB715Nmwwvv8YXLgC+MT
FqB/b/arWr8y+t8OxswVlcmkmd0KXACxyZUvlGmVKGEa+Tb7GSyEN3GxM/8Uzasqypgl0O9m+3fv
+xpvKYZrFrddFlibJ9PD3+sgjYKJ05HsWs+QkUv2Qid7XbRt0DCiwi3FCy/KRrtcgaSTx47ue6VG
0kIEobo5HwlnTBLZEDLMl3KFibtKjDoUw+UKpjFPtoTQJmWzdYf2dUyv6m1dXR6pSZ/Q9houw0wh
Cqw0yZCZdOmajGf3RQH/CRfgu3h6fYUCdVmPR2/C+MVfpOsASUWriOKl+NsT+1HUjBnzQOwaXYaR
0mUGX+I+GHtWleROnZGKXQq9V6ZZ3vqcpMDS4eoxeirPvkj6xLNXHtMaitBq5wknQV7RIJaNDjg/
U0sn8pmOVhcW2zrUfmY7WCB5jwnX0JJm/I4OrwS8DiAAwmeXycWFtLF8/da/JchV+fqQKA8ZZvFX
MY4ghCNwtIy+1MTSaQcB7ghrHV3Drhwy48J1cXaneyAsMR9Q9lm9XxFfG0lj6FnG6zNZBW0NRaNY
JQRBVj2Fc0HJJtQhrnehMl0BeyhOqCm/y59AMZ4REXCBJNyykNL532rBlG1VHdpwWg2xjXwVEVhw
vUZ9O5Yavoc+chqXB6DjK2f/hQLE5YeX1vN6NfFolYGkhutFfrbHrUCcMUtHH1eGVgqmtgu2fqtB
gYrl7jMb/731RMQjxOYFawfb0NCTh/SWr5h+brSh98RVoBGzRsrIRGaxilzmch69UnvCqY2kFDCK
5QYHUMTogsec2/+vRMzyWj+qT/77U4QxZWQi7cUdRopZvIrrnR4zcLUHjfDG1OmUAFm0y21ptLGy
svxkwgfC38x6QlcQmPp9B/uVSBsPhDOtIZGu4Hxy68fGxexRqTQmn0NinpGZlgF38iR1UZMMhEH7
RCjQC0ovk80vSvfwEW9sByHa0JqqG6YAh8Nf9ldVk3Fn4T040gxl3vBbDj91H+XlxB9DlGiycI+F
vU8CBLBxDrxQs6Mgs61odJQVubI2gzJXQ+EGl1EKh/eCH0OcLwzyyByXqPeos1pp0NilIKB2TLWZ
nJ4rbavi/B/Rr8etmaW+T4R2ljK6VYkTdO+E1uBYObIHflbSlOqjO8PrJTdLYGUrgD6cnZlVcShS
+l5cxPsVzlXWn1Nd7fYwwRlU8NJQTuSUqUAjsEVEVDkQIWXfmrCIvGpNR0bknu0uk6etn0t8GDa+
PLat3NjRqsI5V0wb28dU4rV7RXukLNlOo+eXLQFcmnvlU7gFGhqKs/8M4HGLO4juzlzsGjT7eD7T
2iyGhmLi86orPFpwXTOZQmlf0hsPYB/O8YQl9tA8V2ioCoBq5C9Zr+aHAqIh7YZwn7EpyZ0JdShT
yftj7yrifrAVqWU4kMOX8KMw355Ytspyu9KiclIBDfKcO9/zGUZEyJwOeaZAuHvLqTdvyRUlAoGP
maz1eeg1VhNOGWyg5muNzMNjVY1lVohr8L9dqfEmNSjfnL9sJK3VOoZAzMTyyV7Vgx3Uw+u/Xcvv
wTvSFozJctJ1BGLZ7C2NCRcffMTurW8/Mpi9IWAbzVJ0yP8NFxCU/tZL1WO89EqNN5u2CK8K/uzA
XIDnMZLL5D6IlvovBuVvy0RVNnmmAzx4vU4rOx9qg+Zz6C90m4Sv2s20RxthEots19NkagyyrsAR
1QeAo5kcaExyg+K2KaT3/TCnQsmWBbflE6EzntnjTSPzElYQnbTEpEe49uruL+6MegWI0GYpy/W6
91vBXpMFII4xcIck8+TfrOZdW09I6Al6jrCbt578QuN2XLkBK6YMc9oEOPqVWUe8i0MRxc11qGWm
sdriuUF4dNFVW1z449kBTVr5+l6OZZtORAZIHMD2QDtpfADOEcHrrOUwvh99L408wx6pmjifKEgp
bNS8N7KOdUYgEAzmuFI+Gn5cSClHkKiap6Hr02osKA/mbARXzNtPserb6WhrZo0/FSLMj+zmXdP3
an2F4njMoxmJwRaERRLafqPuhM70yoB4HyX+7bS176j8rZ6ePl1o+yALjm9xnrHSVojtR3vJgtjr
7sevkZRacBCcTj6qjVjevdxYEXI18vUnieYEqx17Rze7J4pP0v9em8Ix/GmarnTHmwTgc26Rnzoi
ujm/SnK+SHrg16zFGmwm/6Ce8sV/V9ghd419R5K9rIQ2UOjRkAPOn/9XyWIxyutCYyxTutM0ZLqj
bZaxQ5MckPtHNBTwgp5CHrTJk1dB7BfZYw31lPZBGdOrVSkpmboum6YEtmcZpr94nqm3alksioj2
seWl4/28ktMfnXtDyp9crAoU3DzM4NvVOQz7QcrZYxphASc4XGaBnCk2p/spcbrLkvIqBfvseZuQ
vXzPwruAE90qS8IgYoD9dzV53FsoxEC7LD3oOIsQUY7TZqUjp2PggUNW8Tlo+4HQ3CvT4lBGKYe7
oZN3f3yn0J4z6FaDfHHaSGBLhFp8FKtz85q5biK7dFFpZc49yVBwtJtmBlGBT+N7VBzRVFjCptM6
Pie1dmLPkGzhG1imA0OGlTEFhozvvg+QkFc4IucJ2sni60K6msXI4ZNAK2UHtOTE1DlWBZque3Yg
+BpVYlneQEEdSgMarfTfXGB90fVl/bNQ7QgGRbBY8/pDS/FR/en0WL5rqrkHZRXvWah2rWl59Jp+
8LsG6QfM8X7llpHs/SQonJZC9LPrytvYIADDr6t0LljcY4MGp+vpchoiPyDe3g1Xwf/8d/f8KJz9
+0Vsu2e/GoDR3QORRmTS3MM8N5s2yQOI5hFTTT64uJJ5WSZL9hiVpkN9TaGtv1czaxSXzO/yX2Fp
lcLKtCkGXROsy7KZIsiTqEu2+9/IKl+SVJ28lTnapaX9sfV0C7k8n+sR25FRAoyR0RwiQp7u48bl
Py3Zzrm27dx9sRDmWyGlB1lbWt5nZ2/NoIoL3KSe1UtQIsnX5RLGUGeC1ebUCF25NkWl9p6ew259
o+c6SBXqmMnEPyidz4QoUU0/5NcDLRi77Xb6AxU6JFY2cyTLcrE8LgUDN4wMWS11Pcr/9KbUmgqX
rmzWgOVLeRSHufa1oG50L+QmVwwJ7VOloiljfKeJoffj7DIt5l0azok7uS8RKKm5FzVDtOfVwbOi
UCaoPHMb+bvF7GWt5CNXx1/ErdPYM653M/BArHqRxzqTJyWYkhiGnJqOnH7Xoy0yQMSNVb1/ocFA
+pHQ/Egw/20YMxRfR5tHzT1TSKBae1mWhpGxsMvo51ZVOpzwJztke4lYVxLkD24kFSYe2sKIqGHb
b1NsdkwBLFfv74RPVMn3pMQ0R0UzS+P7hWFPsgzVWF5hf+Cf0D8YJ1Qj5rFsFzKKijzyKwqXln+f
Gt0VopgEgEx4zG7fRSPrTLwFyKk1P9z2GnCMq+6o4jjETjA6jr04+b+ONoCvb4m4pZGELUdN0Y5s
kt0ymaO4/8Xoc8pBbtv4OrJ16/lQtKGMAL3aefzq13+XAZQ4Ep3/dyQENS+6lSIGBswnoxZLkenQ
quE11BsAV5nfZdQyh3D6TzSCt5ZQrKjFqk+E1fKvss9FUYgaAZcapoBMKG2ciQFEqsJVtslzxGU0
mqEpweSz7soPMwhQ3AoXECIVbMccljrYKiBv9RsQVWwhCfPxRcBkNPlUppr2n4YnUHxRFVnX69Yx
2RUBjaNkGbqJup3pzNFbauJTUiy3OW7XY6pm13fP9U7kDU216ZIEElfEIDd8TBZLU3A41017Hl7J
ALj5a+USHla/4A2/gQdxz7OV8Esd1L1D07kaJkUetRN3pGsCevWOePPNXBFDye/VwS9oJfmVzLp0
+66fL/eWjJBCQFGHwP2IzH6Ae4I6LDZRAupCMBeXzn5uL5UKkLnVtgJLCjQf/GDH2TTSx2yJK6Z8
WbRatKwdeDNsXvQ9u3qSUMf3s5IEkPwqbkhOdM4UTuDpbu56O0RRrUfa+uvxKOp3Z8iwiW+KMI6W
j38It9EUybbgHOPjkl0KBbYrpdBquFocNV/yKMIq2d0/HJXNb3th7wDWE3mWZgKWHqaiIG5htGPl
5/Hlptw28aj7y8nT/YjkuH1wJ0TUVMH3hHHTygBYyyJqjgaYj7X3tq3pAlr7rM79Wrk4CAh1H3eU
s+Iw3DZQlo1PZe6xzC6CO+gn8B6pZuO9IMX1RIIwJlfGXWAXSJ05px2rKeXHtrV41Yn3yQWX3vb9
a7fa6QZPYtFYmFQi0n+IGzriJcfToB5vDQChshMvr6oifKUlxNG3oIY9tWa2WvNc+qPkDgcy74nh
mn7UD4kMqP4pq3dFElREu6Ou9zYwnIbo2qnDjsWVXqciv5lvUqM/xBi4sJPU5Khaxw3i0lcbkbG2
FjbkRjCkoiu6UGM4XyUM6qIyekiJ98xcOyan6cENj3zO9tgU50K7kIebTGpk7U8M7Gz6mOFLHRw0
a+AJ3ng3TPVGkaA0icIx9Ad9MVLlBOLCwZMlAzqEekpopM9MVOlz1EL//ByY8b9FC3EOpGwjS2GQ
IyJ5emSQ0cTXqMC1KejrP/9rHjYnLVLH2s6CKieXikTEvSwVDrDB9ObbmQf1HV+JKM3PBG7dvgVK
9PQbZXhTcbEHab32lVodJtPSjp9RBaMdTbOBwo/R+P8LcPZopYrDL+HBLs4aNrDtWI0FoWf83Npb
qfiQHTt4y+Bh3sntCRoxILexoChh+oW8BqMRLgDOBZxagJDOWO7a5igRg5df1tmFExDRbTjlpBcd
SY6QtoJMnR3UojBl8OlOHMnVJOo7XUbEoEUiBlo2JWwsaTnvN3sKLVZ7oiYBUKf9aMGZYXu/xT6s
8hWieDJtqWLPYCjMfPYecfLB+TG0cPYkKEXsZbrpugEpev34TmMQ3/ihuPvaQKN0WVJIzmxbqqQo
CNg0ezL6UESrLQLei6AuZaTgVMipCfIEDQdFIXJaZcUAo3C8/hEfzMpgGf8pTdlf4jTubDV+HJmq
oyN9kufWFOp/x58+350IKx3DZcXfY722LndwNrfE5wM5NI+T8WeGZrRyLuMpj3JjIE8Y/LlVbDnd
rOPFve4NDM3eSIX2+QyJgvmjJi2LbKMEEtOQTrg1MNNMWg0aTImN8SD8XjOqTqh0h6sop3oc5gEc
LW2f/UUngEMiXgDI4hby4kztEqifafdlYAfMCoUrWYLiGj46okyeoyX+6J795gNEQjF8jqLsxXiS
eclwCqLB4cQa+9tbx/HrTEQHtssaYDu2MLwwLwiJR3BLZKdsmW86SivEk1KiSgGu34nZbEMOT5g7
8o0fPrWrD0S1Yrn3xUiQnLlMNdfp3glm1i+laDZ13uowWmixTrA4+GW7QeCi56C//psmDVhwgRDJ
GwGfwwo2M6JXFD0JNV4hIjcolbJF0be/QIRWL7aUS58YPe5wcmoSFKlevmQM0jHDdpfddoqJ/OKa
GAw6TDHKwRw4PdRTXxHbqmyQbxQS9SHmN2BH5CMopZyWAnjG6Tbx3SRqJfF7WtwLY4wkyPmWemii
CNcKJUACNFIQAP1jl2c8rz+fpsiFCwXWQpwvutqKq3p0lN6YaVxnDXLzUgZpByuS8MHSkUnh+BI9
0rn5CfCOVW/FmAVf7+RFmX6IXP3/0KA+9e8mnCQx6FCWYGruDxJy1d5+usCb3iyuZ4LrsN2lfdsJ
oC+3ogiKVx3jOUYycPnXxAX9RDuYQg2TA0gnhd2lnxYg97KqFXChG4xLfcR0Vj8qxaFmE30lpWAv
SaHlJkl6VQy8+kKD3rKlwYxWCxjIciKY7DjvEUMI2Z33AJxBYxO/7ZhsPFzcCtnXbHiqqfyTlC0W
3CpGMWcn2NBZUU/CEAbHjSIosJE5MlH0/NaWS+PgwhXOG1OH799uda/9rWF5qnnt/ReLW3Wa5d49
cCpbPwNX4UAfdlqrcxhE/aJEFJP6uc49R/SFS01IYRXk4Zu9sJk3k5zlUlmxW2OMjXoJ1d+ymmGw
r5kavnptcfqHGiKNymJPvMxPgrOx6coLvxfRpIbMwoHR4wMfKkmVrRZide899QX+Uo694rJHJRfF
nwa+YVoNZ/iJY3lsSMBC7aj2FIUzTOucOBmzaD6RUOXVhi95/toIH7Sb8JF3KjrLTOvLOo3KYB9G
Xgv9Z7uMJBNJ2ZDV5A4za09ezcDNBAW7lMb9RoSzSv2Ml3hI9PI3gcUUf2in2BMy9bI8osMDpneQ
QzozUOiJk6W9shsBGJdu9AmGGJc3JRMIaM8mzepGW+bTo2EAoD0POP92iItsEp3LVXv542alO6sS
+lg5qK+GrwGE7QKIgjKvbiBjqz1xALqZG8pFJQKF7pZ95CRiys8/eVWh4NRcBbHUMQwpcH+OyKAf
plWsu0u75ejokXbSr4vJtb0LFcomLw0TSc0aAGSBJDik9VJc6TPSu0QzfZXI5LS7JjgdlejF2Xbv
6kX54cws8XWCai9HH/8vTd7biFGjS/1qC/WDPDFEBgTuE7sNFgEValsz8cVcYhd7+EjemL1c8d9X
N9iTqNgmvNpE7x2uiRxitBPMTLGK3SgGwh10Fs+j2Mv1Kyh8yM/VKCgw3daXo1y2hf2gPaoZ7QmQ
BCyNyTRR6wit5W+FGLbIuORgMmQLbveEWuPitht2uBL+0n4soRHAL9ViIPA6/En1Dg9CVmRwyH9J
M6kzq0BpLBWi7LoM4MvDgVF243z0Xai9Uhb5xFJ9F8Iw9BRw8F9Rf940yG/rq8vYVSMITRTmRPfE
ZLXVyTYzm0J4k3eWF0BSNuKbZcT++g5OR/R1ffsT+gUcz1ISonPgn4i6D4kpq86SzQ2XaQU8Poqf
RlsplXpCjvvdnZ0JLdfHQN0AUv0xcz9j2sIjHPVE4HxqiOaQv10U7z2gnN9b4BNdi9/NcJrz/G8E
+sfL0psLTPxiqp5OY4A+pBUQDveBhELs3CqdVnCHYqNc4KUhqgEViHIdKvBv9jnHfCr1IXNjzoHh
9Vu+NACgSrwBcLpeUlRv9mEJJ41xISj8XqIw4gwaOLqpzZXY3TEGX8bYnnb+PChhGEyo/DVfhi7M
oCpquDVql7Rc55Bv6rf3LSEp+raM+fmQHgMkw6rE2QwKXVT0++tWeqw6MtlHrA4zkU37taFThJcG
L6TEHwFgZ9joOtAdRE+VkbmCsnLtlx8kCRiavHrfJyDfYhXC6/UlQdYhypFt4kl+neTgVBZbwK3i
dVS/YLiEus/WfnVl+kgfv6VaoDAJju9xZ6E5tP3TTI7+0svZMcX7rCtSClFBoKVHhSA4BH/0MNIG
6QcOUJZ5QsSI597lLrGuVQFpDrzCmdmJE0xvd7R6gdkL1YHDI1f2LXk7nVK/KvjLfWHFS8MQTY4b
4cNzL6LGcSZ0qvR4zc4W7GxpsOOR75+v20nct+vUPfVAcci/t8W3oh7qhO5rL/0svFiuIiQU9Qe7
HG7TMby2UCJY0UB7ujDibuwWEbcWFneewlVGgLf0Mkq6eDPagMFcrnjT0WjvH2vTk/jqHmKHVy2A
TymT8jUJTCrIuFv/HW6j0vVe1NB2gea6hLNL6r5N9gibHgfXAB4dR/0At23dEALuRWdHI5hAeVgi
8FYppF37POUfDvou2fKzYfQ1jmB76xgzEfzf8CRePokoJna4zr2m1y7cebCk1uWZnURUVJiXVmM9
qOUuI4eHgWRbqRHV75bWTwQUHqxPi4SaMKmbu5FcB6YdWSQEOsBkAPH+D+4Hm3kdJoIsQLC/DQAa
v88zQ1dK2wYzft24jEIl5ftuSEdriCdNayjr6YK1GfS0601X8Z4rNg5s/Wr2PFz2KXDuzgjeLw5D
pSr5JSADVeDt1HKvoQeSGmQmIiQ8TeIotUBc/meIXq0P+jfxYSr0T+cw/9C6WuH1+3zSltiocsxn
p9jRd00RhYUpqR3Oc5F2vfpJ+UHAbi+r+cV1aHYf17zDW1FFqIJ1mw0NebCW7icE91UcHKDLMZ84
vnlUmSUvj+ADiK62ml7O3dDT+Essr8HHvxver1+iZwblKb5ZKMOQe4/BVuYABT8NrgzLgbSEsGtR
AwLBC/G1px+yD6SqitKsffBhMTXoVoP3vw20RLeiijxM34m65sLgFL1so3w4tZkqAlwht2HLxz2e
lFBO567SKC2YaJCJNr4cUiDRZ0FS1yX8Lwy5gO+lISD5JKdR+qDuPEg/zKwY3/TT3qZotUxLcEBx
SdScCGInNo49yGRIWabothjSOCDLlAuMjNHtHwoHypic2lYA7bIgKpL+HACkKxoSUqQRaSS7dE8E
cnMjLvDqnJW73guDrPZmA2k4tceQirrq3ysON62HN0+yHI1emxmjTeyAgdJkvOeco006XLlxbZAd
MX8IJzTIiVppfh4w3ToHrpj3emewFsFRUmW9VN6bD1rZjEZV+dZneqCO7/NjrIHdxUBOvidMzcGn
jxtu+r5BMUK0L56vfxkx3oTmDPLSgPWmpakCI+0sDt+HwYPUCGFdMF8HrJUgwefDJ9da6uUtr4Ww
iql50Rui1UnOSZjcUsC3BQVuKHy8R8qNrmkyrYRLxBpTLmYjKaWst3yQp1BlN3hLDr29sBKxLvNr
tn7sZgKi3/c9MJRbWebxrhGlx4kXFJTWp9QjILS7OKdYxmHx+6KWGjmLn8ya2DZz+KYQhjR6XwQz
dyU7NiSGJJF4wccAxnjHg3+Ej1unsCMH/keLh5yDiKVQiqU037Rqk/Apkqv7/qmVR1+vrg5M6naM
QMmfTI9qArbG4wBPZrObdKKH5bTsDAPOUR0sAZ43Q+vQaPrZpLW3+HXmTg4HHnfgRGq0f08FoS9B
qnCwk0UcgUkNJ7JWcd6DhlZe0CA2m5YxfQXlNeGzYBfW+X/tySS2PnE81P3x/v0q0DEafhbauDhg
bodTwiztpVAVnIgfH87kixa76sBC94It1GUA19dRkAsyWl2EzmvIzJyM+FR+AYZlqdlXS2s9dkpf
m1TBmYrCwr4LtihKmFMvltx91Zi4EGQUftW/kfresnmgUCeWQqRVYNO0pba1iX6aCFEWnZ+oH2Hl
HqtrkwdFxckUxxHFo4Lm1WlnFt1C8/9DWE6V+AThvih71t3R54br7daqDuPQufIqICHWfCvua7iy
UdRq7RbJtRaayiD9W6l3Cf6WxPPmf1vGo3uymucb4jryV++MjQtLrFu7ulBlxHfFrXBFG26WpJ5n
so1Os5L+RkuX5LfrExfuYySaGc24wtHAPsNvh4BNtXwawJFocYZAi5mmNSDuhopl8SCzwIsPKuTt
rwrZAbah7fS8YClMRNFrCdfZ62vQP2FFGJ2nudABNPsWy/2ytQXp/uj1etBs//bOquWwGya0DYZq
qn+Wj6mlDgm1onrczfrKhV4SMRc7+kg+IqfNDFV1F8FV/dyO0deZCPl6UMBphL2+aIl7p3Pj3mZs
QS76rJCPJ+Y/pLLwlUglH6oCNLHUWgP+ZgaP/FyL55nVEjqzz1RKbWk5us6jxxA14TF/y2MH3O3r
F84uM4IJeeU0m3BPv5Fkcivjmz0i4WB7oJM9QMiHCAEePvq3acRAKrltINFseUlhhTImhlFmd7q9
IFiECAyiGgypGOYiZOLo/t4tf3Egmx4SCFU+c2xq66jwMeFyz+EFE7/FJlAIjTUsp398rQQDsgjl
00AkvF2+ilQIf1sgD3GV1CfozKW0avQxTnFUBJgMOGTnrlnHmOwV6tJsLwOfJrJ7SZrjwRU7Kt2L
1ggeLsiF9z0oXrz5DXz5L3oNAWuoMLOR5JY9T9D8IeDg+jSZbIPredxmazzA2vx0ELnovMPfLLm/
6m4RPf7pQMat1ZxtIFUJ6HBYVr5Fp8rjD1xAbWsMED15opgLHdj+LTawmgHws+15E5BLBreruEXD
IkbIkbgSh1F0m9/XxGDeTOZ0wd2Pp/RpsS7BLKU2p58XPYbIuB+GT4xz+WjKTc0tc1f6gjnlgGKz
+80dWYpn2QPGCE/DyHz4GYKUlar6PZmHSZNWee0QPL9z2vH9Kvx/6kcpkBrhKG98PfNphEKbRItX
oqDXMJWLksCUAHb1PjyNx6s2K46Iu1EmddUvJxuMQvVTglor3jcZrggbp/xLrgAQe/yA7qAcsNS1
eIllwu+K1Q3PbhfLQ+vRQEbOVfv39hX2Vb+Jf3wJy5SKZrqz+ANCs94wm0y+6evD+M8HwbL3gEBo
YfoiDjlV6OAx1EHG0rydDs8+TMgsSUDfdYQ5UGmfnu3XKfzHuKaX4wvR6HP6c8mprOrdcP/Z9i2V
nnbTsyUVSeeHAMp8SVkWMTG5NKCW8jdGuo0ceJjRn5mKjubTxJibm3Y5tLjX8Amusfz+TJLzTDSi
vO3+D8kNSaSe6dF74APXxQw8E8rymlF9gorKGSHf6185rK+E3G3zeV0BYlxfCQEfq47oxClS6Xrq
D1fK1QYK+/KbNm5q5EeQLO7BjWom4MTJGsakm54ZDAgz7zjTNdZpFApJedbAseHmVsoD7M8rZzco
04lbW95k/wd1K1bz6CUYcbBLRYyywmbzly1EdgG+K3u9RCjes4jElrLL7jjyZJjpc2FzHIWIM6sU
8KbpQlVb0XQRh+qvzoI8W/5XRK5AE25flmhn/1WXDs9v7TWCmRrL6ezt2yFPqXofSWtyTXy1t0OO
B6Pyf1Ce54vFdN4153QrYwzklHUnAATmCP0brjD40yK/8imaCeKkMDwX+4vM86dfox7EO3ZH/rbC
xe3uXAlEdgqOBLkaIntcugYlYgii04bIw+bWvKeyputPFr8yySeZrth/8BX4UWcWjenWgmThPyZA
L/U9XMkNU6b04HBXRiYV0BVBFFYydzikpcFSTKHZy5pnuk+VvDCTvi6j6CLvFHmxYmyPGIrptQZ9
sFLBrBoCLNG0sPfoOY9v3PLfwKz3GQHg7WxTxAlqjViENNhy3cT5UDvAW4+F7ZAR0MglJrVDzdTG
OpNBBEQgNiRhANuArqdqgjR7GLY+6cKZkAMrvoG35LS2IelfszOrOV0oIxFuM3yT0WRk3unC2+Q4
YQO/6wHfhhQjlDh2UzHb1CU2DKxqh2BfKxCDWCASskfbKyLW5w8Rp9V8PaJFeej4tiSAbEgSbmYe
TnJp+9sicg5HgJGR4iQI4q+SKqKPPwBZ32YavWJby7w782uE1WxqiphZmgHiLQfsUVhfAewMcRoG
G8P6tXT0KkCkd2jXa+YaZs0VP/a3lvrsxkCZpq5nep6LOzzEf1PWkNneFlG96HoU6hJFnongKzlW
Uud2btec5xNtnzkSQNn67oHZd67YxlP8dXOKK0R2ApD/MxXmnWdrkGwxNKI1BGX7Okq/hYbNaE6P
oq8UsgWcLB/FpQhSC+Wq7FVVodcv3RsJxV2BGmghX7FKuNFUsLM4GC7cmL+F/xo/iL/+0p0GAIdT
dCgOG8r8NFCz9tAdWG7fHPAK8tVbbzSLU3+l70f/xQeepPVoieCCvpdaF5leqyCGHsIqhEckcMrq
ji4eh/Xv5KO8uEWiFGL3lvetcIawz8FnecHljqt5ZlNC5BNWZMuc0JhICRjgVqg6kX9eyjef6A04
9JLUSKBdVrCMY8JzXmcjCHXkO0UB3v9et7mf3ckQNro7q/4sZYEjBHAWRILFwjQt02mfOshiSFVG
vTObio5aPpojjvLu+wz5TORocki0dYf2HyO4RhWua6k9+lV6ULoQBjAx8xFbMbHaHVSDjHfSYpGa
UXGxh2runmVcR24CYiAzZuaHsmQQhomC9CLdNvySfnLHXOPtWuBokFLVKPJDdTqghU42VW+ZqpQv
f8CoSCz9gg9LiXb96/Gn2yuGkrjDDsh0+997/E3BCoaZbfzh2ONvi8Jbd/RWkYMTf5J24C/TKwkG
Am4GrHCcx7YB82i25LpRpDOSa00PV2Y0muZoTo7oAJ0ewFOyOCb0eqARAAgL22epOX/yLm+9CK9o
poIyJKI/9qhElIgLmc+rwcvWvApzbYMQiTsVTuhruyagHEuXz8OCUUMwwbOY6FtzlRzIp0CrLnpN
oLWi82cqf+rP2/F5D0umWdLjyjPq8I2g67D2liH0BhO5PqLFpPqyua6/kOgLsxv2cA1+ExlciRVG
HMETQjVUhJS06elWyu2hsirzJKG/tJWTr2wFM638naBhjgiCYzEkVgHvYddADfa0LxI6ZvxwcW38
9E0cNEzkIX2CxWGeVqRnB7i9CKgH46+a71X7ya1H0el6oc+FmGQoLFVqc9TdE6Pl+YLpyzZA2dWo
bpT7oc3YbLTPs/s70Gmdw8Whc86G6yoBjfBFEy28w8+4jYQC4d+2esAVAz5pICQDccQcQ19iKQ0S
k4oevVPKJgc2xLSeDOEYoT8BWYOQ0Oseuzmw9knRne5mgl/bmMV3jKUHAzOj9ATJ7uY7GBn3NJhU
s3rE9XChNH7JkKPwNcbDVs/ozgnmvMz4VT1f3ooFdWgZa1igcqP6COhp/VgoleZnNjrVQTl5fNUF
MG1ANCvqyLWkkD+MkFCbRjzGWG2KNYMLO63AXU52Wg1i+TeLCX+ocmRpK3ebbQ3mA+UFfkbJFV8C
6/4tSgJfbaDodWlDr/0NSV2IRttCUSbTFhVmc4QaO5g315oM2bCB7nhhrcRUf4wToPEMfwnUHMPX
E9ZaQ+3tQZbz4FCv4fGWQ6PIbNXelf3XV1hp8eXEmz3uX5YAoaLURLohdp+S//nlRxCH2nebVndN
Mic4nTThGn8GIdAOzwPjijRDwlnS44b/QCwQ0DpZtI4ZZbnhxbB8ejC+qu+eAp+bW5ToVWKtTMN9
F/7CXKtVam/L1w/jb+n94MKxSiFCnBgg1+LWc5k+gsg3GwXXPxdY7gRJ8SJfiPFGvy6VB51AFQLP
Aj8pIzZG1UByegH1RbXkzndLayFLRB1ygkgv4uHOZVE5RqrrsUlt06urZyjTM39a598DGh9hdaCU
PFEmhmUQnJ+AzeFB8PIOV2TG+v2slrFTzEvhbKJb4fmRCD6FRJm7FWkSl0UsB9FTtL+WMQdST9Ho
SGFkgqsaNf9bnFQ8lWUnt8aIPaxn/pGFOFFvd5VBgoFXEct+FDxUDDPuMGGWdSWgELI2gWgesrvS
MBjuaF+7PYAx2uWV8uDX7tz+/iWzYTFXI0Y7iHG+kIkvrfrLySp0Kbs4FcBUIjyFzj5nl4rmYhkO
Z1tuRPPLTdvD4KoBSA1Pcp1XEijVXNaEfRS/WgCG3QUbCuDgcdwTthkgAJ6vmuTXbQheg+G22jg7
rjgip/BlFrkKU8/JXy+HKVGrYAB3NFFYCZXSGMoJfizYOpaCmpOrUWFM0OI8x9Wdz2qpIiCsLo/A
fm/VYoUISdPxmkRrFk31o+UXprgCB6C+SbftJPwbZ7jVOX7bJLGrXnJVs3g7mVauyzN+zT7L1LzW
hapb1ybN2HNjil8XINuv3kFIsPhvzk414DoXe2ckZoYWx7m/0112n3SjvokX1Q+aHMX2F9NdcOZa
x4PRBbpWW9CkDKQWjDHrpgXjKzF2IloB3R6/ZzITtHW9/EehSK2po+xooGkfxABlNRcDffBe8QIs
k29UVXQancTUFdqGce7BqVIZXm0GH+87BodYILJ8d0WsoDpfGKyffceb5HKMToyMlCLYBw1QsZ0O
a3IY7naxbcnHNbMMYNOcyFcurs2Fe7UtUY6GTsoQxdamT0eokn3+CpgPr/Es6KMfyx8yrQ3gPFCN
Ykc99LIda+NrYHNMTQ2XUMnt3dsOAKxLImJ87SC3mehg3LKLKRxnpZFefPMoIsesg8u6OmSQ56qm
ANu62j10JKmejjFStXZI9TxsMALt1F8+SIzrOPUPXR7I1bNgTWcm2Y6xHjuzJxl3Ed9ugCiTCiai
6CYmPUir+kqG9haOL492NoLdu0EsBbf5OMOmuoHtbnAHv5KRoicVCLtE8kuPm/zDI7Qn6BZTyW/F
ZRLqzTqKmab16JUvpxrkfJzlWh2uWn/xBrHuVVlRPb4i5I7YHOBXxaWVu9nKEq40/LWziZ+qGBqv
j9TBamGlgxmK9TTfi0gC0ae6EaklygwNcZ04xtiRxQrzWW5xK30cwvjKZ1Yd9i72QFikQQPE+6Ua
6grnJIV8QN/6OH7EBYlEcv7GArt/1q26N8zoX8qaa3DXter32RK6pX6ox+GyrY78kNrMzGQLNqyy
nbxGRN8sWvbW8DjV4ymYkQBvuoyXnrUhHgFrDptejiuG8DJf9SpSTm574b+iaGuGRe7t2SGTAtyj
BaOaF2bM2QfRxxzofZIxuzQREPwVFb/WaTYKFDkC47nPrPq3lA6w6izDOROWPOI3rDwA9Z6OlFK1
J5Ev7wcADm+B4M9EeeIm44RUpZOPItWR0bJqy0U+Es9lgt0Alb3NO2AmiXigoKLDoSIHtRqqIedT
Q3kFq3UWw14Z8JByUGdMt0PxkV+rcegOA0GMaJJScD0BPQMEsY8aJiqOusdxQqb0dpOPCuLXL8zt
qy0Pq5MjZGFQaIFRg3uw4thKpBmXKObAgGHG29RbHrvXtqOqzTqZKiggyOdqYucyddjde/plV7V5
teYarWOocene+v5LZ/CcxCBbtgCMDtIDULz3U102n5Rgp/8Fy9edRWZutWBkWIXSX405WOGSTG0L
h5yxGl0Ou54QN5bD6J7ALYHArNkkbPQDZD15n/uN2f7vR9lutOACSTTNmhTdH3dqTuM/wVvpI6d0
jmRDLhTELM8MWuLJVZW7QDJCs2Gr2sl1tK8HRKCo95wsFVV7fgtEuUwXOjYh4jqOuOCqmbhC1SzC
XwLqr4woPtoF4ROCLpUrqAcWFCjy+nTO3oJZgL3ZLpmeBGOwyJruROFTTiH6kpDH0X9V0ve5y1KY
TBdzKzTciu8lzFkv4ebcIxyJSce8G2UZlq4inyWrdB5ktegk2/pd3x/Sis+oGHoJkKl7r+28CjHj
ermzbDhQ9lu/ocST8d+TDkj9F+txQ7+gJYPWkLQoCRaIEhZJg7TaFFWUX0+lJmtXyRXg/SUniYah
L6POAC5Qzk8fm8M3FfVgmBsaWcF5UfLjMwWmWY+PnLpqdBNH9fJi1kfgxzXPc/fHQhldVGmYJxcq
LZc5/q0bWKvt6E2ooKC/UchGRKmJZznDR0yfIzcZaPTumFd9CzLN83iOmLfzFjjKA3HhBuR4CBkI
oSdGFc5RTo0lqlCo4myIRkaP7Ug9UldPSaVZiHtMr4IrQrm4LO7cbPJ5iu7otAM4Y+7YDNqYeXll
s7smyvkcC18wMPPFCbGPHBxbXV2IVlBUOxGae4GehD93X8gEw4EujlQsZibNAAkEXgIGdKdM+FcU
0nGWf2BpMgX3at8jPlD42xIby2MeUcnHRvLK+DHETkcTIUyXWovfY8cOOpTcTPB5RclPp+iw7wxV
psQS78knzybTRTObYexn9g5E86Sesya3nRM3y1utOO44kpWplO36NU3ljTo3T0LiP/YDgmKWZnHx
1/G5P71bncwKh/5/qhw1g0z31drrONt+JqskNLwMe13XUFEc2WE09GneBOPqFD+lE+tYfzwvtwYm
Ue+lNqfzQKqRsB+8QLW5CiUEos1ebSkb/AfqHu54boywck1ERkANa4csoPQLGN6BcwUWPaAf0qbK
+3b0VORSFI7aZp8uJlPYs84SDDRLf6PvZnW4VRXWyZQBUb9GlxPdHBitgLDMrOw4R7EFbm479b3C
Oo+hUHsfqclZ0ffnhsE2ejw0zN5FtA6hZpKtaKsPnZwxGub3B800/ZyhsrLHhAUNGaKPF1LhRDO7
pOTc7M5ErAr7q+d6CkJ9sF693Ehqd4Yp0OaU2zhT3TKlslmjMZCyJC0NNMNQymevq60zRa+wgOFx
SevHyNE+s31H+LqzFC6CFeesq/EspJwV69fzpOFE0HDCGzVMMiHMdK6rpLdbLLlbDD2O+KbWYfS5
HeFI7+ikBtzjF5p8Lv/SAfoWXxFLkAtDwtXq/EctFb3Cow1ab4HEXCO6R+f4OaTrr0/L/puroG1T
AK1JqFjTZcrMutxP7T/blwXoELDKWTxhCUeKkZziMHUFLeGmzElQmjxYY4+sbbQXFWQAktPfC5L4
ILIymq1mcJzyhDuaLghaol22gWxhiRgyYC7VLFR8gap3JXYQMWiIXUKkhph1LZxJpzHRL8i1FaQ2
9RzX/MA0ktA/OOkVuAT9xyopuexrjaHTyBx/4+7JL8F//ZhPY8Tud9kKjAGMiZ0NNZ+tSZuC3Khc
xamdSUW5zftxFNr8PSIGGZxO/6h8U+JNY4KLtj+1ISQz3bFxE/QumV0rIJzGtJMq4z52hAH0h8io
wY5IY6Cw6qCpk5j4CnkMcwmbxA2LIJTGPybHS562bKlyIgRie+e2OO40uG2KJrSQXfetPNxQZNKH
JEWISYgqmyJeH7uaCVUaW6DguO5g+jUGnfzROYvrAN5apkoU/6j8Q/RopK5XSkexLiU5DPg86vvY
NtQp91uaEVeodBM/NCter6c3rWxr7V5MbVlOLUF847+1/bNlGvNJtfFminrcpWoms6DcqrkO7tt6
nkWcCtTXPp6cJJyWbke/nXMQ95QWO+C/od1gUjqHRfg8nqDK+x0CFr6u1aRD2GUp1WLAY8xMdXnG
cyVNRZAoPW+BLtDuFkTHdtMzlm4B3YJH1/lCuIDQe4/jqdo4zlePhD/4G8S91CBxeXF2hDTH5NWD
o8/JD/htH+B25OVm5P08EU3dGw3KZlbpvKYBvPR40Ff/BTuOrZ2/C4GwMVtSoWDYLyU+kMS4xPgD
D8vYUzDsLJxURllqj/q3jAY5ZPyudlNzp52TaBPsrrlv5HfAbffoEJpyCRRZ78S34/sy/3dWWH36
5TVoGrSAhLRl5f1Zz4F55YvyUgOSBaEG64/NbJoaE9iQNW/HatFhbcpbVpaDi8QdSZCbyJK7Snl7
C2e4cMaKmkMLNYGoIdDTkShLKIMvNXwJJSZ8KMyszrm4kRZrgihw+jpBl7MYxu7kQZ9ZT3k9K9is
pA4JjbfVvmekP8skFWnmzu/DVk5FBHlOUGVALSEk9TRlnP+szrOtIhvfq0NALEeK7mq29CZmov6U
lSZCMbjmZLi43xB4QhovOhEEp2pBgOF2LcGzR0fBhvdzq3iOoxnTy5axYkd49fNjPBV71IvpYplm
B3BqsBA07hUCOKJmu7K3m5JcYIY1hKnB4Zzd4/nLI9KsGHg2Tr7SLtDi5QYEt9slqRJgOBOJbkOF
yoXAeaZ1K466/M+eQszcXKPWJjYnT32NBEgOWousYW2+RA0jP+d+rov/9lzah85GjHBqpk+oT2Jx
V3PrgkATBGIXrDlD7GCggLIOvvSpmQVfCs3DLMh85mDx92ZIh9PCdQhRhjpfvwv5EeqxTjxCoQW2
J1U8LiV80kB0fJbjJJSN8HPtk8sTqL6Dwwj5tMsDsE4tFaXY+8rQ0wWuMOdvdag2svubEAKPEEvy
YZ/9BEkWx04mHkTtjkScAubUyVmRZ+FrattQ+zhTcLILcm1RbhPvI0PyndFXedd9REQ9YwCyZnfY
C/J2iUR8lu5wHE6N9WjQc8nmR69vskldZsPdVt/NVt5pqvH4dQX3uGur0G/WVwiVstwyv6QXul1q
dJZr2mFsbNkJtwDRsvlxJ86edkoieqroXRMv0T/zHGRxoupRsKRXzVWYKiTYEsfV0y5J5geZW3Wh
ZhZ1Fs0yaydFGbCY+VITl66hdJhH5bTZtjXGY0bJEZuykCBvdgaV790u1EyCUM0RNBbFj7fZ+wka
QnntZuU1mTirsgS9XwyiDYmliW97hgZNOY70yyJBwW44RNVPjUCq4Ws2kPKPdVWo80bABrBaQUgp
U9ytRZXXOoUq5IMv+rfn3HhxwQSCjJi+3tVPHZ6wQafS0JWGLMoQSDy9VsNKhtGDeHY42iYYDZ/F
CnvulcvZMiI0GzV2wn8bqGd5eGMwrqC5Mpsrf3Wtk0A9fe1u/kWP1NAqEk/69c/rPjsvY3/S9F6v
m2KC+WEE830FJ186DHMP8npYsaZrnS59xOwy0e0PaoKEs7/PdcwQ53mFgNr0QIeNGeiajGBMW1b9
fXlR0Enq3a1QzNu8/ZidnfrqB50shquieefQVpxfSxb4QIXbmxAQS8gnaUdrOey2t7l3r1Cm8lrJ
KzJ6CuVzbM/byF1KKc+qeVyrOBn1UymtDUg/WrUVBfUuytNAmqgdZVcGCUjMf7xFBEEJxYKZTY/b
QfogNXrENxqHxXJF6P5eEFz3OeV/jCL079Q2yqPASP4x+9DDZyN1PR7r9hT+jlhshaW1BhYbACIC
9pr/SbSOHMtBD58h/InurP7r9EOh5outHgTCBghZEdHeBuC20XOKall4FNOvp9EiQfdkAdl4Ixa0
Z8WcAKLW5OU9UeP6abgy301qgVLibgopvwFlezSLGqfWghw34XbFpgyJZZ4EzXZBwS8Pqbc4WGfC
hkooq72db8Wrfa4GP4n2dapjvqf7HDd8ZihPKnvJELWf3WUzMLW1beiKCw6ZgnmMVETCCBFHjYw2
cDxg56KwJiKkKLFDIaBIrcHJeK4Xh052Xr9ITNaMBm5gQM7LUZnlcx1n2t+bJMqfVFW0TURu2Huu
WTER7+HZaFEFw5gYn0mtU5oNJBgJYi5onNhQa4dr/wpeKh1efKkxn094V5rFMMrN9G2LBitcttX6
YRO0mpI+Zbt6B1ObvY344xcUM+7eiG3KjIhguKfo9B0gIjG5Idvjt8lbRpjNfnwQY3yeRtRs9Z+W
pwhFF37I1v71hLzvJ7rTOlAripZCMChI4x+OlQAIfg3OnrE3X70uuk/BOfqIbFaSwQsNIgEEg1MF
TyUiVdc+U2cjM4viWpOCYw1ORrhE0nfo8GDr0F3miwoNOvF0hQ838hrmnsdxADfoaF5ZG/sOQnxH
LmC3lw+h/8vcJihKH3txshLhRVT5bJpmIG+GW2zI/X+UbfEk1svkP4kXUmPNWaliO3RsTx0ET22x
W4DiWwD92b3USIeB2K5tyHoxPqWHDcqpCUcz+4On6ldhVDPPyu4k0yHA5SQdGsoFAaiOhOKh9Puj
XyRaN5MM3OWIWvpIaYee7BxY3PYIjq82btr+dskRnj1kcAiokeqeRf5hZgaW/oWe67OOJ2lrO4v/
oQzlSt/bb1gTaXhtxzgg/7sImGsDmNDU/zvLHzUMTqjZvnCwrx3EOxQVl2AayPAHfHP/lVQKGzSZ
Z+rjlwKIUZWAK2+Sib5CXjgQwbjhvXbO8B4uLJcCAMLDavZCp4sks0BlK1F64zISwD3rPmMSLp5N
Q5pUfu+Hj77cgzcn2LrCnMmUMeJ/JFHsd0dVSjbFX2rf40XAGx6R+xuLDk3Y7Hx0xxiZuA8Gda9p
NdBSLDM9pq6Ht2i1GjS1ElPNUdx6d88B4F1FyJaYbyGu6hbDhM1r5DA+kWFfO96t6sDJIyepZteR
cozvZM1Htk6mYnjKlpxnEVSjIk2f696Q4T4u5XkG5nrr7MgLEgRPnXjxEMWEq3A/ekf5GIKVuqz7
9YeAs4V/METHJUQ59IlOtTjgis4gvokC+jprt4lb1IZs7PYhN5D2xwfytTjw4c+CSsEoRc7+iikj
hmJN24Srhp6W4FpHaafOGZUmgVLaZ6iJCrF3uNOsaDZ9cW229MeZLYn/RPTQoAvLdezWMH0IzZFu
1GQPI86Wks6pViDc6CEq3m9pKxiG9pMpErRWfc4yAxDX8uSf3KdRD/wuHdb9CPRIUrLpgFh+a8h7
A4ITTt65yO70kOr1xmVv2S+QsPzBWO5TuHGwK7BUnvpXl3gElx875VWc6JJGX3JYmtB/S6CRJLsk
XbFy92Tu2rqZPQDm1NJbyVEedwv0ZJK5lbxBwlYPEqkRXTw4SRBxPkPxTkq7qJE0j5idAR4o/n20
0GIwAQ55ch2s0z7TI1nn9ZWJngrSs66ndhGCvpNy/C8xhIgjzx7/KWO8aC4jgiDpIj+ghOi7QH7e
cmNs/Ilm7LojeY7OSipLbDQ5pdy7de9QIPeG3rKdEJejwuuxiyFfGmY8ovv3C1NYacBGxwI9ewIY
/3idINMLxtO0qs6FWP/EIO+qYIZ7RZYsa+QvTKFdSG88ThA3Ftx0JeUyrSopXDx4D8cbc3tBu8Ns
7ws10nSsRvnH0z+k00MrG6JZzY8jONsBs4dEDqa9nGhJ0ouDF6hlvxUp+XiEXGfm/V/3BXeEJ3Op
0denW90pDx7KCQTcLNLefN+mUkgRRVt8G68cbDx8kOgi4uxSuHl052xLjxJRan00bywVpZTZu+/v
l6IZdbT+fY4oHsJLyoFFyVuRm+PIJpfmmMM4uWH2vwDxYaBozc86Mclf6pgiusV2q+sVkgsnH28a
hKUfofhM/24D844rK8vi+/8dY9R2ozCQujgG7oqSC74Sw0bC7O+Uc/BA2rUQwXZzqLEONry/3iLa
ztU3lm9hBJDI3teFztgV+d5OkLKvefSGPfSvDBZDtJgagBkWYRXr7RmGxHJ+lxSwpqTgW2/lJwPw
gdO8i1bDbx3+qztI1k+1OE2K16Twk0hUHxeTDotgOiO+uyYPOvaax+EdWFQ98zaoyvMs6wMABfgh
pFFEE3wS0xX1RHicgyeuJNRYnSkvQfNyYOd/AUfpWbuxwC2Qo3gbjEoYGM97rQZTrUobRzEub5i1
jqJHC4y7upaPwx4s9oGNlY+eo/4fG1aXyotsKrqtqNRlrd6nTUm5meekG3LlKMWBcT+SqF1y5iiV
LQf/5+Y3/VWOhl6Fy3PE4TgAeIWapy9Axp7p9UAu/8cvmA6A535ux+e3uFsfqt96wvWw1mL/55az
06BGAYEqxFXEJ6TWmk8wzYWfE15ZLBI1JOLpyYJL1GtbtHD0LizcIA1UzMTZ2MlvlH6jC/pqlyrg
xUo3gaJl3G+XpXzJCerFPaYPn+KEJF/o4j/VKuYpuhwZ2j38nMpAgDMHr/8o0jKaH/wAw3qyPRSt
eSIjmV1NEW74/eNf+KEOl6vJKEXjcgmOEcro+iFcCzndLTptpERcnUpCq87PxY8m5NrxGJXry5Yg
9/ni7iTi8ZT9UUaBuvXwrWJAs1xfOw4PvO56dFpDuprFmWoa+GpD6FkpepzNN9HQIgmMTGkK7oiI
VolSN1CgVtT4v3+3WE03UM0+oyDKAX2i9euEosFYa3h1PXQbu9d8M6R+PK2Kf9NfnpSnCWyf+41Z
gYhjXTR14F6F5cxYMP+frWQa5fFzJwyuZsy5dVOSLJ9fVJQnXjEYYGJvFrlrnV4j9PPx6TeHPrPQ
KpYX2cgDjjeBi9Z0GokCzgFygOPC8lrpy261T+ORLJIxn48gTQvCFVlgHuH2blwRTdqfUPqQDrYv
Ie4oKrVWD2UlCisycJ4nwoLxvlamAC5KqTiRiLD9ug4slCuy/STog1nqTW5InPh5GwP96aUbmOHt
8XoNHuIMnJ3sORvtzLYMPV93mfBu+gUZfNXffl4XxdYeETFV2rEUF3QqBsQkJuK58F5kAmb46FfU
Va0SgcxYqIwlOhBuWnG3rKA6Z/iE2tOeBZkMX4xL7ihZ4trOlnsleiL+avj2Ch8miupgm5Mh7LtO
3crUxvMwmvAtvPImgEytwufMVYpQuGgK9n+gGJR1j2bLB3sebtzfSpgmtFT69IowK0YXMNb44cPA
OKAjyfnq4DhMTfJBb5rLShBAZmIe1YDNBc9UKdefJ90Y4eBfPRcgNVVL6C7gfttsuPsb6b2RoU0X
/2neoeJUiSoMoWlxd2ych3Yhp5r0mTpZ4mgiy7+0fIZ2eYJ+rwAV4JRPgg5eliSiFmEOXfh/JTKM
UKRJtkEeNYE3oVMgdNDUme0jqx7hJkryIGlRvwbzzRczF5bGzn2VjLjsb2oGZgGwGFljx/1kqlbw
T3eg3I1z5RzzJ4ewGa3mtQsxGm8hDH8KSBPHCds3/WvY39QcLqNi3Xczpnx7R4gaONM2xnogqrvx
ev5D4NWqaSKVInKDTjK0rtjN1EAOR4XMWiRu7vGlfdLKjmyO53oT+04nrYdDxmVftT37CjWi0Spv
8p+Ic/lGOuq6O+66lhloOPlKoPLe8txCkGTDEJlmnSfkHAars8YeSrz6XmRwTcp7Pg323Bz6tm1g
XGy7OwO5p8g/V+m8qCeaVwTamjqffbUS83kQiCc51bPUXHZMjjtG9bWiknOf5S9l4u7GCI+XmMLW
0w3Z2zo5TsLMGedylmMT+tGyhb9YuyxQLzA+3RQuDLyZpDS8Qm55AsIcMBp8Q0lZrWvmiKuKEo5s
DOsSlkEMpty/GdRD8kKGxR5leZtDUrvamtqF3vxjjtxx24B8ZqhPwbqB3tBGcParyjAJjaJ7OOpZ
c/9AlcoiDc8wgu1XVR05Mt1NU3J/w7D29t8rS98NeDJMWwQl1TDWv7iWon5SLOs5baW33Bjd8PhO
FoYDDdk1u2jCX08S/MCmvHoHzeNV1DWe5liGpTkRqeioM5BnMERRXFLRGdZmk+uZo7QrfrM1+fJN
M39qLLQiQBg0VJbCuFhhPPU+O9171sthKxGRaRIfNWAq3hBtWdaMqdoN66NLGIijluuAwCLKtNnE
vo2v/uhtnFkFi0q1ew5rTe+48L5/8T3MtVkEKk19Vv1nlFXaC0m8qrQcx1TxzzORugG7bWfaETGK
UcT1P/3LwRvoQPYuRQ+jTkD9EICddZe3R7nZRKVp/hVI/OLstQNfzMGC5OikSqN9b/oZe1TxCl6Y
lXyCsLlAUKAAmTn8NxfSqCk5R3iynSwWYwdSKOnmCGeObDxcunTn33NM3fbjy+Ba5VGzLUJkDuC0
D9Kcpy6tsEcrBO+So9B6KVAUnOD2ntvn35mDYLHE+4O6VsyCij1j+XJOdQ0dK9EpB2gUuc+Qnkl5
e2mJ5Gy5gFub/2VWEgOiwA+UwB+jZjlQIyYpcO/caIKjDtM8fDFCoA49gk3Rur5oN798trL2twWN
xIzKZOQv0bVEclLAkZBQSmlC/XRdRdSlRaJ+z45Uh6Lg9n3IazLAlumykyS/oq20yUrK4dmPeRhX
W358Lch9LoI65BoEXXGH955X2A+bYDgdhI9dEWBuL96GZuqZxAs0+xA3hsZIIMKpAcDaBdBK+VHM
4Y7T4PPO/1TESmnIJv5TRmUqnTZJwCn64xcTYpjxto6NjEiSuTtV2vv01ZC0+wbcWHpUhK+G8Elg
C/gxpRQqip2yMneoDGrf5UIl9721vhknaBAgRksZ3gcGbDHUIsmJP3SwGUzefJ41cPvW6l4iYEc9
eQc3+QjcZqDOPsI7l81onSRCGkChUW2NExNPDtkoOP+p7W8LBehnoTxC5aSl6Cz5M02KNzeLer4k
Ysx6XhtIjTvESbQsbTh8Pd0Ods+cWXNdUTN8YNrLzdZm+e4bAW30aXKRzLe5/pw569dbQBA620AM
eP/QkoJ61eq9LfOh6n6fQcGxnJAkpq8mth2qv+V3Imi1fWJUgXVkHYFhYW64c9kP9LkohwCO14oH
tU0B0Xrvm0tFI8X4aKQMF3I8jVfpSIxrvMMxP7KvZcoqL3M1o+OmBAPkETq/MJfonGtRKVAudvTQ
Lhcn/Fpmx9nlC1amTQtUxhmoZ8xtNxzZcS1N8h73Xmwi3X58YlQ2N1wKj7R7IsNOMeMjf46JPx3w
HPjKKMhQvepH3+8G18trqYuUvCVdC+YCAEp85NYMCHZsoZFsdc1UxXsG0UO4u225lok+vf9esmoK
CMsb/tqO7BsfIsOHue93b4gRz/bVP6sT7+QrXzcyx4YQtu7ZKAtwDs0YqYpf8n0Vrwyid1xm6Ggj
pUowm9W3VI/mzwRgacwmTRPzwRBJHVQ4E1nzeFjV3T+1uy7Mb1bHYBfmmwAep1YppHs8H+XFtJ76
Kq7oUsXQ4ui0iutla+4FI4bxi/UcfMucaLk49zR2RsnL9NMMuMRMtgegbzr41BTOjyUbxqhfbUbw
O35VSyeppZ53s79JJDSvgO3v8IPu4hoF7IniIQbXiP7/1z5mZvUxSb00UyqgeejHZcSirZU9w/9b
nwcW0I329dIzmESrAQcZ5k5bOTSGz2Mts7bfjmkk0zn+LouKSOQKgatLUGdBbK5x9hdW0dWAz3dG
Y9rPmv09fcAoXfSW6OtgOmzg+Qqx5GVSpTy6GSlw9Gk27d62ExqmFslm4G6HGOoymUEy0d71AXN5
LkrwrlS/8zlJSVNkcUwXyIwP9yq/tJ72lnRjzHm09snMgts9lCN7IR3rxA6XXNmCQQQN63fekWXA
lJug24wHral5RTdxBlGk1AhLWZ9PQHFrcOntt6UYRJxBaDftTSxkfl9UeUaPGZv6tKEzEl+AIlpC
SFuK0ArhzXXF12KAp7RPI/+BdNeBlFoFVOPfJ8ejf9lQ0B/nRt+1PKgVBQBygt0PrBirUT87kgzX
zmLNfDddSOvIL9cEQ5NZgvjapf/MpBr3pxfMt783Zn8DtS0BkJD+MzBGpZVpvU/Ny8XihYFQDGdV
LihL8WPRIOXghrp4IoXf/uQtqiVC7t6tBHoZ2+ebim6tZFGbBBd/nDeA6c+hA28DvSmCiIgcpKrT
7h8rOhEqThBrSVvpxLg9FV6Je3SutU7s2QEbOsTOsxk/T/77Ag2mxKp9j+3ViYfwGJApSXYfFaiR
L75pfpEKdfvfSUPxJWL8isGf6RZhFnCPi7w2NMOhOrwumD3XqIUwDn7fDza6kFRY3Dae/wrV1x4q
jY6erQkhnUro5e4aTpetxoFsDQAxUCIHoQ+dmt+GZsELMeAF5Fpt2ihYDSdy6Vc7sHP/O4wZuKIH
sw9Ua3PB+sPVy3RWzoL4x4cp1z01F8iLyxFyegw7nXFuTlSDxnfdSUPg0wXUzdeHjrRHHToxFuYy
bBBj1iqKzZAynpoHEs7/LX5LoD0dod35htMVQuNqOajfV8QdulydG+2jd/GtLFkGp89K2NdD0N1T
7bLO4lxKdQYVHbdM/x5PlQt57dv402Ha3YKGElDPg/ulFhSD/+2N+0ESGtV1GNg/Zwooohu/cFHa
UuQOzZD8ExecbTRe44zjliFleg2E3uG8yfipTBngRLVScIV34bYgGqf+6uR8zxE2O7bbRj0O3u7C
ULEEsgTZD/tGs/mErJy7tWKRLJJCV3AGdjQg7x3GdLO2zsLXzMyBBm+xc4hmAw3OwrdEN/zsGs+6
5STJHMaXbMwz9hrl/Ncs0a1W3x3T7jx4R+eEZ44C35J4tRjl22dv9rVIo+pImqiXv1MLNrHsuyHa
mE2yWtNsxk6s6NG9W5MA/3OhXKMJjupozzM518CgGGOQ+DqBm+CiRl5WLAE3VOC7mItFx3Oyw8UE
/FzRpqjqJbIsYF0IKakxoWvrEB/olNxpkwG5dYHcmeMRvZzRJXRckA+O+aIc5zH3bAXEJrp+S7mn
FFdzY1+qu9Yhejlss4DEAoKQEooM2PWLFinKNtYdf8BMOJP170sruBXSzqTfwQp7lbEZjNalS5A9
koP2OAP1wuwgS/eyjR8hO4WAtGMwZJbsNobNg8F9Jju5NXUfabDaMveYuGhI7VXUlJIrC9X1t4rF
drq3W2O6LZnTHm7ZCE3/bIIvRhZMQBOLkKFE5SOSPvaMId409hreNezvSLA8sUYhkfhOrMYkUEH/
9iMIPHaG+1GIXSJhLlGBRWs9oKxPhO7boRkpp6AagGZK0GlVoe4NIlv+E+ZpB4MsMUoxARDvCKNF
Ovojl7SSQNc2uNEbcuHmo5IjX8ICCijl0zPQY45K+VWWwUVdeXKStCvvENgqKJWIOJgyOd8CDqvD
xYdP3i9+6Yt9sw9Q9zOY+K0sDjpZA8KDSl8CaqKIrbGgQGcSIWydMhsJf4EmwmySiDA9mcMzHVxu
luy5gj7Oz73KbLMglTE53C/JFhlw440CjbYlhYdC13GhnQTjWcM7skzloCNkErb2t7cm53gRqfkI
eYjuDIjCGUlqt919WeJUvH92MSawydHspUdRDo5gCY5qqHBhdptfwpqaQXgJBC5x/U7/PCM+ZL6T
mhS3Ou1noqpxWxMqgTET3CqrW0H4FRJkz/rVVa0QE/vAfLBWvGpqSUlh67SxRscKY+zN0h9HZipR
omY2TL0D0QA+MzF6Un5tRBaHn+AS4WDmqYYvNXMD88DrQMpjzuoCOB2o4gTKzazQM3wnkiA8GmOp
990kItxmIO471jUz9prvH+ZxWP444xZPBtdRfzXBStCFsQwoMhCbk6tUxlzrIvT+1RPmV2sKZmJ1
iP9Cy4kzlfpZubHLwNljYsXIi/XNI6wjISDg3dAfUJFgoSKDX2Tg666/1XkJjOU/BFrRNdmiXQju
CT+BfW73RhBaAl8OJ8U2M3cbBYfg3JwRICfjWKf5MnCCjWp2Pmluwv5GmI0wL0oXnnfcWQSwoavm
cIU6VOQGU9eN0Hv7hKsdRYJp7jf8+S3QJsBtkBijVUwZ22+QLXkW09yZK/JQDHW9q/CPUMjH9DaF
axtIkEd9NF0WmnR1iERqv7qXdp8ytUW2rH3ib+s9sCjVN1kDMevTqyVEo0xDBTuNHr3B3p/xChZy
AlDD0Lg1A+4fKX5raZRKSt9Cfx3C/tnn+fDZ+ySgw/Nd6kBfvbJ2em10cid+R8ujcspsXmep7Uzi
kRTesxfIbNMbOmaOx9jkPUhJD2JYLZAQ3WaRUQKz5LxqKhUkRjtpsIvXJEmnp2wHtqZfVykym7Wv
Xy3rFntsyTss8X1PoQ6idx1BwEqLuruNVLPN5q0I3Yd0RJoEYxoopESrAm9HlNNBusMecuLzCCTY
CCroildW8h/ito88by0CcYDAitEBilyc0MH4fvtjeEn3Cv99fulmICwTZYcUffE3WlR2njTFbPQb
wt/F02JYwd3u+kNcX6WeIuH6vXc4eDAKjHt03z/f1uUFw9jba0yzfQthx5c4y9fISKMXUiDTOs2M
KRnrHMJTVI4uAa/+MhQcvQ7VouMqvuvLpfsXZ24mPy7XqnRGifSenFRHLQYtYiAjljlJekfcd5DG
petYlFn0ipVj0K/kHZw0Hy2bNT5cJ0lSZUZ8RfvvhI1q5cvMlWXwnfl1cCchT+n2KD9gLATRE1XQ
Xgu6xlOy9kBvpVfY2L3+rLkGx1zpWUT8QPwGSeMzUfxmfQzxM8kRx0lmT0fLmPYX0YOc1jeIRIYA
461MOWTfvI61vZTf2T7v08fXVGWUtI3Hp7T5BP/uTVc5DuIf9o1IWFNBEXQcGJZKoWojeIbrEqZN
mxRbwac1RiS/dWnJYeA5LnEodPnLNcO8ZrvOWq2KYqjSZNCwE5OyW6wgI1e0Y3ZsuP23cS5NMlDJ
oe2VMsA/TsrHoOyI6icqwiktzBSJss5qWzaOzGPMOZ49NdSwNfCh0MpBrsFLCeOPA9KpJe70TggF
/YBi7FUAH5JnmuWuQHqhFrVURIbRiZsv/jawc5S9YTRHw/LTT171udTiQiE2sI94uSec5rh/Y29v
oAXhIJrdn9Vn95fUUceJ/7R2BAuxMw6v/qn8ppJn/dXkTW1EW63rmEOO6D95j/xR1klUnoOFxlSv
y28ny/BDUYGkpcH55q/wPKtFgfXzz6C7fz7VdNSB9Z9wtUtBs48FHlOqq9c/mPQScGT3PKZjLlqc
ROy4ilQVkdQt3pXvOvXG2udy5b/gS+lU26LKWh+8FJ4e4uOwwyT3tBPMqcZAsV4uOmoUpf6Dwp8V
P1Wxh3rviDyZgQU5dw1H0i9NO4iG95VjAydTvkP2tM2oeddR93+rgN5M2I6SbsRw/wvjVQ0IUAJx
JBYeVXJAelmyQIACh6M9QKYOycOpeZ9iE108r/U3twqdW5IOzkj/uEd69HR5j36zAr8JQ2ht85VD
CE6V5v0rMTbJopvdjnEPcSDAu2nni2SuaxduFIVf7diMwkANlvIhP/Sd4kh3M5a0NsYTbxXaoQwd
eUlKhbXiu2J1J5z3DF7uH1cq82HaYdyrfZwYbSYWrhv014X+BL2w8brU1MmDJXVs7lL4jCYYhfQ0
OXlBs//pDj5YC/AtS5zsEY6pFeifp94S8ovmY0Y7ibaqkHYdCJEoMP+yHOxeZEFm2+624trkKoM1
/eunY9PIKKF7reUclLknZ3BlLM7uWvV8uLcU0oDukRuXpFys1PhCtDZglxToEOxVxFYh4Ldfctu2
IFpNL+8JcVgytYQrSr1aaJobbA6JOAOI5o2qF2+Gj+96PdSXFouOJJhB7CF+huCXykzNiO80hVjL
EsLucx/crwCRAId1sfSI6rusbkIFlQ+Az8H29QV8y5tpsTsrFlAnOJMp2vRfk3GXHPevDC8sHCBe
XJLbqzhEqcGmT+GwyErat1SQS6lX/VOUT9YPc7S6b/r7yttrLiE9kMws6nq08eKtN40mB/1p5eoZ
JxXoQt44npFCKceLtjElgxIloBLM2Fy0WiDiDgBD7OFOF/RKMhFOsjCuJ+AYPXKZGh0Q0T/kbPTJ
nwRwsiJAUDZtDhAw/zni3zaBPq2EHhwwFwCxaJjUGMGPfKnwGeQQckoOACggEnqoygBUWoq35Ge6
B5ktvjIwXsbQPk4K4oMMBDFH7WumN3n6edO17D9mDCtKFM72Afba9LeZY1j8LStFxZDuO8gaXswl
v60PAvEZT8Ga7lj7dizRSfI/R4wI7lKWKiXwiC6Xw6CGvjG9C9SakjcnKLAhJNdUjcmhZj01rvZF
/Q5iQsy+gu5RHhUd1x9Ndas+XY3hP/Kj/sGhKWobR2cavqAZLVMwhYgEJ2lnBc5pWlbIL+DZ5pYq
406DOm9m1w0zl1kjxO2fU9pFW3WcVJUBsXDsWUJkjJqxqlHanfWX+VefW551JugyY6qBVbIfaegD
rVQknCbppm3PKtTvNTS/9tVTSo0UIdeDB5vv9UAgkbhWxfSju0ChgrvnmQSkxeEuITEHz4+BI6tL
xl2aB9GM0S+Y4WsggGT8II+HOIauAE/rpQnuFJpFlaW07bo8gffXSCcgmZBp1NsvVFdd2cDrHTEc
AnGZKVhZydYX3zIefXsfdObY6+x87VsKTjKuIU2uvtc654mpc5PBlKB2BSyjF6/IvuXg8TpH1ZRq
yUW39E89L7ei6NUOLOayU/T12Rubb9AtMg/Qvt4NrC/bGc0WCjvzwEG1GNluCidmIQQXyGexe89C
KiTnvyOdN2m40YC+l3ii3j1SYZLcNT28HJSCxDoSNO6aKjK3KTbtbtoBAxrjz0h2+yNN9vrjC5Jq
3n4fyWTaImRSwu4JvnHyxalCPZxA3xnRh2vxbnzhlvUvyc2txZxlDWpsj8oLJXOyRwmE0kcGw4MS
IqGV0jcCICtnYmP1dWLzdmUTdPWe+u2u9l9yj+L+ozT7GDN//jHwOtwwcaQPJjPsACY4jQwP/B7Q
jZM4nlfYfocvfHPIeTGeBGtMMTQaid0CNRKT2DrfkuhM9NK6hj8FFGcSwLmaYRnJV5PxrYWJ9z5y
fXXlnJ7ItwRm1uoe38uLr3Hc9el0qq6g554MeIevuWZxs1Vc7iyANHh6swJbO0b2EA4j1eluk5Vi
hIXeYKxJDxY3nt6UncjmTCelGICjLwYnnbNaHxqvK+XnMNcbM+TWDNGrMs+ElpJjMjiStMOb+F0F
r5A9McEXnozb2+VLQ/TJjQw0K1wcGmMcTa+9ZEkQhOMzNjr7c2cDU0K9Wy4pXMIYGUmkBoZsk5ex
TPS6pK7UyUmIwG1oSu+KRHpideRRFRfhGFESjzp4HfYRw6OnJOiW/0kGPS8cewwmCU/DeHAvyjxX
Q/e/yt8Bp1MKJYWL1qx3CJUWea0LXmyf1OlG2fDnb8ZixtqZusV7m/Mg7aV3kQczN1wODCsWTNZm
rinIU7wOcCXM5XkyTrPtS0toW5v5KoOWiMJvSrOrIkDMHkW0y+2F8c7DIplq/E1IB72eqtk92jeq
GjwbZ2cmJmyhzeTLB6Qfs3ZFOTxoLxp6bNr2H7edjpF2UCEse+XhjCJL2DarQisu3v+ZZ0KzRGCJ
y+f0MB3If5+wXJkEG+zXK9X65lqzXpzKSffyipWa2Nt0n9VwWunTE5TMEzbH1uWHXupFZOMcv3UB
LAzxfZxgqnrx0zGrrEWFXtEXx9iOHdiUft2jYqmwdvGrsp8zXncXq7kMVTrGgUUcTympCQ4fCQP+
cOVLvPzSHzbbTnucYnXd0WYcHit5zyt5O0rnP16mB+rQZ4pFyi/FZiUcXTw4Bm9ehIuijJz6XUj6
isz7UDR96itwTM8mszBsYpDsykHn7hltotnRjDEGh83BEryxuieViHhsuKmKR8VaPj1JfyYcT7mR
RiebHkJaZwaVDuYs9A+x8L5MlNS31Wlr/7tZouhmE+B74WU/D4IcOTMmxPu1e9UcEy8jLa5gC2Q8
u69OqGRNFom6tlqeneyvQGYM8yAScqrqwA6iFTB/9roJDYqhWOb+YoL6Kj5cFA9poiFeaBcpCjzT
rAb4zoDaeb6fs9ab1GyB9zxVXcUovT3NTa4fdkXjZkQluRSTZ4UyUnuOQLJE+k3vZcq4Cx2Jj97G
z1t3OxQRHmLM/rNnOjDJSBBVhMSn70mdsw8xKlTqlakRKif7IJLeaeRyVZ0YohsxyP11NCmbB+Nd
KytNe1w/EJthzK1PxY5e6/2CQyFFdOUMCNjg5k6x4f7WodvPhm1S19zA+R5aGYCQrUF3uPMLfHI+
MfwoU6eAUucAmD1YcjWF3uAXpHiQyN7RJryLYpEL0BSoJzL6K8PbX4mSvuV8WJS3VWjGXSMPATUe
fiTiBoEflsiIiH///f7Hs91chFcQFh8KJnF0VyK9GGHUqqa8T9uUqJNGPMxTOru6D7WgmEFhjuc/
2Vs7cQb9GK5W59WRTKbs673JFjpaY4k0jGSfvAmX+86EOgR3gtmMGzdHaX2qgyPH5khHBQVK2ZcZ
tRvOmlaEQP5w9cX54xZcojHhWgl3UKFDLQwMZnRTb5QlGZviplr1D8hb8o/OTQcoRJTISPBoiseb
esE4ofu3b69bDCPpRiF/cwvd5M7sqfjIkfyE0mUY3w8Q7DOyt+plGIebpOKmpY+h535Z6clJ5YiD
WXbDHw2iszbGNWC05i52GNnosOcpv9AljQNycLiqWuAORITcxm5yiDqdI3fV87BmgLHKHGmrDoxz
3ZEtxo72pWK+EqOONLPkPWx1Qcd1lkik2Kw/jeRWPn+JVe7J5B4LYkSupe/dv8wkVPT6f50MQFTG
AbTHSS5rtRGcCJHYQt1vPDxBt68eoazG8SZXaLDVrj4xD9OUnv5c8+/V/I/ZWjptoGLWdu+mOLJx
S6noE70IN8A0kglWeQTk1qUL8U+zGtgGPOnT9Mm4rK9TGnsZihmVrnSj6/e8+3X0ggcheTHAtOnF
GzDlwcl8H173LETupewU1AJ0rovkPST9OrMzkGdkCOAhS7StdQcUJQzNp5Iu4WU+HCCl1M/tbsM4
6WNAf680ByShPAyu1MK/czoz7MxUBAG5Xpl2jdc2N+RaiSF9JHlTJ77CPrhZ7X6IcdYRcNK3Pj42
H6N2Kj22wzV5GucprwM8J3dcqKbYXUIY+a1xzYN8xgWpNSHWPIzXJiwRgyaY3z6+izIjxiLN07LK
/tiBMGqIG5kbzvVAHG0/gXKr2UtbpFuvnikwRSWeXSOS4CBhjl4fIX+fzMaU6tMkZqse4ROoEuOf
uNYYqbAeltClVKStdJS8DRfkQHuapnZAFQEz/7hDfNfoBmh8Q5hs4WyUVPHi8BaXHOyOV70s71sj
SH/gNCW4KHkXDNQ0FjeM6J7cffoH5Ia3EnO18OA0mrlaWsl+2k1l6YDVmffWbEcffguvdItLtBlA
8SmCLRw94rGmuaA0GDkYCFAKfbKno5LyS5I7tzS4DbUurkaJUpy6j+0NF+nJeSEPzwRJUDI8FU9a
m5mrMU5xffkYTltXvzDATGyAPKLQYBae1DeDQ4OVErh4VRVlWFyl9hE7ryL0MvXq9LZAJd5d7/a0
9+lDVR8BJGHwSr4Y+yAMwTrJrbKkfxXtHrsA/FR8NN56xTgueDPP4j9lbeE/mZrIV/xGZkcVeSSy
7CgT5wlPK/R+gYLH49VCVrhASTpFU/FXN40vPuJmY/+CV+oGRMIm0HtZ1h2hYK9vMmkr38c5pR5O
FRy+2Wen8RQ56Yy5SQ3ip78G8Pg3SnjaR8u3xmcaBTewiZ4wXjaNJYpdQHyZlY9MYSJabJpx3VKr
tQKK5ouHGplnwB8TLerQcO7ijkyBb2K5XlhcAFfaEF6jAgo3oBAaH0Qc8XF+3yneHUUgfvyss4BW
QwYfUOX8zt3/5LGAAXOMU1TEZe36jjcsbjG04vSomfz3Z+GlUWiWkB3OKc6XWw+fxWjrwUQe7ORN
9YP5LG6j/y2n+WVjyPUpA8yhhmqzfxkvY1b5sx2db/7cUGwDrdWr3we5/3HZEFyK4Y7ptC34vbnK
rtOoy3Gj2qx0FbZTChRdfoBe0wMXE+DxG/4xzqJG7cYbtVclWLaGAJWHG+HPCuwY48ReotnlOdfb
3Suyq0yztm2fUcUaMtg1j69Rlrbr95gmY5+uD9NU5Lbo/TX+XGuGsq5KRJeppNpjelpcaYN+UApM
+qOsc8obGZ9Yhz0GdW9p4Y7hPRbpIiUOzm5Uhq/dDIJ4QxePQs0LWNl3jTvyDi9A9hwjrTtxKyEj
GGLJxSIVPM5/o2ZIKzedojTyWfwkjdT3YRA7BaUNda0HGpNpMvkZYGcKfjj0qYKmfHQBWwqgB0mv
aLO0r2om3cgwDlvp/PnFkZYVP8k8n9Jv3wsdgTx3WJRU4MCtOVuUdWfOTSkxFCDw+tj7CSBMYsmh
IChwK9P2L+EkGDG08vZBdLlLJZ8fdFMIBS/Ey+wZXeeOASNcNYrUYWmUYbDZ9vSrLvrO1q/l3itQ
n4e0E3+o+ECkr9gIlFyc7JPg3cVZWWHX6YMh9Yo7y8oNGgAdUkpRkNo7ZvXgCilfiPJ2grKgGJCF
rp1J5bNEg3PTVcYn006/b4TUE54mxNFoRclU20iUZTVfDlHdRPHhO92MQQw8rL1qk7P3bCXiUMTE
i78X/h3DAh5eoIlZ4xvSmfhGscFp8TzkRcfEaDUE13M8NQF2t+3GNVoYtlr0t9CgwcWqEc/LPvwq
cHvAyIFnmPBqLjd/0GzVM9BXD8lQB6J2VNzcohiuqQKykjMmuZVybtqRB4blTNF8/ACcqo54umMq
uXuiv6MgeIBn3DtTeKnWfbH0w+/mK8RLyBfR98LfcB5JmGQakyS8xOf8Il3b2sceuAfkNr1phbts
gQdanTPbOBZqxyHiwsNKUZUyhZAzYs9QnwwyAq+4MxJWwZAPYuLX0wW7tnHtSiEhXwdVqQdRGYc/
AuMuzFi7o3Um5XSJzjK/zpi40ijq5VcuZoPTfolo8CVarZoppeKFJKFNeK+aih8j1TOTiSfcGERu
8ZaZXobDhfOY5OkordFjW4MfEu+uU+SGxLPxNQgS+9KLF7xIAhieIY3239XmbfQa2RiYB55XC1Tx
Q5Tp9HnYSzS8ZULttJIeeF8VeV1UWaxTfKlJZnJDvlyjP4y2DXC8nJav8yEpG/lT7cYYwFk7dJv8
b6kamCQ+D0724mLxSVi98rdRJ8h9nxRhyw4QGV46chWN6S52NffDoeoqsMHohseJpDej/WTB1UHQ
b0oCaXJcTajcSk+TJ5QXiSWz6cjl7tOfoRHKsdU1X2QaZBhR/aCTB5IQ1UOBEBCkFQ21TMVdcqkl
hA08O0NlG3gjkWmEKFlw5YMblsH/O09CiAzWETVQnevhSm4YTGgsBdC7mrg2tlPgiMrVeEHo1luc
n68udy6cOd/KogQWlfRP8XKRxZc0IVy6w9wCivHPfSTRm0MjrFhixbiOaRSDkWfdyNG+SDSXOEFX
3RCapxZeNA9rBgA7R6B+mW6b/yNGj5o7wHPmETCNsYnNwTC/ltlZrxKzMCeLMj+IjXbWv47m5Iwh
L3+6ot+Jua2jbtQaMoVLaRODcegC1KmgrFs9akWYaVqYJdGzApzLnzqqNwMMLOOYOOKkh2REBFve
VIpUtZhTQ2Gnr2EtxmOtIU4oM8yhZkfyoMtLoRf3cHutFbTd8L4HS93IiAjJtXgf9Jity2n0NWrX
EEE+0crZmQ+ZrcF7j10TVlL0ubtkXSoaVvLVKF+YWI1HwXMNXUWgIU2vSqRv8QYzTSEED3VlhcL5
UtCApIwbLHW0r+nm9daenltCyRNTVjf3devErltZDXw1QzSLQE+AScoBE4lH0CFpPhNOcO2s0Ajh
G7sGDvZW2xn8GqoAdbEyuexp0Yl7MXGwDFqpjPTGK8P9iQH6uOFIL/pqtUuQoav/kDY4hctYE+br
DqZRoeusrNnI8ycjwxpXdLvGFdTM/EEiBZzeCUcEkLQGrG5ZhrU2lzNUws2FbPgYhdY4cX8gxsFe
wJSQLGS4w3jz2Jp/xQ4rOOtKSyRVqtWTIHTFxmHWvBhCTgZcP08pTkt54Ai7gI/8KV6OIe/FSwuQ
a+I82svWIVDZ13hdVdHiCJeYhOjuftoxIA6DqB3jUWvfUtXjosnjpE4o9UHjEt7KBMpn8V5vjkAf
gdL4QGT/FfNT56y8ujNmDRRXh59yYPzVC16CfmK3zI90ux8nsOhNELcZiVayOS84/J/rFpC1BoN/
Arx82+iUVX5Jvvc7KPDxpsNCmXbsF0SkDGUquKLSfCGgXTtq9WlvRkXkDkmfiHDC4eaD/Jf8yj6B
rEHbgpTdZX3DlFNIKKqtaKnQ6OPWxLbdrcF7u55TXSC85OsfZhKjbT15Y5KQBaFoCEMfqIzOw45u
lgPPZwZ2e24sxSG/132xQCDfUSmndf2sjwkm+tOv6FNdjC37Hr2WMqaPJ5Vi4q9TK9C2POmAYHRR
roHU52s5eI1iAU6LmCZyKv84yKnNoSK9OschYtYOZEm9mwB9U/hSCV1HfSD1LdPbMIk/i2WexOXi
IZCrxUxuDxUIMYgEoCYGhoy2WBtOxzaDCMIkZhnKq5jfOq1Zk0bmENM1QsRLaTQ9NC/sK+sR4GfM
2n+Mold15ZMNrhnu4MtChBkgzEFEPSeI2vnyn0K9u1CHBF94qZqzDtibFFh14siYIfAscao2F5X7
3BJhtlHSVFE0NTW8z2rUhXoy0Oa72K/fsdB/YQ5l9WSYWf+UXXbzmgM546JnbBmK87mJON21cHAo
WjW63YbCB4NO/Yn02A+0wyf0QDC/SR1vYjSoKt5TS+fhL83ThPWXycehH9Ka3s/EysLaP7S7681J
hT+gH6Ul/ox8v8MRTaGIvpeJx4daGXAQdfBShTqYwYxTOxZYXKDE1IFZ1Wb5dkQPgrL92YFPgscM
6Ii4TUNKME42NP6nAKcZYomhcANNfeD2Rz84AuQ/0BqYil4E/34o9kXNEcnUUuCdE3K362lymKhI
yF/rf0VPNnO9QBcprRe4Cq4XgkTClAa2kfLxnM75u4Le0wcbIXQvhHSc7LZ8HJleyvGaf/+gfnlO
Rf1KbFZhzaq1RWVGHkhqqcrcm8owXDOq9R1rSuOTQqFQMMJt+GU68ZZYR4xgit9SPIWxSc4nvLQS
+FYyaAlM+ybURNSQ4gwsS/lAm2XNPQmwzkiA8Qvo68tHCOTyOa2PHzA6edEN1SsRSHVbkk53ZW8i
cPMqll/igxNK5V9P4C2pZcns68FBp7aWLZNPumSnvsQDFJ1yUZ//f0RTJhmjkSJvn/iolqOqdl1t
Tlt3RsO+qIitx/pyWMwN/LfHXrSKt0EUhMAay4GPnjIRf/6YWc7/NaAIIRwtm0S/ZXebtDWEsB+g
zpK4bYf9vLt22p+uLYn7ifqM0yq1z1G+5qbbpMcn1fhCXYP/AKJYiXj/agKcGIhgg/bHrdlG8MwI
EoV55OR/QA3iDm7U9XAhoa6dArnpX3nR3uxOBB0B6ECvf/C3toy9+HxR2YDShzMQ+tAHDd9GFF/r
UKEO3PzUe3Jc8ad0Xr345c2SSP4tc6hNCI+fMvvw0CUJAVCKw04GxicgK5+0R7vTXlSsCQNhT+ev
+Ria8EEM+Kr5cEhJ10hPMKzztXfrqXp82M7sx10sVqQcJ72L37zwRNAr99NgKy3cy8UJf/uLPOXB
t5tZ5pFcYPXQYYSwff9uFS0xr+bPyU1p8FU5aZEbwU/INB6yA/cwEvKG35ENVN6Ahh3AQe9ywUDm
rv7L5JlvrYD4kWqSGXmzP+FHAXkFKQENBDsHvkbJRdVbsPdshKXL+4jABhj/AU1BWftHHxqM+LeV
fz4ClnVaD9Rx7r1Q5D9UU/8o61IgIi8jKmewbXRbOLnClFDth1DIfAy7cZzi7CUbYtKLYgKITdli
sZKJzK3poDKr1EOkkSLZSRNLWKErMTcJyVgW2xxi8qtgaaZOQS7cs5xn+/OYXdqOVsT8W2ocAiyg
B/bPXCtDeijVfZ5yOUoBVqcpaZRhMMm3S3sQg8fZjCqLQq+aXzZ3E7rbh8axpOM0J1XI1Bc+MMwW
zGiad3JrNgqW/cg3/SSmLt6/fC1rpGSsevMxIRS2IyLnVc/Atyl7cpPaYv0Kn7FY9HxZBTSwztJK
aVNWh/oMvGJUBxqQZ5gFjWXtuWk01Eupkl3yuVP7YyJwG4Tk204bhEj8Grt1Vx+FWI0kJBD1KxuE
nZFgxw/jYl68il+oLfn4LGh87IjVYkpeOoQECRLRZh96NRqjGOzLVviVqVSPbX+ZPxz8tHVHAmSe
G6NoQ7NgSCVNPpZbPxrYveGGIRP106bZtKWAoaY9/C9Rv9TN9Su73lqEE1xaBozgdQf0RVj6FpyN
Slhqk8ll1lGZILN6rWqEP4mDGm8Fmlj3F9f4c2kZHs8GMI5/ARl+5TexGFw9ShRVnZEBS7W2+CSf
+C8BWnuK4AM7UHq6vvimT4QNFmscNUDco2HOsdO56vKjYGLxcMF29slUzfwQe4pNYy1Cxn3hHbpm
9r3+VqDbXHYZ3t/EbZQxy4p0DZEBB9sHrIfQxDUm0Q/qQntqe8E/CDYgn2YpKKOop42/ofiirUA+
lY6pYaBqcZQwejYmL4+INw5eSuVkQbxz4Ib2c61zAtGjiZeNTRljpaEvpl5OwXAf9bs4kR9haXMd
SgVjU5cQeEdG8TumaKtg8mkKIvxJv2njOJBKo3SH8YP3hh0Tz/AbTgxz1SRUHaqI6rugfpw+rrPL
yPY5fvHK2jiDpxP9uKM6lziew9cgbGFj/XRrgcvh7CDqSUexJtfZHKBaOLJhkhBPoesnS2Yh1g2y
85SyMjmIABcI1tkKpqQZlmIxfqvsZ9HpJr/a0mcTQq+aPK8Fa1iw9cg5E8Ehee91hVJ6ULMml8O7
gLahS8EVFX9LcPyknFBGJs8RaxEP03vbb4HPmnA/3YNiVwqzI4+Yg+NJV/uD+2XQ+KHInRY6/2Ly
68EVZ+9ieKHZVXt8ACQdaF3shllZ2dFMPDwzwMJdY1WzzO7LALpfjqc91hkG50oLO635fCUbRCl4
vlkPmi7iXOSsff37LbYY5rJ98YK7IP5g27oG0HogiwvpO7q3c8Udxm3RrzzxUxzLgNAccPgfYwQz
F/rzXfjgswf+r/8Dx6Trnx8tcRidNFAMHkjUFmk7zcvVoYb/sCl7nK1WQZfol8+J4jDNJwlBu4Ka
CEdsBknrMIGq7GMA3mYRmWdzOQLDIHuK5g/zf30GhjJ6kx2lqe9+6ZT8ACtb+5dY6ClKBjqQKD50
Kr/d2wwhWX9rz1kkGhO/Wn48G+nkg6fNmUZr+wywIE7/+qmK84sTAqcFUxfBdHfp5JfoKivWMoN/
aoHSJ6OzkkzwYXXjVRnczNS/8d47uvuOGQu8KAr+lxMDl9cV4sOHPqG/6Wv8aa/53Dgsa0ovtx0o
hfzoJaABfxVQcjY+EXs2i7VB4akyPW4jAhpDqfAL5KItHhAWrkeFjT0xow1025O0aTyArXgecNuR
9DCo1vJ4o0ZR/FqiNDzWrvfyEat7HZOH2aw0RgNOsQyrdFTfnSvewwhadKjHMTtNOpCcdx7Xpx0c
j2zXT/XiGv2RIeYT3GqSO8+iHM9POR/g+kME7foJWLQ0K8bPoUZdMGHbN/PQdIkcdbVfeKnLSJht
K1+qz5tCMs6SqdsRkIxvhc8vkaEgSMPWvnpylB3VEbZ4NYLvaitEXtFGtig64wZwSnAuSXN8trxT
O9nTypwtVen7Yq7oxpl52rZOLZD/x7g/1872pB8LF6nHQrEdU4BL/4b7xsUAXgSMi5jk4AioXSgg
78+f8L9eTIyymiT9bpa/vqU+6TFWZhfb5u/L1h5YDFxvfB4DPcMhHQlU+jY6drLcQInHma3lHBx6
tvP/QFvjsOb5C+YSzWP5p4abj5Fq3hsznToiutXZ++IahvJhsaqUDwoe59qmMf5THJMhCy/wmnyn
1CaKEG/WX/VMY4iEQmZDYmPRrVlktScxzEO8JSJc5twFTkCYvhYkWeJ3EfmwqtoERxi3MwYVGZiI
YNxCf4FUfmTZ5CyJ77lfrt1PwGtW4WzTN3h2wt24RtOLSmfVwdrhxKZUO36yabaG/0RHWTvbMXr8
FpBkKlmC2CGdohDneaH+mbb/JakMrEHkOIksCNe708oVmpeAWBYy5stTZg+pEGe5QZUUGehOpCT1
vdXIh3XQKiAVHAXKH45O+7QQ0MOvoKk7oz+erzDO6m+6KIevQv1tSY2UQpjk6DRNs0iVIL7Czx4f
PffaMTwDZSpa0j53Fa3bRDJmWV4Y5/WkKb+vqyPsk6EbazUMQuCJoCkhtgDEMODLZ8rNsxPPqKeE
Wg1MyO+k8BvlM9lFxf6h7ULehPJ/Wi4pgI+v9+CNRoa4QdT/MN5sfSPcZU+kOyyTjIeZLvdvE/wm
M6cGM9Y5C8rmXnRF8JE0qeJ+Jdtw7PLrW3D21IaGKPpIO/x2MKMWtmslxE84R1fz15vYOKBPNlVX
RXiuOJYwpIIg/9nr4PcycIiqM0r560jBdI26hbKzjHUN/5y8aafdAajgybcyBlOcv/29dPH69sDQ
5+hR8MouRchayQsrIGIkIvszA1tjKnmwQCKmRg2VH4L0f8N73CUV2jiP1tNFo/zfuZF774QQ41Ky
Czdb8FvVR4mp9w/o24ghHtwrfViJeR6qEXKvck2RpF0fMux1wl+ISYlCyXXX8QGBafLNMrqOE2vS
eohzIW/nUd5sRE+GLhZBOLCC621iolQ8SeYp+qOiR1nV1quxvH6LyuTlfKnpiiCwHzOjD9WoiLxO
Eujjzz6XTRgDLKtKfKm9Lt0rujtBF/4J5CRUnE5+XDMQek2ASlHTC1p0eCEQ95DaULy3SOhhWyWK
cYFAdvVFeCxH8Wf8/Q579DzLu0F7gt1IwOOvzCkknUMFjfD3zeekGNXHLhi3zw8bt1qVbi62WeKx
DkcwJ+Tn75R/SqQq2qTUTcVmPe1LOvghLQirC78G0QoO3qkNTjBVDkJD/VQpx7D0LHTpQwPr8Qv8
+VTLeuKfOXGQT7BzTByA+eD0gWtrw89jsuMmhm1BuM+2//SV2JGh9bBxJYWJSl5wNtUOkgXIAyOd
D9u7Csq+qd7RdJO6pKYtczOzNnl4T2hcdqcKmQxmb3Sr0T2a9dSL5PYydvcK3eySkPaH+XkY6mm8
NsqPoMEEiIzZp5NHq65N9A4Ww5CI7pCmgdzBcw3E8mKPKLWlqPmZepmpTed7pEj+Jn5eVcrHhm4B
dECUyEEXxQy1kKjKng1DamzFeZUqtgcWq5sD44N6PzWAuIShjVnM1bKzJupeMNH+hodaUXj7LpZW
Cqh21AvapfTHLWD8enU0jR8MHvALqcNnTk7ICQOiVCSVWqZCWvUNh9LvhIO9ALEP9Nkt6o++kArA
PjWiDgCUuNpRKSSit3Y8gxCUdh7mdJT/lUgXswwl8sVFOq5YkPmtCq+WAXD+1JVsh5JnR0OcqFxO
s93BtQrLRdDVEwZWhftM1zBhfsai0ltnJP9AUOy+Jpz2aYC36+yM5eEpLxROyjt8EqTiJcFK406S
SBSfmtvUD5gLa28ldxIUvtL0a6pEmlxjLVBUQXMjJQQUejhm8y7pFga9cyg1zsGuHf3e9EtvlaV6
hC8QWOx+tpFh8msVA8x+svosaRSGr2S36eFLB0hsHOQ2O2L1ED92Zq7TrcOkVKT2EOVpAxwPq2DZ
jk3Z1tK/gQ2+4r9n7edfBO+//qgW9ItunLdpzslVe2uzinny/SUDnjQCaPR/IZW/00Cr0YAANX71
MPNoqXVw9EjNjh2FJCfU9Wm8NSOSMC+kv/XhdOGsWcZ2rutTVoBwZNt70HDnMshbDwyWm/WgI7mc
Q7EshIlvaxw4mIHg5ODUtYv6HjVG+dQi5SoopqP+Ct29ECWj+qkGZp487zRSrOoKHIwmyC6JGCTy
mpFVd/9wJuiJW5Pu0GJdxNOvjWmw3ei074KwreNRDKF3WxQK6y1Uhtr7EHTL9gAF+asyTjcgc0qD
RElU4pv1QDYf0G1gS5fq8UbC/SxxGExp/IPa9aagOPNJZ4qlmv2g6rZfeEIM3b+RS7EeonsTU6wB
vgIIBysDMQ5ZnnIkv/la4chouAFUPYkLBfelzotyftwP7Ia21LRjFP3ts1kaPcA+grJdLlog7G17
yxNdO0NO2UgU5Yk8kLy4xtmicxZ62S4h6fyq1NlbghdRORj8zpwEDoZJMxsJPM8LL3DTGNWH4CVn
m58U173v4PsKKtqK18zsl3UM1GVLKoWJTED3hRdIOvYgccvI9IZ2LTUic0hcnfa1AsCC9Di4ujPT
kcrpA0kzL4+T0NvQ4mT0xz31H++QOW6YMlFrCvC6fm5Ye2xF1WmkvLdL8pHAtK+xPZB08fRsDiqV
2NA9LaM2T4QRQCXo9gT0iWW1cKGeA909p3zloa9p+Ab5ywxndh4KzlZ76tv+QLvece5smSSRK+8U
Wr1jicM8ygLdYzSdrNwTeWi0rrn4kfyKxiXEMI3iKb1/bjLy47AcFO+bCOHu5YjPUvqj0BATQkZq
EOwp337tm6fUXov8w+7k9Fmlfb+vOHCC44DqgVYmhyatovhdW0W1QN+yS/gsXQrTvBwtDWyD64du
qvcxNpZW70Iqwwk2hAwmmXddMPfzdZWy+WpLkF4Jeng/zdDImC6L1Kb5WxTc83T5FCbJAwHqXi+b
Lk+0buMW0gLEA8zRnjGxfNWMimlBkhvOqsmqa9Dx6eavYdG73rYyefJy/FKXdFlccZniY5rn1uPh
Qt/Gk0tx6q/uWD5eSvmfrsvfzPqggw/FA1rT7djNoKvdHBnpmecoYTuQ4Apx1C7PIweaAwtTPIKh
vJNumZGvyj+AGdrcjX7t3zQGtEv9M1/h7T8/xmq4D30DUbf0HZVOXw+NM4R78iwVoIf1+j793pox
AsDrtksdSS3Z5chIXYn3h7kXSnBWSZDpFrQNqEtHwAyGQF/hIWFcgzNB3BKqSBzrLS6BxqbNIGPF
l675dQghmji7gQ+unALnxy/hU0btDDczN9BnK35mA5L2xEnvdJcapr1LuRpqaz5Pcv2RrNhTHcor
TI90aMfx5MJUHmrusFJ/Vhn1aQ4RMoWnqJDpJ+61ul55rH02JqacxLNmgHf3iCEwhDF22NjYZu+i
9zsWdvIuDyt/v+/MEfOYRaQNECmreP9kpbSDNpz5mmTuAbb5rd9U/IVQWCWG5bfvyDIUPMSHlaXo
hmryLptsu5trkCasVsUDX07TC2yGZIYOSjWtYCB9qLAAs4qjtCavpaaJAUDT00lQzhxRGo+PtG05
8ciMK1rh1elydfY0WOeRkupxTDCMOCeP95SzWNe2LzFgcyxyiC2rjm4s3fTzrvI1aWAwPXUqiUV4
CRsbxp6EvaX6dCzerkeHohGx+WkZQfJY0zv6/+B6Ds3mefBnd90AbW6p0Xjbf1o2reJHcQiZa2eb
PaUzCk+OMn9qx7Fb+h/oZgD/w6YhPIWCZSthXMw1vVY0u//3VIJQgDrYBiwgsvPeBgCkSEbxuqUd
vnsi3rTtz60gv84m3zdeJX8dYxVIa6NoMDbZQdTDBEFJTstN9wLR6XZgKQyRLo7axSEjItxCOiuJ
bNgRJwVLRLBf3/DJfLRjg0PFU1HLV8Y5sELGDCBJdS5l0L5fBUsyt932CONSOsmFMzZIt15cbTqe
ZVZEe7IZ0q07ecRMfmkskhALGgLZJeHX/EkWgrOsMSf17Ym8E4HH+hOjl2s7hPLgGdUrt+KzqY4c
nQRPLjER/s3cf/B99Zjpowle2cTeyCqYUTSaZyu1/sjGSOu7WgMi9wxQUyaAF+RBaZBc0hx47lw3
QcIbFMNep4LQbZqN4ytoPK+LMENHbBMa8iXxsHkIIcybOaeRcnkwWRIblo19Ds9mwsZX6PHYFpK+
L+UliY+D3SCW0SOZh9W9/QslFkFEEFq1sdr6L/Jzl4TzVWM7emzc+g5pSzWvxsFz8APIhxZcFOLD
hLYK5coV2bpAnui6jo+l9L5EeXcvHrxvf931P5NyOszGFA+T7TLzucG3/0/pN/EyMFACiFBIa7F+
OopsKz0A4v1ymEAHAkCQ3WxraOcTHCVZ0lO4O1DmEdCItzgN1MER49RLhzUTrIwMNSyyJYT2xeyb
TYMS+NF+SEcEsygh9DC/ANHtjIaREMuIIvPAQGx9sOtY3jxCvdu0/6JA51HCZaKJIcLjlfRmGI/D
BS5RsDdUFrrT3JzLwsIF0xqx2tzgPQGFBpjrtKXsORqdaWxKMxlw2wUDfscPXmGWND/w+ud0ctgK
enjpniDTxc7DeTSVGv7Rg0sct7QwawV30mD5xUEJM3BbeZW6C1LJXpZa9MbZP5K3USnarulGL1aG
iFhOjw0I4b2IEH6wElTN9KEYIyAUSokXc8vFQZwH4SynsVQQ68EyKln1Xe4u5oCmKGbBVrzDyHP3
uiVKtsnKFpxlujem6egGQ0fwT6ttwQWDC8/Yd/9RBEBPWebwBtH/Vhy8uxA13++nMfdkzmSN8we8
l9IUt2Xq5cnCmZS8JiuebBGiteJO9qWUSf6iYAtZ93yoTwSVO6xZUU3b9JpTlHklJZxg8Igtr8hg
40NFkL0p7X9ub5+rP5BmJJ7XZGTqYDeaF2uJNbrwy6KO5ABwCtmIB7KlNxsNmHTQMv4Ktw2Kr9lF
W32aW36XOg0S+e71f/WlqKJhgcLik/3AY9ZwOklnhGo11+bqsFAklbUakxWUIjozxDYPbEZNhdYS
7xsP6/NCbfcL5iPFRG9JDRo3ysiGZiJMof6+/2k01eYl/RMNJyXWHpr/E1BtyNvkkhFTowQuIRl9
Eo1rCTMvEV5B4FA3UzuNTyLI0wtAfroi5Z4n8x0ZTsrr/9Zh9JKWEKjoya0ES0wAR/ULsm4MKOQm
040VmfmIEHwxTptKWVVg6cs/3w1k0r/cTnV0g1+7QyVKiamqPW3B7iY8hDN4pjJBaCcf1UTSK46q
+iQwUrBCAOXYT0U/DsborNjDKGnBR26GMoa36x42nD/qbMnnQ5PZ+o8pbNYtxZaZ2wXScqUWQv/X
ItzUyNkagi2i/7tbqn5ulLhWm9UHkc6ofJuOHeEdwrZvYlqB7JknPc6c3ZKIeVxMQ4ifyxIftxJh
aCVk/nCZUpMdfbnthhjVtwD5J04VbAm7vxLiFeWF3oI7jh30Y+hBJ5lBPV/jgmnGWHtTQ3O+VvUG
A/4TEo5ckACqY378K9Df6ZimwkH7/tZcKn3YuIA50hWR2hXvqwLrbvukiJa6Tcvp6FI2JjbEsGNq
N1lU/OO8YD6giDo9nazwSkk3KHCe8aslqbNKxikDtziX/I/QpsreitITf7bHrC8t0u2doH1noumX
3fLKzqTtzrrhWqxcIeoSX8Kuu5Jpw+/AJR84ZKRYCJI6N/d2BVFijdiOt5/14c7F5KT7L9hM2DOi
6zBnYrKAQnwsF15ewOt9OyvAdzQgKKl0eP5uRIGK5LaWlZz5UXu5fWEoFxOxA1Wrp/4xD+aAOJPs
v8qoM1RSd+AeyBsavbPiSArt/uV+ggVoMs5ZAm0OOZ2zm5qPGcLzdfDiyT+UONexm7Cv2Y8LD+s8
97DAuqylf6/MVenMZb5pf8jN6l9ZkIUUMIMG7DY5B2JO0dFU9OHDuUgND7tW36VzUDpkBsgdlXWv
GYSUe8jjrdIhOytCEvAIh0V00stb6VkNwQ2c7fOOXat2BmZSxiV5jUF2SqDVn4LlDnuvFLvULaIh
6B9WrxnpvN47iDtrs36yDvvo5nmKfcLvLg1HH8H3xV0dPoq15eCxA9N++qJpWqISer2O6P4Qpkas
2ukV4eniToHHhNjMYJ9dkhI3HLAT6ygPpAHYiSGvMaPt/i2HVcuvWh9yNyOgylK9aqLBY0BcSKbV
2ctncz3GBaaO9yuPNLvbH1tGGavi5wDOT+l1WFHl+iz6j0hh+ihMKrsMJSIXIFrmTe55VSF1wFQQ
xxUAS2h2vsUIKz6MYJWzVlZsT5pnwz9jNxBJp7feM+pjjdelV5ZPmhVUBXCSqv873J4f4EylXq9X
U0Lv1GF8qPjyTr0Aqzx6OZIeDRldocKiGpahH1xDDTPmsTbIH0McijV3U1wTCnEQ4k4qnOgLB9wi
izFluylVHcs8aUFSILnhZgCnOoIN6KKnEDi056QfGk2Mqyz2ti8Y+15X1dRCrT833adapytHD3SD
OcO4Gk4csmPU8z2pAp1j/PnvFOvoAWq/MQZj2Q1OLuZi+WhNGMprd1P9i4sYqNTbgvgw2t3QATOT
ohvko3ICJq61wljdN3Fh5AKsq4sooBTBYnc9q976ywRXWDRyC/i949luTcIomVnM/QzeYiFqt0b2
9mUPNqDvZtQxA0+anrKw0PC/6cV/44UHCs5LMLdLwi9HY/95FOn6eScN0mvEnvNeKih1udSf/pZp
rXopiTikKsovaaVaDcDvOQbXeUVhCO1bHlETJJBHCNYspDPnOL+wd/Ci2gOFjvzYaHGtmzaEaOXz
c55ivQSy9IOmUx/0jKbjwR73tgBDukbBe/yP8Jf+8DoEEDw9lCv8ev8HVH51ft+CbrEU+dXlRXNl
4GOsnHCdoNu0FIjG0DIqcz7PEelh/VvQ/IIYwgULbcaiHylUDIY21ifnrplTUKJBd548lSiSpr6Q
8lrT0txJAQjhI6ACaADJ5wyl0Te9LYF1nQ6moTf2cUwXpL0fWrJSmMZylwCHGOfqGc1R+C9yiGju
bL96i3++v7wf7CDpgmTaNijeTj2NN8Cd7HVz1jmedy5SfeNUwlJQN1CZRwY91FVXzMJU0n4nOJ//
AaZTflQtGSauyQlZOdCMcyI4Xs0mvdsE/HBlERdGr41J5IimouLMKf77tsZj3IK+78B9qN+PO15m
1KGJAHgNBVqBT0zn9OyRhNS4NK0YX9cJ+Vx1ptGo35wBLdV+QyYtecHTw4gHVP00dKMRpFT97tLP
y5LTSDt3RxH6zs+s16oF1db0DHE0YSHKZFvfLlyslB4CM5OBWn8R2VEmZ4hvSz8LHtc1iP/lcMJe
nxj0T4RBbIljmnnGq7d93w1J5gYEaI8ZAVe6B9ahfVWVOu609aPs2r/mYEAwH5TtoU9Ih1dwKLax
UNEYB5ah0QY8DG2L/CahJ+C46NG7etT0ZtTXL9ZNdcgiOHE9TdwfFHYIbg5cO8FMKPJYOS9QXTmO
F0+IPSkRBXanzpaJA/mVbkylkkofMgbIO5/1ff0AprVuGJgsbXLNrIs0uao0PGpaH+wgapqMPxPD
FiaMrdQE5dGFjaXyDITHf1cLwP530GYyxXmJr9m0FVmdSFPepLc6RnBygOTm0IAaCCkJLeIYJ8DM
In4lsxpJnkbm+NcxYOVJdBhWR56Qkuu8MtK7lhvrpmH5mywUD5sXIltfKPpP5ETyn8UvnWm2tYq3
ME4bZjYrL7FCZyKd2BA6zbxGEmkfC5jSZfATMAQtubUe1DI13jNWsWgJLBxeQ87nGows/zYu3zvm
3DI76MT55baf8shm8TUTCnnhUrBFzGf+FjDbfjy6frWvMrey7IPdwCgh4am++FxZBk+um1izS3aU
wiAZTrhxQU1xzjniQqcuFDMmVDcqcU6tqW8QrGnr7tpSpFgs0DYLuBMkM3LHtD7+4pOLQPNp+dj7
bNiAVy7cNV8RB/kMa76H7/4vKUaTlvaGJNBG6d4BpEBoz0aiw6yAEePLYjrbAlC2g8E+1wpD/3/7
xtxGEkBZoZcjuNG14TDrluU068StfRqqcphFi1GW88n98Po2J0E+vLf7MgHDXAss7qMrwa8UWJiW
6YYYVb/zBZS4aoAjw96U0tK1jJFCpqtU1kNVsWmuOofSJWK6YKan7FjH22Gfxy4DxU7Mwxn1iVkY
KeiHyKNvVSTPGnSgbPZ85W1xcUQyL/RJLNqr5xkRuLXMeWU36PpDyDmgLxmO4zQWkC/GtsOnVx5c
uNxPn3+Tlem2b3HXF9bWO1dIcl7LRHh1Bcs3Gh4QsNt7A0BqCkQlVjd7OKGZtLwlFn1brDIcjYoh
kggsRxNeNACb2uLwR+p6mULzQXl/TMz9HPocu52B205a8ldAQ7i6hNg+fncCdf/8b3vEgbAwdNo8
/XaWS2JwTTA85BV9PTfszS+OAeYkpt0SzMv5D+MThhMhLCqAWqYig9q5vqVV6Sg+5AbWWlKKl0yM
vKKra5dS+y/kE8LS7520P6AQ05IjE0JW7DhyTsSa6lJaoYKD697uGRIHriSABBKKjl/gwNB8ao3D
fHTIODgIelaLIAK62LSP87ZFFGRAWvYvL3H1EQJt3s2dmj15zQ4CmtOsOr8Iefl32TgfU0PVZThS
n3X+jpMoDPsNu7ARDW8poGZDflx9LwVIhYNUKAyOveQc7a4EVJRaGLUSzYhCcsgO/r71uNuGY5J4
Sji/GF/3++43HBT9YVUnxqOMUCfh8kAJXpCpD6hO0K+oAE1wmk62gJ+e+JaPWNFDb72bLkURCwJK
VL8N4bmCkl8wzSqdraWS7gMLNQoCX8ob3IYqR6tS4T6Xi8K0WFV/TPo/GzgUVHt78KTqaIZoPyaG
D60g6OBMHvqltwbb0ZGUQzhVFuFzxd2WRLZWMo4yiP4t1w5hEheauJmi59u19Jf67KxWhIX1R1N9
KMdsm2P6zuG3xYXvV3ECII0NYXIvqSIrfmwMGgL98okfQzrMUUf5ngskzTA7vD+wnd8CD2Mxo6DJ
kMzdEKcDZUGg05UIPyFwuYxFOrGU4sAwHorFfhoocbybSdF61vlgAvrfe6trJGyJaE+vHwOGIz3A
tXnM+kBCqJ4YsAi/irayUi9JNvQq+4aMSz1an5SXVll+bvy6ZvpxgnWPzBVPX3vHjfQhUjK2wvbF
CLUzZELdtrr2LVUYskDwnL+MUjZWg5XjJIF2qxsuEZKMKGDAwcx7Pr+Y+ZMv7QOjwrRjRjMfpXUp
gyzYMxA4DV5mhFQ5PLKrVMgfmxcXdAumqhfaxy/Yoc5yRyrXTlPkR41XcXXF0InPHbV45TxN9K+D
QSPBQbn4XxOJB+38cLYIU27SaVHJ4sX0Uat9/dMjxFSiVSdQXOMQXc9MZfy4AFfPJyRMBsGeePBo
F5AdgWtDVyhcVkn8floxu10Sx1YY2sRhRGDjV7Aje6T3tqTG73rMyyPXEz9Sp+LyPDqYdhyES3d6
f3CK1P4AcCFhfYceW4j+htVU3YD313vCKaCbr748bL7Puj4DrlBb2OxpS+OmDVfjBfgEhgBStckO
XWsXwy4DHEume7oFZPzY9myoYiEmwa8wyHh2w5cjfEiWkxLGKHD329OVWNgG7bE+tsmClxmkY7Uj
vL61v6hMKJkbInaI4e4F2wrn4MYb26tzjwZHzC/cWtMTMchb/IT336ox5H2tZWmCT156ugfsdO8Y
ll+zpgBtIVZQfFzoVfj4EIMtkhqpqJNtpqYIpBKhexX5Z6NrfOR9F55hMVZ3m9tdKHMyjLNahdqI
kEZ/JBAd8xqxQs02N+SEqoKwfwaMdcgh78iyMeWAIIvA/ogB82fbpZ7jtO82Gwmxudn30IcH0mpS
Qo7Z7hRNPyIR2rNulz13no1JptsTaGdP01hyqvxqb58sreYu77stSn8uAWzVuEXZWpi8jnITAxef
cbRsKateFudFlLX4c0v/2y4KPF7yxI7MmaV0kHOjgTW0pZHMgBpziaUyNDo1WcRaHJVtZQkv1Tnt
Y6QPrkPYLB0zQrNkOF89sr9U40PlU18oCb2bGtY1Xh7tUfMG9mukNsbxot4OHff6DtJnEbykmKn9
BOIZaKOftWgsIvgV1fgeBVEF0CCj34tKhlczjdLZz5LE4vpB/Dyk/KS3T2pByhxRCaUPcFjOktI7
cTs06RYTkYvctweTFrBj2/nOMPxKDCPC2UNwucFgpwNG4dauRKJ2pXetdaCh4DO6qmjnLcDNkWK6
4y8+EnJ9EEIJq2LlwYYRDivNzkzGGD8DOfwl+jcN6qJELdFTbYq6GT7e4EgkX5osLczgV5npaoCW
AoJSOX16G5/Oc68DPyR1Dq8MVCNQQNT0CeTqGEycmhcZHzW5bwVE6E6nfVFiduffEB4B3X1hKlQ0
iFKJ0sd6wkxf4SkUf2k2LJUXVUZRKb4GEJNcjWU609EAMTc2uB4xD4IV+gJpZAgyoB4nYvfPe0Xk
vrl/ln3++eeukdbNegYe4eqnZPL5pLy3keaTjuBbFVjXx9wIDxs0fWjy9fenbOLdAsm/5E6MjVX7
UWShB8/epaKsJXcRCVtZUHOwRY5AK0+eG1WrlAkto6fr2qu2UjoTXTTDIPjSpAbnjycTqh4EHxQa
CAovK8jpM9B2pHhMAJVQ4wmuc78JagNnEQFWhRkCMn9uRaGpo0BobnoQjVHRqfAFC2yYqWyvu+Pw
4Rrsd+ywe8H83fxdRB+O98ZGxyvFqv5R+tXTfiNgAVc+/YPneXCOfGddevNexAF8gPWBrJk3zkhx
W1BFr++bl5zZW7f4sAy/Vbucmip+dbdS+1lAyZX+r/t2m5VPW40QE6yvnIo8h/iMBRQmap1A3fQA
CV81ZBm10wbuZD6zW95CdsgPxE8Y0SBSJL/vazPYV6v6CYJAHUXJAMyxBZ1RsK/7aFZojGG1wTW/
QvjDK972ZgpPosmYaHesES2UzBk60cJ7eKRLhmRAytGgJetiKoqJG7n81AwyPGwkvh4Wsvj+w4Gu
5N2IK81tnmjJ826BRcipBbqR5A25bwaA2SEj1w/KUAjzK2x5X0gXtzCSEZm5owss1O5b5JQ+i+hg
ux3U1v+qW/YtIlvBcn9FfQ3idcu0XBntxF4uAoefsRVOTplS0bHbmhHJsJEVX7lOQMPJOKRU5x23
0fGwdM5q8z4elI0xOX3HVD6sSMwGSg/54cl0YfpL+kv8kEyHnF84d00Y6QV0FH7ZpmL9YS12KUms
mMAc2PFHT/JKrwiBgeCZjyabrArwrSV6dhlIY2cEsx66FP7CpfFwBLJeHjc1bygL+aLptufEKuBE
Ff/achhDd1AHKvNvquIzcZ7AgowTpBqnKcoRI+0invfNXePTynccfPs4X7qjonO9NRGyLZsSENMv
5R9iz+doL/33cJMQUwr7Bpt7VhyhmEKEKk7deBPf//f2xoI/Etm9l34GfY/znktQisO/ADPCnBC0
IRWr6Gl87SHia2OOtn/aXAUz9rltOuR47+k2fbp60Wa7Nw/ch9w9xlHVOK53pS3Titqsq1cVYDCb
2JFZkEeHSa/5bAxag4qhgpLXJsqJe/xCPXuCppOTsMg95xOUgS7OZiCmIKNVRXBldkY2uawjZcod
AHFAMsmQ5HNZOUxOPZTxgZUrHnvSbSrctxHW4TZQ4P8YmsAUS7y77lA+ZFu7FRqQxiZH5caK4agR
WhXFHRimXIe1aYYcRz7wGTqyDeNZF0vkv8ABns/d+k61cQ+81/J12q76JhjQeySQPOBxuFZoLJAm
D2vsWQw1tONXsAobR5qVMW0X9aOoPZ53WXmN7MP/rg9yYvL9SHC0qVugh3z3qtCh9+cGL8iGsrU1
LZWvSodX9qCerGl1AiYyQu4kQCAnQV8wnFdcCwmOVWeR+LsNtT8rQgPdU8aQgDPbcJI1v4OdchlR
++msZ5nVNHMOo06hRFz+TkpeAeBnGw7Vb69n+pltX+x9Oz3eR+apce379Gm9jL4LRDqks+yU2OjU
av5RtWpMMK8jY8SQSDn9vB+T9GHjCYz7dEUBO4dTS6amq7LSuIru6SPUlhx2Ay/WnTiYKBMvVE+4
L3K0C6y+tX73nib0kFtC3A8SxebMe/EVyzp07GBCvXZvRCgUAJZ2MzwvHVeI4Xq2bopy5uems7Lk
zTO0n4QJCP38h67587JX3Ssy4W8IqHyWw0KJn8T0sONVDSXV9ZVAiFcAaPsFzs4C0H5mz/LSPFHN
XT1FOg7dBRk81L0LstEZo4KS65+Zx1FW+Tl0cYGAMbvtM7/Q2TYNDOUjjRSSAJBT/a+3EyRCktlP
zKxk98sPe/gt/L8xcqw/6QXiLdG6hmXUcsAgFHDZN6ETAJ7bZKPyIQZzFsATe4ZT/FD1jWG7nVe8
FqGj/cM/dhNrZcWvgUf8LdAjoTfGTfrwOqskPpVh/2+RqgrjRwm4ATknlYeKPxKcDDrRXDqLHwAi
NBl0A7xOnuj8uGeQv7tJB5yiQVAt/XRhnF0hrYegi0/f/99lfY2J25AjzGbjMVwPufIfOf2FLJh7
HCNue37MO6BzWdb8ejQPmo4fk90+rxL8vHAqjY7XnkH8YfR2M/aZdO7eFUdFbUcLCX0D7KqPLPhW
AVgXnwfqPwxMZmERCIqKNixBkcKQmsMTvpSDZydxInTulkrK4Z4Nq6ZHkpP6VDNK2rCPjxuHkoWT
PBZpcfrUzYlFpy+PcfHQxIh9lavgPQRYSigALTavN9uNB/GLgmc9650JcrBkYObQs5QavI+Ftd2/
Yl8uJIFg3Yez4irbO5bkqi/d5MG4OfXnt6aP6wix+ue6d1leSU0E6zro8+knabtoRBKwdpg/2u5c
NGLPv7Eqde4ohKr3NJlVOoXRoccN9JrZVlwSuqhSA2+qMnmPyw9YLhToCJyUPQvVyWkV+uEJBRDr
gMfHGNQdpZCFlg+X50eKwODluZRyq1mUKw40SrQOvNCq8GHm4M6NbIib8J3cPzkhyWqaMOiqFq78
oiWWdN/cnDQDycB6F9Vz2GzOqMqdSiJhxjVu37DOnVrjn1EnYTNhQpgOWrBgSF0DBcQfFrpDPRno
57y5dyWydt2BseNEArmPuT9dEcgD/N5OSf6IFXqHq+pKCVds78Xv44o+74tWnMGSUSs4pAjGyCJt
Vx7K93txiCPfqIgw+OS1DQwEY9xHEBSsLfrtoVMcBPl5reyM8iXbvZL99tBbzXBb/EGtioQ/CRSA
FIvCjHXFcRVREMUfQhLZC6d0+fYoBHupw63NxQ4PURvf/joVZTGmbXhCEbdWTeMqw+xD6KM+1gbI
HBDg6JJUwWgZT3psHplCiNQn/ubxQpfp331GdMcnhEO1IQ8X2o8EMKNLQr0MTG1ELwiBBFf6PMwN
qVJIuCXfWxyWRZstgTk+S5/K444eTvzQNrcD3135eNkac0uK0tQHNQW/FgzssQjtMdVNFuN2+0dY
5iWsz4LMPZWVUuQltUU6EFahHpSN1sMImk3kwB1/3Rr1w5vR3dPNr4wTvlb+aACsBy6BATcgQqJ9
mZAfRnCPdWA/wZzsd4jG5q0Quspz3KpQ6fCpal/yUOqwVM+lR4o+0zScMaksQg7ooKxgAnxmbOkO
BmHs9uRJpo6Rj3BLf5snDkZYuYnCfGOi6HVyvrhZpYH8w5gGPTgE5/XgvUZebYuP/fxq+Iy23vBv
0DHgFfb5YUfRm3Z6RDklBF3RTBE6ggZhFOKflZEsRagfEKTH0sh7iwoTv5nDY5g8aYvNGehOwcgQ
d6Usr9U7k2W6s5ZBn9UrwFQrv56VPJe3MncLK9je9G1diSrVSh9kkYjxj0NPrbR8lEYy7JnkziKd
35HeqBbBox47JYIeS/rsdyOJL4oM3G2lbAtYzhTGIz4q6XEeqgYqUK0fd/jEtomWH0pSAFJYXEbk
97uW2Tq00LgfcE9nP7fO7ltPz6lm6FoT1HjABzVZf+GglTfLGE8eBkgTFoip8oyhM9G10F4Sknjp
Sugy7Q8H5WoQYWazo00Cq+TmGglkpYygA/880tRN9DVsLItJ9DoIsUHey3jpwAX4lkXPXq9SDnRg
EBV74gO5RC7hFSgjqyur8cwUpyAzSjkSdbtMYtLxRCc+kJ3GnV4udSN/79wxfWXWPNeD2+T7x2Iv
Al/k3jsbF2yuhNtCzm4xxqge0cuqQMITB3c/NcCZ1DK14seMQEeLp1Yd599RF/ZK1hAa3OYJqqs9
D39nHNCUfJK2RbbFkvYU2/JYzXrpZUd1bptHvFPjKly0GT/CvtX0Ecn9FBdAavlO0uIjWs7HWyK5
XDcrcl9VAq0Od6PU/LfIBz8yr7jUro9g3kkPstH4ae8GQocTb+CGIIQZatJ50oMJFxBiJtKA5l82
prEqbDDuyB49U+zkSZX8Yq105Jn/InaDv7+qkAzcWBGYv59FyfMvuolnoLWFbYh/Sv+z7pw8eMSg
vSAevIDYWj5N5y9135SzMz1DXqkkY7pm5XokSusm7n6n9rYtrHR4GIGGiMgoap0rOYf+KDPd6UMt
3CdMny/2/dsXAa+NQVTNk+X2nIOQWNZrIua6F21LdoIfmO7Ha3fYYW77gmFyo8VyHd/6yKHdIo46
irfpR23fUatGmI+uDDGMGuIbUM4VOHjvUEajslTIlW4LexWgei7PmMEAKr4Zg7gpYS1j2enBD/4f
v26tCuFlBvifNkRfwZmc5EqFAH5uvhO1zcxFB3a5Rpa5bQiiyCif8udx6HIX78lakTKclOXoxRWi
/JknUUlIrtICscjn66umlAuX7IMqCucQEUizSR+7AkNN4jLukEQUXMaGDipD4RuTp/Hed37FxZDO
cgkIE6SXdamkPW+fNkWwWZpxO8LEEQyo+AqMNyKpswS6Iy5sWi7fschUwHT+2/+EYnZssz0+LpEU
3hqGxxgjFbAiPWzzxGtJ0iN/tQvyI9YEBJqWksA+vJKKyK+5UIAA9Sm6yxaqaph+gprWZNPEXiU/
sF9tjzdRP8apNA+a/cJt9+h/3VoY85NY4hmnTM+cu5+117Vnfcehy3JEJqT1Fn5YTDK6Ujc8JcJg
7U+8PJlQgy+0AEo5d5kg18iCD3xWE/8R6WXNwAznc02OCKIwZheW9U+0fWjQ7la7I+5LsxIWjCAz
k9g/d2QvKmfrSQDLH6oOGN5bAKPIW8mZf+7HQempKRb4RBGDHHvMhf2l4kJ73FE3laO7DBq4mXfH
L1MKoM6/gUtlk9tDLf/t8/GCr+14ajTZ6k7zDNy6U2zGu8uRrnfPtnylQB/Xsi9gyE+ltkzgQMdW
OSO26SswgqSfcdq43x+XyY++QWAK34EfLBmHi9QHEAuNPjQiLToFt0B5wW1kXp2z1HTlmhu8HZZK
iexvsPLEYIVEDbQV+TXGNVbBfiFT6KCT0bRBm7uxCf1v0rrRdU+7Y00M7YVHaIRt9MCEMC1/ImNY
sz5RH0XQcFf666NucH3nP1BKahnk/fltuPvuXmC8TSe6lEfuhwJJLKg6U6qiRITitcUBHgI4OWoS
hFhs90PYf7J3HNjS82oMmbmMSX0FfOMCm32E4YZRiRZc8wznLAxklEjkcmEjuGh2cm27iUWFwS66
k63+sgdofm84f+jl1wYck2AzmpWL7+6gc0zkBFoCtdgwpQMWJPzOcyLXFcqDzV7UOx1J8/8wpcFe
MScH2O++n2Eh1BLQ8aaR65YORMt4iDDSjSfzEtU+/1hJQvTflXb1AhdIUvziX64E4SPHDQqR+5ks
NqSzDAW/oys8h6gz3btMxq4DCS8Jh5ykbgs+vJniMCd3Gag03KsOLinK/eHa9xBWyWJ4qZP/P5Hl
peoOYtBxQkvxA92z8OMquBIK6Uv/QVcGBicfpAWStLLX4neB8kaiFw5UedR1f7oN5lDOKNuMRtO+
QUgm0NMSHI/4V4058gmTQToP5pA0CKNyvjd2rr52FqVtxEG+uEToYoijXLXDQXq5j12w/eqrn1Jm
wCPDYJUIr4LepQSc32k/MhzXaCL5m8C2G4o5X3yK5TJojCGexEkN4WCCO+DtYqdMAZTSmpjzox3u
8TJDVyxNQFCNEoOQUzun2l/whImPFaWMuefVsriCQxGB4+4n7XlozRx9ZbRuZfQCh7uNdkZC1UYV
h9xPu6Va6imQpilkOPr4ugDtAy3woA/mEEFu2SIq8V9uCchoNCmteFWVJCoeocXbwwX2h1vRIlLg
NHzp8YYLVB8Fbe4B6SKiNV2CdbIScXXdE7zwtR0SrqYG5Jip4cOeuJNlKNko9hUFL+8xn/g/kbxP
fkxAhyNguIWzwsFElvWQVFYiBwFFiwMETtAL19A/2/FMuHdMnd4kNLvF1FY8gq9QAcPzQ9wy8sGy
30DFHTeUH+VtBqgLgvH7Rwj2bKHo0vXfE/0BOLrwm9B80H7TTE8xMFKskJhcJNsrnxwFGq0PXPDL
QqeY5C9O5g38wqlRXEa6Wu2hhWyskK+bcvooEN8ICme8xxUL23Ca72vcpu6TI2QwiekCeV7PhWGL
DU+gEsFEUm0/pZ6BlRMkgPBAHRH4PM5wsQHW8vzKnHKBzt56LVFqWiPuLMV9mVFp+EkjZd6aGLvc
9InwD08d4gXwGQYgamdKTqOEhY6/fbHthItkvm+iH9DX0yRwVcnOuIktuFPBt8nXj/Z38pp9yw92
HwaXXvC6VY3i7RoOVySJFI7AWNb81URpJ8aeIja0R2kj9xUC2XH2Z4Baiq0Pafb7nRyECYY7hWsD
kvBYa0oCI3fMLzG4GCPxfcvR1EcA09XuAZrSC+KxAlUBmQBlFL9IpOAJzLzlvCto8qGcF2QfQuVD
c3d3l6QhHM9P0w4QNZ2QU5Af1ddJkPOpHSX61QF93fPN8lx+2H3hF1GHSzVGlM9Zk5A5+ITO4mqo
xwQkVJ9be+ZiN7hJN52M3+6+G7Anb5LJWOKtnFiMp1e6TILDDgE4iL78ZlQ17EXF5nL2zTfQESmp
EoIHR8+z5/mvryFPcB4PZL3VM2UhSCBDbD/vgR2gd/2gnCXMIcXR0n8eaf3y8azXGd6E9VK2M2Ah
Ob1dt9c3ro7NQzQb1iJfzzn6G9s2SmUlYEn/84hnfqHXcJVB1RovRTJwPzRQsYrh9ax4sDpczL8R
B7eSUWloKpfJ3Fl4mjg0RBBOryFCWuvzQgpPuA+nW7GpNBJW4XUwsfzpWmeHWMKAYCsDm3XyYB+U
cHW/B6nTeYTbIK2Uibq9XEKLLl2RNwSzpqEJNWcfyXM6oMaSqkZLoWOZ53+T2CW6L/VAOBN3llzY
qXIKHqnG9XF8E1riI4jyXQP61Fo1J5w9rxBydnU0e6KsyFg4EzXZ6V8gKgXuXXEXzsHirzq0n6WA
6QBc7TFBrb/LwXFql0+GHzSDJg1sUXLe/IGpCa2sB1OY6vGaRrMZCCwSUJnjoM0RQJXt/LLBppXO
Ck2LrpsJGzC0PM8uYUsBcDMjcyS00PNrj1xxqfMpk+zBCdxG4EEyRGv07cCPXb1NAYUOIF7ATBFb
P8onxWVZl4x5LHkIjWAy/m0QEQtuFyRevujxzQWhFsl6bexcazsq41/oxBnDEH1alkwreg4vmP0q
EibED9nqBJ4mojG7b1dtZsUX8oZKxXVV7M2KUy4rfBSDPjggS6Lx+uB1XqubCansSGKP1RBrhvl3
tNH0a+NyuzUGJOIjhWtouaoGxCSD4L2PgvA89MYqZ0y2aw33G2QvfkbW4jB+2ugfz3t2TbdeMXKf
LWicUnVarQMmi4dXFAGieGxppQcb2lRPg4hGAY8BujVI1CaC6wnNZ2l2vB67krZhD3sn9Qr9AhZy
tvs6Jao1VDy4R9lj0ATtq+wS72Thot6LLlILepyy2yhXiFzjauLMJkz+h8BFArpoAfJH87YEWH3Z
VWZI+AujC8jlUuT8M+/BrvOeDdrFfFC7ub489gnvzFoq5YjaVh70Piic5yX1kgEoR8UkMadnnwkM
ASUlBMTUiLPK+nD0y5U7BAsS9x2EkIyavCD2zV7gmYOcVMaoBKpi3z7gN87MmtykOdGoZkJmZ1r2
9CumK3Hqc/5wGH9jvcRnNzJ0KVZoIq830HnMn95MyZD6+sszPA301Nc/4fQYzBK6qNKQe0IODsNA
NQWVKu4KkH7U9PXjbnu2pgOVmfNVWB8iKN6og8dHYaGNz8TV6yq8p6wm7UvufECeIxyk71yzhSL9
BjVe5eGs+cJs9P/+Cck2/3T3iOh5pXFsIy3SANczqQvvEYVaRD5oc7UwF0nD5cEEB8ui1Ec6L0R2
9gntSP/ddnoFLuKL2pKjErl2j2DVwOD9LqBXvy915iMLloM1Iz8tg1nYuWa0qHA9An/YCspiMUjL
x8vxYa7gTJPHxBsn7jZSBPr7RAC7aSOsgpDX5cQIDlSAigI3bJPsQL9NVV//A38gX0AzAckIB5hM
7E9xl/cSUoC7vx4BC4KROUBS1cx9IFh7BCjGVDIJCz3kfapSsWxxLnYuhyXU03/sOXxo3B3B92T7
sDPdW6kk+WptnYyCu9cme3JlGmvxJW8CuoGdQUJzFAA3T2KGEJ3w+2JReL6+VSreWHmFEkI4jBnF
7Lye0ob8DKsEU1HR4evBE6XDlH5r2uFpfebj3OdPw+JH3H5Jq8VTE7LpC6hgKQ34mrQ3jvU6Cwo4
LlaUThgrJ4s/7xL8MzstMImYMm3pGy/mO5DJAdxj57gYdKkDBjvACK5GqzvCE0rECVwEkP31pmLA
m/pRnQ3dCuERbqPi7urm5l2anIiZNzDH4siPZJRkH9xL0ggS9N7bZLbzySfAz0oCHeoDQZCrLC9u
Q3Q2OJbx9/ezuLg4BZMfs6mrH0dCngeolx085aI2q2e2GPZyR1LrrOwlinWPYgTgKtyCRm+Riood
w18zAZVTlyfZFF6xG6wrcMLQf/pAhBuk4spP+KS7BbO+tZ4npzrSdZlV8PvJVcLAm557a90sOjPh
J4lfYLJSINaO7bAEP8nId+U0tID73r56iSQb1q9vi6qryQ5RRQO3jd/FUCY4iC+8lnJbCv0HLP53
I1PpcDk6rGlZgBxyAgvUJ2NJNeQrmhuSUSkEOsWm5IBNbnN28xqZ2Q3VIVep3U45LbxyjhgBE3m4
sNzHzxxGbLODVtz64o9RG+/Va63Pwbq5ZqiA+DmNE+K58ytJTN2+qPCu6zPjRNtDnkRGh+/3Si2W
mEwrP8ugnCEhLQI80wU0VbFQBg2XOtBm7A5wJybJIc615FjFXv9xVKkgGf72QndBG0dfM300MS7v
rTRJwWPrkpXNa1HjPSsRULnc3tw47TLVOjPSsXmu+AEfYlFwrLRRWPbW2x0E0avIiSYS8Ix1mytZ
fBrlGulUgWZ0gCrsQrvn8Xx5sgsDZpmcU7q849sNUhlXKCapPTsWJ/UHQIpLoWTb6PKRJAhP7qmK
XBjtSKzuaJ9kPEIXmtUZSeaURDbzUbycBa+b3F0AwKoGWWiyCUTcnSSNx4yiQXG9Fw6whTUadgPk
QTDwj52SdRGAMynvrlIpn55b85k2bFA+NNvQmNb0sj5i+7wEi2egNXy/o1AQjNg8KKZfkrvJsFE5
jLwObhqWWd/GAgqTrrrCBaXtrf77zWCvw7BtcInX/66dHUYtciXd3bgeLSz9gSAEseJqPyGTouyl
Qz9AcuhuVkPypX5S+3saOW7eR2TjUcZs0LHI4VGElFwOC9+k5W/+tIIB9lIqcWku9kKTDN1lPtld
gKKWpjWQ/3bEzlpsvjkFGrw8X3jJbN176+5QzYwFFZoZCdebC+vykyKZfC/onpm/J2ecf8PQH3SV
hO6F+Xo5dMLPv6HRfKu8xtijx3S8r3+FtN9YxGH03WgnbLKmeF6tn2n9g4oZCmYfpooP1EvQYQwP
4Ad5jRTz3tC8tnThuDpsbF/o1uL3Qx4/blJ11DhfXuqYze0pXk/mv7ceusTKv3LdhWm58HwVkozM
X6ST8yV/SFn2EeM/O/fF7CDWoIbOtkKqXNFhRvtfIrChQkeRJ9t2PQqtUgDT13218Uih+/N+aQb9
zb4wj8vhr0zX31JJRBps69WJCclliQplQ5CGBa4B8EEhmuq4nMJSQ0nlQAyvODQOH6MWNK/43W/t
PQmv82p8Sw4CvooGRzWDd3NhiJIdwvcBNRY5i5X2OUdW2IeO5YmkV1kjghpKcHzoF3CuUdzxVfPL
i0Fhy9tGKDPpH0UylZknQmrbQ7JuZxAt4KCXIm9jzjb8fckR79X2uYhJzGDcFJxEHR6E8HNAH1Wp
ImAiwK2iUiDlxrESZIG81DQUzSEvGZH4c/PuC5fkqmIb9IIRWOUTgmTy7T8206hQl6R4ecYE50eT
Oeg/fz2s7rA5bme8geLsI2krWV1ohRTYTXZP1xsh3JEigQ6yBI+bPEIBiyN+h3JeakRSxwyTVTjp
C4A8Iy2BR8Dp/MXsp9vzG17sq6TK9wQwiFJPtl8Pndp+oLTl5EGztKnhHYLtzy/QSD+E/t2YZYOc
lZgOXxXOERs6/ZI4fiVdzF9xhkPThaCRag5IYXj9YiLbmVOIiPCNsfp9O4RPnCxHWQj26qCgmuS3
2MT3Bc2BiPxY32t8IfkgCL3B5AN/2yYr9ObaMptKcSlZWiagbKeRqTHWvXDHRJOM94HcyNQ9xsP0
xNfItYlIJUFGlV88reSlLRiorseNkXxoNaVC68CZIFDmG0aG7esSeCFi0YF+27M+0DbqaHQjZ/Me
h7iB3Syv3gEXrIOfHT/uWMd8W05V54sIvSTkNvMBSAhhFSMnBkzcp/yWW4TAYEiBCIJgL4KFrx0b
JSWCqjIR44etGzOFXrC9mCVyL6l1xaBT4Tro+H9IXgohHfaumdKXtyJmix8xdEIt3vGVw2PO+r7G
yrDCSfKArsW67v6zbOr9qUSgNNlgh70KyGRcSSch3RMmPlOOfKFm44sZLeSJUVYo7H1q6WR2Ghml
3iMwg+TWxFL8cIwrw1UWS6ud9HgESBRVdZIye519fXDvhwxVk4dEU+bGpK2+LBa0/LYXZSyWBRhv
MrwqjcVba6GvmAOXbGk4k9fa0QL36txaZFOV9c9RAGDQ3QkEvGbk+dxD2aZ/SlsZcMHBnEeWFA4M
GwwAe4sjz7V+NrGuz/Me2qcsoPJw3Q2gfJaWGt7d1tfo3o53AbIh+MHTY5/GY7ROEjjoLPH3OgnN
QZfu41uLg1r6PJXaegONnr0OY3ZGfm3iEMAZ0i/MqrLSFEQbIDrI/bmNENnf0MX/vqBPWAwUXpib
b3426/dI6Bq6c0NzLC9qraO+tVVW+Y53e1V1suHJRao0JC/kp/a9h/7UWUf/NXcHjEIEeTeKt4Ay
mZ7yumr6OrB2+/Lfd14P2t8QqbJsf+L4rJMlrgtPNCaeabLTPb2pF5BjcyHR1Qjzo+6K9z5UJfM8
KHkpf+4e52SaljfdbuIV/Zsor5eZ51/PFRekr0ZqrzroNa9YQUMykHebhmSzhplcZq8fxmlZfyMo
PmDj3paB9Y6m1qIEoATD7xkz9E7m6PS+8DOhLnvefp+Ccpxuv/46uoAIyxFmVCxKFU7Xt6M3pZyC
YMs+tNV0Jg6Q5zzniqgnC1dKguPJDpBTmNmpDtG0iTqer0tVFxoj0JDRyOV9Iitbsw058aJRhj7m
J1jV4Hy4M+NcqXNrx1ASvGcVUuGwgCjY720goF3A4vlp6BvoN31BhrPgJVVxGF6ACDNcgEoQvlQ/
BgzgIjYt+yUTFrRw9tksDN0qEPl2WkS/qqj0TegjOcXJWGCQdajrL4JZi+QUd+3vJia4/4im1NcP
cDuWIKOZEmhKizDt7d+RWwS/DP28YxpJ/tgbtXyeKMgXl+vaQ1g9m2q94MrE0b4A7BaKRv3jEGUl
WL5Qe7svwjokIGMal4z6sEH5hDSBqPy4W4agD0h8zmkQgBx/L3vKwIGyz7+xiMpSSheDACe5Xq8H
nQOy+8qFmulMQ4cr4KSorb1Cttz5IpexzOEiCwr8iotJuoMWRTvIcqG6mvXkse2AQ03p9pSzsO3z
LUTD/TDc5bibCsQ/mpnTZjmX8YhoGpN3no2Hbw5NVOuhVLIQ1eHR6HAw8FvoSUiaCDOKdMO+81o0
qWLMztLWuCmbNp4iDbbDIcUS9sc8Pjm5MYVFlSJYgra07PsocuWQkX4rvS4jyEJDgS3xgnU5B42L
HrWGV++nSh2z/3dH59XULZCX5zT3FqzJ5Z7X95lWAeuTKps/44g7siBzkjzUBVZ94WBez0W55KPV
YGOdhfO+JLiWOIARBu/f+lY3wAvhHPK9F0kRdxUgbQGZopmKWlWhSXEu6z/5dWBnALWPerz8HUhi
lwG+FVyMTazg5ibF+90/SJMS9E3wX23PiN3YqVlc1DObdtfh0WPVtYp8aFCAD0EZjGLUINthrS5e
b7VlgahiDYTC/x2nmgzXHtLKWhAXnf1U221Rq0wPEpGlVa/YcYnX6BE9GymhagpWuurNidFyva6T
qF9SPFXltr+QbICu+Tp1jCEbmNZFyDf7PH2vSNFuuhTVDMe9uV469+Mcn/OXqGEB+TiX3NOZvUIv
tTr5Ft1lVaJ6vKVryLecOliO2WuTIK/aNgiAWADSbi2gFiBNCGw4Rdu6jZCjpgXffGRjmkouc7Q2
yrJEczgdwsH7ohgL7Po/9E6atkKlkDp/H9LwMY841bAu3lh4PiDVIr7+3S/lh8W0X8QpdmP4AZ56
QabBdtrTVG14EyjRQ08GHasSZ5Cu0iSR3v6NKcuVoaJkBxXMhW20lDj4sMuWa6TQ2bEWni5g0A0r
ecOYtE9e2jCQkKjcon8lkO8jvZu0Fb0z+LINYnlscDhuYpjGPzr5SuBy8PHZf5+3N9PbqgL//wxv
M2ZCAnq6xkmz9jMa2TnRTOL3DODE/AyqzjSU8OUS8xncTuzCDw0AhrI9zFCouRB8dMnXFg0egzXT
rfVA8UrwFqL7PROTbTOnXIIBZbw6X1i1ruyUrQh4XCSjUsy1dgMt+1NcT9u65GEG6a43PAetdwKZ
5Prw30PpNXH22ynwge8FDIuJPoWanl3QwVdiK8uNqfczKgKx0B/V+tUlSsJpYixrlnCHR2kr4+yu
RoDhMNJiRWRYrwI4yHhf9+nlx2y0vutbR2xnR74f4jSJkrkASfYApR0mtOJ/i6kedhZaaZtLr9n1
+qRv87bds7s5doghbS8Hr9FguzWx0APIXoDrM0OcDvpj36AFr7nWz8w4/qJKXCwXp+QYDGxtgcFA
uCI6xRSD16kdo2ydVZGKEsqlDPrm1EMhCJtoHv5GIGyWGWv0ZPEkdiFofvEfrfGm2T7IsR5IAIvl
LpcT5zj0IWTmhH3kh9wOGZfJaM3//rbG0LbIVQQxhudN6hZSIpId1z1eaKRNaOHiDX/k4kJswoGb
PFgV4qXec2szWCrXda5YSObj2Jlx3DrBIZ+vFu/Kug7BIUHlAZu/2lKW+8ceLhcjVkcMlJD0h4hu
aWBju5bV+fjxwUI82syL/ib0sTi5R/xOQiPxHN1TcjHaZzPIhx/yV3PO8XVtQuxLeimeal2pwCUj
irZoAMP7zTEKhHvg7EGy72fnt3E31P0eSwMjLJCO2Sdq/BXvcS9RwuDo4GoRQWpk+1iK+reBXUev
YSexT09AdOGflhh8OuF1wplyC1sDeu99sIH5E4HrkDHMW5iYJaE585NA8t2P1mfIDTf77EsUovtS
qxWo98yL1N6QqcYyyxJI/m5yRdmUBQmH/QXtdS7tt8EPKcxusRmrKb+L2FmxRYIFzY3QpQvKLSn8
Fya8oWBnP9kPRSCOluIeUFoWamtccPFzXTRzxXXmDejaf15KDvZk1QCTQcOML9i/7kH3DIqItbft
etR1PnbwBuzH7h/z/F8j/1wVqzeSXYllxzEZR1VPpwDBECUW8U6mG1mn3CZzLFTdPqwcTt1dI7Jy
isrwFYQZQfFP2EDxFXh5rQwbxl1k+SMnPIqOYrORgX2bv0lvQIaE69tSwdCWecK46JRH1xhFTsO0
ppseYhZG+z9txEyZ5RJ2LzRWe+v4U1DwSGNiGidrbwb376C74A/LTzWV2OpsYpDdFR26A0xMFkrb
yvpUwTrLPfGqeXXTuZQo/DqtdOKMUJclDf9TG+C3K7Xw/eHU/P2fg7RJKjqVMMDZZJCVcd/K192G
TSGQjwFi1puiURPX+1BGrx2MOtU9NwNXST2UUzo5PUAb0B6Drpjjw1X0mplxOiyHzwNzMTGTkG0X
pVeZ5odpF54DkKhoy6weNMa2yI2PN079lZ5q2EnIJ1j4hrybmXmjjpA64gWMomtbUML7Ipxwd2hn
n8DbNCDlKg9CrP29PKSAKxMnBh1FykDQRd728RcxPObUe623dPGVHKMkepakTzybn4o/uyWz3v/m
o17j4i0AcjGogPmcKvnv0GCEn2nKI56ytqxARXit2VCLiYzsp1WfWFyDvA3H2ODMLdMSicxDmB3/
V10UdueVWKk3+7I1NBEImmtNqZ0e8X5ckXv4YxPI25CRtTIUyJdwOPqVtjxHyuOJ2chNhdy+Jcgv
PRvUWnNvmXTcqdKZzf3xgGjJnUUzOLkIzqOqEJeq+DmdrdNigFEjLUXdDsuH99CffEGv081BX0IJ
29obeQF+jEgC6/dvEA/mjCYnKmpnQO3cVag5Up+nQq1MIaEluDT4GBr2lmJHPw/eV9Ksu89QPvSt
1JBNt6CIcTRGVZxxpVAYwI/QbvFZ32KKIsYGBrdNBLfftbHe1AOKItPzRLMARFPdjO3b+KIaX+Kx
r6/6BYgZCB3TkHxHum3dgUONhK60HOj32a94zhTBy4scSKk2/XD5W1Hda5Qe5TXBYGg7ojZzyv03
+cZyweTBKNaZyCeV9qolqIX8/bxz8PB1/TUmvfREWDLY3m2WplACn2+7oUXxuj0DB2srFY7IvaQs
Af+18ezv+tC0cZPXu+7rKHpsDomYBo/VCNVx6VR1QAPl7F9DiIea8bSOx2Oc/3ihcOcM4CcFtpp8
wsFaC94g0usBJ+coMxrMhKCuuCYfPR5UeueIRdXFal09Hc6o95ms5fzPPUTtAIndrbCKN/5sjJtK
rwVlUzPgeE1huR55dWBtbgqzPwtJA5dccljo8dhJw9J3r2qb/nTeiIMUitgdIkIMzIBounMH98Z0
NCtQ3PDbcji7BGlS4ZRGTdbsauVBQZHI6e7vM27jooPrN/mEx74ZYJ/z3INAXMyE8XaY99ZzGRuu
XNiwX7CKhZRCbUA5XsCnxHSo1tf5zzK6cRJnGWPCcivV7F15OqqwpyujwKYE2cpDVXjm5S9FKhne
b6lJdBCcdQNv8gIZ7RwL1JtWzu5SeCEd+7FCZFjX0Cvoc75sB6+mUgTpfmdpGjUQhJBh90NTyu4U
DtxS1TbTcLJy8k7nVYA4Hmi7Zorm9u5/Cr/P8FWS9Pcb3esRRV2h0JshFHkAMYv8RLnIH14RZMkZ
6tfcfVuWwW2JVhaRBKYR6VOrLYTeVd3A9Mz0CHPeB6HWUnMJUyod9VIXpwaw00+ld4ln2HnMO58n
Oj32yDHX2fQ7wb6YG8qHmtmWEaACNdTLHlzJuAi4G7ldBLDz+7XV432E+3jgur1NpwVD9ZF8Tzgy
Ik6E0hCQCDRwdN/wSm81UNjRxiKWav55YgLE+YYYScETr/GNKtNsVOGZ7cxQ39H8V7FS6AECl7xx
0bbuyQ2myCGOb6XV9i7jRYbrzfWlMTfKcgTku/dI4ARjpwvPby7ofMUO5Xq4BpXbrgSswaDz+4+I
HVUuUiYU4QaUzVUTjZ0FDEHH+9fGdMSFN3fgkY1EPrhYEB3msC1bD8+cG4kvf4wAh1niNpCm4o4N
Z52NpMToJRKSjR8mVFI06IWKEX0JjmdAFGCH/cQF1EArKJKqIZmjtaTPuU32p9VLABz55WJ963Wy
mr6eW2tWwv+7ygXOSuZP2SWOGVd9pmX/vuE6MGvmZikdy8jGe2eY8+5ilBldrYLtZSJfuIQvwj/O
R9yWixG1O2a2yea6XFkt7YLkKWOgoykupjhOJirf6sDtxZHAai0WbnSIHSnrAsB+J1CXFy7xJfle
4ltg99jt348cP5PNhGMyod8H+iHAsB8WdCTadksuov3TgmARw/F+g9u3tP90vWlmcV2AtAWzVTTc
JkPQXLHr+f+US5TBYsd/m+qo6v08EurXRGE+LqezWghnO6MFGla0mjjPGpcBYwYPT+jjrqcQd4PQ
VQjDkwxjt5+CCoKQSxogd4K5lrL5VSsBzNgZJmFxqnILjby2jnMyTwLcKCqZLMEugtTIFPMeuqcY
SUOcRvtxt0mNBtkHxDtjgFKrjE0vhSvYxlDPF8eNwJ+kD+b6F4rhmHkQB9p+JbnEInXiT2WeWHeL
mjlYhIb3Z2aEUNF2h/MuSUBhyeWlO/LqNFE/VQkS2yZFyegRc6sCuj+oBwu/+sF6PLl+sbDSscLb
p9ahQdFr7YYYfvP1WGo6pIpezgJ0swBC7qKFHD3bAFblyjCckyb3SYudAVz++igK9NR1ecrEcBdv
DcQyshmeW16sapbTZ7aX0SawtOC6ihHo8e2h2/r2C5YRmG6zH783O83o+auh0nfHoSYb24iFAhN9
6xMQ9Cehs8S4sOYT4HdnMGzcZRWPa2DSin9of9imOT3h+ma/e01wkeaqDP9emXjhkurJKrQ3m/U3
K/b/07MI8ZHkcVijns/oGB2PV7bsMLq0wnNf1xXPGDZSudMLzdH5bw0kBzY1NDZ8U8w+fksreAPX
3Urit6SFfQ4pxDFdn/fu6taHFKIOAMZ7asG8Ho9D7NtiMI5ACJhaOH0jlU3l1Zpy1Kia+bQ6Hse+
zcEzkCqv26Sl3wLlUP4HKNCkgsxsIyTldg5Dud+x04Hdi+2oIJ7YKc3DkowNk+29PpgHkpl3omTg
r//7+DzYRK/o4Gd5QkhdOTviE+TYxxSmxrLL+OkdF/qoTY5pqNigdMjfI1tBIl/HbmtGPwV+17Iz
QWC9MMEvqF+zIiPHhpuYqvEneuiI95EtEmr5RtTegqjjHvvq/O8AgYx/HhoDHRa/Ejab4psUwS92
JL2Bs+Y7jporHM7AEF84zQWzis3lPjddcvDxsLYuiagAmq9MQeEUFjoMcmEmU6u+fr2vPcuJ3hB8
9Btylw7M4smK3JKv/eC0mfvXWS0H13k2oPcN/7yLr2V26Kw2qZxzO941eHzd/5XywBEspahGxHsS
Yaqnpz9OpkwKy0tvKvZ3HW729TGBrzT+46ZmlHMdhmdvR7+JZ1C/I26VbTj2B3TnJKIMdQDQfpsG
jFjxDkDDgjD6DU7rn7fmwb3l+Ebryyfvg1QGvXPK5VjQ6cvbj5QH7dioVhn8koETqHLDRsqip94I
tBeoP+DW9Q4HvrM4w8xWYhq7GYb/BWbw1GjeJba8AC/QYLMYzFVPN6YnjXBHrsjLOLnBIU53qzrv
BhcXHOYVROvZlGuwTH+bB8jX22YkcZHJY5cuK99oKFTO2tua7fUYFPd2fq88XqxyEVPTX//+aLyu
zFbijC4aAZZyzpHbdRK8WHcnJov/xYyHTcOWgIKHte3vlhNBRYbqu02KxmhtdfrjJcrKrSpD50Pj
XADaFN+68QiZOeEupiuIre8U3dZI8AHwe+N5xYx/FLLoSgjyByaFjyAEkzukIfwbBMxkODGHV2Z1
TFR1PENiCGu85tVHhcj2fyosXGsn4vcof8pnNmHnQmv9oVaVkZc=
`protect end_protected
