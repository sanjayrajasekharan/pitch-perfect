-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XDAVN68pGUwJAXZMz4GwZ439/RE8dXVtuovtwhlITLc8dEY/392/nDyoTbmu5jzs8s28yr6B6G3t
21PqQtZbTeQ98b332oK+u4X3kGP7O4o2NVUCtRbeT5744mi3uB+aV3AYnipDpwt92LBwvTqMFcn3
WNk3px4DirYeBAciNdiQpkD+XKs+z1TVqHZXM1LXqKOXiahI2+wODNDwz5hNPddct5JaCdwoqFQp
e+sr2d4DVt7P/9TMOCB/kb6BMgp2V0U1Lstv2WFVE5t776uhpSJ/xO/hKBEOjUgHMoIctXB0HbQk
EP1fkm7dPPRGUz9RwCx9YHCWPco4pUQDKz6nfg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 27776)
`protect data_block
/wn3TnhbhcoGEZnGD90T8ZFtYpbJf1W4BSZt+0vxW1+Pq5T9xu0+k6oCvc9+57YjK1+MHHb5d+ar
qaZBLSAmrBECgMbmAAuDBcoz2Et8ingD80R4Qn5gFwrnxQNXHOvtK3oWqS75D27JT5kPAMrFkGCR
VQmy2DYkpN+IE2pxkvxMTIv9G5AOYs+5zF3vMZe35vFQWy39BR0oWOR4XgyS9VQwQf37Zejn7pBv
AEyFfi8fdhr3a111mcTks569k1drPIUUTN1lyjOhueUVUNAng6QgG/9r1IhvskVYbW3vqpFp5+XK
EGc1hrDKJfgSmfJVEn+RQR8jMeQY6cwwnhguTNSwVDw1aNyyXorUj7/XkAkBXHIukxl2hLfJHXOE
Is9vutM+CBdeAno9MTYQP7rqc1/1+6lvCJtdmp7iu6IxaHlEEjGDmeEuzq+dNwCfJaWn/qZumzvG
4Ce6SSK7g02gSWMWfZoC4D1gwK7eSRq8YEg26nelQkxlBjWtNHtltzEIIF+Ho7lMFIjfB+5FmtWU
tUCt2LGv6aZaykJvHxRv1sS17oi/9+joobdd/21PreWlTh8UuWNjlQz2M6QO5wRwH1JAMy0SlSTs
4c5zeWGwMMN/9FKbgoZV49j6rT0MuSjN/NdKA6k62FoHDoWWfeW+2U//0QsL9AhEmGLR84r2oZRs
Hr8So3okVL4LVevXEawfbWXZ+hm+wlHvh3BthX0VQcB7wFtbDakXV5C/plP/smA740fmtbUHo8oU
ihk+BrA3cd/0Erv4AFrw6K2vlLGrAtOMbE4/e0Sg7ASVCOMag1VICpqbSH6BesBU5Xlw6CPw7v7J
CPj9MHOSOCnMpbDCECtW0yTHa2ze0A/JbmCpHAV6zTmoM72jsiHyAm97iMdfoUwdYtHjQpmBPSO1
VnF+D0zVvU5hsS+Z1Fl6v3+ZgnVbs5GH0YL4PtSRfFOzVRbwL9ERWHJRt14K/+dmTicT4w0C64EO
XrG/vZUCq8Yo2ze3t0zMZaBvjNf/YpqUat/PoeE4qZjYK0OtcMH/fhk2NE8TM/tTqQHLfOt2QEz1
OB7n0GSMUh3NzbIMchmMAL7pC2G4unIJckIe2lgs/7EWbOW1OAZiNb0jpmYlWqCOa1jx9RytYE+K
uK6xNBAlllqk1jaAPQA3PmCnQT7zwtXF/FM+iG44NIvcQy7vap2/AbLmBOpO90q9XeVpO+tgbPTv
Z3kMMz4+pDPfwCiLzgbEFvNbMb/OZ1RMzn34jHmmPee58QtB74nYIG975K7fv+q3Q4kaKedB1fnE
/Kex/460wrCCksSTRWHClYfVEvTPmjkCfztJwxMwzaymNorQJQE5GoNACInXopZWn6u93fbCDmK0
dn8aiwizwnU1nslPAAF9JV/C/YEwblzFEjWwU+sm6SzVgRgUop4+eyXIPVMvzYw1iCwOg2G4Y4Ge
cmu9P+BlGnbHj8Fb9p7XuZn6H1zJtxTC86Bjo7l/m1cefvzJc8Vxj1ik2w8zhJetRokpDiPZNRML
xqqVUx3MVeJ9Jh6NzkGZ/5JPCGRWko2xo6uOxwhhBk/YUw+bzXq2OOAeVPRXWRw6ACmESJwlGfy5
EXLpcqAHuNdrJIRtCuzogFS3ohHA0F1lfQnVJpLnRb3DxOoIt2Dpbc4a9qgnVe8BfgZwDXEaIabT
ahMPhoxwXOkeIQFwuMSciRqYNqVH8WaEQIunCDJ6ClNYE94OdfxdOJhtQrDSq3d2QIPd/gXhfCc5
DUoflrcEUcazIWoGZkU6vnM963lmmw4B1Nqx8KLQsqHggZuCnxq0OT8ORnj14boGTj5kBhwPG2Wm
+M/fNGmYNWcsxsrfwzbGlRnmK/OF6Wv95fMLPu8n7SEH4RWuH5CqGae9u58byvfcuBSNKqjHPs9Q
dF03mUwRC8+DJHbLZwc0JXkiw1geQqW7f7vSBLppG9Adly9Vu72+EXyCfi4lqMOKRA+DC1Mk0+LW
wrYhrHmFVIO2UHaR1jQTXPmYNBu18E3fNyY2KESmiDWNBOJzHjNMKh1/kg9fhM11Wl2l/iTtKsV0
6VIzGv/ZpLV7pI7AnrDuWPAulfH6KvaBGGhVG+DG2+Vq73brU+fnOOOM9Y4JrtqT/ARxPpESmfPo
e9wcgjnGk49GlNEFI2qNFtvAwnybyFW+m8NAfwaB1ztneD+cV21jn/q8/SgwIVCcwmOrisQpWlB7
Pq6uIUs/qP85a9RfN8uxM2oPgoB6KHHAA1iBDvPmcWy97mR+aLyjlFOa27fEKQAT2YJQmhzua4HF
GskHy6UErTOo4QCS4UicPvhYMhFvMStDJTulluy7Gr9QntPeNopZKugd2Lk/kAdACqheZRaTbN6L
wK6zXC9z3UzxICFJm1BdBg7AfdgHFfSY3xv9CQVN9BNzzTBLpgrQz8aLr9nc4Fr2LAqnIMhG24/i
gYhMaEV2lnCN57SubJsjAdWXUe9Zho5b81CRhYiA69Ca2KRL/uv910g9WFnmyQ1xkUiUg4H3ZiGn
nJpj7b/9MbqVpuzh6q+59TV8voP74ETZPHwmJ/9ry0NkJZzHB+u3Zg1jkVn27BExxCnQ/LAUhr2U
yHwdi1Zk7vEWCYsYog5Ud0C2FDi9vyp/wVT9EtdEPmZIOw9da9L+UBq9lyrKEgPQVsl5cxVQZFgY
ckIvaw0surqDAZXGRKzbdRHgC+o2eAQ/6uwSNqWc38/w3v9ZSRk+q+fFJdritopuZyjtwoDDKLH8
ZnOxJ5qRq7x4JVjQ2akPzIcAEkPFPN2+CTyFmfd7pQ+dsckzFjVyZjMAbnCuPfCbkll4dE2aDeQ7
V/qI9F+U8uP4C8zWo5RgFqacLQuK0Ha4zXxGiRRGXzVntvPVrEW0rua1ZTNLgyMk7GvMEhTI6Xcm
arjPwZ7yldH9rL6ZGZ2/tXYwj6RrnYBKcFUCb8ynSz2+zncoICZBtmgFJaVnxNKagho/TvkZTuI4
PITt6JeBMs3Ai9XSJcaFgsbr0jvZ970pzyDcg3Tev8f4a83+HCaq1W3qxSNXyXbyOxKd0lqDfgk8
YqJmXozAFT3xnDLZe9VyWgtNAv1j0e6kg0M98yhWdgR5VfBY5ns5O87zbIrXD+gngR/m/wPKpMqa
80BDdmOJo/i9DHqCVyn3jzeTnXt4xPTKA28IUm7V9SShF0dzTyheeteRqq46mP4z2UIrlTjiHHOh
DRQ3bl4u6MWnvAbNRMPGfBvbsOl4wDtyo6cwrfp7Cv9pN5eOL7RMDEYCDGWMPUwaBAhLDHGX5Qb6
vg1T+Uxif4aZQ9Ksba877PKkwLjPuEiTjgxTJq1SKY2iDfIVehMTQGIKkvc1eA7Sp6OQFsOIzRDw
+j4CX5jO0L6vtCj/C5jSVR5uVZbc8ceyI85DbH29Ww5OBsvW6vw8BXvxvXAxEMeCpKaNx3jjAEoC
dBkDbrt4kcmp3JS423Moss6hiEIfUu8HlLZQvw6ABspU1V2LF3wi6Gwp3QCfzlPR2OHbrSoy2i03
B43mul6PvFY/M5s5J5YOElm6EohEdTn20iKMCkPi2u54cquCTlaBUXUpR12UvERABr/dPca43ZU6
sNPOFRrXS+5u/AQrEiSMQXRzpYls2OQeFPu8Fr7HO3jrUVaO5LBtXfkKOqN/Nt0oDuZxKy1al7bP
NzgGdSdw2NlC3pliuceSDbnY23JEoQbWhU9a5SQJu0BO5g9QQFVhmW7EWAVmMn7ESz67juItvZXf
QOKFb6fP9x1waJfESSj+TJeqO2EMo032d8s3CTgnDCIImV+/CSdL2YHQafL/sNAOq09Zutzd4wTJ
8tzR4jpQ8bzHfwKCXc4JU0kyClr2ixpD3bbSpie12cgk5oo26v/4pOE8eDzhj2yxYo1TH483sx1m
Ly9LgYeipDO260Mn6tKfNy6Tkeolj8BJb3wEfpY7Vb7vElXMF0++TuOw4Ag6n2MyFQIOkQNSSmip
/fS0oqIlOBm4OH2qO804XY/5kVNfUW13NFVB4nBFDf9cFwwMTzx/MQrd1ojwrVHJpr4NBbJAoqoR
kny8o7oO9QqIZmGC1PSOPDDPU3bRvSWeOQxQcsyrxtMyhDkQqqEGcvw9QtR5vJ6ErP2ZdW6EKhC0
LFYpgujeCsMTroeD87vAwWS6j2akkovN7kjWPW7ZJJSrVwZqJdt2yRjcorxJ3/shaQHntol2y9SO
1spZ6z4/pAybM7xHmg5n6vUvdQxZ9dLM9FRwH/NsClBf8GUKn1c9ATVREp9cNTiQKNtOhqOASxuH
71LiCjj+GFR16BsrLIvyH0C3vnRewBYldb6gOnDBIthB3NBrIK1GnN+hwdHQUpH8kr9xAjJ35Bam
pS067tIQVaZhQz9Eu7PfSd8b6rt+nybhZXMkT9+kWjqk2VZAYXLAJgY6+UBfPsZ/SLu9gVslseBs
y72wPRUogdV2HyIYaXbcosLcCF3AAhCGJBncq9lveQtWWSRg6nIp2flDl+BLrR4CEaz3hzdnCjMt
aLB0mVyvbh1SeSEdgRJNYTnbpIUm4abFoou1wI9f6Yufib6bx28fgOJ7gDCIT4NmKrskg2cdLlrW
BHni9u2jjYFaLZegTv1O5b1ANpcJS+CZJCRz6Tspc/eHNpuZ6UK22Xjj6eqh/RzlngLhi1NU+pS/
35U5It3KV0GAr4LART68Re9hmx3yx/tHQxG6B49dlTubPRWIKYTE6ufL+m0EVFlPCNp9Hox/BgkK
v0SlXjdSmsCnNvQeVT+Z3oyiaWk0oUDB1lSn7L/yuK3yoy6Z2eZ0OzaugGQC2c5ldKFaLJ9VC2Ol
x+2h7NkgP81NnUct6KQqrkARBlP+SdI3hu04nL3jhE6pMtTrASMTJKP3Px6NBlkKgG3971s2r5VH
xUIp52Hf9GrFVcDQArqCy9xNxOMIx3Xbm2kbpgNcet4mKUjk+2unO5FKL9Dc4wSFQhjCnmvUPiCl
qggi4skVzjhzJ8c67grNF/z46r0jJv4Jf6tlwDXgzend9LMpqp6QqSl/mL1gPvUGTbOTQAwnrEXO
TTyu/arQcehTawwxmrNQG8DROJkuoHoc8EoFX3fJN0NHQWBetD0b944VyeP4KK4YDxemZl5iMs37
58KcQeO67fY1ikb/r2pjziYMaTqQTbB1Mm8znVXv/vcq1D6m1zLImbjVyRic2IHSkoiPM08xVfMa
biN85lM6/d/dH9HM2eySfBqrCMQf1LcnCa6K7Ppm/L722/zTQf+aaESrhoFW9ucD6rdQ7keCBfpM
UhFsq19LlyGFAoaV3//XyLX/RwM3mMqNkZsDaX5AO3b7j284wKEdIfOkxmUI9chMPQGPiqRsFLwf
24EX1AlDMHMcDGNNoPYkwarejVv+yci/yFogx8douBwK9gIfqPNbAD1hvCgLHb6qRYVa+F1+MOCl
GIuJTy5eNdiJZk+mN3EGuYSmSg6UENPm67zTWFqNfWGU4TAEzPIPH15LMK3+A8IyAi4mXIkgtksg
hpl6lYXaGTBuiuixLnqK+uEfZkCRNiSabIXtPp6bVnyCgoa/Wk3RysZyTRhbL9D3tVCTSt2+45Gq
lrxaQx/3T63JtA42o4348MzxE0fy0VSCvLLjCNW3At441Q7ikT4L3/YiAhrwIKOaIUYH5Zo1YFIU
FOMHLag3FWw7j5mq9gjCGF/dhTDsPeDsPVTdXGov+yEvxCJcYMOirczWgNxewkjqAcvLfBjryYmb
t7u9DsX/2zUYHzY3YwkywhUeBlzl3RPR1C1ALNaFINEq4bL+t8G314bzt74QpTEe+q3iT/bjfgjT
E5ltZStLrfWY8vB6mE9tAKkz/dfJpxeSM68M3VDKdFAvicaHtAzOtv05zAUoLwS8T8o9VVE3iCe4
ZO26HnFP9qJBNWPgZ7ou9v5iNTUa/xSOU1h6gVZst8KTI9+EQeZVMzFSA96Q1xy5j4pFzo2cosJE
OzK+gV53DAHka/mk1dbkP+gUf3uXfyreI8bF98oy6gAJeqaXfZgA6tn+aWxum0BtjUERyvU43hoD
VuAvp5U3iY3KwbiuLaZ5dR7PJA4hATzfwLYxCkJgkBDotYipC649tIia5bSGndYeltfE8tnIBW2N
WC/OBWrDlFmxfkV/khgvPmcZkCrklxeH/ksVNCySTjAU3Jvp3JJS2gwfQl61lEHSxjLroS3Xt90F
ECHlLQFMdtJCuFOe5Q3P4/vp7nCba7QddRrjvzxUGsITetJFijcDPoIlt23ruzwyvvHiTSErvXtk
NRiO6wlh+spgN5hwmExwRiHCA2aXBQFbU+bPNIHnYjNnTE5QIPQSVlIz+RjPjxoxtgZKzv9JkU/j
DK8Nb4diErJsAMslW/xKEjbqE+PQwC9wgrIYik0ogNZHtgiJaWnH7WJVLDDUguF1VZUCQl/lCtd+
hVSI1trcf9GMymXFZ/QU+q3DHMhNb3PmGne5wX5lxrEa3UpxdPToe5TZD85Z/JBoK8lSKHJV4N9g
rsrC5g7NTyGH69WM3fNulWWG6bI464buK+VoUDTtPiAAhEoTkR0yIo0lOkL/eLGCHHYTAZL/BIP2
Svm/TFHKPbfLNQztk+psm+aWSOJabDAyrLh4GaLMzecuJnTkzHCT3GNwMqmgzjs/98UaNzuetWLm
Jit4cqG4C9vDAPwCme7dck393BFmIYD3yLEAUmCm5acKkr7Yr4GqdnIf+5oX9nyZLfsKuByYmNWx
AotoW0/8EgU2sDRvlgwPZfD0V9oUXNGxwQIZaWJzW6GB0CUXJuxI7/mu6Kl1Bs8i6pAqWoE0itje
CwJ27PN2QpNdGQl/bgbk0BI0m4G9Jd+1uHzucJ2LOTZf6XXRk4aZzXPCqVuM/obNxE+hBLR7t9md
HzSu7fYnoa1dZLQHlMaW0wf3hU6/MCZ+Ba7MdwWdHiP59ffJczkCiRLOR4ML/GB42ER4DPjhtAhp
IY8+6a2QdHZZkM8SSMPmpVbS2T2zQ0JM/jWI8Cq3uf27f8644htURRnTHL8YJAli1v/ox07umYPg
Wud5T6CZ2nQsDajxv2ifKp13UXxJecHa7gEKC4PaHCAUMke+2dNgNg498AiFLoN6++xDSzrxpexJ
cAYYyD/cCXYI0i3FnotlTtD1uOfp/+47PSHTUOxEz0JLZW0zox7bUria6qgdStEmJoCJVIIX+E2b
ltmLnj9tldcqK8+VO9ZUk6DnQnorrCJ0NiJWmThxnblBzBHg5qI4UOyo+MSUmQYVK6XJkDp5pjHL
6/4VJ16DIaDosY9rV6G2UzhNrlOBb90pkWtbM1icNyFDPWYpdi3qcAmTqusvvEJSEOP0kCca7Q9W
J6MSEYNawDRkwwXDxTXaoT2JXfQ/151KdOjCGXIp8T6++nnxIAuHhHenbfIEaXsCLC10ABJGSDoq
xtexIV88lnHJ+Xtaar/gwk3CWRtK4J2A1R0T0MEzJ3v/2rEnqwxb2C4j8mN/kfOzU9mSf7UBYT1L
FRYuFOw2ZnEmBCCzShiNy5zjJa+mAtAsDNQIc+RlUar951wOVLFGH+jwLRbGWf6XzMVkP18RVzev
0U0XDOc53E5nlSbZ/+wRs0T8+RJitSO3h//nFU9qcNp2oivckiH4owHi9VcHBlvY+93/IIZJBrcR
OouAY15dyUfrpeFce1zP9mMFCKzboVFP1or5lcka7iljlhwrXZ5XmHTh5eT8RiMj9N8m0EZNH7AR
VjZoSOMR+pHjLbYKVQODYl3yelPI9oDM4dKCLb4g/FMHJvZmjWFjhcz7tZsM45vKDNos27cmvdh5
9Bkf1ZEgqObKbqIDSsoasbRPB8nUY/fMcE7Bkg2XcjyMvopzNYt+Ozvvy+vx/1sP0qD4yydNTJa6
ODMU2ZF4mkGNe8dWcZ+UQ1odG+J8iHGEnONyGSyaTrfYYpvS7cyMDoPA5DQMjIU6F0KxMEGrsDgK
LiM/Tur+/Sp53GUe/xTae0OeT+sylb1kwwPghqxGykXwEExApTSBP+CJhOBRLQnAYXPE4fPIFEtP
i+NOsfcU9zJuUaRgMdDS9tZZw29+PtA+vXwMB1RkOK6iBcngtfBYxBkSAgkWT6+h2aIAQMm+S8a0
xEuDH2DKuSRUkLjTK9VswILa346SrWvNE96a3Kxd0KFMzTdUnW6ZiDxxtWXs1tDiyLE17qW0CBws
wVAGGT/NfjFfJuqfK7tjhQ+R7g/4o7DNIkvAgQQobU1EgE1mr84drQulupWhURbQDK87bhkP8qP5
OhYp/YnhwJzcVtiOz5dAkTPW2y/J1o1izMyw+Tm6VpnMgKidmy//9WUaK57GnjT2NdFPM6g/eQeS
11vPJ4VNO10HmkT9MikJedlSoZHqxSfJT5nx0otCc2NjlotoAA/94od1pBYt0nvE7Vexj7L6sgE6
rKeBIipG0dX2ZIsAuokJJ1DQvsfsPV/JgPdpdxgihp4eeK3YDlts5r20B9DNbYAY83fyYMt9/s/H
QRmVxcrZopq6BtXs9kdmPkKV9rMSrPhEMKNyiaI6urzNOovIotgA8edHF6YdkaYkS5c3r3g1e/KI
WahgkYk7OMLM1u4p7OejrpO6fxwjL/moAyFQYeH0lMkEpmGV+aq7gtZqh21JsIUPIZkIqAfjuZlA
IkFGBtuYIAE2xXPEG9WgBFbxuqa9bAr39GSADLSE8yVzh0c5b4fD9KzOFc5X+5C+9j/5nzKhETVJ
8mZrHkDuS8EjoAr3fnrKPFdFzRWc93JKE42l1CmnpSj77a5eAfAeDsFBeocUz22tYs8m5iZq1z3R
Uk3t9HK9E+mmn1xSu2MYhuWLIsUK4i6vP6HyrNGOND5Acte18sx1SWsK+tDy8m/yisBNSNecb2Zf
Gc/n8yZShPNlCGKV0cGsBHd9hM1Ac32TD0pEzrH+AR7Kc39Nw5CEU5+blO1CentASIIrTYIilBU3
wQtwne+KoVpDlYMzVJj9JrAY12oHbu9t1otBqNDVP3PLnC73JmIyX3eo+FPhqCrmw5HQeYpoa2CB
kGRKuJlOGs6hfRkRe2ulES62GhS94/WnCDRuaECTjm9zWD2BFyj4JTkClacEr3EsgKCVLulNElOC
LfCD384VoquCnE/yGzkQB43HMX7zPAgRZ9s1B2dior+KzI3LuYuZHD/LlPByJJijPW4hpEI3T7Dj
i1PUAgijs60X2kHrRXR+ql5UWE8GYn6JnmkrH3OPD1geARk8R0Y2n1g7oNJDRj5TkudAamDif17J
e5qGSf7DdGP7SKp58emVZNSBQJ82UBAzVONNHYpUaF6nVnbJ9fzxwFAO7w+CyLvjqUYkI7pkMsBT
3IwvWzOZSObOoRC0Che08ZyDaMdMOElxQfKkS9QSpooZqc7myYfLAi17SA7/Y/+C5W411aqowtb0
yypw73jOYFDg4jSpRbRmJEVoyKdRgI7MLWbXZHzI6VY3FUAlCF5h527SM2G2tTjtHWttnhmDUC9T
2TBXYyrQyFW8YDr2lOMRBCXIlYsOdY58dwsqu/nYv0wlr3zGLC/u5/UbB7CTgiJlYD6XGzDedHoy
EkOstPDgCwpFkpHbkXKGV03RsbFCwzSjX48iYsbNUmlDkua7Eqdi0Ws7ILQINOmfooWTlZGEIslf
frSFUlqHH4vRO4CD0fDTINt2DyfeUUZbFXJZG6e+EZ1QgdtIsGA8Vijs0YvEzUT6XL33wy1bKVwb
FM/lOd3Fj0aqoBdM91P+NW3B3tcz3RPyljKYDpGxDmTIYCXteUW9P0aXvaOU1LsakIsHnXkUH7Kx
WxhnLIQWjKOuhdUHBqEmBOZnFc+MjTe57vtUmGY7Y81uFEpg9Taol/ZCYHIo16MjFq9T+0CnizDJ
vKeSGVTZvD018GuI8bDKQaZCpD63q7xoOXlFjcVMvLayKdd/5kSIhohGh3zevu3A+xcfnPdlPe40
hpMbh/qeseKlvfoxrroCyLl2D43Y274Xlj6YSR7OX5qDRH/ybkAXaCdTsROK7xG1l1xaIdtm4VVc
0ZdU/hOCmd6Sg9CSVyY6FzJGkdDNZ4A0RjH32UvUUwLTbb+382LZrlfRNBmaX590HltVnxpUktlD
G1ra1Ok+Ux8P79Q92lBThDVaHgT5grPu8fe9eY3JLgM8fMVJp862jyXfDdiPVsbyb8Ks//zXPq7q
BVXe1hDd8Gq82nXUMgoXjsQ0bOnpuTjQtjqRrkCjCWA6J/YEPSelHT384SolJ5KBhcwMaTguOiaQ
2sWGYdOqJAqKv7LpXFyHHJ+/lmiMuZc6mOpGMbsJq0CNz8MdJP6TyJnFiZV8p1hEzPwFBl9C4faC
eX9o/ZK2Kgn8fhIZ9v9blnsnImKApq0oVNVeV1LX2A12QBy0Exa1eCDcGFxViwT9CWn5YY2bTV6x
8CzKGCA+v6tQ76wWbpt9rI2a1gHZlPkqyReGSh0cxycyjymRdEpy56/eal2alcpnlwxjsux0N6w0
YQX9VhT4Tt5MqawwZA/QtxAiNLH8GRvdUfFLrXNFgYJIbVaueSJLTRrX1AkVFHC1c8kUdvxfWjCw
fFIwjci5Y04TaVmzAEMLBaQyfA1EXAXjZw4gdvonJPncElmK2cxdojWBWJiQSFYBBnL9cMg/vovw
x/7P0NrwXVCcpW3Bi6QZ1IKrN+PRT5BMu+NIDqNe9fALe7iH+Ifb+DNOKyAJnaKEdDyNIY+FSKmq
BaC6D01YzoQjpbqdVU6hmoOoHgTvDdq9IYAG1sGd2LoCpbmjbt//XP8w6L3fb3K1nQtwUI5mGiXr
RLJeK90g6og7/5k1wR0KHaWZiEEgf7liYDvRc95sBaqgAk88jlPJVqxygUqeMXI1gyk15m8EtSNL
biEjB4T49F3c5DqU1VwyzBJttxdg/IaqC4tXZQlTbKSLcGloaf1nbK/8GlxOABVCgzdcwzfHvZOB
rVXwULqu9mR5Fgegy1tWLPqoF3OElCMKUBHxlQTK+HdoaeMMTOwG2AtuCiXSHfY348eZHlnrNfbp
8hlumVdEkDNuqXYU1uqV6BeSq4Ivgz51p8BTed/uxcUd6r+xPRCWaAXfwPIx8NIokTy5UTq2eDsY
jndWbm0T9YqbKBf8yBTUYBZ1HW7QTjhZ6uYhzJ3gu8qRhfkjXn06MJefw+ejLHGZ7eRB/jwPNL2b
dquHz3OZGkFOLGIdM90C7BWpW1exkCne13wsu8kZ3Mj8F2P6qSjY5KP8/e3HJT+nhjA8KSNGq+0M
TbwQO+g4v+azeHPKw1VkLMWcftrUwXWRgTAhlpzOaUH30yKiF6TWyS89/Dk6xA4VyW3YPOiZYMiU
yTajS+X2SfKnOrhEfxCYnivQ02HJRtTuB8KR6mVOoC8O1D0jl+9GKsP00UO1oSoujywO7e+X5Fmn
032uwWgYSTJA2ltcBb+EgLAHlGxHfsix0gkHNhh/MZhbeqmFZZ32Ix6ZmhFqdl/Kt4qdLXys7GQ7
kZZ8w68erFx/gASy1wAwsyP8dClONpXWbMhjO4EUOjADxxATEI8AEXeFy6JlYGSkagNCIOu26e+A
8N/GBh7cM/t/lF0/bpibKCv8QPAP6v4con0bsOjS8hADAfZezh13u587EGZpzWrFsQDLRHdT9hxG
iRvKcElXg/ql3BOPRe0HP3OWUPh6plwao2ffAw0Ihadex+RU9FXPK6lSDiSb3xy7qfSEYmTsuXaz
3rGUthQI2gOTDJDaOQr9qcELHoshxWT3y+J5jk+gxzvxp32xcOg0VkI0hICYkRjAlgme73MDdEAV
VAQKt/qXIiG6Q9o8xGQqgc3ZcjJITiwq8VY3qYSXcgen5BZJ7dnBPoHKohIXx05ohJRhE826gDEw
A1B7PxxS8sdvKStg8GgvR3FKPDe9p7P3CmrfDJE7ZyTFTy5OVPCBr6kjJQY4eN2uUHvDhURenYcm
u1N2GVXaHfLEJJxCWHUOMR4AMatVVy6NHuwXZFbh2C9HPmmJPV+KxiPU35t4LH6nny+/cl3J0+B6
JBcGOCdQUY8Gq7WiRV1NgoX6jUvHNJ3dI98nuiGZ3n02IBwbogeKXDDf3/fw+zE5FtyzawtBcNfD
64Pl/FBz+eTpZ80+dL7q55wZw67QZEBnxncUs6VaOZoHul98eTcupun4RicRibSy7O75gQhFm2pp
d+n5lynQEgxjrKb2zIzZfsDN8/UOHOe9btAE4m4DilfRGSMocw8uNtvq9S4I1z+x9P29jmFv2c25
Hp+q4H3411VD3YUDanlypCHsbe1s1SwpBD2GFz6U9rOrN1bmkJII1Tr0ALf1JpbIAXE/Bd/hQtCt
sLWVR8x/r0nVrfpwSXP0R1O9U56JWrwjaVtyCR2mS4e3n3vO2z0YUB9kfhTzywRb8nxPl/UKVmdy
CT74m+6UN7vTGSjhWYCJQP/wgj1+CuniKkr57Zh7nsYLJ7nL02ZI32uZMURNKQwo6zjkNhXmpEx2
2TfgZL7zCUJYUPBK3TWHYfMReqLnfx+0c4GrNSk+ZT5VwsP83Vk3yNG6c2Otlmg4MgneqzhFYXEh
DXMgIIJQC8HeHxa5vlZ9LKZCX+dcslQIb9qNdkd7mbNyoPie5f1TTeE0HLpjVSt+isCSHHEGQK+a
rBJF5GbeJ09EPBMmmFTvQgG+VPzFwy0tdrgjZQEq1UbY0ZSizu+ZztyEqMIh0de2gZ0BZ+X759Pa
0jbqCP0raSM0K8h1Bi+VGMTQ2BuFmu0lggpGr6jGs0Ca74DMlytv7jk/CUD4AqKz+mbf0iAcrn5U
pEQD67LI3/dLvwxeFuVNrExYGMwIyw0/pr5lrjp87lYxM6jqb1qM1thO12jKDsUdWt286MJrAheD
llyByLyyIMQ8xQQs7Rq9Lt0jYKsVMvq0XIwAuqSCa17V6mBbvwUfkZzUZ71eY47rldASNpFs9vzt
T2za4xE0iqsfwKxAKId2sTlWowpe0PF7NbOi8YyCLoGkcPjsqp5EwbyvNjRfu3HjW/luzLUzQZfD
Y65Ljt8YUtGTUqNC39BV1xLLJ94D8hsRHNVewmRIrDjDC9B8/ptXgREeXwj2J0zECni+S3Tfcy0/
mIXx3BYPqzvZ5Gs5LKdPEwsu2KkaeSwe1EN7OJeoXezN8t1UNhCFX1buD3D0PCS6Lzv9f1tcrvvY
PyVQ8su8xSUAlWDGG+rUiyk1HlUD9u2KC76jpOkRhq5p1C3+0xaqtWhS0JdzdqrPjm8tdm3O448p
aDtgJOwwP/R6QXyc3y2cRvFh+npDmEgj4Vbnv1P+D5186U2ryQlxEPnEGkRL/A9jcfQfn86wgXOq
2z12kvvrqkMZtoczX9lTJpl6lk/5zaTWaawz7MEX3zj5AneeYgryrzLSYc2OceKP7Qdtq1ko+zDJ
dk6jIP3/EN4kABd3XUjJ9DoOT0A8bucJ9C3t68MoNDJYxIv8PpjBOLiUwunNN1XJIEkOdAXZzLNN
c5aJL418nuBO1qqDEMsyt4QyXG9MfWo9GRHP7pMOyPTc4LYQ7L2veLCmXBF0tG3HcFznG/a0gbx2
WZ6wmgHhwI2HF5yEIvW3evPBFjOomyncmeoGibEfrl4u9jgJTFmTb5e3bnA8Vk0V44CfXkn8XFTi
AbogCjbHc8vedlaHEYnB8Eq33fHYGgzocKkx7S8TCxwy8SKpM0peVg5A7p4HLg8IE6085u2Z8RIF
1ol1sbmr/lHaUyhY2UzRwRKfL2tVGBGayRe4OCWeA+e6WvbFoH5e9d30CCoq0kw1Z/QUyQmV3Ddh
BHHhwPw+JTnECLCs8v8HzZdcflVYTNm850Hh2HUAsReQAtlZ53338PrsJevrWvuWAkZkmkykfKtR
Y7OTJDttPDJA4pR+TeFuJIH3aDIlNDRrvnCVb+9PnUFpX/788c/lG1aNNCmxtOHySoM9GL7Mi3zM
5xbYdXHBqVMzcMIOFW6sGONBs42lUSUZ4az3dMtqzL0wPB99UvCePRY45WraSrbVF1/rtUtfe7PQ
FneCaueB+ySO16gM+GY8bXHzt0vphvB/psfjCy0Omq1P04qYV+y2B2MkiTnD0JRKYaH7AHQwA8v/
5/YGdgHmClvfJ3yd5r3TV2noT4d+oGuXrBHmIk89YVyihDupjFNatEC1BeTVYFrw5iSkbXQ5QWl9
ME4DVfI2SNKlrkYWxI5bvQi0WIq+RtyG4Ow8T5W/rSF4jvkIs+why1PFfpwUwzPJ5isHfZ5j5Ql8
Qov7Hv7fqIuaHKWZ3g7cV3+sFCoLxTvgaP2MReict0Ibyi3fnsDdWK0RRK1r5JCde2oDvMWwMZgj
vhQ2A64/YfQ5wb5sIR5uRrJl3itT1jKhpXz9/EPTAOS3hfrnfXXJXP2ghZ1OYXPFJw2HbCCEcof9
yiYA9bHskOiA/HUXkVNwNb2IMlBE120VVRp6F1Bbp9qW3foeTTI9J2yWYMJRP2wMjUkRBCTT2JWI
OStw3+oHrF8PH2RQBwQfL9uwepprBgiriFG41PWrnQ2zDmeEmxWapZc48k5uEK3xQIT0N7uowyJd
KDpZdYxSOYD7ZKRw74j+zZ+LFuHT9h0wQBGPCCRNomCuhojmYfeJmePEOtR1m4x2pjQEvzcgIbCw
zsk9qXFJuSjqGzL4gXgoj067n13a+ivJ4K+Lg4gTriFE5LADn4b7l1slUyWYsP7GzI64+s83WQze
FEghRfvTjiYIcxzdQFQjg5i9SjR/Utjm/1HquMlTberB5DMDQyS6fGQiYwcL0WDPrY3AXl8bJB+1
UcmlkYZWKhtZ4THBJzj+G+2ex5Lbp+8UGQoNZLy2kkUM2a5+G85n2GbLwQGnxAAF1o7fomrYm55Q
UuTws/d2xeMNixSagPdp6sCFlyhrBBAeCuZNkHwZ9oprJ2qVcrRqe4rcNqJpLrLTH/3Vd1YPiLM9
Z3iZfkyPkKFMrSucEZ618Rbi4hXXAIygSahuWGYmXgC9PmUhPxMDWxZfRux4RTpPYZbiF2JAX6FA
zrWXE+c+icgtIadT9z4ZLopIHL2N672CnNL0+8KWij0Jns4BO5+T7AVlnOgNqxWJFcyjU0Svb7JT
6q1BKCdbd3Wfw5+HnjOQ0AS7BcdJdOpZvdiZUzJM9HSgxCVnZfEs+D48myilXnTJYNwvK42KILyW
eK1wbpYW7mOXT1HcTdsjRZ3sqHXlYEVr+BUp+ff7Vco7mj9XYy3V8yNHLqqa7GIONL4qP8rOpAaG
Pv9cvEoZ9x35gvUZ0CECqi02o+ZI73zc7D4ig/t1tmgQJNKsmHnGWAhK/jERrf4qIIbeypASrUyM
MWRPvUtlPImgspQQ30a3bppC6HfFsWlYbx69vKVW9EFffipzuse5vam2F4u0Ub7MZbOy70xRp/xg
xPXSMabcvfqIH5OqVEb9xRsr8JZvVxzXU1OauL0RsTSDr4yaWrj8XKLSmRDbRq/Sbhw4O5wHaWvP
MAOdzLFOUD50Y9I5p5sHoNPy+xfnmxG9PQq+W3jv2gy8oBmpvC/7172ObEwifBAmP8RhkVXYp5zo
BvQDaKvCammD+Rd2R91Z/GPYNV06idzesX+nck0u8O9wVLVzrAuWMWysUiOh0zv9nSClWmwEUzE6
gIVyNVgxb4EzFCGh/Ll+KarHpIlOgnJcUowkdlHGslDrGVqAqIQZT8AyX/w1xoF/qXros75uumot
oaw2iY5/z7DH1uN0S2CavkvXi/elNmUQwzYitiKilGi9HsWXvW2cQ9RDh5QN1ToNUKsS79tIxWP9
iHdOwoSnNAw3L6taOcy3g1uK5MK9fz76pqqVxmsDG+VpDWbPrnnYrlwZ6Mp4U6JIrTbP3NXDRzk3
3+KegLqJTwxN4MNYakYADXTvMhqMd+06D9hsjAMEv9C351sY70/ql5lVYLslz0EGlf66Zgg+PkU6
hAIHhtC6aYQhtZ2o9PpLogEGSgJdaGAh97dccTu2AdU7VmQ7eHFsv3IHk7Fv7mIw/N/BvyDK6x9y
LoJifzyA2N8olQMofLRZ13Oh663zdG8ygMNUo7nISTINAl8nlkNwey6jHHd0vg2DzyjYE8ZizaaM
FgXJ7yzGfloTSkFQu3ejzzpkaz37vptbg9kAwkyeR4wzzzY9X8D0/Jdh6w41xeo4aErGsmgvPkVU
CTZCzOP07l0zm3zlXOPzHlLOw6PoGAAHTgY+26vSqBrjj276psDXSy7diIqh5EBtOXb/eKASYC5+
3ZOhbIhdcTa1PV2Bm2pJqgxXY1x1QBzzxnEB2j2hI+CYpEg+KuP/WL1E+df/z5AuFXfwgMHgAYFY
run3jPTycDne8dPtmeRjKbWZwEHMRmnKf5ZghHpGr2gnYG9KGc90hZm6P+P99SFxfZCePIaD5urr
tOmMg5kyKGAkRRdh6+fUv8yQ6lPT1NXuRLkeaxEgRH39DYGlUgBTA7fg70O598I1bvd2OxfYxxzw
XiME4JSPbjd+v26VBJr+AFCRUB9VxcMaHtIkkceySSKaBOcLlq1M3DKm/178Vg4BOMrJMpXGcPOt
VhrTC1IwgmkCFvq8/7v7gYkyfzz7om0Cmf/86ViWgtus5c+x8OcfXW9Wl9tJy8rH4usaDhHV7i8j
41fazut4UcfRMmqwj9VkYFXKbzJEFd2YyrS1fRvIGGdugS/kSnb7VF52H2hiAbLYQ7tSlJgq0TcL
VIaOc39060NPYPgiXn4xhP1nInd17fDVqcClzFMrGO59mpvMZbcd58G2l+iSQZ4xkD0KCgMPq3t7
C5aLIPMo4TgcWKvktpVcpsmntD40FRjk3mUbKVXBcPyioKnsPA6xpvOBnbaBq5Mosd49QlmEYpO7
dnxOehN64q6u40j/fCBd+aEbnh3UZhCx7JmeZkKrSM625xXCihqkB8S3jJtqhbQIrytqjWtlvWy+
Tdga3Vq3bIh+mgFYBBECytCJ19/aUwP8aRQG2z6QYiEQPC94Bbuc62Uryj01wrwluOVTR20GyTsQ
T4446m58mMod6ozpcfdbdoZOvp/3kNRL2uLraV9gekajuipGDOeNcbOmqcZxdTFdthBDLH+ohYjr
EbF+kU7nNpchfweO9ai2OArE3B2HCpH76yrA3qlzarx3e5YUxTZnHzJGj+vR40zT1qVTPkA2ApTs
k23VH5/ncpySHsP1FYKvCVnXxWImXUYqulKd2cwybRNbnPbiKsWBSa0TLDIXc4LRGcp7hK9JTN+X
JNg5jEwKcm3Nhdr+O4RmwKvb4MH2IfO06kZN5e+qlIBR1p9Bw+orHY1plGrMGntj2IMq8+B1e46U
3WX/4T+RwX8gjqru9nHZUrX23PIssJio30HM2zTA8SKepXM06MzEgT3eoWWbaA/K6fSOvkmGo/Lr
q5jlNtFSQeKabpXFBFw53T7s6KKQIKos2kXufFt8L2QJwJpMMhvWMGq0AxyLKDn2zBGeWlvbf+u0
WADuJcQJdgZBzAlBM66AHRYI3Kn9avBg3UgXqtmdrPok5yL+eq2H4o5ktkRY/UbHyQS+KmDDvkxx
zWSKxrSiEni/7Ks1MsmUOXeHjiElqw5WG4OHKcFBaq0YDnJ1YUaB/mbIgkFKQ+M6VQhdAXKMDJ3l
pnIP22luEugp3cjuI8ta+agH3pXQuCUeLNMCPDDBdo4vuaqr6O1dSEPNBPj0NH46We7fhBOEf7Qo
Wexy4NMjNJPfQlKjCOOzMsWNURzu3rGju5Q6+8NOTvi6cmDTYR+iLV5BCXPLgJ7O2kEBwyGmgC9b
Cbw+am07+o7Iba8byqr0AEBySy/dYHSMIcdpI8Xq53N0rBcpJ+QBZcD05K3y4+Er/kiL9+9m4ckS
3w5+K8Ynk0xV9cZwI2XKr8d/cxAp14/UgAmHphPnYNKV2TMikDw7w1L4oZLM7zUQL64gCGBGrKmU
T8wlN2wB6H4OXxlR78+JUyikxbtB0yfYno3thvC9nftlgCICx9YvzPZ74Nmj0lmnMSLDea0dmkL3
Tyez5skipNlMyR57+uZe3EpvDvyZbuW8ofe7H0YxIcW6m+ZI3hYyowxol+nSCKrr0zYJZVknefAM
HwAwJ1CvN5Ok/kWTmGMQ3S74V1eAvrrfM5xZxExZYwQHN69/VBN1+7Uoei2UIiCA2QWF/m19pt3C
/O9Xh0/ztoncNnpLjTDOwTSk0WCVB/NN5JCVsWulLekN7yfMUg1SXQeOEuy2peAA+waXW0uWgDT/
wgmop68+XFUNLpi4NcLR//ooxlW0Zdf2uBK934R1Kugoe6hY4S2iOoYAqW49esRm8HoqCNpYQTVM
9Dr5C3dqJ6vjRF7nl6d12lukjztTnQwD0YaHV48p+8m+ay7ZxqsjwklB1lVkdjo+NKXpNqN1WL+3
JIyp7P3oZUsJlSsgHThwD0Il4jnCLqFnSqshhYjBh6h38DtsSr+KU3nXWoNduREr7y/8M3Dbg+FI
oQOCqkVRN4npnbX04DzOI3ZZBLeBe7ftb4KgzRyP6PCBvFIIbCA7XVMGbsuqDR/ICCcEb5n2eYVn
zfCwJuWhSjv74ftXlY7d404qyrbjVI2luJXS3bIMs07/Z2CV6G5QO9SxFWsPejy2d94RJl6T1xLe
G8dey2KtUo8c2W+iRtITkAQySTi9EF1FALUOwISQTO1yANrPBkwtNTu2XfiDBgQkXPbaS1JLsHsW
fAsC9lcO+/C/7C8Irzcm66micWYuLKGxeIagAedc0q9T9dFqI3vg4HZFTxu9Kquv/giX+WOvSxGT
E/zNMNro8jZcLIMk1SmPmlJ71Ke/HV5F5X0k8J2Ddxlhn401A2yRcu6hm569RvRusJ8ad56GcOG4
zF8XSvMKpcTzefXo3bqmSouDyFW8yBjLNDo6TK8HImB2iAtCFoKqHJDaxr3QbgZzpNAK+FMBU+dr
ncuncI/aWpLUIK3MxgPGik5j2TJdIfvPoaLyJdihH/sj14X/Iqnp/sJTwVRZmfZCAHteQb5lsgYp
HplwVTUQmtaXAOUkBriPLwOsIM1tLedpi0uTPxFPyJI98giq1dccsNsIcCWtEk3LGx41XaJuoxbL
UD2tkiL3s+OOQ9P5NHOGViY/nwSWHw45/9LJJ8svTXlMs+gUzAv4VxGl8yEW6T57NOx8bWOKV0Nn
LUCD6oHOVGMFOtdzIBOCTwfi95Nqio3fOLdB32lRdWIDiT+6a+KBLupaG8oeGeqaMqTAv/+XY2MM
E2SgBpbazVVYtAmoww1xAdgOtbGNUUMzjEmtQUS2mSGJPS8ZyG+Ip0wEbopzEcyOxbJw5W48eGJv
EhN4rfuj6ZE36Da4/toaCg8mdp6YQ5yUBukLGYvjlZJAcJ5cHUKoQQ1An0Ua58M1whKmvgr3yiFs
/7zHjZZ7v88XQiFzALkEyfDrQFcbSHuGrBsLxfb5BwM/7iCfyPOS+L9IqL30ufXDtWJia5LIUQ5S
fkIre9krzAe04Xqad/ruYOsl6VPAqS0RHyuQpujnlq3lcnbMdqS4tDB5f7DMFWjoanyAge5kzvZy
Iz69WRJYWZZiAGNSMmHy3pjIoM1ZeFsU75Hcquj9l3eXZQkZF4lkSz/U3lQ8EVMKA0ZRye/+H4hE
9vScC4f+3KWy0i4p4U7dOLZSQyeOX8TR16Vh4sFLmD11LcaoocMSkcuVCudPNQBpJmGiePZzdtXr
q77jU5EUiPYb3C0WpnnKpjxz/cNdq+OjdiadoqyNi1RfggdktI/PdcO6SXPWAXX/PreM9G+5TwbQ
KysZJuqynqXY/7rlIOjM3Xi7lr+jq/KPX6AjK/ev+gPi7ZTCvHFfYd1oBh1Avp0HSXMXYb3+C8nh
oYHwlJdbt48VuISurQqajlcx2cxnmh2hnjfmWQU6gss+jmAfGt0w4EeP51093lFTN4ALE/G32qgR
VUTr7r5z6kyHdkpmKVdVMUsyjWg/1uovZ8pHVRJYIuTS5Va6B2sS4TLA3OyBqADFfzrVM6FU9Jpj
3qwzGroiQOfdwI5hDtvCFFns5qa8Pq2llkMhJhjLzVxKsy28kSrbBpivFwnx1z3390QGJ+PV7W75
oOysghiy2eMxRBR4M+M53D7Dr9NF2lhrNv/JVyn6G5sy37nbLjYcRZMe6rAz1aX4n4LkGstAcXYs
hzHNJW7eQJUHa3+PSM+wKTwI1cYnf0mhCHZt2k3gojzidJPhsCMWsLaXabu5FnQZNIDN12D2EwZy
b+ocmkyLAp3EPpbFql9otTpugaTz6to4v1hjYzN3sl10VCtQlcg1fJMDneMoXS3t8+XyaLkGBdjM
jV4BUukPaabwkWXgHyII8vulYnsQd2y95i4wvOtcBuK2YzzJk1u7fcr9QP6JwiNwYZhJS2IVKCJq
gxsbohEArZ1r3WjI1R36tmd8j8I8GkhgKlIroUd0xmLkmhjgz8gArLeTW7jk9JZXj/UTcEA/3VTY
FGoa7j66brqsGQFkTxN/U6EUbmifEyG7EmRV6SC4yLJKjVl3p8iwx1ZMZBBUQHEcETGYoCLzXRcN
FwvLpZ2zVGDsDw9QuaCTwkD3nJvm+MVuNTDpUFCpWJC95ZhKZ986t6NHsTfn6AnoNZfiRxinIULp
GsgT4gMUdVeB0tC9R7E14jvDH/W0wlSk8LFAtxZ164RHdTAoL87DLULyXAn3Jc1WrLQtifmpMAu+
oUwHGUQNk5/rXHh+FgEDfKAflt9ZzZtpMNsydF4heKP/mF9P//ds5IaqCqQb6Q4XdqZMWREVpuk/
Uu20QcmuTKvPX8CViyztvvrZo1q4ixIXJIJ+1mvl5lGMlj5uJKpIvNIGOX7E+iqFE0JUG4tWM6Rq
mgl2bhsbPca4t7o4ODL6p88fxRwSD37I4aY6gQxOCHew2D1EDqw56peaWGqYSeJxyosDrJbSyP87
hEKThWiYktOlhbO3vyZOIPey+xsfYPY1H62NSbwNnMGQtCc/DjTjvkHIpOzqTSfsR215LBVqlYJI
jpeqSmOP+GD5aaTCysnOZ1rqkOIGJqYiv5Md9ce9LpFkKgCQkG6WC+cGnhhvGuXMBBlJbHgNguU8
w8IxWnTHG4O4sexjuGNDTVLGbeX1GrwDn5rzuNSodSOFc1EVLXplhqpGtD5A8RjvjOZOGXKGxbVk
wxlFDvnaN25H6ws4tDEGBB/gKRHXCNCt2E25dgU+Mnlufg033UC5H5wjmpMORV9ThfXpnMshnIvj
m6mjLtmV1MXkdRS84Uw97cndWpAuGxZPHw/pRQBd+55btqEFBiimOyPyCzEnL01LWtQCmeAppSTe
MnnwmU1VKsnp1NovPQRT13cwS1CM3A33ls+2mmmvRY5vykXkbCRL0B9WDtH+OzNNFvz+Lp8v5CUd
MR4VWLIGK5Hil2NPA6Huhx3keZyN2r3ZyhAAhMxQI5IE4xdFTZsIe6JrUwbJwcmnKvFk+KpI+r/J
x8KKv0QuWjw5xeesVytb04bnj0l15FrzxJCDUCpL2f4H19J+6pr2RJedYywk7zhAZWcQDSu3lJnP
LTbwOId32zpku3OyHFMiRMHoxDPvHXxguHVOt7XPhjnkSFNTZ/+yZigoZwPuAAysy/sTTKYlCNN6
ws66wJ6pmoXyXXd1pR3tF9z7utqYUU6wa3Z1ciUFY0HKiT1Q982ChoC+drSRkYC5TJw+8r2Z8VUN
sZrrRVFoEheXh5UUPnKXZM0ac5XoNe8H2b/hWQNp31nbka7FkrNcfrIKiqWSPsmea81/JltTXmqo
kaXALk1kzgVaqXhIcK6tjNwrvzPbiuvv2RbEwQkD9zW4+bthiXleagcwW94ZDEcJ4ycOf8bQK82l
EUKV1ml2hnpSXs6k3Piuxb/7KQLdXqqjIc61a99YocNNEX9eZp7NAI4A60PdXbmnj0vKcY+vi/Uo
SbTh3vmarXZkcohX7vE2wDWhSwwK21NmAd14g5zHhcyc+KZ2suBLiKzzeNmDiB7buCh+3Kib/A0f
d0+tgcsytvUe5Z71IhUZFF3+aiZn4RPSW9HCWQgxZlJDIvEfrhKYX9wjXyAGJ2Q9pOZUvpBInrKc
gBNA2fhxY5z8ENriIzZtfYfeAkpkNvo0/SYbPKt9gk4tC1zTVAO89s7lTc0HJbS4qcOhRzB/V6ig
rPeDObJ8sqouhB9KZyzW+BWJhuUgn+b4n2cdQNQaAdSq/E6cCURUOX04doc4pZ66YVupx1/qUHdS
7CKAV7Elv13YJpNeRj+DT18sMyX41EwG/7k/NX6tbjNES0PfgJOzATZqws2SoLBdXAQJCBL5mIxA
efHuxB8cNmU+/gPmhcpzP4mJrSgH9C3ekbX+V5dpQyBipjAtw3aTyMAKfJz3pZhJgxDLvm2/SHwV
Mv8hkRf2QqumNT7cTJDh/YHdnS7HzJCzD+h/MJRkmyfpi5zuZAhFV4YFrE1S8HP/NI4whC9W5+c1
tJ4sR5o06JmJ8XEHLuTGDdYiIWIwdyxthqhziWp3IWEkGILSx/dTqteT2SSmUrDVwyFfeM+TWzr5
aSq//22s2NT3A/a9U1/qiqKf7+fZZy10+iJQ37v2Y56XNu3UazQ3q+NIFejORWxvYhLqyM3SGecM
A6gIp01fHZpxRLqA5XHCJUCWM1wywdew1kS7TK0vEs6g05YSI45c5GVZUXFtMF1YGSCpjlPv4bo7
KdA38o1yTrC85AFLUOaFOPP3m5pfk/4IHImXXcmBSPOyyzFlUcI1SC+QeBQLJvT5BpePZDpmy9PJ
MixXdI9tMr+GYWCoQkvA6wT5wLHx0m3AhVWg/T9LhF8emWj3puEnp5Xwuhco1eX2IEh5NUCWCgss
+D/B0+Xxp2vdgTqw52dZ/DBmZ+dU5lXw0WaT9i2+eNqbXY6lIOTbL1N7iakiD8aPFEG7zyYCwFRP
Ovw1EPQVa1j9MF2I5h9/DJQnY0t1JM5vUgJqFppBmUzIXV7uEnsB8+55M/YrbSpQ3+QFz/87m4Bf
ZYJG6Pp3Q2G24CVN8wAA8MqZfnWo306SMgDkePLX7wwwCU83Eqb5/0/y4VbbR06TRRiS0Tb8D98x
e/lRWXxXJMdBYpmo3IKnNdQqmMSq4OPyesNwuaAvSqeYYDDq4JpxE9fzXs4Dar229fwejVDMHCa4
1L/MmeWH/uia3wRqlviHSIkp3e3gK8rw6kOBypyQKI4mJ4R+iBY2RmLadbfkReX5YxBvqQxPUdOj
uNe20w9voiMZoR5fSfuHq89ee67Itoc64UQScUnA2doH+Kic7HOx9Zt4WQW3HmU1P+aDWz5ejtDV
lIks7xfdcMWANLAUGL3HWEzpolfASVWg6mI/DBQpWlUdtgSyxyKZevpcOQX7xYizSDonEICk8KY/
JonmYpF3q8VLfyu5CstSByg5BcaX+udSlhTLRrWHrn1qJk0+Y0s/hl5eZ5A00i2+wQn1+xAoJ33X
il2nUKp7M60NopLh8N58A2tTbyORuLOZAOtZni4aNDImu6Zo4ZmYLd7/fvbYPRyQCLRhDO/s7yey
QryZoSGbzat3VHD2uohbE1XDcHz+7J6cvsqTRliZuFAnw/oOtN/aIlMvImmHlACXi/WUkk/AaIn9
AAbGCPSaNqg6ksLJUFM3IBPrtbfwGuVKMQyPG34IPHxA/xsbvkbE0UVNci56l9Mtasv2gwBU53yQ
A/6p0Rbayvnjs2+ubSaQ79qNPgFnuHvCxHJqGdwJk3nZHUMKlSzQZGN+7CPpOr4CiXuDDhRQOtXD
55KJP5g5Y6/03RU+EQosCjVsHCS9qcWNPux+IhIsM3wsO8tMrLxMnuisBp4wT5c15da3C3OBAMG8
9yybL5gBEUZn0b22hhYVs47DX3k4PBZCdi97qRidjJbAmYkd0hR//at37CXmQsEnZ4TfVZlOdH2E
eAue4FMNU1KAzJUTL+8T/ZXHZPOCm6ea8+GYpo+hS0K6ABtsNPOYHp/8IOEu6cMMNWIfJcNZVlKc
aL/dBxSaMMOk5A831SsLdIz7Mmdd88rRfrW2dIkP+svuzF6zvO6QMdQIfMdsjn8gMdCIMgE9wxJe
/bZQzfNsR/jVKC4I/bS4ycMUoASUskXA2WA24h6mHFFwmjT/ez/JEWluiqgUCBDjbjTM3WYsTmPQ
3kI4XdRggOB95/WztacqNoiihN41OLuzuKMNCPNnixSs/PNjKhFRwYWqwroDbbCTPq44VcG5qztd
49z2msg35qixkECoIyDyVnDmz9WcEYd4WYq43h9iX6zypQtUHg6I7l88Gma3Vm681GhFznvvR4vO
Z5gL4LAa/a78VMPnPvE4S2MqYX2sijDbOoQXUfY5EXnxp1qUHTf/jjlNOUaeOc/h1KWO7xFtwqSO
d0Jv1uhokUtzjOx8c65WZGwp4qmsRUhWBmHR2G+NB5yaUQBmdoP0gp90d4g4utobyEVvHuZHXcry
h3oECfu99A4fiXmjN2a+VHyb8VCgi/kBbH5InQ4f2QS/1NDo2CnKcseVlTVY4uhFheq8xyG9+ba8
VBSN+KL5jBlvaU5UCWkpoJ0xrE6eZ4+t3zg5NrlPfAoowlJgz18EUlKSbIug9z9HQ4LfvtuWB32i
Jh70Voo1KkKqHmVQ/dc7m3e+EKqFPsV9KGPbyzsfF8NKH901MIlaoht8Ya9n4Zq363DyGFv5AECb
LIQEFL1q7zr40z2GV64bUzJpvnv3qCKYXJLRzbKORIyhi+y5GHu+R2xwfNZcNqFlIE8EHOeT3jy0
T10DA9cwiqeEQalEU3Q9L9n5Ozqcr1lAVr6AYKflx/i1qcAtsBBO6jeDN3Spr6e9urbsRQkY6Xxj
XLkGyb4GlX7fqEj0vU3qI8iYmjLuoitLxmrtWTfPkUuQzv7/+vLoFSKmietkVresKb0beq6dUS/P
16XpDk/e4WjTmcY9rUv20Y/0Yu7tahlf2X+mFEJtkiC8LyFp328Pu/0pB8peNZfUBF56TSSnGiwM
JTJv4FYXtC0bVWSDl/n+tDCj04Ib3gaQrl+QD74eNYvBbSaO82ptfdxWuB5lMyl3y5foEqhF/Qgn
cz8d65OQMDNlkR/H9HDhTbgrlnaeHF22/BGBqg1gRwO6dl+8DKjtB8x+rB1pKgZgbPAVPgU5PyTK
Q5YtzKK64IOGXtPsEAN8O+/xwxr8Tg8FxRWKP686AUrOGEmP5GsSWH1BDZYSnftoNISzvY8yjO+H
inh6iz8TuuxfwrWVeCHZhf80344o1HCMQ4Ry9E/Iu2CJfXNFTW0fuoQTh4UzxO7UgI/vFyevt3xX
PjiWe1PWXlL9MNHvX3yNllGqcOuxj17v3udY6IVHoCkoGumRWeoTbUluFJuBEDlwT/6wY3Vkgt0J
51YgLSHQ6TZkItmr8K2tq9XcpRaJ8/i4JX2oTixt8EPXT/DUxmFfvrVrjoftX5w5TKivrEUbFzdu
ydGhVokuFvW2CG3J+SCaJGmlonXDmFfFfUg4NdvgY6/LpvRkDKTdjVvNYhqTVvoIByq4CQkvDCw2
8wnyEvSld8fTKjzHG4n44ovjpCXkGawHiQWxBosdYQMK3N2MgC0txnCMTVHx4zuFbD/ejS/oxAol
VrPpi5sNZ7el5aGH37TSHi56cnHxdfWLmxbExJNfY2prtFv3PaTbBH4kJ/YtRQ8QtpgU4sl2P83V
UNKp3hX4nvD+oveu9/H7/D+gcm77N6a/qC3knVGsta5ezbMvnFHEnFtxfgrZtJZovn7IRvaA2Rrd
P5EyAziYiL983vUkigK7heJwUV+1/ScLiPkB3ctS7NmKk9YchR9K+b/qm4pT/xuyXKolJkzctKZ8
GBE4JEZipld5PgKOoNxj3hQNj0VhfnI3p8TJpkpHao7Gwg81uYQD7tfsK5MC+xjxv7nB29N03V/i
qrpAo/FwjAhl35BLCM9LePdrIlCtfwbkE2MEFuyFnq5TOz9OjDRUkyq2RkmoQio7LW/AKV1ybqXM
uss2VAZkgAKq2/YMOquz5CCjIL7LLMBw5h/aES92jo0zFR0eTaflWm6S7mP8YymkBr6Yp3OfW+uf
fCMDIfmgvowNeWgbYHEDbjsFQBWq3gd6EFuIb0TyjohO6jA00DFxr8TxiOR7hu5d1lQ1n48NEf3T
ex/kBm9y6knAfBi5nZdpjiugwD1G5o4Aq0RTzFRn2BOM+QUXmgm1S1tL2RE4MFAUQjynIdPwZPbJ
+or8uiruE9JqraNSGY/D1JUd1H2UrQ2hgUNolyoEWSwrfS2p2E3kCGFqQTpkQ685ObuJAlDbx2Rh
nWGH3FKFf66fBHzVw+ek0lOe/ccFgv7W5UbGtDKgm5HNEjuZLZmMA9r1Ru0qQodBzeclUgwQD7Fx
iUXTUT762tofBMsSH3VTwAlzbY5D1Z946ESkSSCh91gYkYrF/unsa4Y3dLEKMMxQfdwGHYMQIUKo
NqVwXnesadxIUMgrFOJGA5zZbEEtp/NEjSeWSWFteXR0T4PUyaRv77FNNw2trbVV8odBJ7/lIuOn
6tLwobuUI07j8/SJpmchhPc3d0m863vso3Y9qJmMnWwNfhS4w/jCWovpt+BIa0jg0R0QAimbCQml
uo2Ru9XpOcWKIyV1fg1QmMRjlQ6LFTkfAEU5wPO/iaJNMd0L0bDAZfrztZi4x3NZPrcpMAsKkh+L
hsd29Vi8pIaIuIJ+ogXC61JvGMcXHrb7DJwwLTgMCtbLT9ymyBlr96K42G4UPB15S+5+fTuNw+mR
lO6zMSn3w9VfGHBYDU+YfmimLdg7OYehtC42jpNdJLy9oWW96Pd8RW/pksywmbS4TOwbFSr/aG8n
HEQcJLRXJyhV4/i08PTKu8PuMnmsTx3xkOReu3FifFcqNtTBUC7egXDEb2Wtl/HeHpM4a8XB7owW
L/h7eBk1OYLk73+kRxTdZz7XNKuq2l/iKShIwmFOdEk6Ax1A8jRM6UeZq1gIrsuB/6HIO7LdkW+n
FpE8V8T+gdL/w8XysPxS2iNe5YpCmhu4FDlEVgevSsGlJvyD4lyj86mdtas2IXIq2ybSeL6R01Xu
KbTBys1CyI9IaDU7mKWwqB+E9uoZpzjK44JPg1e0GCuDVJZVWpnkCGg3VExzVu0cDmvSTRStd3me
O5FBYk22g+iMewl/KYWxssrW3eFsrTNjq3xgcerWV6SIScXvTZpG6qvOKUNzu3Lbb8tQf24gKKgI
ZlM3c7gYKNDPzkjMCfzGx1WOzWBOP6UII53PkNggRcbmP0hmHKpWeV00hSwrPXwA73LrGIfHxG3U
86MPRWYaReBqo5oftPZ2ta6czzLLa/DuonKKg5w37HOGiMKDafotz3kT3M5yGIbEjaND7+9XPkos
yrS+gXWT+EgpdD515AwQsanInw0bqT6qektngUBO5nHtwQyhr5y0TpF8impaAYJ7tNcg6OikA/dy
3x5cTvDlY3BahyWzf4PRNYJQ7q9rd6aPJMCEe00yZ1PEgVyR1fFa7n4/OrT+r1HJrus/JhxUQclg
YqpHNSd+wiEO8MDy015Q+6l7Nyb5vmnwW7yA5oIHC7DCKkbspKseTqhj1UTqopS/JU6JUbwakBYA
+WS4ip1EQh3ViJrnNy7BvflxKZliLwCjqTYefOWuJMF07wOv6uM8m7cpsli76UjEHDf1vifyvKpx
B6+YeG8YYYY47MagaFIYDVdZjcaUTOqDUq4q/OI1oB5tT/ZHjs6xrD0Xtpd/uIpJuhARzo6U207g
X3PEnV5rlE2A2MgKpLRcgiwU4US8A7GclmMgOQAz4BV6Pe4EvtmfvPyg6JFUzqqHxhD41aZVrqyx
08DM3QvERs+tyO4UUtzihsG4YBGbwtV2rNhcF3k4IaS4UyVeTEAZzX0uNjm/AdkMgXNhpWT7oAdn
7k8MxPuelXo0B8pIqogGr8O3/VbzYin3i7Ptzzhv8vohNOHCQbjjBMpwQQLgHntA8XAHAp8kjMvV
qkB605RclJWzUR/Xw4knfZMjqOnG+O+0ThsEyU2vmdovD3z/FIe3ESLN+oR7WJecfcDQlKjLuP7H
+NTtsOYXXVJJq2DLIibLfMZgHsqBULDRmrGOOrppgyXtdezu693OAMmpc0NTnTbcpUufkt+9G+3S
BViMf9sdNW9KF8VSQKfjtQn/BG/GR3se54/tLD5ATycRwjMxh9S1cK+/LcEJf4H1MgFVDH6825MS
zgZxVPPssUiolbVZp+NtY3ljn7QnrTzchBOIRHbyYtFLr2orzW+6Ckuun1eCjRYFJ6Uz6PPHBzwj
GUEIUwcLLk1EPYwKuZ/m/lI8vdx1ZBcoEFxwiRNJACt98nKVpQQKJ5VyqZAJ2OSv2fC38A7UV8G4
PfwE5wu6ylVlumrcy/nE7udCOc7uhzXrmBU89j8fHW9bCiIjSWNwYPcYpeo4IQyVe2vMxV0P12Mr
6dQSgBVNwKiuKXKtlvN0aKDPtfhcnhCbhfRHzOnZXLtoNfYraJKId+D0P9IMtXCHWeEVzSXh+U6k
c+GibFfpYDzwV1OP03q8tak7NGLZHjUqeHG+TG262oiKECNkC8//rfM9hjxesz+qqnhvPlwB9YDO
mi/EvhutIkdUM43lndcH5hmpvygY5rzoiOpMEltmbiZT8LHWQ8ZczVFtDP4MfQm3B96v1Gq1Ycj3
mXIaqz82MjPsi0F7xlkkJ4BIFtLSTE+3HtW06nzEK//AM902pE+fA3RX5Q21WfH1lD7eWutzw3US
HVvwO5t0EojUPWKQeHlr6zFk8Cqz6m8S0m3QoHZb65w87OYVVQqak47rfArpjuhHExjj8F8VcLTf
uzBz1vE71ltF28ospJyXTuQtMsZe0cqYOLr3iknbHoElNbJV6LxQ9KujYJa5hTjv9slbMpD7tWF6
I18oPXkI0fIO0NTgCn1peTARWWZ/b86ixqw21Ly+x5sMAh/nqO+CgK3aLM+RuwB9LE+Syx2r9uyC
p+mCbw19yQNdkVnbiJJdaKcVUdZqcgqbg49a0kJS4tUQu5CPzzMKZCwdm/tdyS8YeCf1FhY6t7ew
NQq2+9oKB6tJyar6EwnFc91vGJnabqjGguwZgG45l7Vd8hRb3qL+wpoieJHOwxtj7eNfvjb0L1gV
qgvbFODS/7n4kvU+yrFhdQihi7xn3eMcCPMRs9BUst+W494nDa7KKAyYLc8tkOHheNLn1jkSH92V
gHm6dPUzy8EFzzUiqd7aSrNZYDDkofyyxhGKAFeosxAsbevNyM4s81wl2Ay2L5k1Pka+I41zQZMX
GApO+Qh2r3Q7gDUa+uDXmCrWde28AarZH4Fn0oi3swz5uPFccOBoUbWp/Eta50XAi7Jg+hVF26Ut
SDsqZnTETyU6LJKfiKagnv7OLz9pikdOgi7CcPfmuB/AOjsxDy8jSY3aiU6sDt0AY0uL7VpWdqMK
PrqRk8G+TlJwv1VyolIEZh2KkmSQkk2g7SPcqBOnUKzIiiMYMHA5DI2ree4MyGxO5tAFGCA2TT0Q
YbZs/abunTCJhlQi2K86D6l3WU4N9WHiGG6pk4Z4lV2kYFpqOAyAaU+KVMVLT7tgAVqU1D3D2bXb
XzREaU8mlel31Jx+0UAo1zuL7dUxTBRe+huB7xaC7SFBOBWj5VnXgQNZ4iy+3m25qvohT3mxD3bY
vkf7vcU3/L/OQGXmBuSozL/aMZNWO8PITz4/ZkzmmO3sPk0HrBYtLw9UkMOucmWOc1ZXICnCoQEs
DSN+u/r6zrEh7F8iB1+QW1DDXaivCvc92DcV1ODkbKD7XW3L3HxtbnQplFKtYs+5Jcvoj6mV/2F7
CK00qAXIiA2rhF7C5STCImFXqZtTJg/8LGfALPy3AXqByfRK5EU5p8rG2PtI/CV0J9tqOkG/2lqe
UDbO4irie5QU7lB3MycpHU7ymlpppqLuPdLrCr3CQbv3NcU2s/nz94BmVPxeAEd8v7hVHM0ol/zZ
HmVGrjTSY4fmHFrs++dmMO7n/RTTnpzXAMqD4V0zJPpw+lYRa8QnLtKQDSHWvdWIRmVPgcO0QmXq
2ECIwuBh6ZsXa/7jN5anS1Km2IbOxTi2lOkFUB9fejybu4e/EM50eXCWNtn+7qSij+90Cx4lgySF
Hi0zw2PKcvznUlZQEk9KM5kafLLsELIcHgD+pL/bAjydUROGz+t3TXzYoQntDqs6gUYeW7l7BEP4
726d+HOiYivwGBXkpN08k5LwjhIaBqLhK9GhcIiL37Cwej4KMVhYPj1104ed79dsvGtNh+kFxt78
UMR/9tySS/2CC7V3nqrOfE0fzpfW8ha/14yPe5amF7bknYjwOg7FCl64ewCSht+X3NXQ+/ppcrEv
DQ/UD34aokY7MWvNoovyd+5H/O7tn+PawRjDRHAcqvqO4lG3WKsVg0LtLUZzBospUcOqUqe1YdpH
+g9gQmTKyWUiOjvkFKn1x4nh0OkOqXxCHAjOuCVYycWz3kLApWKJpu2iOMjzTM7Q5DcR/nfSIUOm
ut9/szLX3lxQN2o1YwS/emzD79bBCC85kH7aiQByVQfbrCf/8k20kiJRCgUmxWUllov9k6VVkc86
FnPxAYtX378/HADJhRtoMXn72p+g5ETb4voat3jKJC1MKwQB/N3gdodzKikFXbYZGw6ZGFQUXb12
XqiYB5fMpoCHdPjingPmnkXh461z4uY9We606qiPiOvy4/ku5rlGPmNCAz4RzF5uagD//4UV51nr
yFH2NP7h/vRZ1AZ959CF127I30jthWvbzU0xCEEepPzUohX7Las2SRrskFKh14/KMp7egnxXqE+v
qqD041LPoaycWf8qJ0JOSnIUGQPRTQVEz7FntIwH6Bo9qlMGy8twWajoERyg07bhUMqz6OBP2s98
JCSoohHogFI2tP1jVmaPLjvGS6DJXGzrzOaZM2IF6X74doMjCi+z9dteMGm7DwqQTRoEvJe6fe9/
fbkMjSuBqTqqeXRQmHZqOiSXtUX64pvcKSaTYfR/9SnjqRM5CSApmdVjcw68v3vb9hU9Bu4ndvcE
B+Wm5WWZTGniFFgbiOXC4k1/+ePqECN1CvwEMKiRLP5D6aBRLkZgknzokkv6Rx5+eVEEn1aGrrW+
6gdCLlzomHvw+z6ByvaJr13XtVtj2IieYabQ7/1u3FTPh9ciLnoaIRQaRbLLEP9GAYmNBIoLn3eK
zEXSV829x/18E9DiKND9W1tTi+MqOCpIWIwzymIw/APlZ6BKArEUb3R8lEGzgFBJP4JJtu6RzTZI
8I0VweZHGuPeSh3Zq47QfSM8/9MLWMJgkdRJ5miUAecXptwqsNo8O/k4LqJJ3d98NVA9iaYmjQEf
3mwhz7dT2M4wCMkJCpA2KVWpS90V0aKAlBBBFFReub40/cGd2DrlDjOvo/slXKuxe5KmKK2H4nnO
3rf22jd2mv9hDk6TRBlsyoZazWHb/R6H5evuZb7KdabiCBRw0otIbjw0ML2rhfmZIPmssuj334og
uCZARiAA01MfQXCrxvxUdcWvndryN9biGwKRUGiDL09foqUduovk9+frWeITybSP83NEMhdAP0hO
nOcisRkNBlWu/Qp5Drj+sKWJoyY44wJWO1h3obTfT4NpsTlgvvBqKtUNm6MkNqKNTYO+i8Qntyj2
WeXX6CXcaP5fDKCYvLg8Yy44FwqXTu9s0ClnAW50XymqnJYbKKoB+8b5dE/1qGxJLTPn1EETQQDU
/nhCMS7CbH45pkQRH252EqsEE1u7Evd6D6PkosT1orIDlxPFTD9A9ggQI1122KPXgc/wsmb/x1mM
QbodL5hW5LnHgiXt7tbmh6jLzgzi8qtv+jmpQDCG9xhU9JhZAeURqyleJo0jOX1OPCu7KmbpJ06g
Xm9GI0OtULYixLSboT6o7r0v+bAOVig4P19XenXkzWw++FlvDk0waGCsGcNTXrheAserZTo1RQn4
ff30Zn/mmzfl++1taNuhmoLqGKMzwtnHYFyCP5MyyzWB45X98SQXSrS/O2iJvsSBejoQokyxe/x6
FPeSVha7hXtUDv4E8lTYiZiX4cTzx5acXd3yhkly7LGyF92/LEMVAxuZL+24Glwg7YttywzrK1OE
pnSL4B9PYr9pf/TBcjJdWAT+G660lwR3DNklFcwBFcMCkHu4qrv/W+YMd6hedKy03lZ1s420m4SH
td1lAM8wsyYF3BbUR0plnt6qsFRofquslxxf4SoHN37J28CSUv5J84NWH5kOjTWB/RwAQlS7ajxD
v5EdjQJaAd7aSQcGU9pNvRMUfnKoTE22hyb+GmgOEgSgHj4z7VyN5r+CRjYxmO3vBAg4DGNCR7/Q
jRN4ngzAizpA9zu8IXD5FwrwDzgYKeCZ3L3C8Pvoo8Spc7o9VpwrvPW8x4UIVXSycU/ES8caJVeU
qKNnjTD0+TJCf4U6K7E4MpDC2iwlazsYy3KO+J98oHFVs04+CCAvq+lHOTH47gzS0nEvG7+nu2GS
I6D1xNk6oo7Teu5ga+uGcPItoqOpwz5sfYldLvSlDGfYDd3BBVzI4if1fJde5waGQKVMUnhbfwuF
084jP7MSWXHNZ5eLmMPybzKlNBT4YegDlE5osnkRV10E5+dTuudKlDDAmJiDcxWN+Pf0EDA2qJMs
HRItviacYXIyHsCJNrgujZjndjxgM5yvOxOSU/LFlEi4YqGLAyGbBEdyZhwPGhAM+J/S95lqhgR+
HHp9hrdLjEtaa6EjXlyjMZZdYvkyZoerFKEC8mErLJ+asCCPznmDF4fv8pHmycwotZh/GpNRtT4x
cm9awm2byAqavX9TczvRL8ct1Am3yPhtSY2wgddeE+WnBhIh1Ucun6qNu3oBBKlcu+br5m6HVqZT
urA3IIHXAoZYBOpsYteVo1p0ryiBFbKfKgGt5/UcZMsEI0jiN4A2CbsshQYaFaT7C1F75rrUZL2n
001fcbnrRY1AaIVj/d4Ev+5a3//Zc6G2vfEwtVrBiZxwq+ZhX7SxK1cUIpGhS/zmNpNmaVpeiIEs
tqy/ne0K6dY4iQW6ouF9M6NlDWx+655jEVamlX/X24RLYPMqsrT6aFLBeM6gzAj8S2HeBdkZFQyD
LyGUdlrTQ2c6GaZTCY82Vpn1UQIMpkK2UG/npG70ZoH5oSf8fG5sfjW5Gf5cH01lzPIPh0Lwd01I
NAKc4NW6b6/RQmF2AFVDnHhT2PsDpiVv1W1g7itrxLQvThc7tj96ffKEugUBPs5/FIP43VQKHSgM
lFOU7pAHNjeopMtRGPbp5I37hXF0wxS5AHF58pn9EUhiIfNF9y3xfVuUEgARnKfiOY7IupEm0yXL
DI5BmoahHgsRnZinsGgNRHDDL5PTGENe3sHf0EoFQQ3VH7UwoZgwkqj2mhidzxAu6uQMfCm7L9Rz
2EyfMGFJkW/UBOWzQwz5LL95yiHapKqJaBauIx5Td4jU7tp4FIjPfMJC6T3qQIMZ9sh9UcvdDnfn
HtQDq2heQn1uRjA889182ZRXSBSWpKBjMraLQ/G/TsKakbIB5h510hjX4Uhp4Deb5fWpOSqPecZU
yIDiitetlXLh6Oifa1d7jlDEoJt3/A8Nteavj2dUbBFN+WgSACsPBg0SwucUyRC6eEy7pHQLC1QL
2PNVpTUto7PMcNFDgc3hWCONbHfS93X0TUvidNDgbOaUjd9+fCyao3m8qmXxsbwT57m90Ife2jq0
mh4p0KOkMUxPdqQ4EcUt9pnpAZsLyaAbUEAPoQqh+yvRRxK2VUdlChfVOYtL/GzJI3lhIGjMU6Zm
Jgky5kBlmLxYZZMbkguRB24oYJHivEwwv1FevoLcq9fdTKbaPx47NmiCIFDepTRlJnEWxVejWk4j
Uc5kHwb0S6WqRMh9M9L9UceG3AeSQx7kKYkpbRdVP3iVolfLG0LOTJ4OMLTQYL3umPy9NWBFXtNo
QaRZbz10ZzmhVgBqANfCQC9rjeqLxMHnOsEavllA1tAbQPP9LnCx7MpIoT/xf90HWb4jHWpc83m3
7kFQ4y1KdM48xRj7B01PWTSxHmeFrJVpt/NQ6e5TLAV2kq8oUqOr1VENeuEvePwLhF2AvGTB69kt
+UduuioNGxe+iqfLfXkdqH1WuiigCPOYShrDi0k5+IUAiEDBDx4Yx51CfzHGP1NkVJCNcic5iV2A
9DwU+k83qKTyQ7a0zcs/24dQKlB1YU+UxpgyUVylABbdOzEXPUMU1Vbk6r6NaYoOdMgOxTgYKFRZ
4nTqEdJhblK6xlBvdx/EtL9Ul6L/wHNyShxkqM8A7dgAB49/t5DbNbjEjtt14/AmhHnkdo+WHUdV
7oTZMscmx78k60YUeNQG1bGFcd1GvB/moyBjcVl0hd9/2Ot7H+cZRx/A/gczf2bj3yixlst2BCmW
U8ld3e4oeo+zB9e6lq2Hht+c/gzy5HH/WNoTD83defYBG4iI6LNW1RgGphu/NBPHpKftRBis6uKk
eOdpB11IjgVxrcHwCyplgdMX3wWfoYxshgKAabbSlY/ISdToUfPW7GRSzzd1tQ/K2xRLIwfCXMZc
yA5IqBFdQj3IQyDAveV9c0OgLFc6M5VJUvwkPODOCs46zYSF33cM1rlCnVIn4QdRGNK48CrFoWry
rG+eD/Y9SxZDPV9f7nJUUeYqiCkIN8ZAW6rKcTFsjTW2BcY5eyK1UzErhk4qXCg2eMQZ9j3PWDgf
Ko0AThHORpADFHwsP3wOWikjKYVL0E9634LUBF8v+PFzEA6+bHnaF/VIVVskMotRGPBoPdA/GQcX
tAXK9jXGMaWW/9gZ27HnQOrN8UHpl+zFORZlVXUvQzSpAcGhjdq5lPSgUBI0h7MWGiUQVgYiI6B1
avwXC73Q0GUwMQf5v4TfDOEpTH5z/khG+aH8GNCh9LglDSzxa5zuY3Dw89DfusFZ4Q3S3Pi0SjUm
mgwJq9XYyz9LbmK+4OgmFX/aEeGUuh1QQ0hRiS9VtWFGBtjaiNsZpuE5I+Ef5w/Aoni+KmrgxLjE
B+rvM2HlnQ5KJo7oLO871U6Qr3IGojUOBC5aGsuCaw9YFgFDxY4NKcEPn6ZGea7lJw+T+YyDkF7m
0iRT8ab1dzL35aYCzsXbsUQfEeELjXYyYVKhwQYnoiEhcvYjAG2Y2nPaFBnUBI9WsEYy92m30DH0
KYpS8Nc/7FliWR8USmkm0tskuGK/q7/Hs+8iAav8fgf47HcYHE1iFusvaaFb1luGkMnvg72Rf0Wg
QX91NosK5RRzvpl+YKjkdYROIOvPcr4H2L1SXYhsDhYBi0ppXCSEFwUAjtlrLo6MHHHPHDkXE+/w
DZdHJTlrjapPWPV4NCdeSfF2sl2wgBmZUAC4ELqUHK0OgRh/mZcsDOtuh90/oifecips7cyE0cOF
V2r5XBDNHvdxZsxtxHVA554pBLHxFG4Cm55MUnvon+Ba3EyHHPmcROBM6td0UsYrWJz/ubJoi3//
i05GYuG0LyLTqbIz1ECJ6nHxKN4cvHPX4EmYN99AYIUVQvsxClgoffALZgS4u/NnvivLg9USEhzI
RSapU9nNGL8P56lgQdyzczlm1V6932uVc+0FaglK0dj+Gqh/J50FrCnSQr1iCVKH7t8icLH9usoY
tPjlKPnOa/Yp312ziB7Lamu3qMcTdqappordDdhDujzHo48QlTvmHm5BYWtSLzyBSSTexCnhsIuN
o7ifaLFDg8JQN6U8z8xmr8aLukZXhXiQjA9y7w8mj7KsowpVs0hUunna0ZkIqE2qQduXHTvwAJv5
8E37Cb91w7GyG/i7/5Pu5Ei47uOBvdUf1mWrchwny1qZDcah0Qz3GQ97I3YbRQ6fLJ1pdkBraUmQ
Ej1Toit4Et+u1aaBt6smbhHLjfzZX0oZvnl/Mgmpu4qJ1NnS7nrWo2pL1TB1h8ZybYU8Gb71eNXu
VZE33YwFL3xa54LQstrtBrswyGBYB5JQx0BPTqBUgAQ43CrLJUfUgPMlu2PV7uj88d0hsJwKhf3J
G3tOpPbzhRllMby3wacIM0/N3aJ+pwgreveE+FX6gKRrNpUAEhV9QYB76plNxtuOIygqxRStkaXi
qmbN36SnZxvDwPePjyQtcU9egsWG0NBhCFIw6/q+0VRMcwYIPzX27m7IE7fGX0IEwaGL0myCFhvD
Ljss4VST94dXkEEH1dcD4CeENXtNiYcJmG/GJge++unwuP0PvNTqNIId95nk3CbigpzvXPFzLfmf
OAHkyrc8sOzhROz6YXq5VYn3Ysco+gkJDM/3cgRutvG4C/Cz3iR1+Jr0yo02VW4+R2t+7HNVkFL9
htnhqXvty2rduwdMl7I17aU8jUGwv7HoLZtNjnNImQV9yrLjnE61aCxvo5QFOOgIlrsGOkjcHXm/
kQvICEOkrlOeagP9rWHU+sSSJmi8EaSpzMZ1SG2S9BYYAHn3JR/uWckpQRI3VhoOpSvtLQJs6R6v
JadY7ZiXyn2m5tGXixz+ice0XxluzsIt6PkEC56ORK5QwA/1R0/uxU4ZYHDBnnwzReHWGIXZtJvl
3ZPF1XcY9uLF54raBxhJT6d4IEpABZVEKu2svkd8KmfV988cE2xmJL+g5WvxdK0iO7kPHbyNl8uj
ZuGdG0N7BdJ1g/pAEOLpPXXzw/HkwJDjbz7FQ1ogTeBNLSaSrtTbJ7ex8YFIuOk1wqb57QcwfMbb
R9sDqbUW1YDR6ZyJ5SmlBscbVOGZyUIS8U0VwvFVpD/NB5ElMHvbaNgC49s95oMikhlbxbwmtTS2
oMug7OwGoTOv1YUD9sz6v2k1nfEWkMbgeTEgNG9ddRMlzU4T5L8AmJ18fhF6FZcXFo/jDonbqw7W
W2SRHogWM8TdGjiEAvEeoClXOQuO0dVmVMaz1mDkUfsXLIDWVth/rnIalpCIr/CdXqO792K3854a
9s7I4cSWoO/dwzFseaiP+pmk8Xs1v6olX+xLLVi6krXrb/JG6M9v+n7nGdqgNg7zJkCKEpb0idK2
Sjn6aa+i7wpHwZOD61ipOahBxGHj8gL1dtyBQA32zUfyndfxIIKvO41Jq66WXEvshwBHMcSYxuE7
0vbHRTX3Mw/l1w9GYGeJXL2VszkG5am4Y5N4dT14i3r/oNJSvZ0cDak8AdTOv3T3ugCeMdNu+wix
3rqgaPB6TBbbo1jLN91j52buNoJr22l1SG/xtelZFgxTHkepebjL6X9leVghTLqf5Xi8Tn/XFylc
XxpACCRLub/21hkrhx8XBLhw8wKC1khOE540yQYy867c+k7W2Fwyw59afjbM4E+JeUjx6whC2BEV
Joa76OLMALz0eO7XD8diVEA=
`protect end_protected
