-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
IHrDbq51uCMHvZehKdZHS4TCbYUK6AmK1CsI64/vIhtOZJGuPScOja0i6JafwH7m
dFgR8PvA1e6VyD9cUS5CzweOHxlIxsRY7KnmBctoaAJzTCJITlEKxttniK604Gm3
aJbc+LXL01vnKLzZup0B3Wz9wZqdvh2b2VkpRZ3JicTEsoxFnJOSaA==
--pragma protect end_key_block
--pragma protect digest_block
6P4oDQ3P3ctJ3MTE0BtawFFyha8=
--pragma protect end_digest_block
--pragma protect data_block
XOg/uvrw4/huvlae2UW300Lhi0b+Dej1mGdKRkl3QDRreCp4QPRzPbRole6fZK3K
t9Yp/s/mWFFyABy1wfP9M+dlCb1NmW+UpJ/FJLGn74Q2vbHu4sxfNJQ1lsv1shQ5
qU+EdTTnECtHcbNfj9vWXgIt9RrQl2Qcys5tTT+8ESpNTZSTSftcisCAZhUXmicU
OGlOfpqZwKRAWo9AFzb49skvyuoqWuKtvQdNAuK2qiJoOYPavmavA3hKB98AA6Oz
G1fyPEuW9jN/a84tcpjF3tatVfZ5yAuGALrMVaHLwLgUpmSL+ZIX97QXlG+II1o/
bGLvMtkLXqH/51xceDlQtU7Mh5g67zcrCmaxbd9PaTzgwV4toqUe8+B7DOKZkoPa
WXy9M8STydU8FsuBxMYV0rxFiCHcOy0ODsWhekrkpDCxtLW12DAmuid9DCnDBJOD
5t2FtfRIz/FCNQAaBACB7FuZ8/8wjeclAtTWMgj7Ts6WQAg1vy7HV2YmKRQvUXAw
1KwDe2F2HFiIBFTy8C7GDK67OB6CDtAdqNTnIQzTrXfk7RZJ6k73n3Mw7StXEpbY
DdF4CuTGi5+tCrJEjrF49MK+wBaryoQHQUtVAshu9XafiLRP9yam4cj2Q7fsPP5P
Rdz/uVY29/+6qOc25ddeslXQjYFs6TOTLxpTNfaWP0d7BjF5hVekW1Rwyorews9x
eVkHEmVwYN5dtJ24BHsWt92SFEjPTgTaNPMpKZ+eqkHInIXZH2DcVCtmTSZcqwPw
WunfX2K6d38H2jTA+hnjpsaYouKRxUrgItzeYhlh9rnRdOFLgcAy+37HkQRZ99QQ
4tk0IBxMzbPiQXQas3JDsVEbpgWHaEjxv8tbZS6qHTjlDNkKD1e1jhOvcsU1rdna
VEYqayxpqgvWryPThgU4hmRDIb0wDTP99XLstjffgO65VBQl/IaqeL3Zfk4BLn6m
2p0+PvZhhpAYhsfXydkEmPX5U5zJ4E8TLU+mk2EyIKPEb/gVu/oXfUjx6eqBwoUF
HsVB64sgqthrw+RhIH/b9G1G88CUKxgEwy8SsQGO5fFy072UXxyXTIa/WWwbrNlq
srkfCk8Ubp4T7V1uxa6roT3VC6GwJPhalC0m+M/AzSy1C6tTTdG/zd5Xd6ZJ5wud
KI1bvoq3tgby4eCy1JLGP8/RW8GfFC9sEvmU496XfJcNtJqCR5pXdb6r4ytCinV/
iBLmS3PiVocqewQLfXwvWvKPnoJNECJq2OaApMEf/JDTfyljGgDLeQKcj/V7CLHB
g4rwtx7onXIayQkm/4m4Pr7lqJsOT5FvurDxmX1OlN3maZRfNrr8hwMV0MMM1y28
JuZyxVGuN3bsBxS8ZTItf5xmZ0zzn0kOG7R2krm69IhDye3vLKWYgvHk2dMmavHh
A8MAfBu3NLesoLnTzwsHO7HqtaWfWtgWnH/oYKM8us/CnvoapHduMGMC+F8W2YCs
PPJ3ZwMiMjXpuEAc60710EiSHUhRprP8ss+Xyq+H32P9i970v42jZHAnwLnymCHD
YGs5OMwZswiCH/ZSAVhI+8Wg9iY9frvTDFmhTkswb8BeevUwWZCc8+BFPbfX4LY1
P4p0xYg8EldeXDUMubv46w6h6UAx++VEcpL8I2h8qkXPmr4cfGffi6bP5uGGLMfD
3LShclge/PtPBBSB4bAlcpR762oI0RxHJVFAKO7d4pzPaPFzD4oUleQQl3OC+okF
GN14Rs7lwEjlZXRBjJCgIHtyPnYf0houxCSU704Dae1MnLJZTK4WqD/9s6tR8AZ7
lK7Cd26G3gfvIgMImFKjV2/nHkAisprDUDF9CP3PEKbIRgVvtKWA7qa4OiNrx81g
rgMfrgRd1S7DZmufvs7kv/D06rnhq2Pwroj4v2ChvncEFQRvK/YV8XPTFwBgc/83
LOiDEX+bQpDtdGAui/x0bBe9tFbaPyolJ4Batj8KjxJ74eonYCxJ3CjyhuhOv00i
RfFsteJK6vxF/2gLIrzyN7ZZ/QBCNipnJRyTuwqH5WDWqZjci/yFRNSeku3YHy/Z
nDqC8n/V7R81pg9ZdDMu8Xg2jRIJ7BzbZO9+Fll+UopBl9pumviCzIdOguMPmMfA
iQ5ZlUX+gycxWMhs/dMPpV2eEYtzAAFCdEhZFBACpVkdpnJUDFC5p3MLLv88303C
0/SrS1BXYs6wSB21CwidSxPrg/9EXT32J660GQvwi8w/Act5OWXzJ6qqb1fnfJOH
lL1uqbxeY03cpDdFpPiHShEjN3qjnLRghTjWQk0bkYS5HFAZTvYm7MGJq47S7fir
WaQ4pecBCEmq0e6r2MpBKA2UE1tDuBUCjIADsy03kDdBHemlEsTJeHa8ExXz/5rg
UFJoXdQijuf88bDH/MI9iFY++HJTYxYdPDUnWdTRksRlH/FyCrofUvtfyj9wSlAh
PObEsT8cqN8nyS0wKvjiBYo8a1QM5HfckikJPzuh97sEb2iS645DAnYGTVfmj9bZ
Jit6EXU06ib/My8VF5GTjWjR1QVDAKhQMkMfwrb/mPQDOBs+KfyYymy0tDP/m0GR
mofNvDBiCp/oM8ZZOFjKXQCsNHw3jseSIdMVWOZuTYK3fyjAlS1Ewl00N+WHuGnd
4gK8J23XJxU4gftl3SaaMcWhH6bDY2nKn6jA8U4fCxbX5vRN2GzU1QBFxRKb0yV8
i3QBmcyBW+0ko4zTy5dZI5S7134BpOVO2Rj6FcmZInjzrUzIMf9wf9lmctO/Vx7B
f9+jVbWPVK4TYYua/Wf/Qf7reDuER4YLBcfnpDKQA3q/6gFZ89x4y3sqgBOyYjb+
XzGzWkky0w72yluBFjBancw4sZoTA1Bttm/fwQRpfdxqS3m7neGVjQw9tu1JyeYJ
FTN/i/mff4jZbl1akrMBw0dS55rfVahiJlHVGmPli1Yt4ZKkQS1wh/wHRfElb4Fh
jUFl3Vn13gsuReji4R3Z8iskUQ++eL8tOzQlHuO32U+wY5TePODBNcp942xClggo
t+xwd3KpiMKHdu02tU96AjQTZt9MptO3tzg0DAWoAZUvhSQgQJ0SUhmvEEklWA6X
/5Lmv9sFIPYUkBwsGyqxkqp0Oz98bR8M5MXvI5JOoX5jtDvZYek3fhr6Jko044jb
ru30bt2PnfSNL2hcLpIWtZlsUesbVMCjUxBABsKKz46iJB3XdUO/CuMzrvcrPaPH
+VuAk/ETGGLUJTH5GJTKQe3eaMF6IZZIpryoz9Q+OVJgf9f2n1WKMv1+BEYUEbOl
6q8VvLyegcbndsD3e6RZK9RXRKyOqebvWOVlZp02TgCE5qleDjPaJp1NaT928uDb
SxD1SIxUVd/O2UCCN5RhwXhuL4az0xEIUz1SZ+yWMBLbxwnFoLiIIV8mYc9KjdcO
i/InYr4+pbuvGA+jgVQqMiTVs6eCp2wG88Ux8wO882pQ4Eh4Z1zBBp7ifdaA8SWb
1uq5OKBkNx0KHimpF+z4ALz5zvgA2go5XgPK1zCAhJAbDsHB3kkeMvxuKW/8u6O6
Pt8V15WgvFWUn2HvDEewuHqKy9Uf8qsSr9vW9DrRqxFfBD+jhe/DmcfZXT3zgEbv
b4VL+tkr0qqCXcKkcnYP2lHs/OrDlOEgrTdvCdJw/u7iIRZUuhoHc7XdsYd5D2mJ
anuK3aBHIVLjVZ74tpPbimU1pb+QeGjoXLwL8V5GwbPlldqCILRZdYuHrNEgWOqi
HDdXNLKSx6dyeCAQ0Ls8ZHNOtgoJK7sIPMgtiqJxYIl5tg3fj4oiSEm1p69LExNL
HHqUgJ+dzenZjbbn0QBhfd1O1XGoJz3Ksoc3TuXVOSWsab2CYE83iH3ssUOIZfQe
aJ8oY/CxQITlQLwh/ZV4u/1VJ1bSiyBQnIQXWhnyEubTZ/dfsPV733ReVBMvh7M3
9sVyfgjMEAFy+lZaK29zChJIgcvgUt5RFlEi7VXhWzpZr4TqEQSwGBMon4bIvAL/
aH03akRkdHcsQftOJb81Pz36jfNr3O8jU9gaYLNAaU8ibd3dl8A2hN5NMOzuFL9o
P6IOIaOPNxNeukaTNdE5RyycQKCFz6LYOWWmWuKtBMo8RSObjKRBM6qV0IOQXFZH
Ae9dwj1LLT/p+RTHDAcaD1L6a8GkZIjba7BsC8ErSGN/2yrJGCZfyDGq48lTJ6WS
u4UxiUr9vlFXsKKOYvvYFYLRDPbhUH2D2TpUulahhSOHPVucjhQlYTrjPIf0v+ZD
NnBxlkAPTtUVl2gECPcMJt1rLVN3gAV+2mgZ6VT6k9YWTfT14Q0QEMMV+ViW7Fr+
7ubcISDqOLlWwaZF9eRUxataunXSnJHj4p/NVunXG8EvHfBpyOuocZXBIicZ4h8o
KK1sClcsjcE+TXyK1IahSojhcaWazWNhvl6TvAr2vblUEDMuMAllbin8e9jXYPGT
OFnQkXImL2nKnI9c4oYhVIusGHipVdVeKSj2MzMcaUR9saaaHN5cVEwegAQbnRTk
ytQW3eghXKESo6Ae1JtfVekpSekczOF7MZB3ECWVZ69t/sd6ox4wzr1nWb9ZLvdU
SNtXBo89uNOBVd4aP8GMXRq8fy3UZ0YXtE0wKHpsWlGTpDoAm83Y/qhQCXeQyDGT
1TpflkdlwxaoRk+HCQAIrDyyfu5/4FpL+5tIOq8c0RsZT02AVRRvwZbA4qQraL1H
/uOPwnj64MtdyierXZSyW2Bi/w2F6n8igc+xZC0p/ORjKCcgpyjo8bWtZJKfTKxq
lgxL9wWrxP2ez4oHxznVZwM+D7WL9p+LK5RsqCfozs9Ydnif+cZVXjd11xQ5atwr
yjd+w2mC0WvKVRaUZ5eSv8wlaIeXcKr+5YJ/Iygj97zEKiuUbbQO9vIJhg8hhOo4
2gQPAlnSPn1h2qd5cH5lhmcuVe64sK2TSnZMZcipak9oaO1jzNapnx+ZOdaQcZ86
n4U95VRb4a9HGP7HiJi85VsLydTp+P9pDneQ6PyM8wHpkwjPuA5o0VkYEbKHb99P
X0glGN0wNfG7VbXCHNbCyIyF4DwQVKFkMPBcyau0BrxGEIpTcjydkdwhRHHP6dOc
klJGqyewvOkhxiqnEUN8ptmYRo3Fh5lhTrZHDPq3DMSWWSJQU03t+GEuE2As++Gf
pyTbycDJTukn8oAqylDUGKXLNBNeR4qtKgQgy4llOB5L1YJw2sniS7wTvGn2y3Z6
QQHpANa3To9RitD/ECvev+PwPRvj3zcFS7QZ6RMlxTFKcZ64Oojo4T2fvcaL2u9J
YVa/kihfv81O8Zbzvi8z3vc8j/GkNm9eOKgUnua2GQibbgzGVqNOmr8YQ+bkl4xk
N0P43/xPPKIGj606wgrtAunk4igHkW6/pkFScJTbnPX/Z+oy33OEQkobHsF1XZAY
tS5OHYCv8tPP7cmkxiGeD9h79qJbkiZ0KqR1xH5Rg3qizPBbO4r1CQz4qZmJyLQy
+/OmJ9DKl7qZVRjrPFzvbfv8PS6UKqFNfw3XN+WWzQK5uUt5MP5wSRo3Wn04hMlr
yrnbC91HNDyBV3VdAyFPPIoUywhMg2ypAxvvHfqZqHvdw3OzK6C+E1TSX0YSQsiQ
qzWH3bZ5y6qOpE2KMBqQITJ8crA+iQE70PXEjTllozhTLGOex0MM6a4/4YFugTR1
MoyCAXqHIaDoBWrD0qgx/XB7V5cyu1pzIwADtKQ0Mu+zPlX8dg3YNADH1F22sZ7G
sNevYbE7kWstg//INE/ES3dTnNLUyy7QcZJB8ahCsOS+bOF2T6BNnK4dn1n4320x
MLLZh2oaGQV88BftRNNfAhmaE56ZxxnoVRXaX/vqVWDBDt5wzRWTk+FWz6z7dsFI
9JPxOeFQ96DaKyQcU9I6cNM/GlFS00gWnM4w/u1UYzYJNfy3uinzSXjry2m6x3GY
uBQxhh1haTNRNNKqe7bVi8q8fuzDa0IVVIL66bBKZFg77bLfGXhNc193sU5z6/E3
oHNO84RNS5IENuXzWR/bLN0QE6i/0/mc+v4arcwu69+BKMmFvs7s8JjBT6isacPs
cZjHGovZeA/mnrodcwl8p1kt0rlmKPMPVSJs8VwZqSXiICdX/ob1JnGyj9Ru/ZXQ
Eh8jWRZj+9lHCZ4DFi6ZzUMOLGZ3VImGpzgaFF+y3cWySQoMm8nObHR+o9bK3Mnh
K9TreOr2z9ewqqXUYu9ktLW9liIh1cbnvV1Jq5uoV+Sb6JAcuwJF5ggQ8pFQSBQT
E+DQUgLF+3iBAQtESMIQDYpmKlpyDeDgyPdmei5obEaQX4ddlweWSUsbudnFzaff
kb3MlT9D8SV9UWpbf/Ew+jNOYkOXR//M0uR/W/29+693d99nqyY41r91YmBfyGmo
xjcQ3TyO8l6Y/fPUZGpBz4orKbp+onw83cBmu/2yAgmOZiR/Tp+26nyYC2vfu2Nw
S0TWX9Ooj8K4dajS2/pox4zQxauAT0Qb8Jz7DgtrnClVgeWnpnAEKR+zRTiKJQXA
MkLX+yQvmz7FqGkhq1rPSs4nXIhaOMeh8B6Lx2urOjZMTjwf3GuGwuWSRNjHveUm
EGggTkUXYUW56a9LqeJfZA==
--pragma protect end_data_block
--pragma protect digest_block
A0uYoPvCfL93E3SBWdY0qhudTv4=
--pragma protect end_digest_block
--pragma protect end_protected
