-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
/1D+mLk4Uw7KZNAN0SME1keGchhHkcZYdFMevIOGNekXO1MzGd74QrowKlqAwk0r
NiGfnERKfcFWQ+ZvtiOyssRShCPMOW06FqNy5lLtXkRhGzZnygsvtlBijkITPwn2
2nPr2ooFDPExrKjsHnpIAr47l5njeMIumI2VwOpBabDmHp/vAC2Iig==
--pragma protect end_key_block
--pragma protect digest_block
//wAz00YPUWq6w8bnf5kkOSZk+A=
--pragma protect end_digest_block
--pragma protect data_block
ZtRc0pCO892N3545L2ETd5jjDtRqvwbInh0Oboh+bz5XzPCpepDGE3eOdGgJSgq/
d44pwd6DCBpWOEE6sRhsJwt1zSfxxhcInOFpi5e63rUwawgzr40zTsPm1q7Bmjio
Eu2WUsGC/5XFei0efMQPZ9jO3MVogCEDr2Z/OgUpy7PkshrDMiEpGUfslKZZpvHF
0isPKHC+jIUTlh2bZxbUuJuWFzgBoeFT6FiS4PzjLp7DoCRRHKqTikKJ9IJnzBMj
H4MX0P2SCkq+ab2wTXv6vRtSBH7Ns7TQct+tODXT7J5miLG2M+5Flqi3X6CxwoAL
KLxxsDaYKK4dZTM60r/S1aYu9hDqQciv9zRlEG3BOzQhnkE8eOhqgBow+lPZpe90
y96RHeQoSVji37KO4VPdDW4W57k2OOK9TGebfUsxPSWziQPxMVJDcNKZkpUoJMsC
Mwe3tjmJlimKL9y04WNNfjw1ugE1YwG8lAoQtvwHmVoen7aoEy8evGauVbvkTbYC
75mAVAF5wxessrLTO+sIEJ50QMh+fAZjmBs/SOWrcpukVkCtYIymu+F6FZOdAbNZ
dKJTkQaoMcrn9KxlC+z9gW719xhlrTj0mZTkgyY8MCgNh0n27nqQgSr6nuzBcdgM
GsAww9nRLovnlb2FGvvIT+UmGik2jOyTwwkT55mWAOvAFa9x77x5XYqOn44k0i+A
ZeCMSGx/4BWlpRjwMd3dzoz/XNpGlMJkNflu/V07rZHNlle+nADB+BlzQxoL3gk+
3fD0qoEYtv7idlx6Xpw/5fBGi8gKUCDQ1x++KaSg3cS5Ohsac9QFClSKECgdBC/z
V9djwIdJRlhnpMocfQkRmobFYzMC7L40Z0VMS3nv1p17flgAnKFUBNSB5ob0T6+e
ggzArWnYfXrKaUhaVOU6uYoL/Rory3yQzFo3531adxVPfrsOtXyoP+zN02ZHpsXS
QrxfShYsLWH3Jx3Qg2LCLwUo/lbZRFCj0DCTmuaFnxXN9tGT566JR0ZTiSrJotFY
sZsthqi7JPRQyuWREAwPqZoskT4n7XrlsQ71OSb5READS5lrRK21Qwnq0+V7jtts
kLdMEmF2zrROzBAcA4bUj6eIAco7dxetgJ9P2F8BBbCux+xrVNLf4bSHIPgzIvfr
lGfbxB5oagf3R2HhmH0JNRA8gKoGzJSjd9ui7JPTen4uM4fisgH8fPNk3YewRKvG
x3R7I/SUJR0bYfYjsi2QXZNfMYUnnnvuLrDp0Q2e/qUML4t8s6lWHqspXU0ASCdx
OZ9b8zHVxmobs1EAg2eb/TCS3l5CwQihS1IvxmdmDdrywkzd/4N1O6RX+ZXd0iWi
x8p+XOq/6N8J1Jw0V+W0gGrGdVucob36LqOaxf3+IcRjVc06mZtSlX+wNyOgITR0
jdX9wTYLCSXkn3Bc+DjLjlcWOJjSaewk9+FItmon5WRnVvfmZHbenZUHObwEG8OC
7O2UugvWPm+spXmo3psi1G/k9hIi0in82j931Mgb1XtwLMjXZQal2cyyLgiSPw01
JHfRhz4TEq8hCfNnY+vyCvIKRP6ibyOBYtN+FpG7YnilJDEoxWX8zblr0F6mQauk
UnZfUUOL8oPxyHty/FiJ7KaW1OPXP7RzTOZzatELiyx5NlffsJF8Nc8cp+KYfun/
EqyJI3Ovu1mhT25ObI7/EwNzUvPrwbRy3gO0XnobfW6j/qtmxqyhItXZx8pqrU43
R8sFkiRMl6jr/4QXJQz+B4q4n3TkKeIMblCcSJyodP0BFwQmY+bBw2PwIipMU8Yb
1SuKN+1kCqnvf4cxQ022EvsGmZt/rbG8WSS6X8niAz1nok48KA8SFFNKBoXPsKo4
MHN+oaCYCg6DmYjrF8xqyUJQOi/HVokE5pJuMNCci2xlE2THtTdGD+iW+30GmnzE
up81QQDHD2Uiz3770VM1Vin86eao/t1huR3XFbbxKy+81BnameHGSmW5sPEiywAx
FAeI6R81UVqQ7UEeRuRmClBJfQkCYr5V3cG+bjy2UhwOwCiQkV14tKUC6xRleFzZ
LEYBqQH4kNVuyk+BjTmW0vRU1scx6T5DOqjP5CtMMIiu4DSg4nWkleyQh0zv6W/u
w2o/TVFiBKruSheem3WukgHy9Zv0YlQvCB6HxsuVmMUqsWgKva3C/cEjcUD+jNns
tKhUsz+OT9Cg8+HmdrN1GUX/zmEyPxVX3v1QkuN4pDCDWknQycW/YnumCiEDnWkN
H7KXWliafjLV56QIX8tDf6b2hweSLadcbIco4M2YNZO+F3JhQ4/CJ6vy1xmyBiRU
G3ErANDeZdGc+JcT1/OLRL2eqEATkqX3tVZdIUeOk7YxxAg8R5qELnw2GD6bMsJ0
F482kwS7K5gHFxXiFZq3evw1gm0BP6CqbhTQsu9WMhOB68B5zueqr1jXwPLvZe/c
Zdnjw8VeSEQ3RPERMbFXtWxCMONDjFUJiSVCp6F9TWgnOK0Nvpizfx5zyoBH4uQ4
er7+0cO8CRd+WFsmaqy2UFIdGwPaMKvgOVdBT7sQqQonnNslT8+dGnSW4Fslujgf
jOax3suTh+RlsYMacuLTTge+H7e4pbpw9meugORNnKAcitFRbyI4/EJKn5nn2VJF
dgTpcRtRvsunhxdtRNfGzYL3mAVzmQmAyyODmCEM0u2ZGY6F2/W3qiKro0oaIHep
qKgTnTBXypx74m2WYKXgqhD7PpH8jq0uMMyBG/76aqa0pL7ML7odBWlEsElfwu0Z
dZY7wAGU1++MEs4BacNybmBSP8h2TjxIL+AZxY61fAg39/PFCTYHO3q9P2TJfN2T
0DoBEzvSLmG3HcXz89I4jWGKPNhxcLJySS1ku6zA9twSWH/j79/LyZs04grU03Jh
BpSOUOoLfeELGdI+IQ57d/Wqy7FZKsWEbtJel40ezolrKZXUtRRzohzxK7Y+P7sE
aNZ15eieVTSXfvRmBcNfJbWA0mSYiJYqZM2bEpCNb94M+WLj0uYXkquUlbJqUDGw
GIStV6yitEMj5Wl4iUNRI/c/NQ8iNa9NUHVnEtZXiubjRnZ5tS0YfL7v06D4nGV2
wpFre+3ej/54kwU3GdxXbdfxJfEPRAygr/dLcoy4noRvZ1M8binc3Gb1YrOEryYN
WNx+y19aCMOhTbbGyEGlsiAeoEbZde34vfKy8lgZEAlsWbtai9lhn2dzTWZ7aYrS
H0l0/eVJ9z7+9f9UPjcAcaIE9zmQbLrgm12FKXYgXR9a68MdU9nAbDy2BWLDKuKa
mUDML097r5OSeYKzd5LmqJptAqqEaOer1CcfiUHgbIO3wwDMz5oEkp9WwCS5nVjQ
SKEaEM+qWYzVPzI87LCnE0OrELEdxzYh3rGdjEiAsCrsdRQ0ea+vHISJ8MhxD+XD
wVrjRL3fpz2DLBChX/0c9IWKFX5mW9rwSZKMKW0sl/uptObahicYp1Zmr2lc2ibZ
dbJSHo2xeLFMYFdpp7XUe4YUiSuBGTuR0maHfFSH8R3wUixfIIPqGc8cHMGL0sBl
MTeosKEDfchmThlRXsIV59qxQwIRZlMeNOHIVr8GuoiweNQBljT0Hdj0vi2unOG+
8Mc8yQEFgCu0PCc3OooNxaHY8x0mvStFYC8vEiHU1c79g3/y1e34vSDZu+B0P5+0
ShlT+iUYYADWSoqCK0DoDzzKvYnAAW7Us6Z0QbQvhvwNQrb/PU5Dmg6o/Kn+JLbQ
vz6hjbBgt1mOmrQBm4fJVd7vrpZO7xmsYUmjfqrsGuYzRXegLjqPjLh2krRxqIdt
YdVrVCSgQl1TXfGL0TSxFGNqDxZItXZ7t2gh8vitttJ3yaPYD3lhe+fGHct4YIHj
uTka4I29Vpb5Kio305hocz+BFob3kvWP6F7DtNwJo6AkPim0BFqwsA1GpJLYbmw0
D50mM+pfP5ov3nJt9n0ldgsu6syxVE3c7D2n4lDCiw98yOxukX1I19BdAVKmN++/
RzHctMXKRpV3m2wlxPv+N6MDI/iBhSthJWQ1MUd0w+VFRCHAOD04zIoSgzjfLrC+
3cTDIwNxgzsjZc6lo2e5vhxUaDEZRiYAhaQ2A8XE/Uu4V4uCoQSNDMwCY/J6+xCQ
GweC9frbak17fmof36/O5PtKyGZDZk+m8LkwSU3GINWDSt3wUWtkWYG1iSRSNTwc
kWbJwULb/JJNKqeDInVbkTCb8A+LwFpyggl5vfiPid6p+YZyxe+e4OZeiqxUjHhM
bmGI0sMZoS6EpXf5PYFHdQWVRvYh4EFezEyIcdRGPQkeH+xGB8UeGXA7VTKN/cwX
76cHFrruYGpKyWCNQFN7AMfGRqnMgFWCvlhRI03fkHU7OHUEel/H66PvT4Qytq+N
IBD6/YOiZyHr3y31U4Kd2txavkGgOU9Cgs1Kpe2NNJ6+eguztY8/MqUBhO0K8u14
p7L8qBEZtaIJE2FPFDmTsfaPjgtYWigpu7sG3e23/cg+LoiPZxBzBoWsce55j//M
32muS9CRIAd5FqtSiJnkGBW4/dClChQiQX+7RsT4o9xbYyDZ2Kx+Q4WOXsr/+3qy
lXPQ/OgL4+wCIGZFqDF4psis7cPFfNml5gihOVKZ9jYh/4t6Xh/2qW5UhaJrlbJ5
h7j7/M/bZ8OWBAJBgwGntc3SCj5kJzrgCl0N7UtRVco1LAFnaGLMKVUXY0BPigem
XNtgFvHetkwAxzDN7hcS6ujwL/dJ0ihOojEWCzKibgDmX0G+gsk0bgJuVBJjUvhQ
e8dxylnxkiau/YplEVlBYGu70M1xNQLEkV5Z9bMQ9dkxGCBVYF7KJdAa85s4/cfX
ePqQsNNjbWJfb8VzTqUwyD4ZuHex3kInV/5bxQa6XRWOS2vzfgIOlNlhFrkvdvjD
YMEJO/vtgysG1Sy36QXLu8ppX9KAtQmpwwrm2tpwy9NJNgmPGjcgCCUvWQvKars3
Cn4MzHeCqjiaBWRald6QeQBX1w4P9P6O93/yW/B/apbTMTVOprz9e2NXIM1n7kq7
3qPnk/QZxZdiWh8YWHMlNK/ikbSAC331bWw16m2PRFniKEORgdJ8wmf2G9u3QuS8
Yz9682OGF/z9GOggZ+w157Pk/gPEfGMZyEeyqMKTEQS88ZVsvUN+u4bBanHdMwG4
/L7q/6OKg6XS9+T2bXSxFZQFegtfQwzXJ7/kfFS2Q1GoVSe2PRXjCAWPuc7sk/W5
aaRN5PgxozzgoLDP9ZaKNAlYkZ20k93KClAkd/66JfRlycszoRlxXH2eI3lphJWs
QrTTEQYLp8G8cQ03Rhwc8kE1SziR+riY/227mCXkEMSlem0I70NRl50qWa/NzO9E
TbVx0Y9kFXt7lR9jwfRXol3iGXjF0pfEtCCvwd1MboE6ZD3M/MZU/IIcTa6nJ7hb
CVYXz7yBQxHzHdxTdL6HOPz4rcC8b+XFPjg6Bzy0pcapI90MbdVWTb6fiaOJM+5a
YyPl+FQM9Y3nI+CuyRhzRvkwFvYfEaeby12D3Vfu0B8Ha9H9IppOxWihxjsKtofT
xwhwIWq9SVLiIpCIvkY5kcDNB6XDWysUiDulGpgv39rYKAkfMYzjMARrvB/AokNo
utIFiD03+YTJ4byJaBYoGkVOGDoECDeeV11jSDd3rriiDlGQXU2fTntTPPg5CoFa
ZQ0CgO8C4p8CD+o2+oDpxqLlrOvPaNfHnCT7hemskiW7JqmwGAbZNp5tlbx/jJac
Aab7x6VgYbsCEI9rZECIrCpNhDpMeI2g8mpex6A2oQYgj7zZ1sm0C0Sa0OG94g2N
BQVKlx9BcRuAQX6DTuLpaa9/zW0+P7L6GvAyVSyaas9DoMEb+DG4eBOnrVZ39r6s
egh8tTkEMiSNVY8yzaC6oWU8pNEFQyjTppCPmMckUiM5qr6QxfEFkmt6i5+pVylW
xwVHSsMp4fvt0QoMrePRcVRWD4/tl86wL/LjKALHVJxzYOVDgy0dzREdJd/aHNme
n9V817o+BX8sg6WYTlZpQU5+RZCTDJDaxZN7dRwiXbszk08C5M0z9knwH2eflw6c
BlQZ2pnD+R2zwt5F2vLSQQUr3jnfR2pjuHfywFWpjzpfQuG+6BqtXzxSNlzaxaar
qv3CRwaq75WKQ6chPgnSlshdNUwRflr5YpkgdPbzwK2MI0nV8ddsbKhNHl64/MQ0
2nkKLZ6afIkKYK1CnFeKoXlRN18Rq0+/lw7H2DMB4OdwTmdf9xU6SPg1Rtnt3Giy
hB/wWnW3QuiJXqPKbaRO240sAhdlIGfG1wQL94j9aj2M41eoxaCO4KEI6Jgu08kO
6kCNrpEbn8MyRTZfpEJyjnQiGNMvzA4Hsl7BUQJbXF9MVYl6J5vmi+3OVzqvUXyP
Tpv9rUZpHJXhlLdcaufyzwO8sFD8F+opnX349h84yXPBXuofOM6MiCCMZqb3Lby0
GK231ODn3DJARHDQ+Hvml8H2hbIKXaHRvfNRc70G55EH5c5ttYQKbxEgtJFE1YVK
Pj7hV/VhpOd84r49ZGz+IXu9V+8VLh/PeVw7QzQpa/HSubvOmcs1e7towp4QrfST
5jz2nVwqd9Nva+HVLpxe7lsZtQKChWwaefDL6oeQQ1iu+eBA9B4p79rj5+rLenHH
8/5AzbcLvnX9KAJxjlmfagAGNRIuj65uBcglOF3L8Bn5ObGkw5aOj4C5GyzLyLHQ
MizZ5KsITuRa1r/GUqrnfuJwX/E8S1sLcTc5VQd4pCTcHXaCgh3/6zlCNTGRGkPS
ih9Utf+xrE/VCJ8rQUcYHFmdeo7fNbwPw2Wcz660xW7/9znIvsuWOPlw8BtLLdX0
EnFob61ZAWoyyezOrQg+SJ3a0eAPlvXHPudX/m2csqMV81t8ahna2i/tWb1Pa39C
RDkvrsLj/f4NYxqKFWBtnZWzaZWxnj9/9bOPv5COu8BvyIHFko3+gFXpePROSpOa
w9tiqnAZwrrk6RB+I5VSZK15Ct8ZJVl5LSXVYbMY2n1I3I78WLgm4ZwKF1Kd0ugf
o3AEQjVhHuGdvtoUVfG2TGXxqUkAFHtll8Heord/UoKSzYCnD+9vWeDu6TKaMVcn
L3I/O9JINSxcVLVrEL+aTbkJ1sATcfoR27RAZDGAXEHB07s7xyx5lynFLyM5LEFM
hhQp03Q4DjO0K7ne0+3TUUObTJM0IevZCpGsNbe0d3XVCvOQBR8xpkPahdd5dOl3
NN0X/EpQuA5kSCRekO54OxDDjHksrUmCWrBOQonF8a9FgOGIqpsg8RsnGtg2fiRT
R8rQeMaFoijieOKfCNSwJDfNQBm2SNM9iDIuJ1Vyqijdj4QfDLTUe+ra8/BgNDV7
YUWU7sdSbBfSmp6C5EahbZreNdX6sQK6nwq5xa7eZp+773tGS3F/u6loPnkfuBq9
8MpE/y8gLFNjAoFudIHUA7r9Tyu7f5boQXWVkC/oGiZouH9Hml/HvnqDbp4jOGlR
oeblvjQK8hakTg5tqSVlA/tAhcUFquwNlhGk4ncnkuO4qLf6SmVGQv/T4BAwO4wS
fZ3F0GkXGUFoFc+KZ2ysevLrzxEyn6DRKZxRMri6Q3V50AGRyipyP+VaGJIqSLzQ
HhNRThUSZZz8lYERkJfHhtKmMj6Unf9AdV2oeDIT+Pr49HjYx2cgAWeqWwj/aClr
kmlDqpq6W8nMCDB6vJi4l4qFtC/jboG4Mw14KuGVj6aYrTMb50SjAKRf4Ct5Ylmk
qM5tlxDnDSsbPGWgobc5MfxShUvkn5ysu+v4o+QdhFvuTwFRgXCWFPYxvQKA5i63
6gPfKlykfakjoZkp+L/uKD+j60ZPxdd7il1HIRqdlJ/JvCbEgAQMpbfcU0cIHd/A
84CRBrjwTmYkZuA3meDCfCkIKKl8CPPWIRys6Mr/+A3vC/0ieonpTteu0yIxesZc
mqurUUwD7kUm8CpIuEk1HuDMg79H1Bd4SQ0zKg9o/iO6Az5HXc6JpRYHBXB4fg+y
gDTJN8evJ1BBlHepHhFwKQ5RbavRlahDI0xiPMxHhvjyr9obxQeERbTC+YrIIFYx
Jcgy3zLFv81AweZye4/+xwQkNwADFxZjK2x7nflOy0UV4Pk8QxDNV4g4d461cV5s
TEl6f8B3yAI3NPaFpkk5hJN0nGfAmJY4F/io559ZLNTKrYIH/Fatp5bDv9DCRYuu
XFoWFzV0pqdiArOGkNKN62j2P4ZDuAYn9K7+p5fsJK/vc2zdPmoFbKxIS05C9Lwd
j7vAs7Sxi/Cssk/vclXGWYF2Y4InAX1kEnwHfY3mf56Fvm7oDskhcFf1Tagou3KQ
NeMUw2gNwIngSNWw8XKMpaGGs00hu5JHMErSeM2eKCP2ijje9EZQEjwlMt7PX8Ze
l4MtHIaJ0xS2wS1A4w7IjX2eFxw+okp7qLP7WPuH8manKB4jvQGWRhIQer0qnoVB
j5VIHC6phF69A7IZwRrVFxVdhiSt420gXYmIJuwwJV5KsnI6paqcsu9vj++ggaAM
5aIQRT/12gX1VFAkXiilCIMe06XUy8E3ZULpp0lHUfvNuw09Zi8ZNWQbBmYD4aul
CeAyWQds0hipvFcf71vs3M8aLDRFljE2REhIY86kTiRzuTDG8Vqaw49q20OmIXgV
la7IetB+7hWpXG4z2EIk3cuO7UXyr4+EBaUy26xhq/LJ/SlmzpnnBjcuhUbrjRC4
URRwDw2DBAeeoWlPtjMWD6DdpXmgMZ7irtHu4jIqtqnQfsF88RvnyYZEradVJ2gS
2xuh/ILDeQQ9ksEq2MwJJnd98aElRrXr0AC2IYd/K40vVslwKVIOs1AhJ2Ebl58R
KNkhiTm4fRW4dtOGlpSywXoT6Ri0GmlcsQIsOmBmyySppI0xKEYUsO1GjHc5ip4T
CzQQXvB7D7j85i5k7IPfFF3iVtVXrFHWD9F3F/+xvsXGcoVIDHzvOOch6wvkio5b
sVEEwiexfb0GWx4YAhxRCr9YD/MXmtKAEaHKulI6q7DFniLQZvxDAyXVv5w6iNSr
zdu1oX3vPHowUjfIMpVW12egMT4fc1H4xiFS2lqthi5ywaGzZtAvCxxEIcLLyOUY
2IkTI5jP9xl3x231flvGEK50Ikn7qox84d6Oe1eVbf6+4yBcrCFoYJw5t4Ep7cxk
hCeOig3ZSR+dtEa+tgl92oX8Y4IZLWAVTf/bg58dMhaBn/E+50mbep08YAUx96VG
K2m0q3w5HfFjyoxKUVq03nSSnKlBZnIa08t//UoOstFmfPLz9PzFA6iDx1vHWqLS
/6IJwVCZX8QD7OXCOV/Voe6uzokiM2RNDJgyCzlN4ZDLvBYAs0KoHdLiG7g8JGbL
p4OrvJJovJPzEJQRQGPovijcAf/u2zpDgyNDPQKeupMqv0d7ARl57ZXyxBG431S2
zqlf8jDyfUXm7UoR4KI6q7s1cRyNOsr+mANoP4S/Vr1DGgnlovONOOjguf1khBy5
CSqM5POaXkBi43oX55Z9N29NynWzBKqMDeIQt3xddSJ9bVLO7n8MHDzbsLekneW1
ybW27cQUe5dhXXnvpwAvtAJo8QdW/ab6V0QUN3tNOydCQXoyeISLyDfYvzfJn1mg
DZo+B3Ia9Qq5aU8PuZxEEqc1yNoG3MqotopQN58nCn790jeJQmn1NcwyKzeGwSJJ
zGkv4kwdfPQLz9JCSRV+vMUQw4L/K5VPzSFHpOXvk4AqDI9wqZX7D+vxqrNy8Oid
ppQ1lyRCyLy72ugYPF89ZgIvmPG/52pu5y3cGC9C4TYegC5F8X5QpO3gwluzY9gg
dv0mYX2QI9GDOQk6oLuil6k5nFSE3TdTt7wHvmPwgc5L/ARVGfrIAlTBakc2vARE
wUSMsM9jEu2nRPPOaEonEFfC/4zjfme2kakXlmORqEz5+Nb6KvYpyeHKTbVwBgQS
RzR1rx+J3Pt3aiobou6wQk2aXj54MMQqgjON3Cc5vD8k42ixsKHbWQoYyosDsIIF
/w/N8b7u7vRm4px9b/Xj6mABp672Iv2SXvp21KsfM1UveQP1Z1W80iFB74jcHa3G
MzQZW5a/DzLlxQwODn5XJ9QqiYL0aAIh3A9vRRTFdnihdYXQ1mw7/se2UpiUz5bO
GDVFf5djRibLl70etL64BkIg97k7J6MGspjhRxoUlUKXM4PPhtmgDrz3LIrjUlER
jdf9peSuFB2ZHHODWviNcOPYFF3Pk61VgdMa9zYaLb+0cGBc0bSgUe97uCdJsBNt
yo/gP4HuZCgifAq5IXajxphvj5if+Er3k8CQAPHebbRS0N9ShfaS1sh9D6da2/VC
/ibxqAeA6ymvYQORaxM8jB0l5aErbIOZEkR88twmhzwZ1hFkYrqoQ9Zk1J8XkwNw
lNv3ovisBLaQoW5TQgImtO4PZ+fp5uhjuD07C2sh43dvPl5E4hRvdqtL6Mmfm0d8
12M2gu17x8siQ4dJCxU3JFtTZM5GEJQ2nuj1MwfijYmaJlzm99xh2FU4J+W9AJY+
/ISqjdaiyXceXEOguVYz/LdmMx5/TOjMRzWYny0v3Q2yu57e/MtALREp5lvT5iAf
vnIkoM4G6o/0eRt0dZAjP5KvBeU8JrxZP5SguRL8ZmiqJRIaOwaC+T92oFC68mkv
lIlMhNJtzaMXtQR/vnSQfnQ134SLYd768kqvRMg17Ul74o7IfD5MlZSefST3GpLr
2LuByzljCCPhAbRZLMRDXSFQdUnWXufCqORZVBKJCOLOBkSXJPL0xLZjpuJgEgE4
B8YfaYOd964+UMybr6nCo/oX+88VxrD4GkA+79rTto3C86Op1FfASJJNHQKeancT
Svl2alyvd6jun2DUHsUZnl6aGAconNku+aDUGoU4aJCQoiRGuavd4K/5V/DBef8H
Y84dXFZEk9YtFzhC42jIcAMXDrSwR3A/6XPEQ8m/KgqGjioQgDDPm9XQTYUskOCc
2jH7nFmW3hMBOlGhpaXpp7xTxzHRB6i6qMlBzt6xt89gRku58oWauJUVvXmD7q/U
07QbRbezL4bvczKfF/aukvK7kH7g7rIxTcnAuBRNU1+nC5smzDVegPdYD+IsHwcd
Tw7okxPqESbXhxbarCYJxbrLt9dZ0t4P3G5+bdl2jBtwqnpJPDRDDIBfXrtMu31Q
BMFPqaDnuuAWv6MvQXsZCPKPDl6WJlgWP0y4XUTTdpJJWcoODkp7/4wc5EZfF/4t
RzS3kma9iDAUt7EvMuDu7L6/H7xO/C/qN6Mi657CzEjVcf4agIGgwlPySNqY0jLZ
uEvOQ0029jVYZPLxui+lFZE5UrAySSf6dkr4w5GaiAhaXhymyZarMzXdFgeuDIPI
3q5qYfk7j9YSVgowTzOEUc7vvLUbJeRgrhvicQ1wUWZ+xb0HQC70k0/74KOUXnDR
Kbook8qiwTDax4jPHwptfxfxB4VIq82YkiIVaaMDsZRjbp8cy96Izu1vnpiwXCZq
gLcyjY5oe29Pzxuoqky2qy+mdpV1CaXvP+87zeHbGFLosBXeublc616Pb9LSUgcD
FO/bb2Bt+8090iP5d5hgHARzWc2plNZDtWMWf+UgWBozgmaQlTd1oT79KOQrKMQZ
w6A54vGdiXRQysv/mrTd8DCzsIWF3evOc7Ezvydnef/iOA4Hqyf+eLMKwi+8LCv4
rNy70TG+Bs7c9VWPuNPyT4URIFDabjaLhXlK0h974UPeQAN8Faim+qlIipsK+3h6
NS00tDkt4oLW0vQpKMpQemkS75YAG6y+mZGaJfKS1JXdIZ/IZ+5ZYcCsKbSji5bK
2euzgwcHEnNiOX0XWtZ/hVUWam9IydEZlMb/lB4VMQsqYRNsV5l5plEZhRwcXcoD
IpsJMQHuXQBTJLTuLh5HMbc8wZQ7tVU+i3aDyNNm7mp3/a0Rp1MbR38e7ZspPUVw
fIju9L/E4JbIc/vJGwTGI6SWUhKZZEBWtBgKtw3UC6teGKoANDnP32STwteKqHyC
3+xjzKT4/H/JHoCKDGSorDiZtNB3OBX2i5mZ9ad5bk3KFcEir/m8SU8XetkGcNhp
S7BMlJrPAGwPLDOTkAJVxJKYnLT1Zr3psqYd7PMXRkCOXpipzjipUv8wpTGYR42c
JOe/O9OQ+ThqRzvED7Ns8ILQ4ZMkP/yyLy8sfyTjJjLLIlXyTY9scTC4IRfFOK2R
vX0v9ljE/zpsoqUULW2Za/LY0gOQtZONeVb+47wjtGdouauiKZBqjhHTpd96P/Cl
wxIOvVoexZnVvCj8ZjIMM5a+vPfFIFGBOBzVdmSRCOJTGKYBv0eUzHdp7+VW0st8
NWx74E+m2Cs6B5YII7bztI6ec3AcsV3r7WOCtKLBDixlI3/cxNYlDhoZGSwL8Xyn
xPgTy0C1Al1HVRRv7XA2pYW2J3No0muiDYdBLwJvjGQ+kyn/GLLu9d1J9xmEX6GL
ncRPcf/rrfuDEUtIB9Yu2YkBCn1BlC+t68RWBIbXX36zZhSP+5/wBLOrbr1VCWfQ
5xCDsx7lTSjZyoRCc+VWalaefVOhF6kVGGBoeCilCuxR2RZ319PsLmf2hfMXcM/i
UnYMmvxJYkvHllKqYcnLkSWITNonnqJPtMpWdJyrX6HlUVTYDyTL3duBm7c1dHBZ
xBUSX/dlZO9lhxSN8oHJTLNtu2jQTT9lQqw2o7SoqzlME6w2pJ6VJGKiOFDYJN5E
F4Y6PZ7O2pFDgAKbvU7fG5GCVl6TcI468SxxHsUqgvkcvfxFhbMf5sXkhTWcQu47
PJwV2GQFGip7kW5CSoN5Mw2R559ZNq9ZMVMbu/zPkq8n5dqYkKPMb3M7VZrh55AM
h8VrmZPwwz+/KppebeH6IjU1a6XBzZT+tiZ/YP9LHCNRY+bwWfm87b6bFt+Xnwu6
HaNd5Y8e+F/tDAsRfZUbuF1avI4kJTADqPNqRzGtIECJcaiO1NwGFzxQZhuphXQX
EmQdjXaVsd/VA4ALFNnB3vwUL6FdlxzGXhTkUaf9QZu4A8plFfu7O23p0qajZ4om
QDSRxaR13VcTqJMjH7tnrnwmbfBiCIIPrunZdO0505lWXdU/KoKbCMzH0lxgqi7V
0D37XeFPN3FWacrW7Onq5rWUn8esoNcnCC+lYaW7BhF74TpYfobFzIq9QutjlYXO
epXfjqiTkOAEC79WBDqNjfh+XSdAygVSEn7326j/cEx1NWRs4MWM8sACK0eg1Ame
h4Iurb2S9kCGFrxrOYSunCtIQE2J66W3k/EheivtMaq2wfG9IylpZjE/p8mRNv6Z
23dxtRwY3SRbPEJoA6ToKRvBnv+dUPAU1lFtvqPL2BR2xqCc29hCPkjX8+661pZX
IyrYKQsY/1rVLWIfeDpBZ/szvX207wRhlIW30byA8cr3jlbHFXfL9gxq+lTqmcV/
IRanlRtfIhSs5ls26ZbSpty3QbGaN7ibz52wo+GLgYjptYcw6udwWEJuV92djtpi
OzJgwbX+Ne572pFj0Ce/nZoVIgEJDdiTlS6jWZuFNxW5OY7pNKLBDRHrxJjKpTMS
wKFi7dEyfNM2b2us16faJDNj2v8sgpTXXVMVOo/L00zv6/JqDJP18RcrBMLvFC9n
k4S0zn9W9M7TqQszb25YiT5RLGoBo2ERwIwgxpLT9x98xvQW3qHa40Hdjc5OnjqQ
g9zpNhOChPUQ0I+mm4HNjFZzQGqChTLg5GH32r5waBuvzttbxEQbFgLoG3fpMu+g
6IoG64bpzf5LOej6cnIQripiMq5+pICEeLxvVs8u6n1lWWg6BZ5QMCLZJCsycN2K
DWg268xum/zHzSI7nlgkZIsC3S+xLd+Ce9CdjY8yJbM+2wfuM0ekcYGxD3d+4aZA
P6zmsre97ZGtCIRlsy54X8fMue8eOh53K8O9Xi5Qg6tHezGLmacIhGr4DnCV82Ny
VWDX4YzIPRK0uIjVfdhYadYxLDYo5Ieb+M4i6g3creWm3HafO40iBbGbFnSs8mgW
ukrS4nVU42cOZfudyIJgJ96juqHqlXlbGDGf4xBvxkvYd2cBpxKQBPHhRIlaVyre
IBHHM3gg9ttM6d5Y7rHdBwrId5Tfi8+FOcB4nYlEU89pHON/+f2Mihw7f3eYua+V
EiprTtiBDit12mEwFw0FUzjIuI360UbET9nCB+ZuBFnnqFHs+CaslSyCORbs6XcN
ayuWXxxnfzcCdRFi7oex+1AwZ650o8k09XBBo/IPCeYDnKo0Ivp5JxPBTOUsjHK5
64P/10gm/Cq2mQHazjAsJmSyRlYL4193uniiWfEvfi8mht2UBr24RHjLJetFaLid
cmw77WEF4iOx4sC0aXOsS73V02FWaNnj7piVWHZ7DRvA6Q30RaW8nlTt097JXuOu
8tZQ0Q71SaOW+5lEgsoBzeLywRnCGF7EYeF9nW5n2vNaPzAiOTgFXy6XMDoApxNt
llioYoJtfhoVMe+TJcAwGleJV/8APMsVfqJPdN7xikjHPoVZO0P0YbibWxULuJyY
QBlonI081322JwlCyHT+0dxDNQ5U9gsh3/FIiTiCm8UKShaCq5Sg+Nbv/PfRqYnv
bj/ywGSiDYWcgtny6BQgKdiFZks9k/QZbxzpIU9sfJhM3CIJFb4kKxVFUf8AQZp9
xhUUccSRkVOW8MmLkEd2+WB4QG4SOw+mouBvBrugVXabgeaN1Yk4ZTp6YYRPLOzO
4OLVd3CIE8rSyfxyMR4RfcFEugcT0zzgIj0dxpeShdt8ViYwcGDZwNUB0Gn00ttC
kO+0lWTReLvQSvjK7hbtk1J6TCnA/rYN8G+q9hxrDoU70f+68b50/c7lpvFM70S3
NUDBKLEn/XUiaF+ULAM70n2hHutI8Pc6lORfCWjikGgQwuWeA63Vq9jmp2xfLL40
GGRWzuGfqFrm0xrLLWii6MCUALYvUllHRgs3N78O9IgxL5HG9aREy7ZtNPcrVPID
ZAvLHj7bN29qnIyUCmm32mBgmCPjTNhypTqX1z/E8XpvwdGzA0eEAKoTOsV8afiq
BeoH/+MBlE34kDwTdiZIC52QQZ9sjLkHgRC5gyQdfeBfBPkx3V5u9HzCAp39H9WS
JAlavpz+4yjmL2oLWgVTlfCyYDVGXx95x4ajdbRsErYnbgIUi+qeZcnJRa8o9C2E
b55FdHnyPZ4KuFA2kWbNlCEmqOUfuduYFp6Im5vDDHLWDjTy/pocIPp8faFBwYpE
jRbk+XVEcTzaVf3SSoDtWtLriRmY1taXIiX5CQfulkkPKePo91uJBh0ideVi2GZb
/aLEtkND5uVNhlaKrYntLZ6xL8UiHkI4ldOvfjAMffIjlxFJSKj8JO/e1SrpqO00
my+OESlesGGFBXcoSQ3W/ahFpXAovkaLq9f2bKpnqbqIVyHI5xfyJ8B6Ru8HsFlk
O48/rvp6hCCT3xInzt0wMaSK51uq3e6RLs9Aewyf5qoAzfVa+pj6cipiwnUFQ7bp
4Jq3bgbH9247NmB8OMUQ2ia6lzOfksjhxzWMqdaz834vSZGTw6s17XBB1egdRwqr
CFgDtBDELltWfOJ+0vCj86qghb55cOhJshTJmdjrZ8qtL3FJw8Ly8ZQv5UPS1L/a
ARPBvXVXcBD9/lM5TU0jeWGSYZ8qssvboNJ6jn5PGA5lETiApX/9O1EBs0HLcZzZ
VkQfBbgxDMTjzztvEjas3HuuenPYpTXDXciaiqpUxvG+XYWtr8OTBV0TPIzT7+Dv
UIUm1Ln5FXcwJKlFUehwg5KWaGy6pz+0vX2trhwUO3BnwLIJkIaKj+fl4+B+qb0M
FOKiSDi2jOqJ5Jlcw8xWCgbdnzbnadc5h4baOuRXxoQ=
--pragma protect end_data_block
--pragma protect digest_block
wN8PwxLdNw096QmPp5iJZ33kpaA=
--pragma protect end_digest_block
--pragma protect end_protected
