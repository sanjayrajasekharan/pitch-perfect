-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
46ZpQ+KPHKAdp13Xq8Z5jjD449FfoQBW97eNRCWCu7/ZreLyGWX2HIHXz0QW9zin
oJxL2bIisx2httVEjGVMQ05OEPXspXYUSg5/ipQ+xVSxi91Ge194+tEzxOBlZ70N
zo5YCrfxOhykb6LZJpRNGfsCGwXt12rsMxYe9cTvzwq8VylK9vOg+A==
--pragma protect end_key_block
--pragma protect digest_block
DAbQeQBmTqJZ0BNfEmjevDr8mB0=
--pragma protect end_digest_block
--pragma protect data_block
huIr9uYHf4UHdjAQX65vVYrHs5Sz6os9Zb8/1obPbpi34f55DhJHm9HvTqh0GyWi
Zz02DRJSul8QHoDLpnVeM+V9jJuetAsG6EjcwEONGyZ+4dlDV9JLBH0KSNCRw9qi
RaVxECzRfMjzhira9fe196y+3v5jhKUWJS9gEXSQgHM60DrNp9ipjZrQkv6jt8To
mCmyP6mYljhrWXWLBowOfJXJ7lMJv2LfzWdJLguZVBb0k9+rFvmm2PLAy/bhIQHq
JGBm9AqtWevXpZDGfxERmEzQcWLn3FJ5MbfGpvzlmM4NMq24BFZDwiSuQOIMK+Vl
OL9P7NY7Vy5RKVc+TlZnDA0k1OPPZSDdb6+k9hIfgZVzLIvITSmH8l8E/MjifqAj
2JgYu2r+kz055m9GwUef2Khm169ThC0Elr2eClu/3feAQpP/IGcqq9JSz6Qngfw7
3QDcQODpFm26w14ECCCDN+owFTfrIh6hhDuFZ6+99X5LByNSSNdCmHNiOMtZ+I3t
2Y7yiIFCx2FdStSwtOqtujxIVRm/lGCXaArUeSQALRr5HGiNyRPPxYVrL/v5fRof
iPZQSn+SzwLr1D2keIlfe93U1bPaWhne/TFlHqr/ekWhmFOpMmksTtkMnjSsEY7o
6bVRtjZavSqKoSSnYu42YcYNcOnX3hZgdZxeewwIF2L1kwvzIOcYasqqRvAinCk9
/sMig8dU8vXd43XfCm1772tYsJ11Kw0lAWwk/JRV1cLNl8RiSYO+RRGx1A/nhwe5
mGoYNpIO1EmxonlJEUdGF1/InCwdNM6TA8Slqamn4XeJqh/XnmVUKjdhh13O7y9h
Cyk2xE0UDMe9rdHjFLvWmIMMoNCBVe001RebmNuNLOFOF+kElOaH9E8R8XDcdsMR
M0FqM5onAq3joA1J5Eo5K8PFx0aSy48htZTTfp+p3QN+Ba01RKe0dObmukwraK/O
wNbw9bqCJNXBB3nvdn0ew8rRynT5KAgmO4U2H1aoLdU/9uU54HmrqRyfvgufzZyn
3DfSuWPElsTnyDeH2usHby1WxLH5hLOlc3mPOVTBV6fLCB6DPWN/DqwqVTAgQ4Dw
gaYwciIqbc7MR0UrHMHqmDKPJZzDZ4pPSxSXvPEwb334tF79lWi6BNL5xI4sUCuh
hNF4yOYrnXhUXoMitlW+ws3Z4zAD8iEyQsia5mfCKECMDvTXuDzyDMm5Vjobpegm
vdDtTOuAt422UUYIpFSaPDIDKi8tNAyfoPMdoqFSyx/qLUqQKOTqx8CYPy7nR/5y
UpU8rn2+Dbmwo+dZ/s+FfpVsPP76ZX4Uh78HLbSCChfbGCW9E3d/LK/m1n0ldm2x
qM9BiC/3XwsnMdHK5SAwME9vDDeDVMDl+GVIv0hrsawAUL2+x6yguYfLBDHMMpWH
NrXYG6uE5DGBFGZUhkGMNhQf0UsMbKnZDiEOn1Q9cOtJNNNheFD7VC25lQlm/5s/
Bz6jcPZIwS2WEtMuPeO0nUfGfHLqVE46xTwY5T9x/XQ84JSdAu8VksSfYaxpxkdD
ofCO5zxURjmlBrTc3zp1z4a0YGBo6vHm8ZZLpyB/Gwbvm1ON7MkGi6xr1flPLIzA
fFfmoARLP06k5Upjzz29kudiqHmTVKKpbCEpx8grFgYMQJMFyMGgSZcjCdbsgInG
ZGVIN7Jd0X7JSEJzNUEcqhc131dMCXqmWRpTS7FuKN+HMPwRvM7Rp+hbsu01e3Yn
1kbQDumWW47pNgI/IT7plYVCfkkBXnOX8P0rYarKakerU92JRxuIx3JlojQ4/kiB
bO7NpQukOVjSqKTlR6LTUy2+V1AcKdgGta9Qw14UUN0BqkEOomPMxGlqNG4FcgAa
jDdx2vaeKkqZZGEf/WTbOZf8s2Va1vG49gdIHjP+/WW9SgzEDFtqXIkLlNUmEA7c
YfqPZxRkLmvQG20ZyPpuGRHh38M5wXH8MIHL1A1bBL9dDiwIxqlMcz6vZrkhRC3d
dwPg4wbi7wBWf3b0q1oEG6l9fawKAE/L8iPeRNIrOsvWd6936FBy+oRNGfNybrDT
mM+I2xuHv/DBxa5pUcS+Qfjz7/yblB9ja41S5a4sYbdm7/CT6ryIp72y137zMoOV
A271P8fGREySIxxABvOhAbrVE4q4+ysi0afho0zz98vGdj+Fx0+XSmb6UNjNfm6c
tClIrxRG42I0k635dImVxLOxiI/91I3RFykfsSrC8IX+bnXvXsLn+/VIyNOhQ40R
PTAUs2F0H9jHHmOigETSUmPEuoxY1vjgpxY7fM511vSfidZdYCraMtcRJeBXSkxi
5SwJ8YrmDGh9LXkb9cImp+Y7ra01xO+gxkN6CfWIhbVQ6c72sDrlN2CQPbwtgObC
nNwRALG79dIMZZ6TuLEA4FMchQQr7dzOmEfYXQk3YMabfL9RfV1sDqrGgmB7kOwu
fjBy9I9jTEgOKq30qpVAf/AzRvH52LO5cVs1NmM/LKJIsTNyyI1pOFhQyJVHBJTf
pyFElE7uMHlOf7yRdTXqhb9nnp1E5DaEQ94yQGrp8mpuiYivq4G/qOzHJlvjDjCg
q9+bvaaZc75IjQwDueLoafmhbxZCntD/YkHQI8RZhjoAlkRaZomK1bZG9xYBd5HX
/Q3CsTYcGGMgOt1hdRVJs+UJBwGhPJDjWTXUIRYgbSV3neOa1qLMpd52jBCyIDiY
ZncokWMV8HWJiBtao0GLDcvFzYH844W7qaQHiSw8vNsYu2IrKwsXlUlTEYhy0u2k
uk0yil5j5pLBscnH8Qmk5NT/tcS+E+lCYru+n+vWGalgAwqgktiS26vpIY8CpMeX
w8Th1f4r9nGUrBuSPY9gXHinkwu9vo5u8WSH1jP1cgF/3YI/42skPLhn2WpZvCzI
8g0+he9Mfwg4nQB5BgVOZ403U8iPTcrKrYQee7DLqME+215YeR5Y4OQHvFFsSRe6
9kKBEzj+Ks+59ZBZOtsJBUcO5SaGIsTmvdlBE/Ye3udt4iJijxY7oUjeBAlnzXBw
gbZ1KcHMVKUCzBsJY8ybyQ7/LrRnkoeP15TiwkfoEQpMEpjWYNfr8gGqppjMn+fq
UW9t10+b9FMGINfZT/EHr45iOo/4DpJ9dI2You6uHRhXL+1DDkzIEpty5hdvRUR2
wzODHSxZzfmYQsdZ83y/xKfR2V1ztH3Nm5YEjMvXjO82ESQa+2K3xhmtjUb6VpnM
79P1mkVg4WuMR5B0GjS5SloPGGH1Nymx8GKmWHuRFgb+QryKe3UioZpjVus3zy0b
bFRibVF5x8wdgUW2l7AUWXLRNxtAd73h+8401iPVQF3156jTk8Z7fdEgLvk7NUSr
rpes/Lbgx8wth2ApysOB4iUSefZycDNINJVrmhSLjFph40EXDEDGRqonXmu6VXqa
eRyTI6slbCEW1hcPT2WJLmWOkLu048xVrJ1FP9mbhewU4pzWKRs7F9qQN0bk31Z1
ojVH1WxZ75p/bRqaoUd6k+l/vd6mWqCWszdbpX+wc4yprT1OaNxrhBCv2Ayz58WG
gOf6gaqe1NdE6GT46umkwPVIWRQzYh2uV1mlxNfFVZuBLdKBFNUdnSY2pdt+lf0E
YsXpxotyMB6HVjzv2hJ02zru3rUoczKsV4tPF1WQ9E+M+IpZ6E1syHh4ublgk16d
MM0DKQOje6MC2Wpz9740EmZK28GwIyX6j6ihx39BbkIM++eJ8wJm0Kk0HPhNteGR
cPDE3j5oST+MhAfzZ7+ebLTAwZQcwmkTKdko4Bp2RYA3BQfKXoz4p8xB/gUNbrw9
zqm70tyeRreKBRu5bXKM2gR0YBsgwtTVzS80qjMWzy8NEf5CyrreRM5DMDiiq0hP
dESHGhee12HIJzD2eXTc0gFjLh2hYkuWwbWZhnb+X/smU9eXG7z61MFFWBppgo9U
gmjPn106HnslbIt8DC2YXfq17ZBiE/de54NKeF4BiSyWzEuw7+a9fnCzfjnWdMiN
Lj432VF8n8HJy1DxyXJHcNaXK/im2smh8a5Eo78Guc+mW1ferK6TsiIuXb9+I0Ja
tC6HO9pXyTabiMmvGmG79/gbBG7aHi+FhA9bMVneXUuL8iC6kgmOLBcOztKHRSly
Wr4z3KzMZsS+e598z9/J6yZlp6DHzPc6TRvvvBkU/1kTKvDjREpogG2ikF+S32rl
ZeiIZ3M5rL/EXFUknSRw+BOVTR/LqI7KfsJrvnTPvyxWjAzzYnU1rpg/bBHAR9Ql
eEeQru/Ykx4iM+nMpXIFt5Xek/Xx01n84B2ErzZTDNRmDPxhAM0GsEnYH3EodBxw
cAqQQdePu+sAZ8dWUmbETiQrWG2yCu05MqnQCrypGEwoniouBlNTfl1HOC+mUXdf
+GibhiZlMaHqR6ZOA0kYJk+eeHmsDJ6CNUkz7CUK/Frdu12AOZsO0KQcJquZKQkF
ophlFLVXm/T4u1uPdnyCFpWbAnMO4dC4q0RN6kporUhOqCo9ddXodDG4D/7kkZtJ
LXpgnT8Z1d0gDsEVWMtudXWdSV8wnQs5RH/v7I5tiF++4oCDcE0fczZVLYKkQmZ6
6DygICAEPCpavsHT/voRM1O/Z6Lya2IDK+HkGpyuIezyUyxjYutthth8l6R3SzFM
K+U8wTQKvQg1OLHd0VE3QCo6DoD+OnKPQOp5Dr35DTjFGFZ4cTreZfwvA/FNJNgc
2KA4q0bgz0YGEM46q7Ibn8CR5s6JZUYFPblrKazdFHhujL+BpjO9oYJQqOKzykLu
LnNw0x2Iq+WHPzXSRuikfuC6Tl/74Yzsa1gH+fLakfUtlO5taCMFEeyfMzoLRib9
KUGb8BrBBpCtlsPEZZVBqy5Me8Q/v9p42J/fnmd1h6dRpMuJCf+rbaqYl4BxoD7U
haYAgbAo589nhrIsecrRL8hNmitrn4c3kzk1sEnGjNT/qVc3lUOR7E7WHnUqYvY7
nFxsefbJ5nfwXViZD4E1Bf+HbpoX457yk5/vHfD8IOztl3WSkKxfG9vFTSmMWQyW
Ri5dO14JkfT2VpFPDVFKHrBcDG2y7W20ohLWpLQKGuP2HbkeyD1DBpwQf8oS/Seo
nh7SNjwg1qhKsi0sJI4TshCHTb+Xzol8mjDrgCFBVGkDVtTXdfI1D3IkDUha5KsW
iktkWkKcwUY+ZP6tEclfh7dmO0pDulWvuO9GdoA+rBobb65WywMPCPPXguPIy6KV
bT82xHkZ+O3TtDxVs5ipH0Sf5pigyzi67WGB6coESpZ4ttLabKiZORGjnbAUogfg
hc8R0Cq0ivSkZj0IFWIXnUJViz0vjjo25CFFyTZoy7vj9JXkxfrIc56yTKQ4vFeV
cWMpErJA9BnqiLkZzRSRnB4wKzf8/BnrvO8VhM77ekjoWJVHKGHUZOOf7tjqQ0od
LdzQIYqJAzbZW0oCcS8nWJPtmdnANmy/+FdJ6pKVhxFYhA5rX00AcDNROrbRMQSD
b/W9fxbZvPfxp0PJWfRClmTQSWyq879VCBHsvJm3mkVdLi4qjp0Gyb8mGWIpbwUu
LkUPNb6UPt1+gAeRWgYhwyPH1wdXAJSOa//uBApqDvMCGAQ4Fza+9OUnuZjaNOxE
9X+6NgrZuJxH1kaSZGVPVzvSCDnXSKBfGNDI9XuoS5ccUTmLf8YGC7suU91SSW+x
qmDvp93do/74jfDq0coWTpEKpjC4b1NCDmfEKL+FFnYeRjELi96Z6Whkt9ExMCA+
0fgwrQC+fCcjq4j5l9rYmkhzazUTNzsz5JGnT4EbF8FMaVEnWJBf4/jYKfk7r8Vi
4vOCaG3N+rrkGJ9ejN9N5r8XBMG12gjBHb5pumVNpKzOadceshn4Et1jpJvSt4n1
iOGfDKK7/nywQGkfJ4JVOebb/wCv7qY5EaKyz06VX4buxPGVheebYM0jmjZwl9md
r5oQI1Ag9M6gXPNx823VdNtKBk/tzvgBcgFfl7dgQevNDr3+lGxe8wdk4qqUUTCx
hq7pYtRRrHTGz3A157ZuEss1PxbHyXaPI6pdO1MQ+tkuPZ6sOb4kjV6nSpriVnO1
hjFV+vkQiKUnQiBo+VzuyNw9bEL337ylXFHOPwwSUHOjSv3aXJwC2qZUVqzKX/Bf
o1iHGLVXGw0+QM3S0yfYp+Q3ClhEigbYXePO/CXTFwtoeVpuJBnTpUOwXAyddcK/
X0BVbkNEpMSaTTJd7m+rwY/geyF4X/GSY4UsC21xf2bwL/viKKKiLpgGZJMg+yq3
82QnSDCeTkhOYWNJXaH4mXW6cgEcfmffa+ej0muaKBsUboIsYS2GaGC/61AojG+w
XUE3KPB7AIJJTeTmAqWrSCV2RL2hi3J++bbAY3M1gjiZDuHcq5Q+TIWdQFtIFaE+
7SdZdDYMsdupZ1jKuw5HATHIx/s4p4COLQnuk9kVM14StXQ7YMdxY63kffjs44Jc
Ds3QxobSsUTWmWTAHfktLkKX8pwepLx7qDEHmiaXSMMWP3Un2wip7YOYwaCgdx8k
tahoeDFKE72cKh4O5NJglqoJL/zGkW/W9YUYccqSsUirk3nf0wr1lr32IcyfdB4z
kKKZSCD9SdVfM2g5VJSALgni9YarlkBtjJA2Ny4LFh0IjoGG8eTPVHSCjm5FwhWM
xcj1E0z7Tcm9GwfI3wP3devRBFsuoGC0g4Is3LNKHKHEqvSTvF0QdOjJGqhvoCxo
db6JeG7HmdtjnsIAnRLwkNaF2bvXT3J+gN2HhmtTBnghVxCOwE76Uy/7zu55vawb
ij1n1u/qehIGh3GPZr3sm6xNK5raUMSBk95D9KFF/1uZXEgZ+sPOscdLrD6TiF5Q
17UGM2J/15gGCRDl6D3+VMih2Y6NiN8J4p7zvaNuE3Jm9as1g3lTYkHKNDVqy2TK
CDjAIGfwV3lT/1xdqru4Ja8wS+jdO+r1O7ITKSGCh/y4unupCN8GN9sKGBNTvH1Y
dYVXQ9q+a6ETyHRPLBAr/mg5f4wXOHvuUXPtqlySTkPhVAs0YxPNb3R1yzQbmgjz
wENuxbCVDlsC/Efzl4rHDK0ovBTYGJSDdiCH5w3kOHgYhmG5dAhVXxD14WxDcvhz
GUSLHVO9UNsORPRlRrz1tkXk2T92htmZKjegUXaPY/xE5Bpe+6CLk5vdQ/D2PDCa
l4Ck6tK6wT5UjJoWomHIwb8vco3QvguzZ54OaG3n5779lW8+0k/Sbd5AvlfOgiVe
Vi+zxSQFiYe/dimvDrJVLtaMynBvwqeM/TOT39a7iew6j1m9Ob8YXFpqdAJGvkiX
dTs3U6rN4oo0tXjj1TOThQZvE5ZUTYKPn6evhIZrp4DvREo63CEjweZS3zlG7cNH
HfipuDD5Va2k6kICSuRxWNZYjOd0rUjaHjRv3vfU837GmfOEn+ytjmvMW3ITTw70
e4PTD7+EQOUxi/rrnIM5aPGQz0NmRyeSY+yaSq5O9akrqve0GIbK48ZCeFKYSdrQ
17Q5APudffNY+vIgHkDoQLHMPrEBwbHfErmqZmqL48dRJXpOCW30feYq3/SSAFVO
5g4R+AM0HtLy8n61iVD33Q+BcYW4wNyURd4sLm0Ysilvfvr00Y2hAfcMWIqAwJsI
rMCeIM++PVlOX14Ikgy6xodY/UiVa97J774DdOZKL19HJqnIogDSdm8Z5WJQTApN
CuYCqQHwrHOtmhJo/ObK2M+4//0Ys4yhLk1cNkvCJwyAmEARA9A47UIktREO55LY
dqZLj805xVxez68azJfbPkKF4euxtFXSTS51+lKq+4ccNWnhNC4Wzt1wgtco8se5

--pragma protect end_data_block
--pragma protect digest_block
InGQZh5JjmCUIZ7jSa1C2zZH0kE=
--pragma protect end_digest_block
--pragma protect end_protected
