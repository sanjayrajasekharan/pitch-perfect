-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
j4AxCIu/LlA/38CuYaQRcqfR7pYCBhp8Yk9d2vr5iuSX3REp5tsNcWpZ+FB+13sW
pTBcw9uXjfL7+zk/9HOaHjJHDbU6hVRgyUhU/xu57vYDmSH+1NOw0chACKJyc29Q
ssqdHnhaPEgylUGEko8dH73iFjg4F41xkdkhpZEWz30=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24684)

`protect DATA_BLOCK
ABL6ah8yUsFf4Z7KoxML05LQL8z2M0skFvkK5ojNLiTzu/xHVQX2R4/jrAyNzHFr
qmCleifmhPeEPzg81XPi7LCgzVRYRs5F1CDB/SFsKsEsc96/IZKZJ6Mcp/akQxPB
y7LgT1d0uRU3PaExqHQE963F9RU3kSOKO6J/zUR1DrbtG0e8QU045lwtj4+hGXLL
5g34+pnXxwv3W2grB6OTgbo2qtJWOKXlm76ZtxU2cNjeG55xtEFWNiAX/K9MxPr7
0ct0ydwgRaubWq/g838CPBVQHAoBdGlbfNnejc9x+uF2myXhrs2YdrG/7J0R4L2x
HSypwOm5p1ZpAFU93oFJIy2+b2b4dxsGFDBx7fk2wv6QzQaKuB9AVkc7trlh5ENW
mBX1keQXHbfaT2sfBD2OR0VYr9NYvSV3gpLbId2CjrOITkQD2Be29Vix7PiE+DkP
XVFwRhEvds7QpPD36OOIauuZFk0p8Rjv4f91XKYItAfuquvq9vbGoiWtrHTkqoSj
dwwpsA77RnUSCcHAoQt7zK2qeTzy+BifatPW+JoLFM+Tc6KRnVve6J7Eqnh9gLSP
ZCZwQv9a1QDhEYO4y7VNoyz5jEn3++GTu6yhtks1T3pseBpQyOZTZzNQpZjjprpX
CakPDXaaVv3A8A/8ByQbwo1uXCp/nri17EAzlC4LCcWlrJ7JqWHrNjoeb5br6gez
NgzeAIbsF3WMzjAPpY/J3d0U1bMdad5tqInA2vZyQNXpimeTnQ3w1SVlkU33Yw7a
vQoZYUBVUSKDgzLzj642hl3pHVlqGUfc6vVQa8HwiLQw5K61AeuJCuosTR0z49q4
ojGFCLz8V+RaCZknYWRfaEWkSZZ2d3BURBhm+khRB+LntdCiVnqt3jN06SGZZ/Em
YPJdT9Pdv638uCBJ/TbIqsyoszTPC9G/A2Yih9aRouCIBqYUKrG0xw4m7WK8v/HX
rn1ri4uGyciDKAK4943aIHFn5RLULYdZQPAqGDeDD5fgjPAElspAdfsmHfoRkVxm
I40eePJ3s0u8wA9OzrnaX9aLFS81mrVqXbrH9lkmOoB3Edv5JbPNpCPK/UcD4IdR
f7EiPEA458Py9WiincSMhW6vH8upGlH9Xinn9d4b+SiS0eK96KXxJibPRhY0x+lD
PtwxhkNPoT3cScSl9zEAyNhw2qXMrEKNvJ3xnOJarCdQ3txXS5teFeghIKsVdVBb
h16gVlq9AYj9bPYlZuewE2gIdFEKjqEoYDc7mJu1OVA/yqunVcvvbJrYuK3GBtmv
L8GqzJa6vEttgSACWxKMEHlAed0YY1XuplPsoVIbukxb9OMx2E39TQSmGLJh8+rX
c0fiEUCHCOyAgOpQVNs3mM5FdsmGxfK4QS6ctHSNQuzAGZ684s/9NP2rDMEvVrh8
0Q1kRACRUq4pmczND5jVqreFaoD0xSzwjAL/2TqMegDGzC0vBnzkqUFgPnOKyhlY
hQwwG3XWr9NKPbqFdxzstTnv9AdEuva9Sb+Xa9J1tyq35Jgmx/EYn3Cl4cIeteJc
tX7EVoK3gMPEpbTnxJtAGDcfMtEQ0ngHXNDasQ0alIshUbK7lavaiEwc+5c2K0Ay
evrIuxWKAMJo+3H+ZWlQr6QS01KaEG7Ex42JBLfdvsRjlwhjll42Oes+T3OHG/+7
g/5MzCCsDyrqQQgVlkHOE9bdQniqYPA7Zf3UJ/afF7hLPtJqEoDUKGawKFp/piWS
2/4Oj+F18toE059FBSYAaMqG0v7CIac57l+f/pb+312Be6+bI01/7+q8/DNeH5ku
ZDfjBS5omBZ+/eqIO0u5mAb2LSaPRIuvm4n0RyXAdLJYRuSNvAC30/Y/Eoqc/iPk
tYAdslCna8kctKi16gs6YL1ALCzwuOwN7MGtPc/K7e9460meJGkws/M0wqxWfMf+
IIYQPE246Is20qjLUKrL1Eg1T64d/J/CcIIcowxLV9dsBQ3kmaCqfTsW1VwShPoB
3kCpANiQBzmh5eb6rGOvlqKlEs/62Jpe/6eaVBAhGAuoV8/zmtHrcGfvZVKFm5Jw
EKO3IbjfNi+BmrFzqG1F4OrlxTlLNeaWjc73JMtI/6oQfJXZYlr5GtXisk8olihI
vDNKDtm7qObQF1w/1x8XdFGA5S1VIOurI2BLtCgKHwG2hE/wmLDMDjD4aRWf2REu
jZ2CcN303wdgRcOmMnQM9ev3nGOjKvyMuN8y2NbxtFr4Dactg3m6JHU2ujlEZvi+
qpIDL5h81mzPentUewn/2tb1El2nwcltr7ZPwikYrPWsUh/Td+8N4NPLZKpITVNn
v6jnoxiMEHYf7kBvWyufN2l5CSfSIekHAOZ5rdcxlV2cVb4urtvgp58EICWIY4aR
6vkWt9E0/bcuqE/9Av/v6Vb51J8KlYzH2CaIpK5FnHdHnUdkuwOlGalzb1sIHv5R
WG2F4LqckWA6VlqWhSabFcTEsPWeYwY8N9BrYn+VPjNgdntJSBq3+aqkNVSYb4JL
FXYQbeDvgoQR0h7vt+YnYF3gJCl4Iz7fbjI3nOejr+l17al9fQNSJYgRA/shhB4w
Auus8uVWdc1EYQdORlIRnKhQtqtE4oDlsUGS5JieoZcfd85/QeJpojpt+niA+CHJ
gRkoK1bFx/Ikn5zVp0qmg+KH3Qssl9DoEofeM7svfg8ZQ77HXAFzelZlbM3Rk6Tn
srBT3ywqGDkpJQUrLbryz/yhG7B2ocMXtgX+9C+2kQ7GOm38k526NGifqUShrFn+
5FhMqxsbuFO6S1XG7nui/lJJLjwY/1DTkIFg7NJDne5+EElg3WVHoWaWVO6/o60u
XgJkrHItZ9vKQHeCYBVrT4mH4ujvUQ7IGg4lvCvGy0ieKIwxGyEfbRnjPFVo5FlO
FdHAM2OzTFGuO3jGVXYUGDmyNwJgNXasKZb/n7+K/gKbAdzmHz3/8+K6bPC9NPk7
tBDDNnhBa+6MefMsLxPyMDXWdYRXDNR87O1pH1h8gZlYiqKsjffInpva9g4KICvH
zHlAb/pFb39ay+tmLRboCv0scepTIeejJ5hku+ku3q3f4zbZzvIkTYbnlsG6+SdS
iAt8dMg21be1AfC6T1oYCjTHzCr6HqEVLcsIpSYv0KVeG4LqqjEhcvlmA75cTsuo
Tj2/RJ270VdYWqQPJIWMDIrrJ/dD7MVs5lgu2NhtiD9oDiwu8dr9SKWBJWMpFI9B
vKTKCmBH18FEjvP7KnI1NtK48wCkxxYKEnMMhzYlUHkhQ7/mFHnNELzMX1KBSXkz
patOp2TDtMJjBkmnKjw8HM0NF3NpH/S2QF1EyhbbVjjM/ndw1mSrSoc8TRYxs/tU
V3W2t5SH+oKR7qwnG93YK1czykhQ2zNw8FGxCnYnQYTGGGO4wH5oAxBzVwS+ZBFA
iqLvaprwOW15/QoRPNxzDC+ocV9lMyJdMuKxborMeen9DhTjP66skcnA2KYSmA0/
xLttOQZGxlAzwRzRg/3rz5R0YDq9mF0OuuNG7tW9PvidF5bHj8TPG7dcVgw3drmK
lnxU1KhIMU1c5WR2jzYltr8+DBiuUrKlWT6i3kubGySm4pQxS3rUCaQfChuV9KZM
t9R2eSZGjOYeJ1rFg85FEWtQGaIq+A1wt4HqQKWb7A7bWznZ697OXFqCtPasGiYG
CWuqlT3qcDiBvwNsDcr2r9QhyJRpjOZcL+CR2R0aY/n1N9mYtYBTibxEUCjm1KJ7
Mx4GiUuBVXh1o9GkITzqhV1VVWACj5rTvhZIeV8qLgoX/V8X1FAKg61Isu1NXskM
T2/afRKAHHKWcVGg9g1rCUiiORsEpRob5cOxlRT/rub/KOzc9ZXBDvh9Gk5PrMh1
IGJOr3qky8B0wUnpHFp3cZ9pDlj0kaYR6HlSs/tpavfXzHzEUPJhaVpi2Veltm48
jrZfFmDLUGIyZfsREnYpL/hm9CuUPJBx+pfJSCAu0pMV5v2ZMtI2vA0ft6ZT0hto
RNx8wr6Y1xpff39krKLsMtViCqV0YppPuNNUUK58nyqBHKkFjDf8txGKgMvNAJ7b
VCcxbp8eDYDtQheeNsM6OzWgwSlU5X3m1Hb0Hk9zQX6RcIP3cOScnk28+NA+E2rR
V/uP4EafTHjjvLIOMRxKtA815A1akIo2e+KON0oCLxKBFj83RNUj2i0VdFcg5yGw
4F5FrSms0+piW2ciL9lUHqKmLCx6/E9r3hQfdj9QcMTwJQdPn3k9MouHWGHeq3Nu
jZnMfY7f6Ppzqh6KkuedGRmpOZ+fyvbzDtnadiQuIDUPkl0ZwtFuIxiBL3M1EjeV
WJ/XYmOKEX7tULZkL2sJLVuc/bQJQr8N90pr98VFi5Rcp58brjAyViCEVrfwiU/Z
Esoc9chscNW3R+sQLccJ60jrFrdu3gBRbZZRNm1U3huE2ZYNkM3t/gzb147TDqjF
nKHf35jA0idTklWeR3PC1GiiCpNtB6nTfsXhOjmYBv0Oi8DGI/9nwoDaatRaQ05Q
FxLNzm/fzUdLkxnjPiS2W65R2oaWbTzvTQeYq8voAbLvCN7Fnt/zK2edRYyPeb8n
u3V2lUMuCDVmA8ZhgJRcwbj4KzJjY9QoXMcanh9NPEYKdatDlm1PD7D6HVcIYlrI
tobu31XSBkXJRsYqhpCon3qGG9+oEc0qnKhm7bhA1aG9S+CCfIqsR5SzSNclCZWZ
kOG3GNbD56EPxtsxOtb0ScedtH+7YBnnsLaOoj2H7VxlIxwTLHYPhXIqhj4VLnxr
GXpU9lk2wLbEjF2oxZpL6o54c+OZNVehl77s0QF0w6oozVFEkxbH97rhOZ/ZcVzq
YYB5E0Gz1TIBnPDE25Yv7ouDfpqrMRT8lwewvLs157Wv9WLfiYSJuw2zD3GnhtGh
XlJxx/xY4SqFGVM4sW05NMIipRKvWaYRjApblb53F2aIdmsyPmuJR/uX7euo7v+9
9d8ttqb0IawUA7i8d3zz22xMQhr/iJ54SMNx7G38lYBhZA926zFxAAwA4LRZKA7y
FjeMDJUxBowbu1k4dO32ZR5Y1X9n8nBqOvNTJqcuDufXE5LjsrnuVTpVfDti/5Gp
6zOctuvemOSMRRDNZcFrKRww6c1alQPtIyC4jqBnq6Ii/cKQRDvK/cW6a3nSI1HQ
uwlRufQpkC0n9eTltfAsv4IN+SXFl6G0rcHHvvFyxxzMR+JmU2Q2tuHMWDNHqPfT
Emkx+docmJ5Ui4J0QAAD1/CgEFr3H3PXbf92nHjY+Vvfy/2vsc8A/JGKSko8pslP
NvfqJEZIvVjyEOKu1cgeipYeQcPjrHiu+Yeb6UK0GeHjk3v+tNQE1y/CbaWG/FBB
yhYsTvoKWKbisvoprkg6loeSeOTN/L10wGr4/zZhpsWW63F9ibdTKSX8iqqEn9ck
l9FbD1qgEKMWM2KkVS8E3FWhoKecWyRet9nT0/zEq2GQAUpyMOTP9RJJro5POB00
LotwY+MhFh5SdYQoqOpv55ERTS32DzC9IE/7m75OaLpaS0TIVXv92OMJxqjblJj6
QNaLq/+bil0SsATTd+22CRHEdKT2lhjuVOJAqGa/41451+QSvsYKaebkQ1CoZHzN
dK2st//WM4t/GqLlHPjW2w/cSL41k38zgkk++/RxWekR4RiPuoF1kmUOyQv83R+G
K7QgZsZK4Ksvyu3c69WB0YC0+V1sLmAatAYccYGPNAjn6wEU989JbAPfRJGhKcio
IFnA1lBUaUb8yWRPpGeeQ1hU7BuG8pVPtezGEkdb5bf257ysCnxISJ4adZWDRZke
dm6ukuqlyilb2IBMMHzgsZ4FBuMJMi3H56S+PKKoFKhKcvH9CwZoa62ZkkOAclsb
INUgyA57Xt2Pt8lc395yU0fnstNUEe0OIBTB2rUwWHuicSFGbhs1ZYTpev1PbNlA
tuL1C5d7x6X7qkKuG5Zh0q4egaG99nw7VaHDAQMxno1ueL+8p5YLgj5W54v1Gju4
GZvhM5/1w4x6R9zNIc4YobMbuGCB9vFhLcob2P2O6H9MYzw6Hgsy0uKYUK6c4aQt
BGXwFO558RStjGFu9Jz9OFvH8Q5a5rWM7GUsvj6stviXmmtrrR+KfWd4QqkJ952V
MMOw4LTLXduQMk7kGzld8lsqcz5gtSJfdIRmQ0mEyb5Y/ovyELxZul7eUTFCftz3
IMuRBtfbjzhn9lFzDoz6Cm7POT7ER7R+zdgVMc6eHdaR6VNjnmzXSyXhV+GU8grj
mJ8PlrDbgT1Vhwn+9cxYp8EHLI8C/NR1blQQkJ1v12hYZX6zvBuSXnznr74eZqPQ
1ZCusptZ1LvmqmFVS5SqHRjC+lgV5/ejorAA20877T8gql8V4oDGHNdX/snoDMVU
W/BeAddUQXak6jbRg16oofICPBVN+qj5b3LJPlPQdBNHk1iw6nEcKLEBI1FbWbrj
2RpdwqgjQ7wD4C+HgybN79WDIZRapgx865S6j4hp/Udi5MmAcDz52/76C5rQBrS8
fzaStkqjH7Q5NlV1Ls76v2YejKtw7oVTA0J7sjkaCjERwbiDM/cGsZJreo+fOaz/
dDMmEaW9Akbl3dC/J0izN1qwJUy+UAvH3WMDW+zcJRYWOL2Y5/Z96eAXeZUbsSh5
mi8xKM63rEoygJDczh17khshsVHhrm6YxQbS7jzcul27eyxf1IBqhnuDvXSOxLj2
Yz9/jmUZwtiyRoeg5ABho9YwcE0ayicCZhN8QANAm1vGTv1LOa1KXJPcnZKKF7FM
Zegsdb0Og7Kj34epFZ6z9slcjIAwPkTMVl4UNOdXi2D7VM235VhdUDST+Hq/hwet
xmD6h+JDVElw1pKY0WZc+AlgYgjjsZEfNjRgM9EW7AUkukN6PS8ZpFjBS/dPvm4F
wBEsiFLUXFSLrMk8ftbiLCUZ1T2+oyIIMAxQsT1Kac7UI0DFIzbcCDyMDCt/WmyO
cUAqurysXYx72tX3hT5My26CD0sdfn5M/nYunanuGZkRB+8cZb2Cyt+tS62l4PaA
5ys9GrxqSPS0Pe7W5aDQ4KbmaT8aOM36wotxR7pu0+OR+BFanYTI+9neAn9ddVHt
GRfJB32P7lYdmftRI+qVSeGtUw5Qn1jb/TP8nVpwHOF/pemaTCMRi5DL0nMIZR0k
Y13pOrz30J3voCUf3YSHZBGK2OvJVOmDzxf/yzJyQ15wkXjj03pTuj23saK7Xfpf
eABB1iG+foXo71Uw7zl1ur3c7PBnCk7lwdDwGJQbb1YkJ+l8gqP7Le4Tcpjfejgr
mCo2AdqHDmBwJegQg1IrlZaz32rVhc/zLwW3repjSonxiJ1nB0EZiJ4B72NRJ8gi
2YhxpqClXcBuqJiFLiTy+qtgBjuDYctPiH1fToqSM6dOmm7bNqkiNlPZ2EYjOe0r
e3ZFOo14bfYkXWqIr7AjCSPf2wrM1vbfSMTPsuagFcQEjnmXr6VDU4qpbLgAPkRl
e+wPDciBiu3Ck30PBCiGw3TVxbcCqMvAj9kohxY/QsQaUvhZEes6wXpSqgHmJqCB
tJrsbEv9pWM80kMRY+e9r8sK3i6Se1NmPcI+eE+1UxbfCyi/za7szSbmZtPf79S0
PgQECJDmcK0cLBMjGKNTrffbdaSwmNAFwsKno+d0VBsqnjI27qEMHj9ykLvDoblt
TiP6Dg7y5tbixwwdEIAXxJMTAJQopXJ+Q2DytTFKJ1hiRND80K3/S13/DCxoGDMx
IwX8YWb0Laq8KCc1QYXEGLSdyJjklvi8+frolrvJ4zNRwlUWgmfD4ibpEpxjRXoP
htJFUOuKuf/5E6vJclFspCwqC5litxQmPckCELVPioNUqPAma38Fv1NIWorV6UJq
Gc/va9y6YBKOOcz0NrEcIHmIjyRx6N/bQlFAaYYsx/YmZ9Qq7lmtRmP+7JwS2bJa
VUVHRhOumsmFSir/gTiOox9uExtw9yYfqJC7wWiHUtWSRU8W84pubDKNeYC0m/ba
SO0jS7HAl8Sq1upCT6mpPQvy4qf3yJ99Q2uyXaqwbx5eurNO5vEWa4cW9HMt9hrw
lxuqqOqJuAFCVe2GNkC+PsbJGj8iTFz6g4tg7OlUXpeyaieJ1UVig2/Qo84Viq2I
tMjtkivX4JjaN/fT1MaSMukmGAdeobFSPQ5lrdL7zD1I+fIEfvMZsL1ErnQ4Y/aU
jWui/n5ooVUxgdXDNCd8sDZmQLef2qo7O+caxbxFCSoUkz+goWtAkHspZ4eNHXXA
HRuNrAL8YAzuzxdkeVxI5RDZPPi/G8IXcksNv9gvntGaOfc+5e7R1+qrHjPmryTD
W+vZw2k1SoJUNBeR6N17czKNrr+XWN5aCj04oX/JdnTwvIKyGMh5MFVeNfWm6Oh+
88YeO1Qyi3sjq323xIHcwYX+XGuNpeUR+YFKaKD0VU19corWe3By853458t+IdH/
HFZN0+B5q3S5eT2hQqHYlNwWJ6c0pLa3x6pFsNzd162GBLidfKB7PU0ptE04oq22
FAQ9gPLENht7vmmFPrdEDP5DlDWebrXbO9EG3oelY03aJPy61CyO0s2LGCAuAQ8j
w+LaoUxMnxjc85goCQUihJVKFRDWaSwppDfKKGBQmrmystXjtXR5TA7w6dPJJqDH
Hbp1NIF3CoysC2g56Qlzg+afI0LGPk5rwrYKVwsvX0JJY0Jr4Ej7sIVqG/qssFI5
/jVx5CHs7Dq9nECQFVMYaEweH1k3gILbDrPq8ivVp3hK7u4r+25MdJiH+buD0oKJ
zBCQ0ydgFavZnhimLfagzbYL8LMqiJNKjSPRjCjxeYIfMLWXbzaDdA8Xwc4X9yF1
CO1LVcqiP5N/dvcQa5h7zJE23pRZnqoOoy7EdmazFfh+nJujPV/BKfr+7Ts+LX4A
VzRhUUYEFD7p+0BwDeITj9+p/cKKSLhEF8nlK7Xl1CwSdta/sLnhBx7NRGgFfIL8
33Z+pgRFZIjYafgnDHTlo75qw8bWZqhdzF6a3sZOsHnhJBzeoY+/y40J4tG4UDa9
osvpXLMOcSYcCUix0bAjTm/TuPCuMy2/IKZVX543nkQtF3GvrNENhuAOX2zE7TIX
idIjURxvPkawBt3KReIQjTOaf1PIxtf8EKTM5qxbqfKoLq2BqilrQblEF3QSAunp
hxVXtKVI1Cljd0yxcSFLWXBAVMG/K7OSp5IQ57dN/kPCMnlFx9qY/edfxqEXXhYT
8w/D1eKffzldvxUX2+dr3zsx08qSdKHxJ6ra828K95lyR2Rz0fSy6Gti2+XQJvS8
m/tOdYOHi44AG1XbC+GjRR83+4xyY7ua857xdCj8dMLmqrjs+yFud+Z+iSUldJ1H
W7RGK4xqid0DldM2sOaiGTWA4WjlB/hVSQ52DF54yYe+L0DJjufAym4yvhcYVDdy
8cdTvJc/GDy5MpT2egdtQItU1DWwIO57URD9lBOjp0ZzgX+VhtTXs3x+cXSpSSNS
1lyyUwTl0NR5xbgSS5qp5BdAyhojQxiP4K82jRiMnFQRe7Rqh8TXLSL5L/c/SQEC
PmLFNxp354fQ6dDuAcCWpG+Uksu+0JWZDEbOeFU2p5tEQ33P5RJ119iHaBbgtPHM
7RSkP45IHYDwf6wnAbdgnsj07f8VEusY3ZC4usdlFkiW6kX+HtZ/eGIBp66qMRXo
Tz1ETaO6YpLiYpKcNtuFuRaa4TmXbnJEEGZfX4ZsqVgfCWXLzOYblkwveMGU0mdh
Xl+euuoHCmxuTupYGzOjm77pzVi3pM4c+kxlkN80/U8/YqDAybtJzV7G63MIx8hh
y4KBMhOFHu0OWztDQt0zsD0d1+RjIWQsv2ng/0G3qQpaocFSXDrSHV0Jal2gBM2k
a7hqjKSeo1DMJV++5HTdb24zK9jwRyYjQLtWccnMjaacXCFG0KVrH/q03Zm1D6fn
WRT7txlBsKrkqhuP9Fvn5hm1pcDgSaodLkMRpHkUVZhhGTMR+PY+eQEA0SAdLN6a
jpHP5pkN2YzyvmAw2XAz6UJ7SBRzT5hwzoFbnfr9ZLfoFirs+ay73dfzm85I8Oz/
y7QADIaZw9LuFiLT7H8FoHTkCGsiCQlyb8TK2beGeuEOkr0G65JCEL1wIWQ8I9Mu
1mKH5WmpbI0y7L7ezDNY8AmFGuDUoUbaQkztk+oe2vwYMxlQLLE+Z+4guq01X51o
4Zo2UtwHN1sEPk5TYBg5+iHxf16vvn5438xo4qEWL6ECSoS9Fw4MsJpM4tSivZhd
C2rmU21kxgNnHWYap/5OfeDM0XvgurlFVBp89Ace4+2JVqJ8qxztIf+h2a9HKDgV
WQhW81uo8hh5R7nGbyEmYk8eF9+P7HZEYIh967OFFGBDQrJCDm8Qd1o+4X044mar
n0sVfeXPz5g0WUyniChHU6198hBsMqLvKOq79Q0lHqX7B0wmxd85S2ip06no6ITL
mnZMFCwT51CfUlcwDUVCuuNI1ZT/m+Gkn24JWuZ/PbsZlKXeFhIrpf+eUeCf/5Rq
QyrJlPcV3UnAMon3+Iqy664ShEYfnWVTSbaXEn63+hfNxRJG0watLleOP0AjhPJY
4MCY7VUXq4y8HcjXJlmBENf538bLxbKRFIeIdm7IwiHqpkNGGh+DRqEomLxqi2Hj
KmIcZVnSM0us46oZ3+HkRTlAJpTxSdSc02OIkZkOdeZX0r/WyKfNCs5BTg3JN27K
IxLIS09bfbDl760SNAt9kLpGPvd2k80E25lhRBA/iSzqUVNgrhfy+qSS8IOd1SYL
pDKikl0zjoFFD2AB6kEV0GCfaUI/SbOrXz//LkXxpTwuw7WEDpxYu/ST36PtAP4Q
xGmrzFPskw6IthUhMftd8i9dQGWdNQkQr+NwuepFIGDrgM3H/d1AJo1a5fOHoCWn
wE6I3SoB7498cNQuR6VDTy6ogNZHBfXgTv6DqLt6N2msonOSRmWT8zoqU3doXVjR
yca93Y1sD+q1U/7n9e9DNDvXf8KjUkxlykJ58MHL2cRFGoQ7gbE2Uror+09XpMye
Q4Kd7DMfNf16t47ou7F5P5MYFrFKHjKooAcRR/aDofF6F25OeIQnUD/CPicwXThU
3N/0L2MtigEkzFyYe/EPNjXV3xn1bvyKmqyQkIRD21MsH8IC5M8YUB52CgPJnQ6m
TT/mnlTdNltPdw3q7srJqyQDFQmVIESSlw6AUd2MoQFSwJffMic7nQlxNK7E85Ux
F5nN36EksYV+j/XphNBfibXBdgvof4yPF5iJVvFrh1EWlNTCiqaZHwfM8hL/rMgY
ZKeBX8tCSPZ6YNXWOfyUYRt1F8gqAaHThR+J4cBj0JmYRBe6BS0fg5iZuW/1fvm+
7Zj7tGqIuV0tJRpHvCvTJCVERWZR0tFrIHd42UN2b1ppo4QqEXL7vrA6JUgOoG01
0g6wRKRBNpak2jYybgKMXnksbj24TiTyCHPaAoHnpCUp88Daiozz9+z5U2D5p025
hJ10CeU9xQtPUn2UgOIFr45qzfx6+PoOgbfBQwUNwFSttYw3klVuV0+hEFRJuWGh
gGhCblOn2GDgf8X6LTn63sFIv4sV7O/4tYpn+w8JvQT0jjuGjtXgI+Eo7BPBLKQh
a0wsCVuulUY68CZlq+9iRoXBaAlOmF4nteyZUgEiwOmfC3w/SMHMVe5UgNVr1vP2
+ifmmt2TMEA69scAGtFMgUkE8g4JYsw+X3HZsPKo4gkT7Nwt6TzxrpmhV/CSVlyK
M1rrhlNffQIHWIKVPBBLAhQZOJP6V/J6qg23Uh/COtEEOCPzK8NU2gcjkwJzyHN1
MgL6ersDTJ2Lz4E7VqI+TICWJRg8CdqofUnVdKu0L3OKkONgL+hZNsBx9nc03/tX
8tMFCMXthpq+OYY01l1x7x9yEtGQFE1BHWeM31HdrlEEkbOoJMNg/GW7Nc/SFpjd
pWXCPCudJns4RiU8r1/T6HmmPq2HOJVPDWAjPjHS8GtqQ4nLFGFh+Q9t5okyBr6a
Inisrdc8mYFZxaP3Z9Xhvd2jeGG0yOjhKmxMBnJhdTP81Vbj7EsRaXSD+PYZ4cCj
X8fyY2KDfybikiIccTitw824AnuvWXtoDXTkjv84h7ewhB1APXafJp2swogHmrQ6
f354w3p2LgItzwryA4xsiSR868KKaOG+cmTacc9D5hr919es4Vhc6SnK1rX1AHXg
a7c8oWPfomMAAmnTvTf5xvSYB0l6GaervBTlq1sTkvcSUd+nM8COEBXwIeuQK5eb
sOn0oSexm8nhKMg7/dm6Z2PsjAOpuifOJRmB7YODtVRDy2bP7LLKMCa5xPgZlLIo
WAe/HoAlJVxDKPI3HjcFCaRjLYtpm1v2h14nFCul5sXtUzxfR44vKgiiIWVClpri
t8Gq2HXtAbWDt7ytvoivSLDCecj4yXPKf+IqjcOsSFXdskCNRkz5XT9uJm65qNiL
xkXmEJMIl9e+dmmgYG0+0r6MnZTswsZA96be7IFH20Isifx8DGqLbsYYOH6X4uGa
NLGT2f7XGJWcU/KwU60AFHgW1H98YznsUMUYZOemcnUsyJos+WjQ7y4UFtJktLP/
P4yR3xz9wCL30N5J/l2ZWp3h/PJdEEZIb+B3/DQeJ1dlnerzxzBSnaqu7OrB+iHn
qsWzFNri0I3RjkNY4FjdqvBr2qlsRHOSYQk10LIbzkj/PPX66hOEkv4wuAJpRlmO
IMHfTGG4Zf8dpF9lypte9SkA0CLMHjSVBSOtvjAZsXIKVDQF3QfjCpgCqIQVgVFL
nb6v3rVoRU9CkxVDnVmXRp0cEYm0JVrmNOnmeW3CcOp8wJ/k2l/3FeyW1WMFKbwJ
ofOOhuC0k6BKaWVrQMMTSg/rlwI+ShSmVYHXxdtZxW3PdIEtw8BAltOgcqAep2t+
MtFx0n7gwmYl9kXkbK7hcXPbsP74HWnoNRpx8hGnInRNqkGb83W4kuwg3RZG+VeJ
HuaMB7A52E0shIMgwUcg6s5uCMUcvSIleQnbhzIsBfxA/9TWOabKQReQROtEdWPh
6tQajFkzEN1BE3+mfnW7DoN/4NbNZldlYX01IV6XA4bxV74RdmW3cXHV1u3OT8pw
7KFZ3chJ9FtV3hnLLIueQa1ddZXicXyA2dGHxCB5QMAFyt+PYHI0zCX+J+p3zdsK
Kslcypz0LBTe5QeGhjVPRSxRhyzFJJSF8VXQ6B8hnOEXHVIdVyVeSv8yK5On49Px
7kOWAFVUMmlxTenyUV2f5yGSP6ExgsKqjfZVgzDAX1HMu6HV+0ciB7S/j3fnKsqz
6v1oN8oG/jzdzE2xa9gXRryt1lFU6iRmFTwKLZlW6m2GcJGWtnAHi8Oct3FimKx2
d3R8Z96Pavzwn4jWk7HGZMBq3r+RG3TVZEaamxlEwuuP1p+zPMSOVKrDBwOCYaXv
lVSizZMpiyg4qSep5ztbqiwghAHm4vigBJAmwkGQZa+j5aSuCxk+3WTk2+QqFqdY
qGwaxNAw/xTK/qa2RWwI5wDud+8dT4pLXO3u/EqHk+N+tkJZiU2eqLmRni88y1L0
XDPQWnpdFrqgYyTrnE3/Vyivc0r/IEaBr8ho0OINnuUwP2pXWvPPe+3emIpYLqVd
dKtI9jBUQATS128ZG7TSa5QzASlW3Okrb+tnvwxxCmXL7UQ6H+UQcGfKQ45q0SYd
Q2oq59mSOechjR+g1ix/a60aCzlErsGbXtxq7uMcCEe2BfMrG4Ll/3U0d/78G3TX
YyG5KUALXR5jGmD3E68YqQQbZ5jnOpaESEo+dA+3xoL5Yfub5hgFBQAvNzqWvwmp
vXYiTuBQaQsFzTmDaaf8E7WJvpuKOM+1H/T9eFjWrSPNnKJZwSBTP0kjh+Y81Jix
53YjI2NQMmYrKzVirLcXpz2szeYuWDeTOCv0ciw1M2d78JGB/u+X9PfaCt57ToeN
JbZe9h+UyuH9CkxVS0hYtOGaTPm6j+F2ndF46HsTVPuX4tnq777xedR6bsHMrj+n
8YYGxNPtzmYIbqCyXLN4VOBuluW1NR/eRcs3rmY0DjP2K9uHBTK8rFlVZj+v16kO
8gXG6zhIx5cjetRSpekdqPqLLHYcerzYSpGvUkyEs6SldFSLnNoylqVa28uXrWer
4YAWnxRGCbHdKl41SJtEbB+xRTz5kTPlJ37OMs0WmSWYmUmHzvLlHTp54NHZKK+Z
OX8TUC/t0gZxhLVZJ7ovL2ukriYhhnnCELuiD57WKqwfK9u/BsnIuR24BvkmCIZW
OrVFxAhsGj2DfNJTyvVjTWorJwJRtHamF7+swmSLq1xFNeMvy0mkDFY7cS/jilTb
H+WCSMx0rZ2NJfdUX9B0TXcpmVkVImvC+h33OCvNiPcv5iL9kX675y9076zZjtUX
2DeJU3/iNPvbsNNbWJLei7VDrzPs6NFZaq7VmEaQNwNKaTFvoLA+dSIciHrvPu5W
X0EZ5WQnu0N5jMbaJ/eyALJI6WS+1BahAINlTAB9Xj6OwuQA49q7MqTRzCr7ASn2
gcPfxjXqxFT7Iys53849mIKOrCy70+cAMIiesd6ckp2/3em2iSgLvoPVy2Nvq7XY
Cp97jljihkQT9Qb2MvHBWMqfaYpTmhiXEaIUY+5GJEwsnUw7yIs52MlGVK4jQFPi
bdazaUJ8t8rlDuaN9UZhe40KlQRcUtKmZVzSxE8hJp6bWDICoSNMm7DNUkwaRXzX
Q8UmhAkmayDlmXWhF6GzVLRzwAW91yRS8WQ8Z3daj6FazPw9wGObIt2giGsK17Lo
sR179krWGb+Pvx6GK14bciRpPy9hnuPbAKP/z2WyIgU9d4XzZHTWB2HVyOZ7uSgT
dYV34Wf1E3uvk+5izbKLX/s+Bh3EWzYxEmYuoqKMIWDKA6gNhZKK/g0ePGjYQfYv
TUNkqSSZrIs6oPGlt4YsxNQlGOaR/+lwTMf7ZkA8R4YFb+DXy7xkIvkPrB7tyiny
8uJ76Q7KM08DCIPdf4krN7Ny+vP3gZXW+m9ryfYj1QD5SFzOajvDZzY37bt/Ceye
CsUYVwy7S/FsoKJx3J9ciyTcbS1EeycGmZV53Rbz0ZZsTUW9MGl/GsEWPjCQdD9M
FQRm4i/sFucahzLGNXiIkgY+CdKZKqXCNWAzxrbd3PPtPAKVfkIm4wAwFZ1buxtc
5CxxRoZDfT4/A/FakBO+MQ9D3qDtPGkQMDMVoNyxQhThqaIdJMUWQnC0xy3kH8oA
O8wyQW73SyLqFWSSH39LOQF8zrnkO/bzqpKYMdEjrYwHXEHHROc7E0G/YLgGKKfP
J6X8ZcKlOUIwX0vIAox1szzqP+fznjK2tqfghAyiEWlPCepFlmIJx1TKO9jTlWXV
X9QhwLI9S2BzW6cAaksAGRK2udvOFW0Urn6eW+tFJe99gnYoKcd9Y+xHVPRvsxZ0
HeHanySGiwSAGMk2cVKpHB+n4q25LHL8js3DFs3DKLwLgerw1XjfJjY/zd45d9xU
O4FDorY0DdP1o2qRpy1PNwOtMLqsYAHT7coJfXO3bqB4yk3jrNncYUCxCXxA5tvi
7GrDYWujtliT+Q0DfB5YG/Fj++VgvHn6H6VXI6LovGsNbLE8HyzkBpIhvewv758v
BaDOwuW7zJOd1cP0RSj8h/OCUrlK8tz59WhZSQRTL+C9B96ZCyoONs4SAl2jm6Ci
bErAPLT9676zEHHak/TO7hX6kAuzEKsmNwGRQfeNHZoBFxlensKxrMlINMG6XOky
GVys6CI8LXXHnTVKtib+D03mM0ST46VSzOptTAe0Vuz5VwLO5ema+vDwTtsgZS82
1KMTc1Mny6m4Xg8cmBEJXLEg7qK7Mz70gJYjUCgkvnooBRREZPSEdUI8vE2VlpFD
4IGttGr5l3LkMP51ahzcKlIwl1wcxf1jdNAhBG70A1Qsys+8TEuST0uT9C/Q3sev
PydUd0SP2huAvcM/ePgRQuxy//H+v7y7HARY9hh2TiB87TdfWtoIU+MSe1FCw15w
6QEHp4ZljwafieK4I6UmvsVq9MU4EERwZDB1siMMiEu7S23rvjnxgplRDG/gzDRt
ZReoHvZYDebbc9NsHeUqvr9RAVUdHicEy7/F2Mk1JZWphT9YosSietFYty99D8Ax
BNwDBSYIIwWURelNsc+OWZSEjMG5bf82gJgMZj+b3x3I3ld9QNIxaNnq2FhM39MZ
RR+hDZVFswBvj+zE1u+W6sk8f8cBTBGFSa7byiL1dEcc+n6Adu+dQD0GThhfTulI
0W/1WHcWbSG0f8BnhbNefcpY13cdy4ygxlsS3/uuh3Dr5dzLgjtSoKrAU/+1pdPa
8zrRLBkU83yJ2QyjcQ5O9DqmsJnC3di1Lo7W9s/11hph+Iy4BOOScKTgA8GLvnYk
h3IFX+vQGOaU3sZFRNLLahBZCj3iv7l1cf1WW6AAFNcfP3njlR1mzp+sKLJE1MZq
i6v1hcMeComPyIVpdyzuHfX2RxsPLjJRyKzip8WUAVGZPg8d5Zavzcv405KhUZYj
P9NwyuUMm3Kd+KZId/ivSNHkbk8gbg8KUhoc6RiOsK8XdTD0f9dBjlzpoA6W4bP2
pn8Kb3KbAc4IpFLyESV+KppqCp0FthE2ihIHabH53Shd3Gb2aK14qK+sXOkA/BGw
WPgY1/itpAtg7rZDEMBZO+qwk3pxOxGfDxV7MGq4ZEv0O3RLaGpuK8NkgKOvIFIC
r/900TRq1SLIzP0s/O8U94nuP5R0Lw5NI0v2PpiW/ncqSjbQDzCTPzenNY2vwWZH
W7e74Q9ZipTA1u8AVEVj6+TpJ5fMJX6lGXhsb+FAh4gKjQo+wfodceytMqaq6KtP
zYMpt5iMNvnAJM70BexRBP1DbQZHzJo41dtymg1ZLuY3WFy07U/TezIqiiVKgcx8
Rz/zRBYSMsXst+xLMY8rrCs0e3+/CNlyHr3BJXaB879GLuj4CweGCDw24H5bjAB5
8bRXgkNpEXUWvgZ5lb1DsmWDxAKk7krepchPEuR0ntHFXQdIa+Rt8j5KEha7X5eB
xzbvWYIesBO9JwZOb9arcDW8Z49DxLDeZ85Rpsf3u1UKDE/LVc7OCftZGQnXmOU/
8rfIFhFOXYwPNyWtPlyGapTTHMAict0wRkTpiJ9u3TLkIBoyNughPBQRa7Dgt6pz
XCwjLdlpBKJykzvvyiDqLitrI7vv4pKZBEI1HPJMPsDGCFzdp5m82ie7H5Nz3YUn
cQ2EmkA7MV6m28nXGCUocxKb6qRYk3c7HgVEEWaksJ9VQzjwh0p0VOoE+rsP2sXb
Ux9gRVy7MHbnlg9jvbiKSpZzKZZ+TU8agU4sqbUrn5i8Gm0CGtpQ0rlT9QmGtU5w
0YnqS7iwl5YB4+aoji6frGUFfWUK37xQqvIWntnynSzNovAKQGeXxOsJOITSphed
oNnOUl3CGvetH/N/IP2fVKPuKLcTSbzRwl/gEzGmG9R+Z06ryPSX4ITH/aoUVCql
XPooJQIGn2yt7Bov6N5CdgJ3v8dUzotGtwENTK/9LlDlV+Uq5GXhcXcQmrSFPsrE
dyPywPByX213EwSYt/JkD/jKDuY4+p/TtvzcJgLaQvW4l8JabcV8cNuy3afsfD2V
tztZmoT9jCIVMrU4IwgXI9OoBLI68EXYJ0UBh3DoOsUWE2KGMpUvjnQRwhWHWObn
yXruqwucVAuHBl6UURP+8Rvk04jAfJD51S4+zDoFVgxZS7PnJPfB6tJkQovYbJHS
xlSF1pyi1c92RXXNeew4nSDHY8iKpSLULIbBA52AxrQrL/OTVGhKfqHQRB6oTEQI
r62pot5obmQ33lwZU7hjg4O2Z6c5LKk6qAG8lkdSwajUifwFmU0mXRZDc9oEW699
wSVJOMsUzy9x6lIwhrKoLDH+fyg6KmVXJlk7qF7yTyi8v4nW7HGu9KS9CsZ89ojq
m5q82e/okZudCSg19xDm/rW4vULJKS9+rVglWOzXRF3LQTGRmLU6s21twtGcBWv9
8IZ+DPB5hC/U5dRyGsrWsWIm8HRf0a8X9lFfvJeKUs/QzGquQXn802rkrEGxy9lJ
q3c2bB2DY8/92dqkc79lm0c7gp/YRikHmfzB/+4Mnpc3GOiKFznKYjnk0f5BZIY9
/AqdBW6QqVcEw0B6IyM8lfrmRuiQQcGAeYkBbNarYTs4uUyYy0ELSPhHrfKsXPKq
FjTTkLE+GE91xZxVm7XlkQxDApx3bMPUE/O0Gg8nNNJpadoI0oKnKQ8Wew0MNFKH
7a2axrxEMGBND8xdf23b4APzPBOuKBo2awOGAkibnsKC0H4JneV/gijbMx73Bwpw
FYsQBd6Pinf9p2aH/wVoXUGo7hwwMh2nfBhR3bb1ySb0Zar5+ARUy5NPw4pSN3tn
Tis8L3xlFsPyRdLgXleJaYi5CQEs3WIv+j3tQCX2MJtuuTU2Bi005lPKIHXDE+lo
nYrWjobMcU+UGf2kbfNlLW7Ds1m6C5IdXg1qL+lItFKFDoYTKwLBfg412S4l6785
03rZ4sy7vSRB6drFu/JqM6K1Kyc2PKXk7qTA2aOO4DIu64/BqFicgn4OYiTz+DLG
EVNGNYhkYr+vWvfkz4cGTxbeepmRcMN9mRoTWu1vf1J716Pw4dYtp3kaPmfkUjXH
XpqzhpHkpUMPlXJ85M0pXHCEaQZ8fyKIGLvQAumYzJNAyKR79X9lSFaRFlg/Qdbm
i1Yy0dxgIFzbf9omPrqQn7jhP+PUGu/cxGpCWvDN4h4Gd1MMFPN7gu/pcsUIDro4
m2lZUn7Z3KKw5zM624A1Xnmkk0UQM2hmsf4b71QZFob00jXtbWwXTGjw8crWxTHo
8S1AvkUc1Tps5wmMcEF3HxM4iDYTnmw/PYqq1/jQVfZXJ12o59IflP7kfAhFRtcj
jAB1Xs2f4x4AMhmFinVlk7CJAcpAcaF4p9UAFJ24JCmVnzWXcJNRSPPuTbeNMyU3
nqZlbQhNPvv+hW+NYqxJY/wbpg1iNIruCCfqRHQTx0KVCTw8XYJ4M2k5LuwELb89
/wEkDK/7dLh0/4WRabARyTod9ajTE9uftgNJMqwI9jaMYiFcpt/r5LNg3yjDu9eD
hWMbJM+p3u4TyREF9bLKP0j2rgCRd6ayTY/C6x5UXQRSCTvcpPnFg8oNjze4Bqna
DBCqykh8YHaPKnrJDgZO/4aDreKxpch9Yi5bldrE6WxACsVZa2ivtyyuXNf+vq/L
tE6Ny0QKbRIIqysbV9Eubi6CEbDBvmbVliJHfLyh3BwH9lMbKeIDhFzyV03sbS5X
EX1b5HXAFE6+wthpcnu2Na+ugSNtcRVZpXOadYhYVw5+WG1t/kkRk/vqebfpD82C
5QszR84+H0Ezif9q4K/WIVNcM2cg6RFYfB5eqLQYMHtAv69eODwP8matWMI1uYSQ
Owj566iJuWnFiSHvS6S5LSe9T0NKpmWyqqOLy8mP/Q3W2pvbFI80gAG+87u6yzIm
zlRVmaieJZCsN9SESL9+ZOVN6r9XJIXl2cNOo7bM5CUARV05kExpQ4K+ndUGVqxL
TKCJPEdqm/n0k7CeguA2da3p6B439wWSoHauF6zl/FBkeFicLR8kJ/rW9ao1JLpy
FJ1/YVat+N9MSLPNShwfMr0HhUk73fG1cN3B80LvEtH4rwEQqaVXps5vgtRp+8s1
bjjGHfl3+DW+jqwn9vjdwaZWREohyy7i4Xujh7gqyL2jrSMo0Mmub/kv8kdfDdcS
x8HJQD0sofjazjOBLLZxO8RclYP/pNoD9VQ96XvClLj0hMKfC/r0LbK63PlV1h0F
TCHd7XaRESY2E/bnWs30480ri9kQH5i1SeamH/YNd1ymVGjJ3ps8hGxiMwhpkode
EX79JHVdxp/wUKLNfFiPGCVWzyvELmiwcmByNaPS7brHWGB3Oexc+S0xEGunSnSa
iUEU7IqpZp5vGLnRAg//JiWzOnta4tq+KVEm06Yl4sNwpLfEUFFGMa/Qh1bd9aAx
UooCDuR5u9Mb2g8IXWL0WLjQsghldVXa3BDpWDlAnVap+0k5YR+1EWnyv2bOPxlb
43wSs6AjId+xgpFg/Ti1emVO7q5R952EtfbpNe9p06cHl7xBjXVLbChhdDIVRW7Q
GeB/CZdZwCy6J2Sz0fwEItddDIvnH7wrFeYHdhIVMd4qIEgL5CB34EvuJRlkjuXh
rxjA98SoS29JKF+w3fCCczWwJGHstoPb4SRsgQY63K0Or6z1uCcO+VJgTmazhaCH
KtqTLSmJrxqdt2b0Vfm+0ohRCsMGeD4U+l50PDCOjaKdDNPtwfer3/E2EP9mBG6l
VR8F5F6Z0zrDidLr97xfO81xcOsawoQHb+CHV7HQ/4FB/WQf2e1UrComqI9h/Gqm
dFjiJfIsSWHotg+w0lS7jl0dkl9iesQ1bGWy2tTp1u+EBJsZQmm5Zm7EHk1S+eXs
g92TKebfUovbzCodEgEBraNf4hOshJqCPaL2IjcuqvM/73rFb4frtdDz+3QPYUkD
P499K30HTdW+h1At3sOI4ebrYtA32W9r0nnkwlEsPdsuzyRoYQERprqyt5K0l4rw
/W6rZeMsxwvKEnpBNfjEA5Q10BtJGpHGTkxN+IccYfd4HHvpkXoGx7f97OVtt+ML
oL7Yc/H/4tPTs3vJLFpSdSM7a5nVjsAKh/t9vSd2V6P6ib2hLpgWWm/rW/sYiDyo
dJwNOwYyRbmYUYTitRNL4dGyi+8+Ixy3XcDDHPL24PXJE5dI5RwaD4F7BRwu6PjE
qe4ZqjMGa1OwOS03k6jA41at2qPL54v7UgaPkDowSzYxL+039+o9/X2IlycrUkna
YRkZxHBHDAYv1FHRLpRjK14nRPeutM8+XvSxr4V6LhJEJNmKa8MjSl8/V8ZK9zOY
UEWjkVUIUFoN6/6koZZodmw2ACUjHs3VKN3/firp2pPLr7ccrCcUiJLEeLyPqzIG
qV0LRsmS22i8E9i+UVgIHlpJYcR5fd+8SvgYsuWpysHQ0cwVMtDm8n6av0IGgX40
YUSLAoDLzF86eZVV9PC7sxtWorOQgz84+8SWBuDb5pkwoJhlI+RLMSi3Dkg3WNo/
Hgi0O15ghiXDuWdqGb5LkCVyT05xiyOz/iUj8p8RSXEG3ePPqOGTEZzaIBZxZ+xY
tUVtdpHPm2cuQv1Ybm41UUUkBIjtcKwZPQhtHaglxYPmBDfm4SZ1o6PsWraQN+kN
QZWyBSjmhmWy5V4OYUKruVbMA6SYTQlGveMiFQyPqo4L8nMiovG5v7kb7KsJztyf
wltGIxvvpQbRtfkRTZul/f2Ru0clTRH93TfkSmpv0+mftWCFQl+uYnTeyP26Xt+Z
5/LsEQ4Bo1h3bdzIHhk9YkITzzdnb+OV1p3a0iK/CEH7743rnGWLQ0gV8YoxJgRg
mgKpoB/dz+KlIInpxVHwqIDnZLs91x8uknBHzA4ofd1KSGzrcfYihVeojb2IX9Xl
m88EfwECc4fl4iMCOuz08YuVJG8j8/3RmgSYDshiWqWuKOIj3ZQ4alRqzbov+bIU
dujefoIwO1Jklee6hckFleMkl3P9VdDGmt+RJTyDvq9gjHlw9Usut+ilLjnnzLGB
wPY4rRJCrno+EWDJjDkGcutt/ggdsAnMAxr8hI1ZG14sBmYhTwrnFdP4h9aO+Epx
YOdIzNmoETr3tJE5cS6DQJ7IV02PiNpu6w9OZKvtQN8YKxdIi09W0AKP+4LfNi9g
zlhvX8sqiRAqOiO/rbOL9acs++Qr83NQm1A5o7rVPnq/JqTooCshJ0VMyaWw3JFF
ZA4kVCUAdGhCShXq1xONx6dsi8pxLdEkAUfmJBw0nXXH0j8xUAbR9obwAvQEuQg/
ZIolhWA/2oox4ms600qHTsOg6+qaC2ICgoS9SOgqsODwBx9QGlXAHLOUuqqxzmn2
0mtofOj/VPfNmC/P+q4p3+ObTWpCdBiB7HOTcTleMCxyV8Uik6Ka0gtZPXd9SgwC
l7nvCxkJ2WcGbwTw3DcEsnvOrbKm215TCTl9Zm/D5LpgvMruqBSL5oI0C7FadYUF
lxYXg1qkqP4ZfC3lwphv74lNOScukCqiNwfvnycFCYdJ2jvdT2RfCgZkocoGb3sA
lmfwEhRQQn46tK42RLAeZn4ITedIkQr0uY2i9w8jBI0C627S0lMz7meYZwUxotgt
y2JYrX/PNpqryypJz03C9fhjQbchyGTgTsmWl0x3fmHmHWwGER8EN/P+b6Wm/GiK
ZFx7Ah8VDKi+Hqbgol3oKuVqmf62HY2slbWcSdMlWbltzolTUM95vh364Bcblqgl
a76VM+GeJ7w3VElGFuoKfL5P0Zr4VWGOpiCtVCYP5SiDH1lKK3K9zaLQ/av456DA
qMNkEjqOndUPD/n8zwDN+8b32ivBhQDAMa3xN4HgH8ocTzJ5Bg0OebJ+BeiidtoA
PL6IoVbjW3DsigMn+pvX1qUBnbb9Tn3RIfKJACHZojYJ3RTXhVk0wraKsvwFe/JS
onKxYfVGBQ0ogitvNquKKH7HWJnwNvDV6jqLHUjGLtcXbR+ghR2eD8hwL0rzBtFr
vtdQZsbUkr0oD8AbX3vSoAdmPZudQDOHN3EkUOcvprdUVJQ9VcV6zmecp408/vXt
ZdRX25I+ffaXUzukK1RpWeJFUEuyeTsbedIazU1MfVygSpxbXQ8XmvtfYCrtnT5I
sOxSZSWCTx8ynes+qd2JxjV2U9cmpG1tnbDdS1SF1y07pyssl5j6Il0zJZzhtC54
GmLk4uoOl5KiJj5BuE1a34QJUQ3EH43kmyFaboleMLBxaoOw1Qa7vxpQtRutNoLl
4e6QvSMKgQzsv2/ddYRFwfxYsiDhzd5P6Zw+2TXvhqi/WABewaAIMyg29Yqh3uDh
4xnewChzS2akvCkZNnLr7TAcksw8jy+6CvvmZivhNm/zu4dp7RMlZ4+D/CXou5f5
vgrhWN9wyKMC+zRTtI6xatXjfqxJ6LIePcWcHSbNxYamhz1d7htXjWa7vBA4Y5gN
3FQ2iuwRwggvAOn8CMdfMwQoiwrUtNApWe7SenIVbvuByv9d1286xAXHlBy4xyrH
ZF1a81+01uqeWvfqcaMShp2dA70alrNirJoNUY4nvVig41NSrRzWf6tjNSUOAbK5
GWKMmTTd9qgRiRAYd65+LOWx70Wvu6dk93ODUqEODBKY+Aiyfn9hKRX5YnlTRkBP
/AlZKB+SjEqKZ775y/3B4wmH2lNm7oaINGOdj85f4cO7fqMYeEQJIxSoGqVFaKMy
0VlbKd+zJLTGnADnNOxjMmSTECnm3+0s3/YkecU+yv3HLKc8j+VHhXG8jlpgrf4v
tzIc78fs4rUhxnwMNjWTs7jOGXMi0RBuTXm8fKiRXsvMyOKYno9SOIUjItU9sLN5
tOqRBlnLHNTEn+xh0Oa1wNegno9I1flTvgxwHUkVRtnfCHqna77L6yzbgeV2wP0U
CQ0rvgDEo4DCQDBJu552uE/W4gOJVRrE4M/JLNmFEyOmwu163t2NkPmds6mPqPs8
+JfL36uGd3nLUv9JqME3dSWASxr2q1Ky8h+sLcKBtDhwpDm+ngNoTpiMcC/fTUQx
+fS2OHJPaTNE89HFjumpRFfKqoeWD4e53j64ZgjdQ6hsCw9RcFxE4MkbzcCcQBwi
7z8LFYRBoRuo0RSRMBJ5E6lNdK3wA0GdcZs0shVy3xDlX8Brt7TQ+diuUGZMAmoP
DKZXjxTYsPt0o9gAqzhYm2lURfvZ4AZpTi8k6ZIVciJ2Jah3DhfdDT8yil4kH3tz
DNf6HT8jESGPiEJVY95ubqagFJMocwE6+e9kzNVM1bnyeQKxLTK7I9xi5qoDdQ26
CvLhdvpUZHmQv4K24hPfPOzqa+Bfyffd46fpSGNa9HpgA2hHyxwE2HkXEl/XGQhO
JW3rSU3wwuKFNtiKcaj2kJS7V3o1/gIlqhqvQOZi3K1oNaHIEHupl6Yukeo0Vp41
/1HVKbz1Cxc855pfnWM/maLZE/ECUukoN+CLcF6djKWwTaoZyWJJYL1Zs+tX0fIr
FsPeu8eyQ28fY1H1m4ZgjJbxPgX2k+gibviL46dj+8KKV0OR7wfO/SB6qk1LgKnv
Sqb/NaDGest5+Hd01SQMQh2rx2uK10H3H3aUS1wMamL6wbYwQdTiYNieR/IidVOq
Vaj647uOPqUxYKATV+S7FAw7jqz9+CUOmIaOgdR8bNuDT/VzqtOCQy0Q+7M0YoIH
2I6APNIrQMFYvMCCXCAiX5Vrv2iOIyLw0MRYD3sCBsRs52JQO6QC84nJUzNjD06X
HkADkBcmzJY9PNsGlAFCguylKEG5fOdojOLoizjqVeXca/OCSpWDCoTTxjgmRA4P
o7GzWb11+0jCMz370zm53xOUWcisf7a0V/0Bu8I9h200+EYbQEKzvhsWweVSlYko
BhFjvj7MpW48LFzYUdWGQqqcI360vEhA8EhbWo0eWGwtWYlfw/QNk7DPJ9Vu+xoz
W1vpUfyA4DSst9Vai6XavXAb1sWqGnhGnR1kHbUcufS2j0didU7BB52O5X/aYUln
eOGgaOEC366XH0McjhFHSN43uvOTeiSNWdKz+4Mpfoc/lSCh/Qkx14rwBrcXJuNo
97YisJnDrSi2NYhp3WvGNX3aCMjLK4DTx/HOt/ql4gxodNvP0GyJF8RkY88/0d+Z
4eG2jWkTW0yi8OKgG5dj3zZp5MlmW+5b6d28cLDCziOlmzi6SoCHQxtCIdX3h/X2
/5ecPT/6HWDJE15/Ax4GQ6YzU5k00SbZiDWLrRPT9Ol+5oQWeamn2cPCaq9d7Lwk
e9CtCZNZ7rvipaKRMg5eBLXAXAGpvqWQ6bbYNEFZ/uUpJ6Y/SXR43jClTDWdqvea
qMTH6cNDQcWLUiV/Z7z9Sz4NBeEwN+Ev52ElJu4MSMHgETRtNP13tnwTCK5DpXi0
fxReIN9nC6Xh5K1JMTci3zM2IUnXdN9f2NSqdhEA29tNxuZ8zrUtGXWc7cPx9njD
nM1/1IPp95mYMmDG78KxsY6tiAO8MVKul7u2no10Vzo8SlVEcPo13tl3hL3S2qku
TwKQANzc0OdZYGEzkk7fhGwAouyD9wLqQO41XiI6WglxzbthuR8AFnDpsR254RMn
Wai7lo61cS5mrXP+s7paFh68So9cViyd5FOiUDaGp2YKB10KcRJpeN2/AJI0Ktf9
Qe0ZiVsf4TduQ29sF6kn2a7uet44dRJh3+C04aJ5/u/r7EXEXz+ysTU14vQKMTrb
5zGHFdvqrLV4DDM7OBV1IFmTOG8XHimlZzMlKiuBUlk/GvmAlUu+sgNjq+8PcYVf
1tPGFC/iMhai2DIGA1ORME88T0ZztO/SqybxMtMsysfMsb/k20s+4khqCB40+gIJ
b8uws/TJeomSm1K7qZr7LrqjTG18QBz1vbA7wymDE6S2vpDUZAoj5OkPdYunCejw
3NgXRr0UXDyCiRwIGU786E5+C0CSqIlYw+/PSVgiQofhha4A0LNtVZe9XVfo9Xqp
LhOFl1U2bjhOlwYY7uz6mTQT9kYgsNQ2L0JPYIunpcvW/6VzxuV9QrRYIW6+GZ0e
7eH09o647WLB0HoKyqFCtURkBXQvoRsdEZwZKI6h0bf3Z17Kxz0lvtVDrUSGfG7A
vE4qierQf6I0URDl8Z9Lzo+u66D4Eq3WNpCv6eVX0JdtNWTyR5lJJmoBmhiwaeOG
f/NQIVEgP1a2iCT+Gii5RN6FscbmRNYJt/ckVL7RAnc/kfmVi3ef+rttsO48XPZ7
+h3qw0jGiiFBUqDfWKaLx/eBY8sn2bdNx/NLTwqB3HRm9Yiytw1oqVoJB4yvpZmo
q3wWHU3c2+DopKmGPwH22SUileLpcXAS7qrRVwgcIqihlqVcF6tekOG1zplARRTi
26FYYdnq6mrrNnFv6cfaQ/wvjgDN0IMDWNm/cvrQ1xz4yvC2I3zTIU+KvmCIboy7
Qi1BPB+oDtNbVBAR67RF178rioDhkpYXDgRHRMM9D77oh/UVNJSpSrTuvYF+JTu3
7+mzb7cqT7bin4EQHwc+vW/TJ/Ltx+AQncRdM2KoYvW4SUvqk7DyvHY5tk0znXrD
t0aFxuxCn+D5EywvaT3g4wLkK/jurYSzVxmPSx+5S0Pjs5+IGhE8O0J4aCYYW9lr
LcZusSe6FR4wjKdzyvGpNxdBqFZr8Kb+fFU5hdQMb4JTPv+ASWAxgJqFs5/sBmoy
AWh82BllVfN6/7b4oJ3RuAXZDEeFJgzQY8NHN5K3HeccUmba26xtk5wgPgKXu9an
UEyRcVF1QIs8EIny8lsSq2v7hzSSAULH4k0jg8Ws9PQsG64gCVazC4TV4RSUgAD5
SiJREXHYVgKIfbQSpoC3eiIX+jqCdA5wf1XrMpj8tSWbCBVqM0JNyF1R5w9MTYXB
4by5kn1k4NAkpn4Gkz9d8xXpL8S1uAApDKjo47QAEr20yw1cqIdrPYKEvmok5a3c
X/rG3TqHVp9cEne8QvXtI6jzGI5cCTgaNYDbzZobElKLrbVqQEfSbR+TbPTCKRF7
36FJ3Ar4G9Gb0hONqEzLcyZI58FOoHz6irOjV+/puNGCyphnA2JA8BIlnf0Do8AF
xe/6BZRxiankJMw/FcOQYb8dtqheo/WvDZA4zWksSVa50wpFv0JKM6j4ReYj87WP
gwi1TmGzECGf06Wvie4zP7b8IdwT74mGOz5dsXab2m61zTxQHIkmMfdMFVVvjxCb
Y2voqzaFVaw1Pmv7BZuzuYA6buwYopt2TrutPaybrEmKSPofdGvlwy4QwcnMOTGK
/uA3V7GX+0fE775h5jnOauN62khv65vfSLa65r/vCK+8tdxOW+qNxoC/gx4j7E8W
PQzGasyp03tsIS7nATY3t9g75hqv4LmoNOm2VJFG1KGxO/DiW8ILdw2Fv6NDkB4M
XstohvGGqR/ZCciUi38SUaByMmGuedfTP+/PC9hQuW3I5/17lwV5xck3vO9MsVAr
0Wh5xaIA0AK7/BFgEACkJCQplHOkyyWFbXXIFUTz5wfz2SNfvGCV+7ZbY78YLLBh
O25ekisshnz3EwULqhmLbvjTpbbiwU//cILWXbqWmmG06giE0AIPVdDRW0eZUZTE
em96L95wYu3lEvSVt7PiDHXY14Lqeno5M5aWGNBYqiQb09Zs5BHTdQkLgjKJbe3J
Tab8e1H8lMFEIzuRy4w9ZO0v4iR2CPWSIQLgVU8zVz6xlT/0bLMAtDB+uUwObcQ5
RpusgQghsqgEdxvZgqLdgCQOXhAEd+7Fhrti9C/SoQmTkWxlxqjFh2oGOz78zN0r
iWeRljgQ1xEdsdxoLjHHQGIgpd6Ju+Olsvg0yc6YoAFaQEemkI5ZVT6uof+JLhDC
OTugXnp7yQvZooPx6euw2IW4HQJPQmWMK7najHGvrpvl2C5+AUJOmTmR/kgwZlJ7
uMr705ht55SSbQy6gkt7NgNKMgsaHdtb4PnRVuVE+l1lghudxvaeCMewn9nrqcL/
MotnUOY1ataGvcY54kpkvc+SbYqZ5svw5YGCl4i66l8lgi94u22+we9jiHDOMp5x
rj8Jxc6JcgwDHEKblGLPG14E06c5zH9XCoViOTBKBEWhvFb79jVmWlBV5NT95/I+
od1hY06F+WVDJQxQky5gr9yQiqPSBv7h71A6sZJLGweOm5WRTjTOrIsFxt2A+YZD
Jil/awa0pynmDgHLGA8goDV37GpvZ4S6UY3LOARlNy/qdPxOslqISOXa7U7yPApK
Wd8nprrN+qeYwFG97UUxmoVsM8zuuwkJwW2iY6RNCYmAD6/MGoEM+V3PZ/ilUvzo
hEKn9f+EUN97Hj8m2fPZoWzYmRgzUJFJ4IZVMtYe0fK3DyIdpHMe+V4LhRi3ujws
/9UsyFADAJrTOfgLfEsMmqzz1R7hH5u7d2+BDgRgQWU1b31KaLkewIWKDR75N0aY
rtJbbB+UBhIqOkRNTtW9J39R01PgHp3tTxEhce/RyplvmzSLa10whI2OUjgvg/cM
VdROb9YFq9trGv95dxQ154RgkoFa/IKvuvbeOJ96lAoVh/zMbSszB9X1QluuZIna
LXbw0w6hUnCyLzRxiovP2v55ENirBasiZIqaqwynWmPqi1miUOl8AM7R1WSt01Os
M02SynoKFONd3vNPFo3AVBBW7tLPGZn/3fvh83BrBB8ML+UTjojMu8zyI//Cptv9
aOyYTQdWNRdUyDfmt+lmdv4WP5NkOVnpU2ymR1pTT/WaR+eAQj8j3ZR03MdglBGK
SUBN50i5veQasX3w45zG85Z018qxmF7HEnPfqNHctdLF2Hd+LH8N/1WpGW9IexDv
CoJmzxQDEj3cBheq3C3/nt1YEigcMH+j/4NSJytdHZWZmqXWvcfY6y1WN3PPjsUJ
uGt2JnONq1jfy/DuqhQVAUGfJd9/S147m2/uw1S+lKmxptAX8I5p+7KNvPvcf8jr
CqrYsamopf7I2TTe4w1tT4KGcLTFlWmEPCDplYgC+5p6EHSjGWOaavT2Vtn6FR6f
zpPpBw6cPZM/TbYuuqN4Z57cOkuQLbRaGoHzSwf5RgxQNcYW9RLAKW1UBm5bIesW
fPIHf0/Av0BQNTkA7XV2S3t0fWRUGHNDspnJkEje3X0yYoIpKGZEdUAET7LyhM4+
m+6v5Nak0KRN460gpmsbtSFPXkl6RVq5i8Hqp/+/cmZcCscnJeahZRfrg83QIfb0
ubu1tRhAc4dvyDz/0LQyD4V415sUqYv2eQI81RcZ8Dg0cmaIAqAtKII6B3hgfTva
pwEud+Jp7V744FBqzEVlJqvy3yHO8VezydRBnmW1ljnEpc8tsVFiiGq8/VrIOqrg
+z/fBPQb0FdyYkPGgrHBxlmMW/o/OeZwaNUSvMhSApTVj7fGxc9if0YLsrmFVhHw
TQ+yXTv8TRjJI5rKypQVvyuQ9bILycQJGw9GQGukv+/1XhY9QieYxFC1dp8MhlVX
W99IPVhK9pvvhRaoZ+Ad4qKBF9Q6gLeWuyFT1h5wSSbqGF2zuh7yH5QgH4rVxj5V
4U65KBGttpgICxnnK9O4TswMtpAj5Uuvnf5DkTFKYJBxTMrg4VAuixHUAB4qjw12
UY1RP2PQjJviv9Vd3+MC+7pSMey6EwI3KSGo5NwNlfwnHmPgktHzCXxbtqwDkroy
Az+z65ES0vJz5rlJp9oCtlECguyNNwTb6c/C2pJILk2+DOHSGlaIU/p7DwuJTqQ6
n4iMBQcIKPcSGudqHv4I63PNYdcmO2gqHFAm7an/VJUcygK5cbVzYwszDw/US+Ek
MLGfk3jmsAgSpwPG/6oqF32LSFk2TFVAwM9i+08gQ7jYWMACyX0Kaf3RRKtVCgdm
eagawCKx9ZPV+R7DfP65uIKrqYSOjoERy4TP0qlEt9Bv+9ZoIqKLcy+jfE1U4LiP
kSRw4GpnAKiZotE62Ps17tGYrpeWMvmKouOSDoqUGCdTCOBXbT66PiSsf/PqD1s4
SoeoiXOddkLoL9gsBn5TCQt0eZ0cAzkcWb5CKFjHDSi9sgbiWC5x+FXIDrwEdIU4
n6ItXX5Dh5tprIpatz3HOy5lD3YnbzAS+dkpt8ONw/4zqDla/Pg7stDokS5NQqwN
cFAaSmuwhjY02MIKTorkJpMBenwn9WAmn8w8CPmnGYxdHxuUkzIKZJ8R9GzqW45V
Tvomaz6OLjv5HjKJMSwDLe5e3zftm4eBywPppfu+9sr1NXP/1Hw2vIBo7SvRQWl5
UEvNJXboKirasBatgJK9uN5MdQsLgdFvk99vwx/wtGHghsf+JMz3XMxx1GbDTn3g
YaibH4zIn9gC8Gw+mvIw2pTcoztJEd5Pc6FKMpNrJxNJWRyO+UM2jC79Vs+Q0B66
FS9R2CBgB7Bai2t+sF98k72D0lTxeQ8Qd6/aZOKxk9GTMoxva37dMkGI4z79ZLZR
OiHweK1SUcw48wBOpb/r3Z/B5cEe5tYSe3fLewSTcr2Ppk0HG3i/YhWPadyoxi79
AA0FW+6KdqRJQ1ITUokK0x7OoVdOTcsT+umYTIlUrz2KowC/Su2dKDtFLf3fgi+b
xGkFE1ed0MU3nlslXCebAehi/0Alk3wsMUx6GDg4h2LnGBAXCS1bc3ccqbxYc99O
2JotThRRKB87bqw5BEGE9TdNjyYA+nlbWK/mdSvtIJUUm/p1XrdvD6Fo/aAxSL/3
Kk6lMgujHBwi2Trq1q42s9OJSYQg8s+xPBq4f9JZlHbWrgyK7/RF76S3onIyr5FN
AAAGM2u+l7NVn6wGmOqKm+ocB6deTohw0QlT8RBOlbMR/SxfO7tpCye0aqpLC2pe
BCYFwnaYuig3djtHttwLw2psIPh+TvO2U9yJhGXzWsXVOyEkLikXeh1o5yoXgM1Q
2jpqvJJOWgWMR8WH4n4IH7x5SiycvLWovfkfDxBjIuMt2VVRlc0lCkdmVarmWKsa
vsPvs4wNHYMsdDA7VBQt3r+WSVCWSOJyf5HA8Mg+tPM1AeyMbwrYvu152d63zveV
B/GD1mp7IDIAjHRUhUZAqs7w0vHz/ExCVq/lS7MvCckrJl7zTFcnRIP/vMKEfC0J
EVXdWM065HDWG/DEgNdQ+BfM7FgMdkRqXNXeuJj+QHv7S+9RP9BHQrynaFIrrSNL
rQr456qD+GI0bIEo7Ers5DfPCP807YXyztcXbQAQxqtYAnbbvKYq3McW9dDN+8l4
u5hjSeUUfzrx0cBAZX4S733ZLxu4K2ivSO/xxbdidB42VBrOW/HN4LtABIiqZVY6
mdZbO9iu3vLW8k3mjbpCvjBwtypWA/4O4Xcz5b7AzFYtb54uUyxYzlNkWaNZ6aha
Idazb6+dYuB9ESmJxOqpI+7Iew22Ucq57gqshUBBLYJ9lA3bUj2Gbz0Peb2kTYX8
rNfePg701EBXzs/DngcdpqRzjgwLWIF6wuz5ZqDvAeOlKUuPH06A6rguvZIbKrls
bnTLjA6y51NPpevCZpYFittJrXTq3kF7ijTlOwAWc4PjKLNBN8kq68plWZH5m6Oa
t8Tmq6Q8cZyYfQ3KC9VjLWtgJHyc+OMU0DRPV7+JcxyD7dmcGbOjhvXGNvzK2X+m
4g7ooJ9l/PqoTp+o91jcv2sScH7qCNpcF+GRmZO83UVD9QeSxMEW/qHcoF0jVDN1
ID7Y3i6THu6HtiusVg0Flv4Dnffo/MCZjZpq8N91dmyzt/lIPKohrrtpQ9h3Pr6q
hf78EdVVSYDG2CpdcVVirzEHU4PSbPng6jolBdBSnq/hvo7Layey6LMxdiUB0+1u
2dk6i+UIBOh+bOyURJ8s8QISurGtOaY/2QdaxcLKTyM0EaXW7OmjTWYiimwuBAyN
GCJFIj0rpzN8+m0xHrg3FwsTjughNf+vQOoxI9wmT7Kopv3QjIQY92kjcSsIcoWa
yK4F44mv1iADqJ61yVYfc8wPB1H4WVqYbaI9zCivxBy/sjAjb0UZCEt9nYSNO0i+
WcDVVB8Qtxgf37TV6CQ1u5FVac+0nFNzdXpGG7v2y4zC0spN4CDbm0kTQLj4h7Y/
Z6US3ezYOymmJqPxVbO4ZXciMPjw2JQvuZB8a40/adfe3AckrDnqHKstOkq6GX7S
72UXVKRy6mZglitz34rPLcf+kr0yR1Xtnj1PYtvosNCrnuoC7X0O56T9xACJyP4H
2KjrQ/nqTk3Ad6QCADyud7RDSLxXRm23+h526RrpXff0HdPYeqBL+x2tpEb4sPjX
3W/gMEWq8vRu7mdg9sevZ4ka/KVLE7ze/Mf2cazJBR3hOj9I35EYc7CYOwjgSA8g
WPVoRw6nTBko57z5YEJXB3k/BfTrwBWUvLx0dACdhECiu2XBYEUGmQBO5udmXdZD
H3FCAPoCzEJboRdZkalb3nnm3ihDOhUM3iy1SwwHO8Omdq3KbgyMuKQzl1j79fFi
wRhgqb1swKf/wfNvSxE+0UDs+DK9RYUrERExWK+IhzOypVX2WvJJ4PE5jnNwzCDu
WJE6MbVBwjdFruN+b0O/viovUk4t5vl7At7WgUmHWs33x2q9I4lnv8nlzrWg3mY8
5rQuLRZaPMuXgYfmFtdyITZ7I+S+QhOFQO46uDkx7LUKIyHkyqmDeQNy8vkVUX40
il7/CFS1lwczEHjqp/6etL79JQzef7GqKtc3bheI38lF1Qk1nYY4+fqZPFA5yreY
znsXwtNh7EvTuVhkGHnuWNASsPWFaYtAXij5RXLvsp521dui128vF58KmOzgGNlB
tj7YS2fs/mtIiillwcrzsYUpn6u91gkCkMNMjnG/cXthrd8NTzMTQf3WXkg1+H8a
rly7oxSuC0TYYRH/xsYq+vPhid82+wjl3b8yc31op01fkixwS72ev+qv7HXoKrzp
gaDylJI4aW31yCLwDLKc9AMi222NLr4DMGTAySlAY+fHoYZrwzg709yu71BDRVuA
oNzV6r7Y/y416XIkPeRN+M4kdltVxOjvtYgozpCoU0VuikryEqJgYg3W9f9/+q7m
D4owqvcrCdrcC5zuFA6HKj8iDQj+C3R3lKK0wsEdILNJ92vkhZaeXqdJeBIegWc3
IhBF9WxmA4U0vmD1E5lVe5Ku9pR5rtIp1ydyzlSb7P2hSFaIXCVge5F+arw+A8gi
mIDyCavn9L9SN0Xp2oZuR2a7YP/7UlqQJ1+yrE7c0JiujuGKg3GywB6EM+kapBmW
vyLoVQ7VwkNlPZbZi13VBhpmq/eWZq5/a19Fe7HUxXxtbiXWbuAweg+QDKznSP1H
xR6QU6bYpU+rnTwE0IvCbeajq5RNCC7g6rOKpVlg318CU7Y3oBhpgjVUt0aVBNnD
06AXIIISXR90Rx+OZP3+rK7V2GMN260ppQR08PfKQGzB+kKMABh3FmCwP2hp6vya
mZ57HFOXsQbJyWar6ZgHUTMQDtdXTgR0HUxzO8KIeZhqTM+7Yr2H4H+SP7QnQbxc
7SN0TS/hhKsHG91cGfok55ociiCK2796BEjwbgIY81hc4Bhh+e9HzPtMXNJ5je9k
W3U94E0PExvRpHJAXaCN1MQ9jHqXz/0TvOB2/6ep7IOjgqJPwi5kolWnte71lR1x
HUozu1ZxFaRCjqA3FMgXj+HK8uVerCLtDaUf+hYzhLc=
`protect END_PROTECTED