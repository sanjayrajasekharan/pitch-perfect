-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Gq1YlU8an/lyGBpYmw1139yfIi3w3NJtN0p+mLdX7heuRqCqqH9GuhcgeDB/sQXKYfBV/v6gTtXY
wkr3qYziZcA1SmxNdz6ktqCKxO6YnUw+dgG9ZutlelRQ/hiRTprotZwsv69kdjPjRNCVvC5jg4fi
p9dksJj31jJv0eiZlEj3NUbNzQq/ECK7lLacUHtjEziF6jerfFdaYahVF3aDhFw5dfz0X71b4ty6
AB9VuFAseVEiflJqS9Au/kiofU02SMgguoKIPLx+CFVoaN2q6do4IjSh03FnmOKkATBfBFtBSbhH
688jXEluvoaaUKQtTeDmWZYKikT9TC0NgqBdjQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10048)
`protect data_block
ZBnxKom6MJ4zmC1MdFp52I12VAhEP0iGzaAFZHqUXvma8A7U6JWQjHqdzRdQE73w3jJtBk+AfyzG
1ah/lHav9gUg7H+p5aIhTA0JQDcJuJ/qMvLypNc/lqzUbyEaoGWE9MSYqXvgvc5xgyy6n8+7Wl60
TjtiZWANiL9Lkyno9jjgoBm+jeAUiaqV1lj0OBBW7PecQcIGYwMu3Y+uFZ2nv/ktV8ipH70sxwt1
oVLW61WcJlADd3VGtVF1l/l/tFLWgZum/0SxVzUzuNKYDcWuvIgCEN701Efx0VOdzsg1p9tEnXWb
9Y+HqwIPS8H+MVuMZMxdNh1b3Qp6fgjFgUoly9cDsJEswx1rPc4yqrieCpXeBUhC6Z0MS4IT2gkT
OFuN5n9tLXMW23QVJn7cNgwyNtAtDWUU9gDQH8SorbmaexISU+7b4aw2mCakMtDJf5ECYHSp5JWu
eQM8nzR39jOaM1AH41kHrevHKxBGFgHGu2w8DFVxn+l3bMaktl4mSmGpZm4s7ZBzr721KDj9sJh/
rWOwBcItECNOfDxohfw2OZYxA0m3mrVX870R0GE3lHdU9oMu9KqdgDb+tGHu+9+9hG5iFTBVfnMq
lhxrf2n3GbaiA3ltGsH/bKRSWXUnxgSIhUgU6RA9ku6w9t7ovxH4hVoevivbP6H+VHU0FqcFHE8P
0eGn7zyLPHJfzIzrzes8hjTitnJDxIiVtc9niFwsnjjtecjlSuw/bpcMFGUUL014PbIzvBUjdfA/
Mx0X1e9yhshwmT8hCwdkAabZby9wa3sA3wSbn2ElSffmYqt5FRhhun4Sa+DwN9a2/2iRsIZRRv5m
55ihkrCDeVJX8gB1aPoXOtvLwLBmo4RN52dNso0tMitCAiONWO/RtLvTygXB3gxLSFFFn//Oerhu
e78/czr6Hddo/a+yyyM5+3iu/sQ3pTbuHU/Si8YkcSbQ4HeosmAIFaeUDRVJRzvq4XL0zyx9Jjwg
xzH+9XKPat5OzJr0n7RLL3TcH5YktYNPdoGUGUFeQRTsrkn+qS7VVGS0AjbQaE8kepycYBqVuZxf
bXCw4TmB501VYOcg5iDBRKuz2jZ9A47csl/Fsle59JQ4aMUTp0Ych9ia/mqp15H1BAWW7y3CewsN
bPK/WK+WguqrWJVy/7g4nVAEq2IXK0VxFrayqQmHFoSxmi2ZXO973HLLW4okoL5x1MuGAmg1SoIV
+/JpQRDWbS3Im93MSl55tVLNoAWWAxJvXRvOOgC3ESA7uQEXqTHGJQaIBci8nM1hHgUQ3f1YzKxe
SeT4liFDSfXLhXZ/rVl+ALJBZwAJDkzjP61EPrx30JORwR3hEF+63cNydRqdVMZBbecBL+ktPwCf
WwJQZc/vYR+OHOCp+2ZsIdz/WmLjGy30CfLZLDVKZgPLwpPPpZ0CVT2N+XW6/fC+y5IG8EFU7dz3
MqCZK0YiDjhNpkkQTifG/RuzO+1VxhGwVSDW8TR4w45BI84q8EFXgAyPkv3c7AJ9WfvKTcHjOltI
g02n5JDqTvkgwuhuwLzU+wQBEmLSlm6E97nuv0swNnBczbNxsa29Ii4bf12siL7KXUwtdlTSpmb5
BdqMaEybJAfR4LqL8bw/zPuZ3H8KDBoSbIuQSwXQ3ctOKB0m3ZNEjmRtmNh2cbibYjcT254V8Kiz
SjbsF6M5Be2uphV26wG5QGAtPxd6aLzD3Cldcnb4P0UKeApJ/jxyHAy8w0zeqmbjMwXpD+vF21f1
P8EssIwTsjcheCLTS/4+4XdykFHnmeyuyQHm0Q+nYwjULmJseVWoc75fG7w2kbQqL+zcPrwN418O
QuyiWdXAOZ2JBP9nDOIYFb8WQ/LyowjY0qObEde+OvTSnthx7zo0EJPAXmbLky482z+Ef7uFWKpM
EJnprH6Nw1z1bsnBvdS21ISJJbE3hr6Ke3eHws8gKnibN5t0NZGNeUyWxnzU3Ypvh6ofXTz6RJPG
busir7czH/AbmxZ+hvBotYf/WCGKoNIHsYcVAbifaVHT8oDtITdb4wbxi4z7L8KsfTn1945Fxb3z
y0WaCVvG6Jyz6FU4OtoNAvc0EQi5A67ZwwlI1uEleM+0uaYxx3Ll4KbuG8OT7bXIF30MSsbSKQjE
DD1vQ49zS8M0tRz4TVHkfYUCE39agFuDuNROd1XEutYGOihQZ8nc/Ww41AsS+8wKW2sAAkO0cq4y
sIIZECK4b5n/0Ri590KhWA3xKNoh6KDdHh2Ne6Pi3jpufn5zKEQNLf2ODm6RUWJoDAemivG6nEpx
wfpiKWQbAoDTmAwOT+PwsF6Oob2hMaIqHT1MsJae28klQCU61bG0A/QghgQCzk3PgeBpgxT8IIbw
84EXQJBS1XwAlaSCusOcnfbfWQxGR2KAlP4RURF+lPtlEjMhe7GLSM73dBMZ33M6r1GxEhTySYvJ
sz2JQy6QJybLqKVUiBE292NtpKE9pkcCdI8F452LymwlaYNtJDdUsrUthvag2xKAIWi/SWutszHh
arJhhObyHmN5KKN2ybYcCIuDygdS4dy4+V2GIh3/t50KnRoMGlC3ICaOxwCq93XHCnzbw+puN7TA
tPT8WwpUQwCpOyqYQ/7Pps743xoZAOLzvw0hOo7T85hTeOGR/NJ/KBljZdzprzhxsmbicXIHXiNs
lpIoB+FdydYMdbnBUWtTryliQqJlIidxxFgFRe0kF4HOo2jUkrrHOF6bBbUDKz7UkwaFh/S2M1XW
MX65aI5NvbxnOxGHjcNAb2KqCEQn8u4ecgvPT8p4ss/UYYTcjD2b/S/To8Y/EGzgJMDS7svnEPhY
04Qk74u1KSBbmQp1ZzAYXmwPGa0ZtaZExs9S7zHOKQCP/ErELZt3OU59NKSxdqnh/sAjziiYlaef
JmF79o4ade2xNzdFJ+dXiXLxYyvzCAk7h8b4sc/IWYdhYMR7QIyoukgtcN+MWPlHCHlNhEeUZvY9
2Y6ipNRVAbPsU7GNf2E2PQL7g4hed1PERV1icIkjVI2xEi9gZBAVponYDPIcUam9gpJnIcB1vZpK
3gz0bTSX8WCATRQc5E4m97hz7WxgJD+oZOBMp34BhhHuxDz5/U/CMIFA19sBlb6UXXvuf44S3y2s
5P/q2oc+EOgM1lTabvQhO3F9rtFjqGYBDxrD8tnpGkvntwIghtLuosS8m0KZC5tSZaL9C5KJPEHg
oyotLsl3k0A7Cp4V0kKx0K8duvsHyoFwHhilxW+WW3fDnBo8TTzXKCSFR18CmMbJG7aPksgad+py
Oj1zJRc2FnTOl3gP7JQqN2B/FOiT87AQFaGmghMJTsSujgxJ+RnIGbDLEJoAmd/y6/zzFd3wEZg1
IAFtvKifcYjgyFJ6Yd+Y0iXdhpzndF0GYdBsg8t3TP6g7PRQoc1dXA8z1jJY30wRy7TBZ/VjjXS3
gcu3pHGsWfyi+aNN4//7MRP5jfLasHfbGXoM/l1an6hV/KDfH4aX7O3OqlrVcJqFtF2tYMl5ao4A
4A+1L5o6wgZtXtbz3edYKo9fwjhVu5j8MUk+WxUdw3GL0rkDvPRte9WED4dPklU0lYlaMloSVXdN
dc2P/YTw0JPIOfwT/aRLzZ8imAaSpP6ZxdWYBqgZx/8zOm0P9yp/chBxtv8nGI3TfjE118BreueI
KUTVDw90zCm+JfunyFQU6VKTJh0Kze//JNf6Xe9ZFGYW+EVrKhzySooea/jBSEvDLSzRdgIttw1g
bU4XRhTCkM+lq8qRnRjn5+d8VC59kGYrD9d839rrveZ01vm1YIxSV6ZucwHLXA70GeSHSmi7/hDA
uh+MYb7S68MeHQ1XtelzwyfivJFK7l3tXJvYBLQsuqJM5JSDIIgN68O9hiT9OABdjLpzXeQXMvZM
RZVoRjctVFsC232DyGJUoN4aSwi0enenBwkk/CEAt7dlUnoKyZtQ705+4rGE3SsZZHLUh0mUx/eM
JDsu9aQVNmTH2FCFrpuopS+CW+Yyqnd6TNJ17p2sUgRpWgPiUZbVv2Py8/EX13SPJkb6LVHCJM4v
ZEcRHmYGgfePhvEbsFSGgHKCSLyF0rKjtgxK2VV2jZZxl4utkM0HxPM9JTKQk9z/6G4DY2TJgzQF
9zZLU3b2F4M3TW/OClj33Vel6PePPo0sY4iI7NUgQsgzrgjidJ6GVCYR3rY1Cu3SKr8kZXUe9b6y
M8qUD9iLsu8n0cOWNNo/4bG5oHIzJFmlwbTG9iK/qRgyarplCzZi8yaByCmT3PDb/JVNdbcY30yt
yWMC/QyrmplwyWzyHuC/hgfqJP54ZJKwAlBnncPo0Uor7yCoVPGolG7Rdnn4hBjd2Fe0ThxZEfii
iaIspcMoZNs30Wlr7CB0ap11+4GtlmEZN8+zbcUwY215OBKuD4Z8j/7uORYPkJMKOBxsmVn5sQ/j
l+uitm1LyUvcocgBuB5oxGCTGaFXrtlDv6f0XqBRJRUoGXX6avZ/n2qS1EihiiuFsb9Q8S2vd58V
RlVu0qz5c5plaW66NJva0KQos24ELGVgQOkID1hLy1tEqiPu1Esw0EA8AqvzQIdXUvIU0yH9DL9q
zw5j3bjWebjyA+VJ3Mx/5cPq0229nvzYSDUwcnGq2ZnrqS93Rnxm9vXHFLiUItPbJHvn12PEXq0R
TtVMYnKy0soBjIMayJsloase47/16U7uKrvGGBygzuxiIRDJNLkiW4MFilYOZ/w2MTTp+gpIW7vR
uNbRoR1Ovgmgy1SkHKBSwjm8KLyGhTbO5OvkZn2vhnSOfaMPIkmWdzBwclJP4UGGEmAzVs3oLlOg
/V9KZeJjhHVaozU0RNKYrZGBxEe1vgIcDeQ3RJvtumGf8hvyqgHlZ/fx92SpbaMCEWTUgrVrFUu9
9uoj14zjuk5vBpcHWZVas6qedOOWGUXAmD4oMPmklRRP4uJX2njikHEAamzvsgdnPKuTAWSJIPdt
d7+wjoyuALIFiRaLY07TivP5xIw37ejXil8xhC+22/xZoPos+wmqBoBLqfHnmY0IDU8kLMx+QRqU
8gYb3IUYsm4mp492lx6N9pT69BaCDwYmrOl8htd/2QOlMHjWgBY9eu7me/fYtwPf1Pmcb4zuYbfA
3pCUe52p2FuAL51V06a1ydIPNjS3Tp1TptuFAR8ABRDwCdVPf7lvjJ7oh9arETh+5MFNTWTPrNy1
f2pwYJDOl+uXofKDY0ofFlJxZnawrCiec0V6KzkMGwKg9HAohzOupYunvsWNt7Ll1tf5GmGSWkxB
6aR6jL2zPCdzW0ab+NEFaWz94AQwy+0u697oObmG7/xbqxMqC7U/vu24ip+Ikq+2VaNW/u+YV76Y
i0kg8XGSyf+2jPlrCksO/5RxsF11+HqRMroilvZAs1gzxfP4qB4R6oaF/wai2vKWnt1af09Xp/Jz
wk5VQcOl/M+lXtCxb4HLbJWKmf/y/s8La6HqxfJHN1xfNkoe/q1P5GCPQOpt62s3owolfyIxRHn0
c274rbuLXC8Fq73MiXmmAVYberZk4Q4ytnGpvdvbKtheQEGmDPT8Ac/xIj/0+zHO7I9mfZQpJphx
9iyzBIOIDXrDQ161+UoABXC36CCxEtxDS+UmFzZJcXcW0MHkAV38qCz47J6corxVjD4xSRsGHT3q
sGyVqIE6x+S75aBeYOOYrWAcllusj7YKkMxbm4GIErU6GMEVfyVTkHVIBrNSoTPHfzjd37dYaHC5
AwjQZpqrY0UQtlW7J8aTDj4UhuA6JCXkWkVSfYa+4H5YXafbsHfUy4GY0ci0iaIwgGb9CdLvnQuT
j+c6Uv4c/J8zGD80kTMsgRROSfQZ9am3PBHxSYPDySddd6LoD4OmY9P61BYQkPzA7HkjgoBjk3+0
PIuo+37htLIMt8feKOo+yg1srYfo9ELyaVhs/3nsiAsv0cUmJhCsMYAUPDtHiUTP6tRK0HO+RDZy
uJUUn3DclT7ifVf64YOsSPb5Mr/+EZMpBc1KO06mCA47OyQFCw9NRFzZKNqsREPtaNH4lNxnoKgM
agyzUVDC3PNWYjE1yYztYBDxJnHpBEM0wzmXGu90z8/0YM7A5N3hSAnV56L8NS/XemK3kKyVMwsl
KhSm4wt3PVIPVI3MgjaaLUMi/H/JVnsS+eaCNYYi6PIv4ifOFy/e5r0pLGtkpd3pjpZ+MFp+yzGE
I8yAGgXUj0wslx29//h5zz1Xgw6Xar3XjWn3USulKZoru2dCs6d0plCih1PpeIjyssSdaBlo3ffu
T+gP1AIp19IZgBlWLKydtZGRp7I6x/lLMsUCW+u4CxCByWihAqRhryh6lyLUkVZK3PqPM+Ym4V64
fkrN1uMLhPoEkay+jrCDJrbdpbJAYEtD48U/KAgVQvbEfotuJYnHgNqgw8+SnPFcH6aKUD8IEZxV
yNjFLzi4IEB5NE3zkmVILUt1rR28bd2QwamgeANuIvpOHDAlDwtx7q9aimforAfGF1xrqVTEFUFz
T9/CIJZY1TQJ/6cCGSfaLoE/xSewByFmg7gVaVlRQ+dwI9jzXQi002MkQu3u3WwSJ8PxyROhiVbg
J7ufRI54Hvoc5eXJcpsfijj6r5+neNP9+G1JVo4FTz2UgmFwOfIj9fhZo4mKZAEPMSmRiIq/CZTu
TddPy/SiYwUCTCLrMvF04UGnL0oABpB4W79kUAUSAyDOEZQokOiQsjXgCjZ5wvbihEVPsFgpz2JD
RBpbcmwUeP+Z88mEqsLwJkSUSHSjBKbLhyTkZPUnAXPx+VzCETmMIPZrhWSU6BZ0AgzHDUuy1hmE
tEiMJPPsnA1mBgJt93dUuJpo+evbOJuw8LK52i28279D/t6KI6OTBa0+iEZhtg8Ojlu/SkMDB09R
5TL4rk5Hza9XyeqvP+rSdSnD6fYGhYK1f5/3A37tWJd1/xxIaKKnB0BW0/rz/uLYjlNaK4K/pBO+
k+0TtHvvp4s1J8ObLd4D+G2plI0nyzeRv74Q9RtYPs94zrdfefhmfb47zvP2EAIU8mDhOLvgJXBW
AAeKi6cxMfcRRIJWUEBScLUvCRIpFNo1lDE4IF1fT9RSSe2xnwCBEOzWeLvqODYSc/xxrg8uaOtd
Z6VAn5GbwzhMUSPSbwvy/RKm79jDxR6QisZ95q9D/vVyS5auusV9FqJqAEgd1zHVKFKI964h6bkE
noHLh5eYnvmQJzA9Yc/iEswNOySFnmt6ZVFCWbrFN9IaweiLrQf4KXMDaMWFJ8PezZ0u8cNzkaRR
Jgz2bR78k5NOorqtCNWXbForzPAPsvY1o4G6811qUH6oYb5Z/4ssq6vmEC9G5E2mGL9y35A+Ah6z
VW+EJaHyLfGlTtQFZbm1NBavQjSuPP8rqDyVIHfPvWPyoKhVxYxUGL2QWDLDZsGB8E0TZYqlvn+2
oEJo9zsqE2mg+GRQwdYNWVUFDslf4DsdNbySOmWYej21MMVZu+XW21lveFJstpMjMhq/Qm++/7Mm
i7zht0l/F68CRuvBmQCTuLomBxeJtsSJVmAvrAYKNicT0+hkY9rQBbVcsD4xIYuESw+tDDKwh1zM
ryJ9WVZbNxMHY+A2aKufZtouQa021w4UL24EjiWP1SH+x4b3O+Uef/swXIipL1CMNl2lQU7V5ble
C0XmxD8EOykl76NNRl7/vcXP5xl3OtSx6pEQMzn/nD+ptqeiXyBhtIz27+owgWc+qg6R6ek/tiAR
8tC3TXem0x2QcaHQQ+zaumFfRtknJoIqM/1nxBRZ2rU6zG5AW2l6EM1ffNg913+rINRL6SZiFexe
8GJ8uOoMP7jaoBgQpEq1ZMBtd6xPWjYDc2ZSiOVg5E45gA7Uo3dmWOppgjpn6XZqWxtFTbEgQ/fe
/ikt6joCELjMilACjJ3N3f3GdMoKHe7DaLYa8/az5WpuqzBvJN0B5PIfgFTDcvuj6C4SOyFx1NE7
qgMevctfrLbCQ1a0MTN8ICqC5FUvE3O71Wd7fQF9G8jJ61xuy5bOFlGIl/hrOnzmxKOsxzm46Cbw
FTlETZSfoE/gEBtOWaYdOKd/09xGgXOFrCGYOwi2LE1dfwW77Lz2XtEl7MTpWdBvxyCzGMzT1GUm
XQgxdUzp5zUNFfbwzKCDYsBrgM8dyVIxDiB2EQHq9YVvgOK0OzhFhlSPq6ST551M0o1+1n0Cq9RW
SzE4O5NoYZQ19+aadL5rJfxoWxXhGbJ7uojeA+AFiZnEnwcUS10fkzK2W9mcRZQbvhHoLLORb/TK
vNiZs/49NqbyHHLp8Qnl8Uikw0utcpr/rrRFcliOuz2Ih7rYqVUKhdVpzBmvEwEG6gKIySr9aVVF
an4IIe/Y/UTpsBJMGt89IzP0IKB392Id4r6hloFOkB9ZGnedDjZ+pIRu9gPIAV2syk/howYkDxlW
Bp7CJwD9sW8G+dLnlVmSeaVqN31pKteVhueoioI7JsQoZ5KLj99QqTi3UE3QBGdVSILmZk6Q8JxO
8fVBmsbCVEamD26Ean3Kty2l1jH16ZsUtkErVkHWa7u9OR89FNlSz1EJV2Bt5QnFAHr8r626yRF7
g+EZmYSVVpjlgfgE8lahxtzIFyfLgZrhmgIwVybSqzi0UXnMirw403eOtiv5WPY5Pkprso5smS8A
NxHeiDGtICeZiLro5tdLXuBieOhPvGaFKj+3GqOR6aK9VNpR0O8TqDIR5rMfX13X8ZPDNs5Rk+C+
dCbGES5hzesTm3DGsBuTUHypsPXlHJpJDzENlDTLw35ukQzaendEFSJeUWshUyVexvRCvTgj3tB2
RHb+6iv7ynBK0vhc7G4bDLuCbr9pZmpaxJtlWXd+BtrGr0BKWQ0aYcLyDUHpusZJmTCfNUUCrLEL
SZeZXUgNJHCE54O3m8DHaGk4b2Rn/gxCcsiTmheq2r7FsHC5c0yuzLIBkB/pS63ALqRlWc+Wqf2K
2aZQbPiKVwfbN6+y+l+Uyf5N3Ig61/d0ULtXFQASNCbo+5gLsgJfO/dr1vYnNpuvr+mKuXM/dhIc
ZHqZAFwieXi5gRdbv24TgqBBWHFQJWT0W5uhessQSTyNeRv5i7LVUzlK9X6HUKtMAFuRbrZ6FITc
hvyWXzVb0PrhisZZWsbOMcbllU8xXbPhZv2bnufQj/8KVVYqSvNHSuaTBXSsbA+kg9oB1wIxsVwj
xAjfLawHMhya2oQabqRKCb5E76l92LQWKtRpLQgzVVVACMKFxwiGeCRq+Dw/luns4ZG7XHEDDXnb
kjHXRhRP797fnYeIKAqGlwFkhrU+FKu5zZqli0lVP86Z3i46/QLG2hwpe5lxLv/tW2AMEAUAon5i
dhVRmuPRMPEiFdUiULQGFNG/yfP3lPEaUymtHG236nrrWz8ctXj/TCKnlbLZQDyt8M3hUHIPvIhl
nZXDmnqDAt095BxRxoEYeu2Y0U6IN4ZtFbI2BMcxppb59dgTZh/tvQKO54COG88QNZRx6+8jIV2j
yQ7dEMlr0of5YG3ZMzPBXlga+AM+o4osTs7elW1UlA+QSLL1os0Q+kULCFG8wtA3cuW0Scc6UN8Q
pJLb4hvgaQMCHCXxkrcd9CAflVCpAT7GlyHhLLl52heFa1uEAbO8m8vhCXMlKMXA0Y0eZpuNfBnU
0zYjr0/KOGpeQqGzP7G48TzbBuYENaPaATTlqnaH0/9aXoLv6jih++oQP7LATJev2KJ7amx/7pKe
gPsq9uZyOv7AJEA4AM1T8SvBuDxKRelUyccHTZ3BGayVcJoHyMphFBjsAvfa+ivn6H9MNS6f11KM
1n0NY4/86Zm++Jek+HTbBPCb4I/pMzX6u8S67ctvRs40X6Jd8NIU0BJ4JRgpFLNmVG4j9kvV6F7p
w4PftxgIkJ0H8fvrZO5uJnIXiXLgj4znvSf0BVp/4OxwUdoXMeC8QEQEjJmXuXdGQCCVtVfsERoz
SbnrRldU83/dHjajdZ7EyDThz9HiWD9K4DdgIaXANfmlA203r2dHQmCiVywz2puDSvXQmnH1/LIc
H1/O9N2yOCcmSM6ql63to1a8QNXZ5nUPM8ffe+bVo0L6YuAxvbFqM+6l2iXoK6bC7WSTPrL7T91M
hF9+rtysJGRWdJoJZNgqrb3ChiebTmoAOFYriSimPiLTtIxYRWoeKkVOH54mk2pGPoJAm5G9R8wk
mhwgbjIw357ypA0YDPMXy9024J6ecgmY1qGYpmpnoxBGb/tUhdUsiPyIen6wrdr7acUD8Ic4QRQy
cKkSyIX87+nvEvxlMi1S2AocJuMyH7OTJojoTVSp5JR9VzJk9PvJxhXluKjgtkUfncT46QGslNfD
DqqnRn936QY9KFydvHpgjrldqYL9CN9gxkiCY7Tm0Dcp0dbodn71/sTT+XIDfhPLOFegDITnHUVn
JhTqK87pykj7WwYP1p4aaZkquMdWC701RNexJJmpQO8FuEfd1fCIERz399SdfVAAjQPl5o22tj0a
N7POcQveCnliDYPcwfeKWJycOimfML9GNsyrs5in7NZDJbiKllMal6i487dkGbgARLu3uFQG6cDJ
ecFzAcbgh08gy21YOt+XGez9+Fl4qns4cll+yCl0QzcgW0zQe2e4X2PGCxsmir67RS+k0JDNd7JP
a45v5ZYUZ27koCu6O2tHxzgbLHFCEt2YN+TmPnxd5qX0gdyMIKgRh2zlXRLG/r1eLJ814z+abhvU
xZ5EkUYvLqzZM2zZpqueHulDbeHxYKTQDqCwveU1H0Lu5JTH16N1GQLs+3YRDXIZbnSx7+fiJQTL
U0EOPmahl3XcjSvM9vDW760MMUOfjGKFYVKu7v0/fcLCNdUbloqztRC/pgs5OJleMsr8YF4MoLYV
CktbK2V48q0nnZRCRr2RIAmfrp52tI5vGS4zTFZ0mRZ8YphV45sWA5LScBsX87nqkll0QOUdx2ef
Lw4AszgqqCl0p+L1u8DBi3WHKNwOGCXQhhqSzn91MoqBXo2j7PUZ4VQs4UfBSzaWxPXVBRBTCfCj
eJIdi29WIsU9iM0V9t2PtF41RkeJQYzyGqEqtO13JMJYsIHJOYdOmF1z/5SaFAQnutgJSzSXD8F2
03JWyCKy2XEgHsfAbJgMcuuY9bQ6AdPB5BA1zYvEkw5wGYmfyL8t17Dc7WGG+3Ianh3kMb992mqD
FKf8HPn0JC3/pg15sTs7Pi26ga+3ALxSm0MjDRA8aBn/HAOUw41BPsfGmXZnEVEthPYS/WMXif3y
8YMXj5yvZAq0YqoJySYFZsybvc6tK/z4bALYe5qS5LXx6deWzKDTeouOdKUvvNh7b1O5b9PYJqbx
Kx2RD07GPY4w+PpdMUYjBjRgAfcHqRyL9tNZeL+Mb03japDOeUIrrmPYljbhLyNwR+JgW+PH0JOC
Nfjj5xdrvBJpj+nofgJWJCcPdW3ZnKgtTaMcyUeIsUv7wFcQQFP5blB3Zn4oazVa+DU8IZZx1YxB
KlA08L/iBbKcd6F4+e5wSzPeVV3zCshekvsEqZh/mLMpDyLBBEuV0inAj/QzQH2B0/0AfeelL25D
vbwwfxQhZIq08IHolWov4qEFAQnUhuJLAA+3otLaeyfzADRldjWQ5WlgmIPHB6OhFzSRRVroollO
NldOeQ+RMuo5H1tJvPVHFPlfyKIS7t5qgQZZ3f9EctmHuaDOib12ezJWTD9WxngFykOEXlnOELtL
fjB4LpHmOI8vtwa8zweAVxihdc4+6G56rgFWC0H9E78uJF4Gm7hx2nWlYU4dk9lQ/RvJc+nO+xZ+
2/dhx5ORy592GL7E2OmuiCKKxFEhMnkqMY0ba/SULE0863ZxvgQZnGWF1Syo7ztDaWUYIRnuk4KI
H1JjrCVbA8O9o/W/h/kF/26VVO8MopFZJGKZjbzfgNWrJ9oTy40UIYwNWANk8rCL51+SJF9oepba
kuigpye36knW2HH+9L0FoKxqYeqWaK2DVyhLd7Qt4OSAMMb9LDAqh5mDDwg3qxcNd5nhWMNDO3Ng
HDZ8BkFxdkRU4Yfrp6PgogObB1iNOYrLaD+bQr4VCAGHzEoNPu/hhgm84ID9H/tlv/dNVTDQyZS/
RNeaVKEckkzUGpBtutcm+CZ/m3LZXo3Jd8q0bBTTT1bi9JARc1iU+QVOYCEnB10ET0M3qmdttfx5
NKzLiVNFudrIQrq43XQkY8SSAxsKKhNDrPWogjC9rkLK7nIXsArEBwqdz2suvaLfJWM96amZC1B+
Im38hvoLqrogJxEDl8+8u4Z4cssH6NYCcSz/nIDHixeK2R2L9sjUmpGWhkMjgJi8Y3Zq+gLphJ1k
hq2HU6I4mkSJs7wg8fyI8Rzr0ARJkSy5KUa2ZsFie8gBiDPrlYQyXbR4Xwzl91Iidiz2ncjqw7Jt
gneo3AIX9BCM95UdkuywUHCgRPD8YX6XMI1LaucSFyYOTZtcFz49+zck7gvEf4kNnzO1hlw+eELC
SxHHonDdXtOdp8y2tAppD32I6DHz9NLqs/WtqGI0kEMr/81E9qEx1EIi7JaHuS/+6yzGGs8P4jCv
lrWZdkvMUYZ8dbvtR+ATaQMgmGkaQ3e45RMt8hv4RYGZwjintxY4DP7VXnqFok111wYGu7fQR+Z1
XwCMXReet0mAQ/X23+UFdr7Yh2+mWRxcSFcCvuKXNfs9QJOZEUAZfBrkITiOUwU1+HMaQZj9sf1u
udB/t9OFelDKTv5NLqUNrAFYMkLgFqs6zFR3igl5mDB3OpNM2X+RFJ/4CVlAFS2ftcuNcbyV+VbT
mo0x1aMoQL4AMcAhzeqIAkDDIlA9l/Pvr9u0dx+D8DbLqspFiAcWYvEexjd4lZ2Ln0fudhzc+Ruw
DUEo9EB5fykNTBvpLS0OOzcIf1igsjKqgeEWazXV0XqwMPD/+GfzdHIpH2W07XdFsJ5WzNTtmUll
3OfvzPsGOQm/i5YHxAxPiF5Q6xvx4b6QadM3ZwoYhEER6DPzcBumBc4Ux14WmmuCvLPLZOVOkDdH
mMberOqlJaVFjrcSv5i/GG1PfTgvI6hJB+3AtBozLDW+ItlDhrnWxSP6LJ5F3/AeJ8kwoRJ+iCL/
c0dxg9S5QzKn2u7bMD4m/FMIUCD3P0aziaIDo0AcrBoSTgD6//GmfdogZ8Q46PukG6t5sWlclGod
ToXpTcw4hPUKJsbPudNBVZk6iCWOOiX63w5pxZ6fjyNnI24El7jJhs4YaYAC2Vy0FFUoPi1T8/5P
ml5Wb/nHjpEVIj5sjRZy+NS7ib8SB7B2z0ZXeWdZ6wNd5kX1CZNheJPAdZVe7DjbbxuZK/2m+/28
39pudQv9r79UnS0pEgYd44zrWlAYrGr5sCq6n6OFrGDxZOwC5vYtYnzXh527Vo3+rPxmqigLuJow
ybvIUyp5yzTLXY1ftczPbWZGW5YDuhRLCCdWszJR+SlfcjrCBG61U8FFkeEMFrIbKDGGW8Sd1g2Y
f0KD7+QefVMoagKPjbHjsg==
`protect end_protected
