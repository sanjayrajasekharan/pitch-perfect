-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JOroSILy5Pr8iNsv49BMzCtQUIJe/k0AZxl4lXLeG5HkmIOvyvmJoNdJOfRASPqo5HA6GfccXOOM
qCGC47XNtYZ6+zn2x421kOAzI6gCz6gOVXWpYhmcn+IZxImnQC5VmbwIo0lsTDqgJFwei3HqF91C
FqgrYnQ+lmk5w3asqj4D47hJc8DocNvSVv184r33qpJCPi+KhYwYuUyNvsUsl5hPI1E0sfvhd8NP
hnMPUqjhQOMnqnGVD4HiCQ/bRCe+rStxUPvJckNzy6o72YHOZV5Z6tg8jh7GKc/XnOyhJvmBd7aW
heaF6yihTCdV1esngWo6xpDsNQNOp+W7hsztZQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13056)
`protect data_block
C0/52SLya+YhJyIBlS0TE8FpZe7XW75GL5mx4rwDYEETcoAOR5B0ryTdWNSwu952r+tj9q4T6gu9
mbXLqXERk+jmDXqDUXSoYMSTstQwxzs7alSCXEuXvY7LCOZrClUnBHJRx+LZXfRpsrK9FgRxRD+5
nkq+c2RqkJiEbMr88m8U+OaBTL07ES/VqJaHrMBoJIwSNTMgtnfMJd8eudz+gYHQgsiMdAme7OiK
b7WIJrmXooh0EsKdIK4jTY/+AS3WctyQbygrp+HLjgrTaD2V6vJcyK/BdWlj0BbGh7kIjU4V9hSv
9rwRht1ZTodP6UepWAlgivxXW1Qletmt5YYXJ4guRDGVpVU/qWVGPC6JPT+wHLeylW0fL3dQNofV
ozKUPx4pnqr9gbrazGmOALMJhPyEgXc/cGdqxgoFW5BbaD1qiYddMQwPo9f4hgzssaEmUIByZQS6
vRGBu8RdwU+GtmEKeqndVpN3NzNvVUm7MhXqZ7GOXNxkjh+lBgrgLEqH3ibwVi7t1ihf/UYpopUX
FQW3/n5GFVfdsHVkcPPilSrYFoM8NQcuydjovCQdvd2RJSx5jp/5FNFkAnQbZGFj/YFUHA0hyK/b
STs5PXzczFMO7gggbZuGMSPyWrqdLEZt5Bl2w7XPOY7g35lWpYive+G6czxlDn9o+n4HMeghnP+f
bJgEHwT8rwdEwtKJvdzmlFRBZMP2wmUiH+YvJn8pDj6enOFWRsR/gPtPpVrY3xNy3S6salGhTT71
6Fi0I/BTQIkm8BzZpxf8ZogTqaKxTPZf4j154ZcEEucoLTaMfSu/fikX16pcorikHdA7gG7oLIqL
UB+Hez9drVhtfQ6q11LO4cKrCKJDVBEvEulwWzUbElls06aORDlcIh8XneiEc+eP6tT1w9yjr2dG
qVmQ3gV+SiBC1lKq5Sk98De7goXpjLL74e47SpSl+rFh7RLlU1YghNeqgnlAGmnodeCa8xLRoeiq
i88bMTPb8jISMeTL1dS7B7ZvGpnkz1eX0anvfW2l+c1JmK0XlhGm+h3vcove9LcSxwAcEPAVsamI
0fZfS/1EYKh26eOUA6L/W/eMWwZmCx6LOOMXo3F/JaSNihhssb+57JCIdyWSJP5yEG9EZI30SyY7
DgXLTEsv8wh8nFB1kw97kL71qr/otlLuUHLkQ+VRuVY+O6bmRfnzPogHUjpx4HeEYtdw5yArPZCK
0jRzj/c3Q4qe/pVCfrMjNqXnf4btDGHv9wt+fFNVw5vTcCWMdTV3EotfDQrYkA7dtwUbwt2nld+E
48f6Qg3rOtTPyBx7VL74Y4w95YLuc9ZK/mHxYWjrZ5IR9HCxSKv6q7qTeTTzgXLSqMYXLPZMn9Gg
kzmwMBniKe/+heeEaOjPi5t6qpVcqEb1JbzFjMngyPkwizQbOKD1LPyHpmymgJRtC9sDbbOagDuB
Dmam3E90l6PpYTisWsRHyKjQlyrq5FawfGSerpuk1MGCI0JiOheytNpwNNsxNZSt4mqEPl0XeNPO
/WkCbTe9CzgIFyIU1qOFGVjbquh0pwZsfervWZ/Edr+r5PI6YpaHiPJNhIJcwnj2cgLRWITh7bjS
OUnOBJY3yfNCeeupmnRQ95aLcvXLFOhlHqyqoj436eG4X19SJ1wvjLPdoBfC30DfmiyEjY/tnNHa
0NuSkkrVWMJzTlV7ziCcqm5+SacR0QxBZNwct+sZwzxeHoGO4fOL6NOsJN/nam7QRPCHkIN1dnJd
Xj1eSWvnvBzqUGRj+VjkscPROAZziYm+ocjWA4eMQwjyne6/0J2OQZDjm8Ekl/o5Ij2NHu+NF0jL
FfsWEtNwS4PGDFgvB1R/Qcurh7TKGnNNXjbw+2masdaVk8H2WdicZIgFiknON0rSZrrGitmxjHaj
SLHR62pHBh/+tQmvo7nn80g+Ro6L0BpZc0bbMIbFH3JA7ECxieTPjx/wQgPTygxTyGCdzTNXx8yJ
JlvNIThNIi2r+RJnB6/yK7x4UzqNXF+eJPsJBsubzxBxkykPccBneoRy6g5ITK+TvGglQhYFQ+yS
FEtMAqe0iCQWplS5bpQvBc1uNAEKzr1ebQmPVNtu9uHWHtrmSekERba/d50ISMrNktISHk4o1Kmj
LqxxEzRjMH1w4uEf91hlVUyM7hl0m+Ae2aIhqRae4Q2c5TWQRB6PwJWDZkcCiD5AWjs2zxTlvGSL
HzOzAanrB8GdMf5m7Cp1pWdCW3uA6DZq7cxQ8RVNQeNhTmVi24rb5GUGgcpebcKU7nVn6ruEfrVN
dlc9J8zsjFIRKIX6wVS1vg2KCBzgK8fk8KdbqTyS3S+4XwD+21rlLeS20OAmyiPFkBiwhwIfctMd
gmXsmWgxTKVLqgv1Q3qi50KBFy8xzc0zrDZok09eLSnIPFwYs7qw4F8g5jzCGD/xDQDe1lQMVGZl
hp5MtsC+E9ZfCeZY8YQR3Kk7w63UNFeffEAtYm8d6jjDKZBiyX8BzlmbYa0aGkNE6EwK6mJVMhf0
hbA4jr0EoBaNkqyiRcY76nafVTbt5jeHMquNrCZKkgPhkiQ856ADqDr6sF5q5jsBU1BCVDZejdV5
Br2rCMUgeTiM5heXo/KrVE2n3Ky7aZS9tVgO36nZBujNc9GQK3nLEplK8XmT18WX/p2o7eQv1n07
eh7vCGuzXfsANsppZv3xt5MPQTitOlLmpAJy2mdf7t+1khdMjAbN1S/8zKTrnxi+x/nrOFvJKTMK
jW30dcaMBLSxT1STHubUoFdWFaeMTmfmETKh2I7KbKwIJird1OFqxuQJprjujBJR6Dk6nuHnPwad
JaOaIzedQ9ITBXFDQiHuPTjq7Kg8el13A1YWK1pgeq65Y/Vev3qBcvbSOj0NUJyMtTuboIWNB+e6
QVvmtLtIrgt+YyIdyOTPJkI1wEQdP+nRf6T5l3Lj9IEZbgJMFgbr6wj0nRYs19I/7ECE8VMv/G5J
Y4rpy11GA+ZE/QF5q7yFqTa744psKCZmlZ0E71Sd31MesdfZUh+Tp6CbJQQSYXtibIIglrXX53Ek
+kAXYzk9iV2TKhXJbO2hRXjFS3SYpfEOKaEL3RhjcV5stKvuvE1LOCdm5NIxXVppd8xT/jNQKIPM
Qu1/JHEufPW1J1X7IqhQ2ewwvwOlzeHXKuN/wSUEns2G1Ric7S2Q1fDMrr7FoXtY8e/rEm+huoEC
cSP8EtSsILU9JRdq91rLB+fKoX0/32bC6hBumEuON0NA/uuoQyis8WRpadkxN3V2rGjEiGJ2/8Y1
osyvHp7In1wZw8pbdcbcZd3hYXUXiCJsPY+0x6ajEFLUZsYnsmKyjbeoHNc20YnllWicAEmppCfh
aM4m+27WKMeg+PiMyXCx56Okta5V4XTG2gZYy2gmv9J8MHA00tRxCkSPoHIC4HciEraAEyDeAAAj
ist9z25bp8KGxR/ZMLxgSPP/RxZGjAu9eBly0C4s9+Rbpne/6TxEIZObGKAXmdzcn808jW86EP1n
SvTi1Tg8IixVFal0KiE2vBgxJhk9qL4dkQajk0IcQWzzIgTCoAgZf+XGNQKv+zEnqOenH0L6KlbC
bZKbvC7mNmeKdnW2EgKPo3iHDGwoysd2ML6EMfx2CcsWzKlKxcd3WREWkTsuBgZ81q+9T5TM9NFE
8mf70uphSxjMTSfMO9Np4vMC1JX5ljcOMZsTNzBhvH2FBX1EjO4SFPB7dXqhkEun3Qjpt5bYeP2Q
I5YK7VWQbRcV+jjAtf/0IKNX/c+Apl6cKTqp/ANTx0mcw/tF3CqScJb1nvQw+xiz2+qd5La5WjG0
A+7SJvrJABF3/3R8/qIMo+Wo75A7agEo8zHTG7sR6G/Me7Vbj6F/XvZUpUvxYepuJb/danZIzIbn
H+4mB33sDvkGlSN6hD+ufJaCD7cYDa2zUR9RBuZFe7pwbtO6nyvH7UBYg2ESobxbmN0ntykTRDPk
Mj+UtiWqqVFc9LIIGHtpKx5M8JUWe1+IBZbsyW95GDaBKQY9AoOmyGWd14LO152DFVo98UHQcvBO
F/3RcIrjRjH4h+qf4ZiT4/0Y5ibZp7GEiL2YG1C+aPpDXXOE1CvBQ12tRdGQYL9lewO/NVN1eHVF
3xGYB7p4m0sXp737ZanbiE/Xbr70uCp5JX6EG0Mxf07gcpaKBrj6SJ0g7n30IWQiuc/bNS4fztq6
I/8JZrX8BEAsS0HOpfp5UP5rMEyqJTfNz2aZF+FTEw1mRc3w+mRTtMVNha6IRQgknftJwn7sl9w2
IL96wJ2jswRwsFnolFy8AJ+c0ZCM2ME6hlGb5lSgrlX/lnxMU0PggwZfWGVq5hLqysDIIq0IxNjl
XeFGrLXNMIWCtpDvMNT09E4NgtrlPj04xLXTMeBSmUFmnkPKv7KoecYp6W3o2Mh71mk522PhKN1t
ff7yOcz6N5kYTeBDtX5DpwpWeuAEn8/2pD9g34EHPNKeGsoA/a0I8ulJzFCMwuEZtnnlRu38xICr
hIE22kAQMKlsvP/+4tNz6LiO8SJ7ACV2wRLddND3ozfKZspaIenC3VUVFcPRRmAimpk3wMlQ/LUg
syd0hKisyzKtbUgXSBSojo0e9rRRpSO7TPcgpIs7EHOoMFVV1J8AHr66LrOifvwERlwglT0VagNk
NvWeQd+kC7RT0Zb+WfVQkSI6kOjdnO3tK+jacvQooTOKOUJ/wDAvWF38Uun19wQB1hfAMTUg5Qrn
WavAEkJCwMO0d/MizN+93MnTM4bbr35Y9rZi2DUJ4cowOBwZ0Vm164hIqlc3AmLTqKcOo5QHQ/S5
rl95aoZDbodSVdeesjxG/y5k08ITHajV2Z8RPiY9JHEYGxSdCv5o7zNIljeggKo6FeBtJL6aS9lp
hbd6wAhnkHeFAz2deA96dFdoeaIRqKpZGV4VsS0i/M0szkomVtgpC6xn0n09qZvQ/h62B42N780e
/5tK11yCsQ0Y6aw6dCRBLul1lIwbR5gErty/3ErGQ2cUENV8GXZ3k5pOVJKSKKeUxqpp2Wy3/M0B
ZHbMX2fHDNWkrGevKocU7ognBXQo1qgA5QE6oWChAP/VmHzK/Z58USaxkZa4fP/V+svhd8WqmN9N
ArXSm3xFTJww+YrOPowbjepYT7jQjV5pfyU+Bpr2s97FSf8GFM+bsJTo49PoHy1GflpUx3J65rcO
YOkZ+fcX8Y23E7R3R+dUTP19gZyJh1KzLA5fopKSAfhGI8P9CpKAhD/3MuwOrBc8it8acUGnhkJw
nA5mD4MJuUepPkbsbfKdPcdyCzQxZtRowcapOvzTL7Q2IogLLdoMwb8ETMfRx+eQ97ReZESkDGx2
CjqNZnyJmC8y3rHRb+px0oWGE3tk0+Ks3LyOV2SOVtBOZifSLCcl+TOV9JJdbiBI0A/e0AhcK8nO
qMnxamfAk0i3WGk+IBwplEdv/KlruUECMV3Tl3RWURqaJGgwKIlm/cibyIokxYHTCvAxEHKnu29b
gs5kXI6oq/aFk6x26ljz+W4h/QVHs4gU11TD6pvAFkezeSYkx+2IvoqK6AxMRcZNQYOcoAuQISpk
NKGHzrOc24MZFFeM/FAstHEzvANQhNKvWIY+0eTD2FZBjgcJfQ3IiDyQ+xFInjBswFg3Mn+VE36W
oFj6VQELLCZPFXPwasdgInWXLjCEXpEH0ddZsdDDse/9SfKuY1l/U96hvJABnxJq5PqfffKWUKeG
4JFISEx6fWV1J6i70Xfre1psku2hQiYbWdklyk/f2bJG4CN+ufP4YjR9kZYqQiXsC3fdxPS+bsEg
BTfTh2aneYj16j59IF6QrUb1ytGcLXVIzC8nAAZN/kwr1OJ4HvQVYeVhdLwAd1TXY8Qirko4NoDK
kD1VhqNdBGWJYJa4Ix4LCBPFqpJmyrF0Hedw7Wwg3PmfjGvGz93rLgBLsKeIpMI5qz1eDjIEWrfU
s8drq5yFubBJr+Blk/ZbSDol1poQQYdSjHecrC08TM/iYdJl+wwo0r/QbyP/GViU3xm0i5y4Q81V
h37QlRDRWmV4XoTJ0eRY84w8oKDlqTHZ9rSXwT9Lnp/dDYL4I++jpW05GdDMjjqvFJee4x9hlRwy
+vSR2iSI2M7IYgkdxqWYhKaOXWpN4LuldaF2rv2zjHkTRFG0X5RSZ+UWbj6B7xyf/jpnCbhq7Zwg
G3ySidQFExYw29eAn9fnUMT6RPVqxSSabX7ZWY24YENBjUVLg3YwAxg3fKzZgKBjH59fEEIccGNR
MOR5XXuIYySM1RprXMLwgoYSeiuUNeLf0mmvgjiKAOXYKWRvE64KHyneok97bN53EaTjERRa4x3K
0f6qGuVpWaXa0ZYMx9Pua0k9ULZy1ht2nCgIWeRGWWSilHjlUy/NHbxxCMBaqcdd+KFrYZlUCRIA
EhKisIkV9YpV7FPGkU1b4NdtJdY2RB9yy8v5X0Jh/TbP5hU0cLiR7jNbJM5byPzGZcVx51nOxh3Z
cYqnOT2MGb5bWo0I3dD4/mb3fA/uIuw0jio2tYgW0yfxhctGdSYLyUdHq+kWEZ43ZsNExYMPPjhk
W1r0yf+ETpIB/suduUspc1TAmMkRios1u1IWElWyZqasvl3tZswpEccfhnXAkHM7/n7ScbSccrBP
PLLrZnl9HBMDEnBdFCDqd4TTsSOxsNrjmxyDMQtT8s7E8vEelb6OpRbB4yw7ogaFoGSqcClBVFFe
BRRMQ7XCqtBonCRa64GsDGiSuvLkR3AfgrqJbP6QYZM1L2/WRn+bMsUr+tCBSZCV1jr3+bkUperJ
9Sh1xbY6xce6Fhf/9Njc1Xoh2+Z1/FyTtqurSAwzTOfJPrzDnikTkI+/tIEEqXSnTJVYVA2dQnj/
IObB4gUuli+oDgJ5jHEoR33Z1On/8XMtab4dsVqqst6VkdtdCnOtPYq2kyifEh2v7L+3myOxS8oM
m0e9iP4DBhNnpThvxdwcAoz5V+RRtC3jUVRwj4+09EfPMu9qB7/B4k4GG6eo7oOtTRn0iZg/Swrb
PVr4Zzm/AKqPN4OUtq7gTwgh8smUr6aCfQFr6vDjfU5V7uoKfTfYBdY9i0zl9iwMYVzvYMEpfzVm
rTmGXePJQ2Iq1kB4ZJ/4e9W15d3jmptr5LIVRC6gZLVslUd9JLVFbjNIMmEw4/p0vkYCcxygXCFU
5HGamJDKSmLS3O72E6DaUv/3i6Jxj6GcCxf4jd4d3IGyhuaYle2bgiBfEB3UdvIZxbePGK0UN3lm
GbnZr6+vnSS0Yu57zDCqeUOh813Do6ZFQPvT7Bnif+6NIyPwzjySUnrmAIawzeyjtWo7wQ2oKS5O
xnsPHG7aNlTkm1hhbvs/iAVtaPLbBAxxpWElsBQcJKo+BVSI7gPn3YlhGIia5UZFxhC9D5olkZRF
YsNLWqwL2IFcWcGipvYtdG3ulKDelzsTnqfMyzm2wMWjxind6PBqtJ788a4KCJwy50PO7gNindw0
4VvwqgWVlsKrgnugz6ltsMFlyWN+xy9Rfz5dy8fcmmLhv4kdlGwyzs4WIAwZw6439X5lZ4ZSOYI3
OONlMMaR3uhVHFOWtTJT2LDy9cboN/ZqSh8YvGQZQxSjnsctqMkBbseb3nrg2qjlFuTZKS9ZffH2
6y2p2adt/vtaliwYXJPKAWslZhu4zx7SJt+PL7bfz68YCWfYpOxeGNop/MVzCqfLumigNcns11mU
VND29cG6L6DDFrGwo2FnCrp5Cs11ZlZWZkKm+633J2u0MD6IucXz41yO8TmAK64x95NlUBc6soAV
tC9G+Nvs5rwG1VVfexroSUIQAI7gF+okOw2K/WG7+9c8NygSc+IMs11ZKD3Lh0WVITVDcDBd0Zdo
jOtIQoGHxQmo5KRRIHj48c6xFoVALx9Ln5/isiDHPSpR2aflFcqmHWQIePorVQyF2SorkN8U5pSj
R8muSWElO7wi5p0phVaS56Q/N5ztY+7Vk5k37vVxBIFSA6EYwwz/5VPTHoqtPf2L/cJc+Hh5r2UJ
eemNRNJ50GyfBpEKdJknzMbbGhEU+IWO3KIeupCrnGInA0pg7SluslHgoDBjJvVuc/4dGC406Ii9
/M/7HbNNcHLohjmW12pRBcYP5N63SxXPOW8c/2QSfZJl2S8dHfvzWN8wqSKASJ7z7xI8DaLFrrD2
EZbgn9Iv7WqfUuC32pyemT+Ss6KVhGlsS1XQAzbaojgaReIBB7ExqRy41pp+4ftflM2CIECpd8e6
XkVuwclfqX4ke5gVi1Xr9AY4sIlF7UOhPZ20fG+gsAI0eMGGVl9amenqrGBzlw7MPie3TJTM394T
j7JczxO6+hibuo7egWH51GqXaImNK+tQNWh4vOmnH1xyDGPRoB7be/4z7IcGNo4T5+C1gpkq5avI
50MKhP7zbup0lzju5TUfrmjzCet8UAHxcYG7E1rXTc1rq2q5qGNssCIp3nkenT9umjWOl2dEyn6X
HdTBYdKRqSGtmTgm0fEfeERWw2tpCW0oIYTRYU6Zhy0sg71hDoXsadgnppxNOdeNe6NCsxLvs5EQ
VlxlAYSvFAoYkmpphP+gydXEJ9mB/+j3bIxEeecimB4ZBItnvt1WmU2e1NQ4mFFsJnIHF/DatpBf
/yZYmfRyKtzG5R3JxZ339YVvjY/6Z7pKk49yyVzdhR28JrZFwB96Y4WENDjxOYymMWaFieHENkhG
qHnz40VtwzzkQfiB9LYe9gKJmOPX80URwVpqGgt/5Qci4uvgaox1z8An7X93UYH1InbVkidt37ve
wMJrB0I59fNeBAe0SnW5GK2H2gD+Z6QDvWkGbz4EetYd43aYQ555imopZkezlk+Bq5e9XjoLeL7H
PstSsTm1+a/XqY1OvBBX7QWws/hlE8wN+iWLje2ry2/dbiGUVxMjKkEnTsJytYoVoXAala7t151N
+YjS3DW/ogLj0rdN92sVju2i/bKyZ9Ie5lC7/hlKcFQxb7ZqsdJXNsuefuv5NAnT64TBOWw5fmRn
X9zGkKNSWkM2NPK9LxAjN4PNY3ydLAp1xj8JzEvZHF8sg6Id3Wl2tAmQWoadCHBGjAcKdea5ZALY
02XagvAtt7xtD7zxDJYqDeOz2qKiF8MlZUEp8pu/ypY4IVhee+hnCcZCpkr4lNNV2YdnGyQml3XS
wdqAqE6rL8CxBbGreD67w4x7FrR2f9ejqzS18XEo92LGKTISWnDLe2hRUOnbTwS12bP71ZQLViLE
rtWWOZ3z8xueNV5JHPl1iTeBW2ylKHntCccQ2blXC8NNkK4qyZ4YhHxuFX+BI4VgIWVKOGxQ/84K
hP77BwLR7hY35qz80DM7vZxTNmeqlCMpw8Mc1yNdGul2t9ig2mPxrKxhu2YhRVPAkPPl+XORuD0y
FxjRxoW+oSs70Exa20LuUjfkhicr3HtBgOaE32QnjvzvpyGwzYiUO48YZkLFfc2ZOk+QHwJnK6dm
Y0wHmJ/RMxL+Wg1PdnfoTA/i9vSr8Fjf7MS6Een93kuiMfAvmRfM6osTtASSC9K3N+94Ek2UQfb5
H/PmhVde9Hmr10qWrO6Lxfd85WE+06dZNmRjV3yZcSvVMOwl5VSH548TaSBnyDf37/F8PCwbqDKE
x8BtYnLNSh0N7fuWDtMyMwSjgmZpLbJ+7o6lZ7XmraN0/RcJR1GV9QJgthbteC5xRtyi3TElbBZ6
1A74UeA9glRaS1WjirRRBflILi7x3ZLCgky1tRn3x5LU5NhUFsa2DpXdLqCBJQ6PuH4gm5uTlGql
dGvjGweqXmgFriw6fdQIXB38RzYEKuIuuAZXEvxZVIc9DMhfrbfg3EJTLR40U/4V4rGRyfVBHUTT
7X4YEDY6+1BWYD43uhFrdWpbHtb518DUxnUBk/2jrU7VpZeO8+UU2hCBf+DUJ0W9AqvtFMPQ8YFK
7mvhj8I4LNmJ29xBn6l/qi17h5ALnzTzQpbDpY+wyWOkX3nrJ+SMT8IMwMFHc7p2SUjL2BtCm0g3
kdJluZ6N4nTD2YpyvhyI4qaD+LLYKhz3OZl0qU4sMUBs85FQCxfrGMOCzRXgV0/5sAmKaoTZRmVy
iMuQgze8NM/sjIC6JWX+yQaMH0SRJvnCncuw8TR3S7S218SgvYT7gZ5oBkbxWri38+xFPNpCDVXb
wYGHxHrCA/mA4QjkFeXYujqrioP/ZYtpzzoa4wPeIe1crF8fjUzAv1k5WIpoCyAgmJ0waAp1JMMU
6dlSA2+TwSb1uOlvS8+MPOPJmL0gD20Iuho/5iQxCw4pE//hXPTKDi5HIApBGasWWp0RQEqC43rM
xKQr6qC6ndYMe9gbF/2d4/Yl378OmARNiKjR2SIL2ehE/zrF8XNvd1XimUA6bG+Pb+dY8Ss0/x3R
m74cso2rI/QQAsAjws1QxpwNuIWVL1HQ1nYo0EkpSZM/mj/Xjsz5yoSj/BzCzSzta1W2X1Pc/DHv
uzLXjqNggHic33nFOTzOmyzjEQnw1dP4LX0au2TXZDe+6JJPWHK6m4jlYXb46XFsXs9X/DC1JsX/
nomgG9MwI5xZnncf4VCk1jDBNnqJkXSeKMCZ4ULJrkGa+l0eazGrERxxrFXcPGtVBDYmNIYrpiP3
cl+uDR78nZwjH//MzqTdX0Wy7mXVkCOKUN0MbqiovzsZZTKL2EPMlXQtdSOFrolQ3PrH/ZGHGzim
q7ujTfu/4Y/kbAwhB7aM508rTNUKyMIN589dN/CRGtSZzlCSIivfG7fQBQJQx+BFCbiPOuG00O3B
SoyDhzO21z2gOrFxV6BxmbX7VH52txFDnnn0mjfFu/rMWoWO4PFHfLjH20r/GGGBWBznNbfhZ2Z2
OQfQmHEwGM5We8Td2EJ0uIKD4t3BGDCK+1GKCeYwm2q4RieQQ7+eUgDUMqIKhkOQSj/Z/1QATeBv
IdCpu1KsmU9vzTQKq/C8IaV+/Ah7Ghc6vMvpMilduTUyLfDlq/Fn20lHRt592XPgOMaK5R5wxoAH
h8xYYE9tBgrt7WsMe3SPKro4M54nVhlWxWrfIYViNT6Dq0GwiQMsz+C+DJAKONRYFm1xOi1RpMRA
p+Ir4zQ90e8dgxe/em0XFoysvLS0pMbsbds8b7MpqGBCwVUyxQQj3xJ4KohNbY0/HlIEyikbDS6W
NZD0+L7C+146IFHPi/w0rtOtKiEy1ZpAyIiVnXLaOanvvuCjCx9GvlnES1PzV5qDxJWsoOsEPxO+
owKC9mLJHQL3wdaYrmatoD4V0JAFIkRbDtvri3KGKT+fMYoOaLJ8lQm3XgbS5ZLMsOMfP23rFNVD
UZsdtXSlBVbHdvpq9HNqyLoVcIW90chiIVmsDRuLHyElO+FYbcc5OaDXzGf8cCeDnbjwqXutm7Zd
78c7EZEnq7SWPk/kYba7YZe5pv1wYgizWQPqHcUW9p8IDZpD0KmuTy1KTnlt6pJFoKPEX0FSFBjM
yMFJuJeWUyGaTCfsvlm3di9LlRHgs0MMd15k9QNbK0ufn0+xxW4hx9EdkoL0bk3vh3LL8qq3doiA
PtM5ZX56+uC+HW0BW1HLEECILbxty3OHqB2QkBXmS83eHi2IqXJhJPNgQCpS9SJWbKyKLvTv5LKO
vSJsJWUL86cp7Hsg6B28iChW6LJ2s91U5AgXhudVQ3JW94KsKT+daQu4qAXVc3P+1NAnYBgE9qOx
E+P31L6yQo+ibfJ82KF91l9fpQPo2kPWqwaVCf0QPtH/vMLbs9R8VmvdKxQCdRo3FXKa2PoCoLI0
lM/CAA+utgMnr5YJPXYpMl1HWdgm567EXPf6rumJQVJo0JJ8jT6WySFYYyAdkr3PFokp9X8xf1nk
BYJEU7zEGIjgmyPyANskqRQKrNxKon/0D9e63Cgn++kSp16Y0x5+BA9dmq20+stObQY+n21ETjRU
fJ4FMzz02zE4v81wrFPLjnSy5LhJTUlCySV/1jhZOaNUaPGBf7S6cNaHaZcAPaYka0Ksd+EEJtz9
JDzZWxlRD7xuFB3BlLfP9j0GeZSLBis2CDPXbsHqdAYTUClCZ67V7lcySge7dqoa5x1mDJCsHwLw
0ywAUgRHF/ULhAhZyRqf3febGv3LfhKTuXnlS1GvGmNAYYUTtwbMWm9AQPYQ4XSDbIKBuKDjozt+
YBm0NbcEOPsQH13/crg3eMn7mz5TTcbxpHpHUe/R2kqvBvnZVn8//TIoTWI/tGxBaUAxg6B8kTGe
42ZN08bIwVgfEcOaZePWhd3noOIDL1397u0FgTOrTU1EIWmYVxoHQ3qzyea1bx3WHIFGC3LUrMGX
Kunq2G1NdSngdwO+eUqtvzRaGJl6kXJ5luxbx0k3ioINClCPaan/ihA0o1gsy7HHtLgqvX5jL8lt
xZs7GEb3fUxnGJZtBoaqhbfgVSUP5SqpGnSFXZjBeKJdnbNtO6+zddoiwLxfVtqD1Lv0Iirr9osN
Cb55aW4VCmI+O9Xr/c556jFAYkJD3bn+YMBBmSZuV/8zusAGXXzmhlgc2is0DIHEAVFz8m/Lr8ZD
f1NVrPeOTnOKLQulOsMadP9WlpZYB8uk2jgc3o9/fA263vFwqKeXJP07OEqdW1oGRgAltnzAyBPG
h1Gw38DYAgVw7PeAHsxC/plySkjhqgi5CdLXdb/fMGdor68iGpmem7l3PNxI9lOj0OPJykDaNBeJ
Xb4Ik7bI+VOETyAtPxn8Ohwcn50ENe4U0Fd4uhAq1vY5WPdbyRifxTikkx7hmGxNcd+iLjUCs7Zz
Y11JGURr9OZQwwFBk4ANoFn/ThBLB3SBwMtCwg8QYGsDapjqJH2b3UTUiuAtPFgU6jg9wUQmNv9c
XP4vQ48B4/QdXkTIu+4qbVhk6lvhts5MDDg05Huv+JoC50RzQSEm3o+Thod+ZUfcpjS0fP+Q51uN
vU53fwQ8oCHAw9Ow/jH1NSPo8Uwm93NQZHrf2LjF9ORAFC/PDuZYS91hUsy1ubIxqu02lGwOM7zi
oROaAI7vCt3f26c8QHbJnICy0V7md++rrdMJ8AERdEG1zFS20OguHQVVF3/PgyHp98G7c45Eja09
5NTVAikWc2tiavJcHHm1CsoJP0sqnp9nYlrCYs2lurU4sHOCforwQ1AktYH7TdZD8CU09b6qnypd
3S6cVe+qo5OfaygD9NzQgXP/V6RcaYaSZTjXm1lH4BXnI7DkNag66RJ6ofYI/HGLqxpFjxbbU+dA
BTxtKbdvKrv0LeVtYTwek7O4gT9iDJgUiiJ77iCAVxsx0WSQ4lys5ojNvbJMa0LJOxtpJRKzdF+s
kFOHo2aMlkYQvC87p8/VD8ZLbGVpp25DivYZbotL3EYZBZj0W/23i6N8iapypKQX4t8TGiy69MJ1
TVxowUFkYqkjHbGHDjIhymmzfZls12Y0tNNIdtv/mAr/arZ9Yfxx3Wty4F4L7zAo8iGuy8Q/hwDf
jZ14fh1+9EvrtnDc6HfD59V6s3fXXNYAhgrfWLN+QjuzK5+FPLH/V0W+oDQ/UDK+y9tXMeAUj0nc
dNJPo0ah/Vs3ComO2M+4Z1PNiyn/yFkdC4IfGMrq2PchG11E1to78q80mkDqYcw48KrIv3T3BfRE
10a8TVofKKw8YW3pAwIdQyMqQkmrqoDlCml6UMe22ns9jUmR6yMXL9G2+XY88Nw7u2sPZPiTlfeH
7tlngOF3E0G2P8kmZwENu9i43AuMXDXkaGBHWumiAY3oupnNuTmyvGjLf6lSllj+cwTayDnrVOgN
9e0yDdmCBUDri7Obiurrz/ZDhcW+ba7RxGxwOhc/v6OTF+ZgmBqzOn69wroHVrLwxR96Y9qjzpH3
Q0Y3IJqj81NnQTgwzFAwNAVte6gzCpQu2kBjLTIa6WTt1BMc//4VzH/pyP04oWlRAEPpNkDyPm0N
XnMwP19u0b31tRX0QBbl5xNzvWpYMDCIoyMek/hI/u46WhMxaTvTWMIwEv7HpTHhAD7IJrHCLm8j
9Xccu22AFxokO44efU/0Ze1DRrYBLjF36cZhO6zL4Ym34zYV1JmeyjMgk/P/i1+xjrXCulxo9q4u
1Ank/Z09PH1GP0EX+hqhMQH6B2YS2ssnuvFVMeac0z6SQ2fUT8PdJUTlE8MOPiNiptvM+2qSdYT4
NycRFmK7Z0sPUqqBCjmp5Wpvq2sEMLnca3hMHyxEqL6PToweKO+nBtawk0jns9dt06jGp+o3h5U7
BiTGsW04hvaqQObEj6D4XTOPU5TYPFvcX/Vg9cJ7uu/3A7Fn4YUpJPyts4UXGE42o7pmR1gpjo8Y
MQsCrF3Vjs5UrglJAB6y029tg14nLOAMDmup9NOV6hZAW7QSp/aYtgfOQvoBe5cL389j3FIKuOnP
wROPKeew7fltsEkDw1rfIYgvBwD4zZc+L15AX6+KvSRZbYl+u/6G4KhSjYp1RGn4W341sfcbeBv/
trIs2p+TuRgLhW2vNZaeZ+3q8Fyy+5vgMw61OhvErtxua4ZdHG3P35x+E9C1lPKA8/W0TL3kBZdb
UdTIN47T0ZkkiXxUwNMevn1NiDIRORWp9ix0y+REBYA6XTZed//v2uhaBXsJYVierHIzXHd6EF0c
ASEMQlLdDxoKxVJrYzbQIRTQltISfI21dGPkn4KjUqV5tFcWOOUMclKd7RY87kE/Bv5ZUPAAIM/k
436RBwDkBqekm3zW7d+q5BHSFaSMaqzPZIvVHSCH5KP7FVPv8Bqq3ipnm1lTH5+2Dx6BkFYljLSy
l+iCWdsHSig3uzNEH4zC06qzByZXpXwTLckD+C3YAn12BbRQYaKxVGuRzKhVQA+PzUf/+kWDWLyE
6lt23BiVkdGbFiUg2SMglmODvRG09ZtSVa7CinpA2Qj0x1fbJbX5tzGGLFl/OqEPHSaOICa/gIlS
+rMeh9MdLxb9I7o9XGo6JMvK9eUH98tsanklpfMNrDFzQ7c6Eu/p73I22dT3X689vIOsN9tik/52
RdD5fVErcXRoi0nj2cS/GmPVZ7T4frvETtZyPWmlLKz/8xRl8xS3VLhu8Lh5Sk3O7vXY1N1S33bJ
2iufey1YObgBnWa7/qkQpkj/OJl19h5VbL1+ZGZ4pIUKdDsRgoANSpTrkIToP9Q9zCbfJWDUjNgf
nfISun6ej8Ypvw1ZlVty+kW3SKyRrT3Ybxog9lMA2+zrvAeXPlnprzJ4njsCCkZNOfw0mOfuM5tx
yyKIVT/ODAD79WWibsa224IXayWYmJmvLz/tAlIeMvSG/KTfq5bWuHW+nPHh/vfGqpTAaBpx5tQL
AeNvCe0nVPfuj0WHrKjaxgvwi4LmC72ajevtpbQuuGYopYDKfNJMxnZahown6tFgZOI1YrGxOULV
ktOEWPa4OllLjLwToGCpzNh6ONttkdnlLmBqEw3zxyHhumubeCCSSdRHOyKtZn1tjm1sU/uWpPH0
JoUI675/BylgbqdAyRGoKCoSRgx1cjXkZ4ly7OLVucLO8tLeHPFcNWYIGshYjts/JODFGM6zuKym
lnx8oN3Iyl6J3fibG8LfKagKvGTwFLP6vZ93res1vAWcpnV438FeboKATOqWYSP7tAHc6YbHi7rG
M/RIqWHjaiOSndKIXdWC+BuSlrB3b+JmKHJWqMT4s/J+7hrjV7iaAYpMOxsJfWdAKNUK0HNdsjuJ
uXOrx41ML1Vd1TjE3IFz9W+3k994U79Z9lZd5A9Xkz7gQcL6jkD0xXPrV1ZSm1WHe0BKt0j9er0Z
oAwF8e2shBsH26UyVDUOR4ImMykPoBbet6J4GS/c3Ue+oLgmTAJvI3tHimr4ICWYtEfmSTc2hTrp
JSBjeo5WPzMePxjo+PTM6bJr+iZHp1L7Bg1JlyqOrx5YuJ9HGythMoc2WLsw8kTMNdy4nVCyORLe
rX7ylTz8LcMhOwn0nuR1CBZ9s4qePIDjM0XdE4Oypmawd/6j7CnofVSGOUKW11/WINdnNTI8udnB
dbqgxwkNzwFlC77aXFBZvl5JWcQH6BS1Na0/SGey4Q6ZMafHn+JcOiFD9gCoEwCx/oE+q+dthxLY
FqeiQHqKcEiPSm81rZKeCtAeIo8wdKu8nOWhPk/dtSAt6J6mTi2d1845JscTFtmWw2LqgE3slLuS
ImDyUytE51f1ugz5hPT91tTDGdJWTkfFeaGKUc/8Gcp24962ceqULHA0ctuSvj9KeJhm4EeoU6ex
kLzeEMyiuOceW5PA3K+Q/mZm8YHR+pBmXPeh/b36NL1w2vDW8L5ht0xhRbmzGKQ4dOD8BY0MXrCE
w8n5LB5S7vnVM8vRxIizJ/ukyc7x7CpdrFdF1XDi5zp0cHpEQhBrDP8OnV/mxbUB+WsDgLYwRTqa
6vANqIKUbY11+KRWrSOxestbOhqPxAWS2Uai3Eai/z3+v3p+r80SiUjNFHA7zz3U3PrUfp9RviaD
dZXpFX6Zc+SxDhQ3+8RJmXSh6g8uHuvL6ova4lqcGag7iTrQ5IGcyZdTWLOtq1GaVwgWNvPCIRJc
74pIvobZeBLXSBbRGTpuZbMl36F1YtW7DKlTBcgXdtxFgpdJoLLTtpTHG3BD9PpHThxNPpaRqwzO
YGNCTKJgM8anDOxn/nFOxzNAxzgIEbTIDdS1Lhy92PlL7gX2K0xMh/ofOYDVuRYC5/gEzEjrZ93X
A6sDd8im6rFNV1CYwzYQ7yhpPu2kDTSxuGtsH0qnTBZiVl1r+rtlZhbjknBin3LpG1PQMv1zlJ1l
zS57vi2DDJHTjQEUxoMeWGCyoo7OGYixVhCAFJYHexVsnn46F3Vb9fnmaDMY8a8d35IxJguj2BHb
9IyhRVNsfujAL0K06dVEH8fP6Ha4fHYRmJKicaH8bKYT8tpLAKCpfAoWo9QwlkqQTUUNIEVhQu2o
GgPqio9xN2Ga/wAAKFtYNSj6WBb6RNpvjWJ7wSRaoFxOb3d4RRg+hGeYoHVlyJYA/7GHvNDRvzjs
5gOYuI0mQ/ZfjO8K73JQremU8YL14cPH4BhRZckbKVak0Bhh67aTu+X78ltayRIwLRPaJ6XS1IOI
/8/raeYIWj3zUI09d7u6QEU5wSmOl6a7t54XSnHNQohOi/2oogqNqadNH3Z7MH4SlRP2YJtiOlSe
jMde2EAFMf+PwHNnQ2h50fxI8N7C4PsJeVtAnfPP2Ts3prBTkNE0v+PWLGgVMKjKWx+4KTPGxfj2
fYJ2fipMTbXsISX8Ldht2Jmur5uYfClf1hCHJNxmtOuKjlJzQTOBF/107oCxHFwSBLqHGGYn5DTY
jSaH2SJbHQTOmMgp5pE+A0D6FSilYt4QZM7A42ssTw/dnlzOr5zcAr4jnS3xqEdLvBbO6daFZ85g
iDCZpZWOkMOV8RQFA2HigCwNv+u8ay9LoJfx9LOo0LAQTW124oICgM8EXdPn1IbFFrSISmxNnGn7
sUYQ8Y2YKUpOfr3aHZrixMwDqlsTijl2guexnR2SRWIzvBEYNizp73OovhAkH49H4fDMGnFwLLQI
FRUj
`protect end_protected
