-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
6SqWxNwNFCbhbCXiv7a06rKa82ifqGRqAZQp6BRYHT5Kk4u2xT42EmAlkRDWv6fP
tLqpYkjnO0ij9R4GlA+9X2R/P6zB5KcK9yFimx0AanCFsvDEPG0YEaKNWkrJh5gP
LTR67x0TRFn7ebv2ywXpVIrRWCrGVwyBT5TJa2scRXNAIwB1goFYkA==
--pragma protect end_key_block
--pragma protect digest_block
XSRQmW10nLtYc8GiKu9/rbD2BYo=
--pragma protect end_digest_block
--pragma protect data_block
e/JCGXqulcWKm0bx1JuiPoJQyax0NzPTgn+1tOeasO5M2+kcI+y4W/QMgfNYKp10
jCoeoCR2iYwLCzMgN/gmB+5noiFe1Sei7yniclave2tQZ9oQ5VPzWmy9zZOah59h
6fw2EwET/oU2MJ+1JrB0HlIOzaRtftlIG6jWNW6Xbe+fZ8zLa0U9Qjp9AHBMLMi9
ao8xncjkp40Ugr6J8zxluq/tm+qX9zwtdz43bLVOaW91nSGcCeDrygp770JYwNQY
Kt+N6Os5ubO2d9uMQvepXDB6527LTC3EA/wrL9hL1GAHVEaIaH6wddFDEoLVLq36
PRPYZrSdatg0EjcI6Mgal+9jKsRWCTNgEqtd0kGptVQPzyXEJneyq7dmA2u4wQGu
f3esZ/xxCqbO41Esz5R3g81Zet4ymDQEe2e5loXEat9s5S4J/JOyq/Vek3zn/rl7
3A9u/VTK8enKsei9q7lLTghI8CyS1IoTxxgMTsns6t6RoQG+Bk9/pR7ky6oa0sgz
0Dx3/mqQEuFp6BpSaMCPxr/H9+ze+DIQ35SKbOOIsAPeRojFyDHS5g1Xq11TuQAC
AJJwdyiKUPC22QTU0OUgv2Ocm0OFlV9yJCQBxHt0isyLKz8t+lImQx82bjUq5nIE
HkBVgSHL9n2R+xOIqnTsWLbcftAgvJkFFfKA3cDRv+iPQ14XpeLZNiQuyDXyQe76
d+mdrYKy3Ndo5bboZEs5h4ztyvXVLVmJoRN4jP0DdYH2Khvu7pgnNRbTB6VjHktS
P/dQjU3hHfHsXBQgw/278O56kNzalzupnlduHtWIcp17GdPMPpSmsrlTwtPtW2LK
LB8wQsga0QiTOeSWnqEifHVNDl+YxPE6xlfJ7lwNtPTw43MdSZS2fHKAI1BQ5nic
8WoaaiGGX1Ua429FCdu6Yfyt5U2GeYvl7Ssdg2eOKSu7oD7PAS12e8Tq5v6T/Zdw
prHG/oBY++sCpSr8R5eDbhlvUSaNHpQL6wFHqqw567HIa2f/zchmqQxcEeSOpp13
DV0fJyFH6S08p9PiMNSqThNBzOmMsEXSDGfuiE0IdFXsj8dJhSx1Kse9V0WYwZ5X
E/U9RU0rbPhSuQXq89XSXDmaM4utyDIRP6UuiHAYqv1UoJhIMG+TKdy9KMfCT4nv
//TCtAZLGKXLY+iLTtxeWHT2TTo8diwDazunAh/sw59Jww1Fl1jTUhJbeTh7Ejbe
/kjmxcH3rE28nVrPI4MIHM3/5hQLzw3dqOQRKyEjHNY9dQaAajqukMwbgaVVFN6g
A1NKHZ6z+Wt+/UIEenbF8Emhgh9AjWpUQ8yZHGsZGFrFGeTkNhLPt4uYRObtmiWz
DjmQ1dpaNNSEe6M00N0Y/GqX0GmWaxlxnWaf4Ru6nnlYQoMCdEpOUgAgJU0raT7V
+lGIOn570HHSpAQ8DZ9NPGvffot5wxmXRcXXwQNYcgOen1ZpgHnrz/Sc1HC3JTjF
oalOdhzlS29rK9Vyla7X1NepETE7H2Qq8hXo0IleyKsy5Xo+serHhJxNZpSKFRlO
DGicjJD5xxSUzFbOiRcd0h+nU7u/278TE/OVr2Pfx3hHl1EELiNNFZ2hhB/3dIqX
96UWlhUUuz0hPJ9nkmyvOPji2kTaRV0IPSeMVJrEE5Xf9/rf9Wvome7rDZeOkjyk
N5Qef9l4AMZTeoy1JY6tuw==
--pragma protect end_data_block
--pragma protect digest_block
eCtaKVQCAI6YFhlzEAKLJBCy7Qc=
--pragma protect end_digest_block
--pragma protect end_protected
