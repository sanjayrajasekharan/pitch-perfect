-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
D+Nj0Essk3RHkwYmLK1uaagUqKbHbwVYQLeDEjiz8RfFO+sHmeWa1mEm8xP3Op/q
kklPxLdakD/R0VzzNlJsmNar18eio/uSMyOoCODSdIeOZg1HBSs+AlVu/iCVERhZ
j1mfcEmRprn+z3d3WLpMSBkEZJuQuxPnGt+JoP25vCbn2lQaW4MOKA==
--pragma protect end_key_block
--pragma protect digest_block
HI0tOcQMDnt0OJO7LUXeR4FxY90=
--pragma protect end_digest_block
--pragma protect data_block
tcXJPfrFSUJNlGCrphVqJoI9pAKiwSwPx3nP2k4w0AFr8nPPnuAz1na9W4BzragT
KApz23ucblOgBbDVgcFryMWeKpC89wQa9/SG4409kRpN1EY8EYIub19MWzgVqoI0
jPAIJbiLObOaD/qtjFzxvRbqPexbhbsz9nCqE4jhEPEnv4C0Bdo9xCnnxK07UqkK
ZUH6qTEvAZS3/vwlWrSXMNckBBRCy1D+3JLLBeuQFzZ0gwOBweKm5cKKenHZqqMW
roSVjsbX3kozljL9HclmOh/cEBcmKd4V/bGw7JZZWJPKXBxBZv4cxnVXRjexBgdj
Lu6ntUHEhaFoY5TaDkul+X5u2eVazDmTn9zJ4Bu2XSyAp1aimwB0wU+n50WWyiMf
VoxF0s+4rFcir24YcyV1PqmSAXhaSGGf/JiG+WRNzO+28hjVDROY9E/7QUiabkOZ
dVkmwOmWGfHmH4QOITVmcjyT3YRG+Ipb+sbxlqxDP/BnUHaZm4ELEWxC3vJfF0Zu
qz5Kaa0li4IOSLfsjbQw1PyMse9uWL+WpxPqkHGivR5GSIqQOnYDpLSi2j6nIl8C
qiDg2sxIypvmGtk7tF4P6q4YxOUJFzD8J0Lmha9EGf2Tfyg2kHTdAF2DEom5UJir
kzH7AEBvZbQxdJrs2XXEaWkMEwKREDwPb1btPkv3GtsZ/zUZo6MO5vMd9DvW9O4N
UgiKDlSKLDo784mcgsIQr5wGrfcliKEblgSmdZXDb31eA7b/hm/wd/cl2fv9Nq+x
f8vC/JFjFUflJrRfV0lS7xfb/6Le++gliW2tnpamtLEEIFAfvrCSp8ZL8j8gQAzn
yGvDN/SubIf01++IClPvUksc83TL4NNUBM5w+ZaAX3vura7e6jkG+kzSfhYvPgQU
F5t4syxjkFa7k8LCvRSKduNUHwt2EPPWZTTuGqDNQpt0vVWjR0MdyK550wNhiFBG
sAXj7v5q9KhuA9eSJqFEMj5li33JV/jWZRukX92mwnAYCfsu0n/CqWFYmnVzTyqa
Pz4jVZnCkV2lBw0X2qrcwktJ0IG1yE3J6cP3nW9QvFQ6Q5226X9XKTIal+hZSTsO
nQWX3hSjU6ztToXwP5igWDzjCuhjjCuQBEFOajLi5X9i13+BJIX83MWTQP2ebNMJ
0pv+9M8o7tXPcpO8PL0BojaluqtLL4I9MI+YVI2HYD0r2LCZCWTkyaGfS8h7/jyZ
KSG+2arim8Hr5bdQOLlP8sNmgoK0rOjHldnuH8z3SlXLJnLEOleXX+t63PcKS9HC
B1ledOKU1YL90xQ40/+vCVBPDbjHaNIxRcy/ZSy4i3RAWby2Ki6e0GW6HWVDSXzW
8fAVVDtHbOs94V+otaieMnJmqSQ9vZPy9Cp6be57PheaTfwyPGtmswQHngL7PbG2
iGSGyArfFZLEQ0nZNU3IBJcviWPiJ+bAQs8Bu2wcCqc+qNoAv+mG8KkuzQ2pdb3e
E9RfeyN6W0w3oM+oCWIlYrSrQuUif5VhQFe92ja0IMC654C9M0kGNeVaWMuGCL+s
VwpH0ULTT3VvfbG66uwg9wabM8fPim1A2WSSq1wM2/DN9PuEHyW7sJ+qCNgk/+iB
JMoFC6AghBtVwLDsWH1pT3RMQWuAGFMMBa3x5pkz4tl4AGF6ftrFx0INmVD2IuX9
ZKEtKpMn9Bvb32TbSyDiCivdZoAzUmI2ANKHp+FKVQ6SDB+I0TQ4brngInyFTuSk
Q3hQ3bgLTYeqQOrzEUACYKlJdEOM16/I5bPSU7tKdlnd9vpJo8r8LmgNtIqN9goy
j3FdMCJVAsb7GguKQPOLzvETrfJb7H4nQKsyeGadikA4XUnafXF/znEEsmLAlo8m
Y8isdq5DuKvhUUEt3AfbDarsFbZ2zCtjsI5kIYyQllZ2Ii9Jx9NHTIahQyN+sfCy
fahlEvpZIlUPYfEFpdIA2IQrXPVOLAj/PYflycI3WhytEiJ50TQSmOPy2OnFoM9U
r2cjJjJwShgGo/ihGrRAh9VvbKv6D8j2a2G6zAtxfynwgB4avJ44i9w5l2ltdva3
/6Lyw7KotxodWAcP8/6Ia9q0pnVRSQoxYks6zEK2A4iVNYzwU9urO+D7s3HOgL4j
iEpxYTzCt2DS1UZ2z8ys+1n3XBXT3pKgps2OR1kXfGf4ad+KtSMSqX9kUYiZB2vL
o9UWfO2O5A1egLnKr/aMD9iwCYUApYC0esra4Jscj57FqaZ8KzBIxvJQqTrrvGYT
18UJNY5MaJ93/VlEK4RTrcPUD02BbC+MTU+FcCK65/f/o+yrJ5kQC4yQbEAfl0hZ
JAH3khCSFrsfmQQHHBme4uBSfKqkBBXfvRWwc4v56LYJ1YBV59ntyiXaxfIzW6Kz
NXQouJy/4Xx5Vc6AsbaMlnZgq/xjrEnHMoi/wa+jqozC4HRBE/Ud9VhJrmgck92V
eTULUbd75D87qAu72AhiDtFPP9/6Wje3cI6RyMiuDI9iX6Z4bVxUGW8sgT71kbNb
jiwM9k/muiihejOw30sXC4S68qmEQsG+WOKZYJ5xg06oCp3fdt65Xq2fKvNDRwTJ
RC+CupgncoSAUt57iJqWKeLbwCHpXyN0SiQDNH1VURwnZ2RXov5sHGzKHHUD2Oj7
k7ukiSkmZ6vZ+khFvs+Wnfjr3R1G9raEf8e7CNUanAnpAizGEpfOMB1qgP2rZdj0
tte295L877pUGSPVZ83E0SZ8Nq1y+4LWTDs8wB02zdZJVEH60aiGQeyBLe26QX7N
oAQqfOoxZTvoYC84pdkiAJfm01ZUpKeiO/oovdxHQ0w+XwFI/LGyy0PLeKfUePWx
EunV24xm6C4zZ4+CjD9kzRw7BIxQVselRu7Uw4P6AnHa/10haIP7ZZ6oZOE+Ts86
qEpOJg/t8pAel2TBBLzXzWWyB1EAYpl+/RhR1waE1hZAzhboC7+xaGmR5eL4uJPR
WHbVpHH900lBXg8sBrnY29TXBb6yr1SGCVc4cB5GqX/Y5I9uTK4KftMRSmQ9V2Xo
ltyRoQVwFJ6pnFkxW+3JsHYlCqK3mMXXROQs3voLn++dKXcb9vM693/R+eD00Q5j
INYulhQQTZRIIxWLEHi0XMKgFA37Wbzi+zaJVTmQ5f7i7tf63gSS7nfRhBM3+sIT
Li3/x4Gwm3IK/62063FXE37KiDVXYqxQ2WC+00QTpXBv7oL3CGBJRldLxU6FayRV
l3WE5UaGa2nb3XyizFLYS355lodpMSk6wOpWS+acmv7KUoMHc5XxJPyc9S13CMb+
EFgLeSa6nj0rXrm2CPis2+s1nZLAXFG5mv+XZtca0ogXOV2TOb4LnmwOLz4t3xWv
4TsKRDKepdLBHpQZdVFVxeuIwb+RWTYf3uuOLEc0Bnhdr4R7wriv3QiwVQcn1UDL
EL7jvzzoF5m6pXTEmqt+/lG84dDcyFKLhUrE86XaFp6lZ73me8BvXtTJQ/IGAJoK
OzebeVqX46kPB3esYGx330ggyhJR8XoZoppFQdmZ8mjum4ftXpme8d6AAZ8KA29d
EfxUfIwcsU3jtjxRt9gF3kKmAwHJNapg1UPUl+7zAajgWVVRM39n2GrWwJj8YvlV
FrBH0cVM/2EDQLR4X0taipkTuJ9HxQZmDdesG6wwtwVxrlxoWhwIQRBdGA7DeJYu
MOGFe6vRGR+lGk+DDqC4KvxgZ2Q3vT21q4GsERbtJxO4rxK6zSCcjdhXLReM7Dch
e2D72RQm2jAe0egWqz6UDrSvmKE+aL8sFVkvUq1oIGjttD4JAAqzQygtf/A3w+Fc
9/OaJ3VOIHdZd5iRrfzMxdlqsIkF1qn6NFZF+PVaysw44br+Ca/5DdyIcpEcS6Ue
zDX8JKHp1NphZkhZhgF345skl0v88YePRVZwwc9EqKH1+Egqhz1AN8xTAcHbxuhJ
71daPLThI6Gbec6IEaznntxZQFWx/gFuw3IEJMv/2qXuXAXtMk77glKcMzSig08o
Wje2Hg0X3Ul8VakBx2f6ehlidgE/iKP0AZLLbsJ2OoqA+r//JwdpXdsY73ZTyUu+
yGrH30Kg4celuavFb/1dUZvX/HNuBUUQI7TH1lUijN76IsPXh4HEPhyd4p8KsE2x
eVo7dyRArQZKT2E4mA2Kw2okCTmBRHsGHj4hYzS6QcxklNhuuq5kEF1dTu+zueef
JeEGeEBy2Dh+1qMcUsNs/W/PyQI3R/TzjsaAhUWJ7/rRZlDj8IzUFRQ0KhrNFhYu
QO7Bpi83yFEelDLXHQ0vLZgmVYiX9ktEVFVRQmnYfXKnDHcl+mUKtIQ4np5kX8JW
CIrgurH4igQLu1CVA4jYV+NC6IV40AQV+km20LrsZ6NUKELjP+Ps2ZST6yNHaNRH
pz4JcDV8VyNZV+8qjMXIx16Gq3ovEKqSJHdHOt/RZctDJdLlaFnl1glba/8qKJB1
cq8/00U032mhLlaJejNEeM4xWbQvkw+ytPH6IuiKuwBcVS4RWU53bPN2HdbeGj/u
H+wf59JPWIfo8nVIbfp4rYibdlamoHeZAxypds3ZQiyKMYHE5rH3snpd0PnvZxKl
kPH6mLBIytJR7oOvcCQbuX7T+yTUizoQOIdoaKOH/e7eMs+4Wox1sjMSmp2oGMc0
75AeM8/hnO4q+sGZzETIbARSiPrjCTaZEgXp/jWo49pE4SZrBFc3h07RfVrxCzLc
tlnP4QUe/9T2T5xs9Z22wMIQdD6RlwNn3uGm30OI9APIittykLE/iFf4armPs/dO
mbrCv6G9ImcCec4if0hVAKhYiBulKTA8hvdLREKiFC1ZUpPAh/P0/wm+hH+FhzQ9
IQxhg7TYQ0WuirczlqQjmZogJVpMkk1IpfmWF5bj35n4IWC1D/hkFhA3a842wCEl
Ue2bSkn94tVfy7FX/V69HamlSHjKXm47T3Ik+wUUxqIS0tWpMXaFJW2RG7xwqW/B
y8TUD9oWD/eyqrn7d3lZGyZmQNJBPKP3YX0hZwQnyls3OpNlEpwfTpvPXOocAUxH
2pyZOPPSvDXcuKuQIF1I6OWqErelwdOW5veJcv4gcuVD3oGK9//7JPLmZ0U3iMCq
3DaqS/iEOS5ljMmLlozE1jOPk/sPBzKMx42QvKVBy84oiN2Q6WJ1hGi1VEYlEotu
gs/qOQc243wEiabl7OKcuCtyDEgOJ7zC34CPEJkoJAa5RJJSrxYnO7kV+F5G5QuR
/l11y29B2vBYohXnwX6ujrlPYuJmjy8s7QmfW3mBqDcDgDbAz86xBNvsEc5V/VaC
RXAGsqPI3miTfkfNESKu/4GhmekyvJ3ChlprzXRsC7qsYzMV5TDOw76ewO+W3JVC
JOwmqt8VerRHcWkkGHy0SWmR+muFNGYpLjC5N4A4sQMrV6V4hx8eX3ZzYV8S06x9
DN3O50YYGE/4QFZkFmy/NPQbvv3Bwb6cFuBKbBX8lnEdCvY0bYOFooLzizsgEbs6
Xk+KnW1FtATvs5KElkpZSMKTPeJbgKPeR6jpieRBlKUdySSgflnaSEtYH3APRiew
vNJg0ekN5LtmP78TX6LdTDlL51VLspVOnlFzNYAc8ljF99KFHXJOjNASjUEI7kMu
UViJc3NWFw1SURU6W1ZkdrFWHCbeYw6RoZh+X4EX7UpOy4ETJSMxiDmhLx1pfZ/1
ujE0b5AFdX/y3OzQY29JObuW1sF+lr0EunDD6XuUM2wAaI/nyieCJDJn/Y/u56ev
7fBW62rO0T+y33AskoDBmGMlh3T4DT+l5OsYOT8b6qgRF87JUQ8vpxr70SErXgOr
3+spBZUmrx3JCe7SnmwflCFyMZZ5ihj5RQTLWTGmZNhoeHKvFEiSpu1clVEq18R1
jEZeYS/26CnTJ34sGzhDNlOmYXOnJbyM4p0b9TZonoHQEZR+NHOmfZ0Zd03T9uDT
0KiveUAqcDWVNwuND/xC+fi1A4sxYfaG4v2PhvTY1uoX+mfoOb9x9iuxzjA4eGbS
m325f4fVMwmOf+efCWiVMsOfVMaAuX580ZC+Oo8jZ18ynieMrvFkCBjJF+B3QtOc
jj8Nq4cztTR+ZKoTj+ClMN3G0ApfAPhy09L5D2ArWSBT4bB7OJrtAHdEDM6VknP3
XAVmSEZMFb23HI4fJbemd5FwrypqOY8+O3aZh38a4w7qSd/DsDdyjd0TBAFm47d0
+gvoaJCYMUWvAgEDoQKNKd1VyHQQPkPSaXYei0jGdtVhK8yERZPL79MgO00THZ5C
Q2s6v+6wdgXlX2ZnL2btsReeFPWp0buxTeWU9BvT9uYSt4Fgd7UDtYc8CVUhuQin
Xv8mMyfyy9XRseFXIMTzZlGV3tk0h3d1vSZf6NIaOdSwB0FdLOO8vQE33D6kwIh8
0E2c6NTfyVYETW8oxlTHaysd4IHiIfvDKA0/oWATPIPLNJHi5sUB63mRJfW7HD0O
j64NCzFsdvWy9FYWZgEH7gjJhSHIx9jb7uRXE4kfUZzd5rhGUw5FMxYeH+LSgHaP
9nOYqwVFtL9dlfBKlcNR2GZ8Wq7H1IPWdI7ZOLlAIKtfjUv2auxp5e+G/KnBEE6J
jud2HhPuHGeUGrqqiLDKhHzXKCwMSRtQB5Xmm84wZ3CDkroRR9DRiOUNAq52TizR
B7bUJGSq9XTD8YL3Xs550osWlpl24rS5lro3r9q+ppE9x4b1GGo6GPI64G3AvfQk
wWZCUPuxerLW59cxUMT1K3BZ+WkETKlcXCgHsnkN4pbRtLTedi7MpU9VWCste/82
jXagtvn88Q9dKpJWknehXixUx2DWRXm4qPqmmaGgsDmgr3trxa6ZHPSbuVRKRT/T
ejEt6RqkBglEM/t5dMwibiPIbEVkSUkNYwMV2ncyImUUFx+GLGDdTR4uf2yCu3PT
DKN2io/gEt0cbaDKsZCkvjz9a5Msu9I0RgITfUmgzxUd5C3tEayYQwO1gex6HHdh
EpH+8EopoHNNDbnfILfQrZ28ypA8ocRyk2l/HK57lAl55YSqapsc/G27j4FTfFPl
xn2Axv29N1Tfc/TTWCobBIPHMPlyqDW3bYVvBgNwSrKC8ACCbSC7eCi/ELaFhsEc
i+zSKbtStyRlwiVo+m0m7aMzqxdsYe8XK6jpGNZerndO9uBEi9V6GePqJbkP2eAk
JUD/0jWaAQTEvL+ZjgacUmdkak+Dj2UypE1HvCq617XTHDhc/JxaMnlrfTvpBe6I
UH9e8sVlinnNJxKXRfTzLH/hkdZHblEH2eQUGuWfucz443hSaqucb1Ib2XXrtdMW
dIqD6MtdqY7fsIyOTSSLBoTVwjjO5jBIifvr/mhk7uYsNfly+mAvg3uC+hq81kqT
s3ICX5aMaG9qRyEB++XN4JMWPrnQ+R5v8Nsz4hBfyLEK19XKvSG69Allsnlk3Ow+
VzaK6MF25v2+RusGMtxW9n6rvgHmTCCXc4SXCp54OBC+DAjkO+75puxVIiDJVYAv
mrkrs4zrP0Gj/E94Llj83B+u+JcSvUqpSZm9x8TXPc9m3/kE0NeuQ2RM1L78WUWt
8mTbIGo3SMz5umGcbjYY9Rp0PuBwiY4HO0BPCbxZGLriiCO8FPdy/jzcDvchWXM3
CWG/F0seN/JNIvsVSpC8oKU51jxpsWEjTvml4twQx0U8u4Z+GFrIVTei4aC3vZjp
l/JNOqgUj4slgnDaUf/BO9g2n61KRYdPEj7VFrZ6ozh5wCC8osWiff2CUB5/XWZ3
bReZNu9tycvc63n1tznfdiGwDB4onOV4VuasS988IhgS+mSYHW/MYuHbEGE8qNFh
JYcGA8myknL57RsD+gfWMHbLA4E7Q19a8x9K4cDhDWTBjclhdfcH17qufz/5/cUH
cX3I4u84EsOqKlfqmJhKBal9/gVi4D9oHRvKw0uC+73v1qc4unM+c89qF/SVKZNR
DUIot7/YUp5oe/LoecXJYKrTjL9hegiHDbIUXliaNXEGdufJwy58CmLiZGLoHDyk
idiTJQsUYxmuo9ATHv42967ikvIltcfhpkL3iXCWBr1CYcTfZ7VHRmoI+Rsxl3H+
PsCjfRoOEjUuSnECLPGUL7hFbwuklsx4GRL6mNdpWhAovLnUzJIUmHvi9boOQQMe
Ng7fCUeDU99EA6mTgbS3FnrOqjVDCoELXtqHQ41pluJ1w6hKqcUsf2JcJNBfdB97
T5irb1yuH/WbyAFV6lnxMlxAf6Mq0PgXPQql2pBmjJNRcS4TUKBJhO0eoYclEHjY
cWF2PqD0vCHxcA9Oj0/nUO+0MqXccShwyUSGHZSrq5fA85Q0kYofPVvIGAy3qNrK
Yoze5ddL4VntCnLuPCCN67osXnJQTrg1Zc71VCXqUdAFr8QxIE5eFemVboBITrcf
EibOagcgwe3SyYwT85LMEWu3XAXphk3qXmk832Ym3XtYUUnKNF99/60xXa5LhjNC
9fxxLLL5oA+SL09x6KWRxi895BJjAtxRoIHYXPGw5XAvvEoweDScHk+xGnys6LKL
t6KJhFEqJY6MAZVyAlIDw/Q6TA481Vaxod/BYsjCr89nZAiyYpfrMCBWAd4+2GPb
Ahswv4WbTd28vw+BJksqpA0VTUYBsCSGjWC0NBlMNa+IAsVforAgKqbwqvJvt6Ya
Dx4qvs2E5jO4LauAQHqIuFKGpURU5AW9G6/pV7c/Fvl/Lp+LVzBZW4d1TiBcK8kS
YggLuLAmygpcXI29hU8bX6zvbD8A2neRU8ZZmQkAYVOLgVpbhPWbVtXX/bmGgeAO
yMOW+9DC5A2FStwSDt45Acafv55zRyyMhGnIrDUAP6SndmyVrK7H4z7zdAWnIoRR
xPS+BVpabUnaN9PlTG/dM4oaPxvYv73YtWlF+1tLcVa5sCwj8/oZVCmEjlXgoE5Y
L+l5yAoUvue4pbQsXHlBxzuGjeM2Spuy/YWtw4C+y1LbndzVp8cAShwxbtiu12+d
OAZaVgeMCJkEiATstBV4UAjG4VopCS3+cITOq2bKc5bUvPqjZQlikhGonRxFXvAi
dtZC3h+1i1J03yFylDWTD95ex+oyqFdpatF2iAmtWDZLa/I84tWZVc9Cd5orIHO4
S6npg5uqdY4pXbrGq3kguJI3HO/hSY/C4xlrsnZ5CTuIwden0sCK3KH8aGMM/3Si
sPNJweVEdR73AcpZ102IQUwGp9cEmUgiw8mtIFzncldpnaJUQYtnhe7o3xH5kPOM
99DNR0a+6hq+yq3IJsFPVGChf2Kzc35W8/PWXr7oKI/VkcUY8XX5N4a5xlpSeEgG
4T3gP5TfaLNCBpIyUrW5jD3pM5d0pyt3peGV+c7RIPY9J5x2akBJF6lOSqZrcDQT
SQS8sXhk9RZs69jFgecba+J/OzIiXIXCz70dKdL+ZCZbVnuyOhIqox9VnnxJqgV/
L8k+RONw0OwgMOlCQUDyVzKfdRrBj1+6nFtyUgPONGHopQ5D3Av7gU5ORn4ZJLkD
1diiCVzsSXp1ts5NH6fnyScLKOF4hrG/OufRKIW3HpIIbEwtDbFrydjcS2HUWxtq
2nqQDQeo8cveexvIkTwCP+ZC7m1W3+LL8VXlWRYgWWRpJi1lErKsP13SXXhJo6Pk
tm00xlmEd1SPuyCPKWT1RG4QqExnK6unsxzhyyWFmG9uvT0bhAY6ycaX2D0v2aXw
b9dBt/ZJ9zwF+cikuZJuzF/MBsNnxFfEQ44xP3bh67RTu6DWBdld9Gldwl3sKiuU
vXC7/DRggIkf1LGuBMuSsbkenV+NfYwevEc+QvD8lLEpadFjdJrkNGW362l61u9Y
HkzpJMRRJ9i3RjieWpujNYyJa2mdusxFPsxF02Dij3kRgYI0Qw5kHF6YXU9XmVs0
k8g7dCbj2RslXW/WKa+eAySjDdGesR7KWEiS5jxEIlr4il5wnaRdzss5QGnF6HsD
ek+7VEtKOnyEiR5XL3bvtUmcjvcXRX3QKtk9xM8R/2riq/Wo2sp53ZzxxoxWYh6S
Nx2iYCI20nf2ehLQxVe2h3t1gUk36OldgnjLx8eGgtapsQu6ZhDij/hw+X08TUar
+CTj4geRc7GsSJESrXudMUBezGJUxwLvXmArtGw3tMaYwnCsanlhhXK7kP9TH9vx
8L5Ezyr8klIZneTBH+POtetoTzxyG7sRzxY1OKhBJPGGmsO49cGCv1SpX5g1DxHd
V4HHuoCL/wzc528W+Gf6MJkvdCvfnU+mxJ+lTu8dQotXGWVsH7jANDVp3TgXWrry
fD1oOn7dqwb1kTe62Oo/LmpyO6HfVpUXK/CiZXMdW6HJLEIdsG8ezauwrXsPBNia
I0A5lWsOKoWL9kJ95zoMru3Z7jxV4+cOE3VzKCVfRSl0PALNDiW1wSWo2EPi8OIs
vUQOUSSkTv3pgKnNGG0HiV+JPS2VdOV2NUMQzftYKqexPLpAwslvXKitaNv/ou9s
DHavOLtuNclIresH2MD890zVVd/KDhnNlmjIqriuYDlJ7B/b467Rs+LQnagIMJJa
PAzUAxGS+cECEaE3Ar+ewx+bSl/p/CiwzT+jhOPgWC1ehnuUdcBo81OzHRQkMli3
/BuMz+byHeEFquKvqIyzLe724cxSbzk/Ldyiqx1ehDy8cMMWV2Q7M8R4rF8xaKns
0VGUeveuaq9IH7dfCkAPcgGfW5KHh4G6xzBV5SrWdIGkqlD7I7LIsCBioi+Z6f8K
F8hA6DO6HR/+pBIiv/E10+cIZNVefWNaMW/DQNbtQxAH6KDL7neQYnABR78IDNMr
SMfXbkhZYL3THjN+NhPHyuExmi4VgOoxgp3dwOvcu6J+FWJ/hQ+JEdWP+5O1ROp2
L4mmgoVdmee5VprqovCEVEsx4GNwgd//jMx6JQBcf+f06aOIMmXx1zutRonm1bkf
B+INe1hGB3p34HF9tXobwNYdXN6JmVlksD9O3xjjyZ4vjT7suONufBGn/ZZ1nt/F
p/QS61t5uZ1aNAFlHkAf2sGVK0JUJ19VHvwONktf3KDPaT3Fk/F1/4h+LCzSEpBA
8AaO5BT2JcikcH5E9euSYt958T97h7uxGL6ZgJQcrxkDFZhGfxUy63m57N75+bmk
2u28gIz3LkZP6pjapxqTCH0ql6USQRsQAye4BM1cOQBQ/48kfpMgNsFrauZ3QauD
Sv2oCzwFzWEPt1AVWYkEMrSWZOG0vAfH6X6DfiM1soWQEwqXZMAnO5Zb9cFyZ3UN
OiH3MhSdH/b2TMehABEuXWcESeg4G7K4/lPuYOFMDJEqby3YSxUrWdZ9kBpoNGT5
eTLxfx2Ymv9RdxqkubQ3KCM2VAm70FxCsdt3gKI6aR2Q+wksG4E8ur9agjbNrfdu
V2pvhEPAyKPssIILDEo+hsvITH2HheJxCVsw0Ch/myjlOXkG5/bEKpIOlJyPhfSe
kEmEXnnIw/df2RUgOPKtu5S6QKjGlngiQpk7lzpVhSMWBlI2qDSVrJrzma1fDmNh
H9+A+vBrDwFnf5NUHf6mMQzxCWEegWZlPFtrMXqVx44WRieH8PO3pI7X+jvLNmuj
iCxipAxMwJQKKphuNAjMI07Hyf8zjzCo1bHqSqqpERqHN/EA85d/wQJnJOnK4me/
+aEhYubfU6vzFZaAKpji5NVYJm9RdEIiIGvqDkkPgnUZOu5Mbsohtg3ulkhRlfE8
XGZ1JeKSvbeKSj00CxonD/1cMU8rzpOh1VF9GkBJHAEseMGkNZY3hsIyCBwm+BjZ
jMP4mjpF33Ib+kHJnk9bYXh+c+dRk5JEXtAzfBdaEtiBc9s1b9jocyfeXbTwVd3O
CHaTIWZgu3Woo0oRm0qO3CdRk+XUa+Gh7upEquxwpdUHxQfKwFReanJhQQz7Gdpa
bRL+V2zz6Ih/xEvghHq0KwPJpsA5z3+CAZFjaj7W83Z9nVkYB9NQHZ6SlRp7gTPc
HS9D53mztDGIeHcqtmHiNy+ViLyaf3Gdvg8amDfcRcQ6YrLKRf5wA5puvLLOLuw3
c4dQC2H/WUmItO5/5ccnYz7Chht+0KH+pTtns9iBTOwrPORemJfhqZzRKIRSVNCf
HUgAyGRTt9JVkgsMtDmmRjqWcQnkyW/DOpbRpOCHcqhzmAWlIi13xp1Y0kVEt5Nh
gkUwxpsJ6GIb24xWhLiWOknFziMpxuND2pzg/EKZBDyIZdrC1+ekOgB4/7+iqxK9
fQyFj4viPjnLnKMGh0ebJd1f/atk3tUsrgBu7tbdowWC8Z7oqi5n6fpqO1eD538V
UUjAUohgcFWFXSopnhXD6fjJ7KkYDNylSpfny/7KgTqikefwX+swb8Es/eHfsl97
549eNJa3eJdcAnuZU6TIjNpVTQBEErxNtFhIv+x54fUQONK1U1ViJrEWelIMOxRR
p09NKG84h3SXv7AUZFwHOcGegZcHh2/fKW/tMyZX+aTmvub2oiO8/PeuBMxvi/Hd
9fH8pXbxlrmwUwe/Refn4QWe/B/aUw/UKFiKG5rz8I8Bby0gxQkRRAs50chclNwG
p3FyU9rknxGlLCecLU/wb6AVayQybjgKoLnLTSdK8xhoZiijVsmyXJpyTpl3jzSH
wamUvzhihkDe85flu1Jp/BjaR/fL0lNTZ8WiUjlfjJWp/qx7ElAJO0iMP2+jbZ1C
DqecfSifqrz6dwTWZH4RIRiGr8/F94h1rW/E94LVFYLiJHP1zEXxKziOWbFdPKNC
FajTgJuLuenY+n7Syx951jhXzt9UlDG7EpCgp/R6S1+5majI9csM8KbatwUhAInk
WasOU0AUCBKUCaFObzZvPdMx0UR5eGu3RNRsLQV820Dyuo2PX+0OHV6dzyBEHmpq
2pNYi2smuH1SvzS44D76FC8C5RtvWG0RhqI2EZUeW6cxjbNXfBGtEDXPyDZk3Ko/
uzzuGI2kVF2UAoUHuqpc3nEZDH3F5+WnuIeBDNsWSaA226ezgwtG50mGlYBUHLwn
voRpi9d1YEB4zDIEEIwn3oPkfcE+hEbgd8LEqdWb9LMKjxP7gKHlMA8/A8/W9p4N
29UxwXJsvIq1YCZW7LKXvVX1b8q5BuOLvuKV15XShYwY3k2zvubIR+cayKouFB2J
0naBWBqTC447T1gHZPgFz8s0MiIR96GQOSFSohTIr6LUdAdu4gK+xvVKX0jqfc07
Nw1500RYwjl170UhZwemTaWwUEX/OjWjXVxW9JiNnuwWWJcNfvetRohCSOIpcSUT
Eoc1pB36Trx16akQv/OliEAWcO8ebGm3uO8zDop0KdnZEnbnGLEqhJZuUxhOW98+
NuGxjjUGfjBw9KkWrBg6WIZ2WBNr99m3qrvfk5eFDgZgSwSXK399V45AKdBmJW+y
5ywxUW4nP0NPT+O8GylpIT92/zxJTf/+X+Tl9X1Yh0oZ4ZHqUMusJEI9SMBircw5
lVCsXCMzphQlyyIrBuFNrwcQg3NdANlTgQJSUmK8bnZRAb0+2YFXqqsFOf98J6W9
UZBR6IHOOhSD5uo+qBKDmVoQb8asrrq3VcFYXMlAJfuIiSOaO2DwhqcYEcKJqCPz
DpZMuvQuQJjcWZqhIbcE3NAs6oZJPxNLIqc6a6zA/klC7GRC0QpYjMreluIGNPop
1MzmCDEoxLTE+gaZF87gOr2YLVBn8etjrqRP3QPpObP9ofyNgXuW0M7i+UjA2cb1
NpkizslewC8WwfCdc8Uij/PXCkQ7+rLbipduxDDJtIpxlcaBuu0FyJFQQJnd8XB9
vBc46B2S2YfMEu/rr1SjupmlyOokUR1z/lIsSVuA5ywGJ3+ufduAvZDKqKQXT5tv
oZZqAifx2Dr0Yy11E7jzD6O1u3bNEW2QSnZWD60Jr+x8kc83MwxGgujCyfXoJbjH
R/Ro6AaMU8z5Ev6r5FEtjZDaIHy4qSsYFYJoNEKN+Sc5Q/A5FRLGAvXuE3xodtNK
ORpg07R0K5BOKI9Jn09dbgouuysfvJZ9ppKZIZwt3e0syeVmpUw1rBb64W7gbppI
lCjunuN7GJ71WQP0AyCsHlBDuZPmm6o8y2AAvUv7IS4L9BTLM4469c6hIm9AaYEs
uGiUIDsR8d1I2HMusECAM3hsT+Aw3e1egcc04QTlnPPSwFooPf8cAly2NmhbpOJ+
jPYOMMoSsDl//ijNA+zu5E1moCGcvSVaaV8LLkr5EfWm8ojkiICWR8p45PEMj3o8
hZaIVTPvk+1fZegyGrLCr01CQkNhwlWfBFCDLGytBBQLj83zOzHdkrJ0jcwq/cNt
lhfyIV3hrfbkYsFgasZhWX6gUHaHATbUOYEBXnTNLJi66EZbsC5uBe5IPJ+6PW9r
lZwSt4UROe5QAjHPr11g6QEKkdb1Hy+k1JuBbMU3kLM1TjO/K30qT8+On9rm+5Q6
twFv/kAPyq8g+XXDB61jkfYHoz0W863iJJuquyFJqmOSxk45hbAz+F0ly+TfqEji
TJD4+gnuP8zjBD1UvLT7Ps+jbErZDw9RiEHKKF0eWxPSET8wjDTq/kp/wLOR2ePU
CvmnZnplDi0S+3A/O2cOU1Von+iPf5K/WIAUIuXwQugB/9arBmISv+I0CsdSFjBa
cSrmuxP7O8CdPuCdr+qIfEOOLTKAUmEXhvxF63OG4fvVbZnkQyUnYf2o/YfaM9BZ
mcmmu7UEy4KBbjUtwyUZlRqnuL4JCLNMvw45LKgG2crd6b8BY9LVW/HK/SjyCG2p
PH6AHuJJmLCdr1jIIUrMNWLEj7xMl+OSsi8itQcLG5OUhUd7uTdHd+jxQki4rzF5
NiEjexwhkdBVaW58UbMWwDACu07CZPRhY6xgPu3ybroNLGdgabfxgFzPjEKXeoJG
5mYIw6tPHGkb7Tr/EFLYG/hCUhtgCXrDhq4+BDhwptsusbmDCddkvWsaIHkJAESR
PMVQvK5p0by7OB9ww8Gsb5NEz/b5gLli2jzg7NaTKTir/8hMF+LNsmHzQ1q89Cxb
yh9QUQH6+JSdGMTTLou7geohWYiOpNOe8RDsXbfbgQBY0g7Y4yBnRs7ZmTJoqkyj
EgJLNo8h7/O+SaGN5773CoiRhr+rIGrw6Q+pUjvgoi5P+YWGmBNMuiSv0Mievp8/
Wzvzf9d1VFY/e3PD/PPzCOWkoeGYurkN9I4WClKeyfnvEI+FDOlWQb+QKkrjWlqi
Et9RaxAIYCN2q6dr698LU3y9EgnUEa4o+52rkXMtsjieplY/mnjoZYVF3EL48zbh
e7mI3N4WUWEbOb2D/i7v6jegBGbCxPLzhhhLzua4cmt8QlsAuXXPXKbqZIxHynso
/V8U2ajgDgv9OQIAcoTnDzQQADLIoYc2e9wn/lUIdPXi4jWklQRAeyBR/7TJe+gj
4kWo6s0Yh0kGXkkQVRMe2PzfZ9EfeTU5nCgeF4DWzmI/kPQbIgT7nCKPmbkBF/lz
KuSCwS4cuf3VhjK66uxcNsJy4+1gTKk+DBytCqqMb6PVH0IgatYKOWrc2NV+SCk8
wZNyWy7kWPGuU2gzdt2rBd+Zaw/dJ1H6y9R4aUwi+Uv9Gpe9IRyUjandxiCy6M2Q
0sXhcc3Mv1qAr/HKsr+8AWIj5fN90U06L1YASeipksxDXAqTJPrpHPeiq50W8nhk
YdaaIMvQC7kU+/9dmhyh7CB0ENlKqZ765KWyaBugMeEHcLQxPMkTUoZ0doqQzOe9
QrnpCc1Lgf9GwdtBt1fNKVDfUHZYxPqlrH9xVCeNy1U02/v8s+RQ5LbK/17xLfft
4cyg4DIsLXt40GOJuNaFJnWQOG890Uu+IRkip1+YOIAcB2bDMc7x9kD46tq7LIbw
l0qV+3LOOsHNDJ0gsjpzGWKIxy44FMnUdEQB6BY7gUiUMAP6Q5XfPtt5a0iQZgDK
4RrJaR8WW58AnUgr0whZhLiuYDLhFEihzff/3+a0Srl5nkW2/4LPCd9nhhOQ0EoL
H4cc8HRa+M4alI/MPRNxAM/MJI+rbtpo73N6pU7IcIbpRSi/uIi/TKPtBr9TgcZt
aehF1pWF3D3OzdzhiJu1KxuuVD4a23PL9P+GUisA7t0zoURE+ak9mB3cgLak7Dqy
J+XA6habzKBg0MfQTic+1yCee8Um7Vhd1Qu2mmx/usaENI1w0ggu3zAO3I3xAeIh
8qRfD6e0q7WNxOeFALjD6uALcgdDiYEVkom868IBUI8+4lBYGo4AkxdrOvNtgDpR
bBf+fgdMT38OEHo+tqkSy76XDpoccZU2yb7M4L+zO58VByjc7mbID+HSecR0jdQr
W79yYOPmCtYWXAqG2ayVKL9kh/a8bYp/5LuFaK2+GCKmwSYF+CwN6IFQi4D3bCiC
2QZpe+zEB4IUxrdSKORgw8otXAheQfnXntXabdGy3/TtpXYtZ+cybNXF6hu4x6rJ
z/RvCY78g6E+D9UQpusGfsmz20lKKYTWIHkgHdKyUWMqMkngbZp3XT4ZOFeHr1wg
mFTHHhLlD92ptIKqqT+ttKE5bJvYJ9FdUOqlIUmJDmeiHMp3gfbaF3d/NzKcRYmb
d+wFXUxrVYqdOMV2x9tuf7Qx2mEmF53M8DYP4+u3XlOdtOS09Jz4lR2ImGZIAi5F
KCB4B2MKYRk4C9mpoeXA3WPxEl0VYyLU4rQZQWOZbj+u5qidJNc0HPDmlVIMCpwW
da/DtGPO7vZRAI1JEQDNyRYqWPSo6EABUtBXYAqPdiiZZvKe8A8usPbD1GIxdv5F
t9eSw8QjAG7L8ShMtmq/P5jdrHiS9RdAVIjPGd0s9BkpQiJAwggRy8CQFKpTMSj+
xK0R0bjGvx4HyaZsB/q+e918HUCC1DJ6+bJYOcCgmPtbjkODjKp4KSx/KjSZitW7
jhZe2CmTZmfTtSMU0DN1+c5W9Uy21KbWuSXaJMpBDZQwfW6qVKwVtfzlNgvHyMzX
Rf37GYPB1Z7ENdWHKTFRX7KNIK0NusU2zZwiONjkFO1KCUL0qBN//v7a938Lyz9V
NGS+UGHOQX0f+dZqpmeiwsDaMwIUKcl0GCz1SxqVyWmevgsjZbMoHfXGWdfMsP7T
WnhHR28h8t/nY6Jxf62+yXZXAMYSKBAZ3XgUcZnl80N/M0hv5uId60V7jjZe0q29
aP7PfdwN5XXQw5fJgyw1xuvcCKNILhTYCuIyjp+S1K5i08sbGJmcDadYh+oZdDwA
rMOEQc120e6VnesICUWCPlINunthyFMxBp17PW92L+779MQpk5z6X6G9v7DM2qcT
UYUOTZw0ydVCD9aN66rmDkysYtw3oC/mzT/1PRWV07XWEXx7AAiP8lKTaAaegZeu
PC3eEEZliZ39th2BZK2xclyhscIrQdqkqkarXxQrzDlrcTBqkXPE+2DTQf/A31Ue
d4a3PknhtzMLnPcDzsdnsH1EeApiEaZjeTZTrMtioBD/qHZ2+223bB3Cq2+Kkdp1
vU+sGBhvBEzQX8ttW1IRLkA65uVplswi4ZrtaMPxHA5u6uW4loADC0oG6LJk9eVi
JEm+ARHCqfKoddbGio84rBbBgDtR2IsMzq8PX5Du47Ei3YpOBg5zo4Cvc85yMJ+0
TXirPjcBhiuTzcnD/q0NsIAq+sDi45mwCH0gAxb7yFR1rK3jh1E6AY2NgvMdjpi4
sxDYl+QUvAgtFdETocNH6Iw/IevTKkdaLI82Dy1HLVmWOa4ymUU4QBleqLj98QIi
COTxuNjuiKPVu07vW8byAo0jghnr+r3bpI6e+LfVtgdnh9O1Wqc24Om9eZnVMMC3
x76sL2ZG6jeLRFbCm/6T/IDZwikjoDQTbzk1aGAhnaRBrBTGRzpas4zvQjE07uph
nO/Id7Y5XilMPXJCCLzQbH/VpopKc20ngFzzyknmv32dGN4Spgh7pLRNgpinFWts
28OPcXY6KX4RdxsmvA7nqAQnjXVUDJ+rjl9XV6sRw2XlNmA3H6CPreFYJUQVlXcx
VxmqE9kZZkzUWhxr+eVefy9UbENKGnYsFRRkQJbjP7ZbqShVlmMephf0FdtvAVXR
qBYSzcRAo0pPG5bjQF6yCMIpa5w0TvjL8qZaol4C4V1MdWLyld3qGFrHO8sq1C6O
Aw81RbeWTK+km/zWF3ou/8bfSSD4KaxdqwaJ1Gq7Ldy+B1aWio9JO+RJG2ikqiMa
lsgusN6WmNwDZq+KYcqtNxyCtgyzliO4J+813jB614jGYl63f2quBB3mANxr2gT1
ksvobUd/zfMrajAwwYgPg8HR00C7d4lXgBjOyOuCaTcIymPg1GwhK/IypvE0BU5f
MNjGvXSgbsKt2jtnGPmDD0QTygQm8nk2s0D0mmMZkXJi2gDxkYBCOeigxUhK+l+T
3ezzFCo8KoeV7KMe8IaXWlLhujYCiYcSrJyfg1y+R2DyzK9kD29CbLvEp0rRG7iS
ztw7W6chddFITwlhtfbwLKJ8OsgKEC9CrQhNSqncl2VkpP2j9qbvKqXtvNrWOiKY
geA6A+dZ5wmWC06CZr5K2G4AuaG4DNjxbq1NKSaOne5RbVFsaOivucApfdiVpNo5
CglSmNsszETeS518FBWASZ/nmCoTutB0y1f3shTuu2TRmSa9PKer3h45jAnoNHty
DO9zS45i+P4VVZvdBEmR9Sf1QUV+j5VjaCh0zGWkwH8yNma5nLQUvtK2PpaY45BE
aSZ3QMaGaa/7xtuYNLIbi0N5inCvaBXJpoI2mlCy2GTz4OQvSzLFL2bcX/njzBOI
qIS4sFtC8q5FTkmd7LuU1mRiS80yp0FnjjM80BkBZBmbzPgPBoQjV5+6o0kcE0s1
BuDx8xIgtdhKMM/nhGHi0RbUmBxYoAbP63rIlWgPruOWR1T4anZk+MJT0zHw/pnH
XqoBWCrNS6rNYl+DIMgIH0jolM5avp830Z2YsUiLrCTUzrFMCh1XKru9dP5MOrtX
b9VYdQPibMuS/AAL4fzTVsFPRvEm+5ldK5i3sMWqN/JzXZy+TEqQ5cYYJNXCf6n0
vvqQeAsNJ2zKR2iIbBFmbft4XXSdLvNCrJiNdhpCi+EvqayPjcJO+oAcNzpMmAcc
CV1fGOiPAgq5xqgNOyv3Tg7EcJaKF5gma0WOFaCU8glFDVq0HpwgtuBwbCu68oCk
2M3ZFHdEIHD8ZkZgoi5shVXsjLu3lUwwKwbWO12Wv4J1kCbrlQnx12+qclVIY2qe
BbouCAsBotBZyN9Y5tS4H1UnhmGL6bEI4DQ0NBBKCT19rxk3QjFhCDjBLB9Sbo3m
T7ZPnGOKwNQwNfb9K/mRhFhT6m3qhdVsbOlqtJvVvZ01VrLfiEpNpwBKv5q+90Yh
f/TLkdHf3j8BXfZnfHxBDlc8RU34M7vhc2MeGwyVX9X9SysySU38OChB+fXAcHiw
uQZPx9JRQiz/GsbNe4lEv0wGHSeX93QeaiW76b1vbDWh9YDhY47sSbgs6RaAuPKO
l9+FJZ/6XC45d2SHlz9zmKK+mavHykrJiQrgIiE8yJkDcHDGLRy/XBHcs9Wo7B5u
6iKIrmFVsFi8h89+oTN300DLvSJF/V9ppfo1QVDWkFsMcewGYoEYtkjlzhzstkPL
LmPwVZdVijm9tT1C5AKPzGr2ucdpuoZ1pZOIoNgnldPbeoSuC621MQ1Xez7T25HI
GUXUsWqUPX6DwOPq1fHkh4NMeHmCK+q6KxR79I9QWsla0CDnIIEh6u2vHbM2G3oe
bDQ2DMoS/Fs7UMa9g+GTFlaUxmuNXWpN0/LwZa65qiHF/j7T+xHaorBrOCZmxsZC
iVKSoJVc6ZCyWAfhG9I59+EXfJNEQFWo3Vc1RRSFFX16OGY4dE/Mv6wSLWIDp+Ig
2/bNwMubL3rcU7GjbIiuNl6HQ5huaPmD6F0ZgF5+spkWGBDp5h3gCU6HkiH19m9t
y1Rt6Rg7J1LO/kDjrEzOEreFoQ0JFoZAH0dQ0jlOF2xgjlTYoHAcwsjdkaPydvnn
benN9RDXN4fOHmvNhMRaVBIb3zeRLAo9lhICddii3HfdnRpdQMmYc/1y3s2650Fa
d2ojwyAQO0PK2pJpi4TmxVH9JVQ8NkYWdWmDikB0phsjIQKhQIwmrcgh8nLm6L7H
vBxoutM4tfb2IywcpkMV2Dm0mqukAGk14q5DzKzMCh2qyftr3IHvjzIRIkeyD+e8
OsDAMJeOGnc2wko44n57zfuO+EnL5Cw8xQQdUBM2pzXOK9InQSlRUXqEYx4qCWYL
9hrNK+jwfyZZgVTNu7941TATQMYoaQJcPugSXi/l+laoCN9SUMhPyDi2m2DtRL10
rB0tIyDe7hE+QQqj06VISpZEsFs+FymOLQieOjyN+nDW44zdJJ6wRi6P/G1QRYs6
XX0pCzpfn+v7ZUSerIBl2LFTDLXuz8QwH7Wk71uF2NkZZDNgFp5l1gYK5AkmFC6F
ylG3BuQIoUDrzWqThpKLS1QdSJ9RBoSqyGJFpV1IfiEjdb5WE0/gx3eSjrbG46yo
m0hZwQRVEcfYwUw3nV/XAgDVfAnWgK0HkGF75XlawWHaxL2DcrUBRTw0DUk3q4wC
X/8P1IR2kiOXnvj8EAGDgn/LCNkpiQW1Z7KRsolMosI4yPrS2wnyMBhHPBWu46g1
EqVFin5hi0wBYkOZaSR+/mx9+5fhMqrBVYXr1V2VL8i2r4wwCpOXzhogfG1kHMm6
nMUA6Ll4OZ6HLBNigaMuKUtzXJtxFIyqBwAi6ja1p0LwM41M+46xqLZ3fUvNSU1p
4epfWnQ4K0JRcgDhxCtNe8zTii2pmC82AbghMhXoqhHvkid1BYUbj9R90kSuhblf
PWyb2NBweDB1PwalXzVyKVPvyqYMB7xlsVIZVdvzq4t2bAiNTlq7ZOZn1rx00tbl
oe9z/OpcUYrLxVnhVGNnA1dKo/mfUJj+it5GrIKt+fk+HARUyVobe0+F8fhBQp07
qgdyGapXYcKxHsb9ZMtMuMx/IBs5WaFdDPYImaICSiZWbHDKPfihS9bptprvkaVY
vF5a45UgufwTAXK/8lSnmByyxI8ROu6g0GjdLXtL0ag0+CnfTYQfahFxn+DVNvW+
PN2zbjzcZoMq7qDgZPZJYG/U313gYtfABuXknPxMkQ8/KABGZ2Fs/e9ce3keDvo9
MaxYozFp9TrtSaCjOvaKfNeiw9GzonzP9wvzilz8yfvgpDTfJwYX80weHxV9xEY4
AX7L100GSTxGH+VmFiLeV5tdwbtu7qdVsmNLCEWqfRYFjKKCEQHArHVeF+u+CEqG
4MS2k5BYuzmpdL3cZEOMqxQ3U1lAlp/wk3+ed6217OTSK9l6D9XkDSxYrkuGEX6a
FZsj92seih254oTSubQSsEzAHrGg3Qogjdjiw8B75dZQDeZHtm9TwwOX3YTqF8/Y
Vtlx9HFo+JUswI8eZyxdQmVh8Xj/eSbwUwrHDmvCdkc5CtTMKy8qRXDV3UxruBYf
pVaRznh3XLW8AYtQ8jFydm6tzoUqnVFw3yOyyOusLOWc9HO42eOIPx0GKyjZQnf7
WqiOlJGrvPqJls5aP3jjqWzlBQdgsLD2h9om0v3ZrcWX+a0djV7DE4kTIXfkqRY+
cTTXTv+9CSuGl0vd20FyYjvyxKLSyUhI4FK1C8BaVbwm+JQW8GhqG7Ji8g58ZoP2
m2lbYV6iCF6CXjtwoQAZS2Dfh9/Bd7li4/dIJVwVVleHu5dTjxwAjUOSySEwsrXX
+sOCKJOsz89Tgcr6lj+kLAm96/djAvGfQPHeRt8nTYGC9PnTUIb2kCoj3CpiuDPi
c+HLPXEHBT6b/EAZ4Xfg5CIekpMGnLuOO7GwzEUoHik+cJ9BGCS9PusP1LoPFtUk
gpM4KGZ9cOyz/nbSs69qqZeRh2YGnP4iVlgKXsumWF23Pe7atQUcuoFoRSBMguEU
k6+O48YtPY8iPTbyqOShX0fRH57AidHzP/+tlDt+qHIcuz8HXRyakAjs4CU4SLcy
/NDfeeG6dQUzubeqxZAvtoANWTBpnLgif7fBy8Wp4qmMCKdk4D6Bkam5jkuIuS+X
euzIEizx7nI5AT0xs7mxucE3IRWA3Z/MtOOzFINXZbAHKZg5G0Pm3a21drc2vKG1
21iLJC2TjWWsmu1972ulrVgCKQ1bj8DlySilEp+P5TBa6Pfu6oALgytR6cpwYEz7
rkJPn+nTtDXzQB93hsxmvGSsu0bjDZpxLCuXLfsPksPYokt6tnHbiec8E6HQoplG
JWex3ZyN2Ywhd2+xTVPEZRxxyCgm76q3dJfrwc5kcAUTab8Z46b5VGGgmKFRAM/s
u5TUGk5uf6exGG4G5DGnEt8Ms+rh24q0uvnp7eRB40snNZQ1oZE9IM+4H4uRqy40
p9YPpwH6ktekwcadMcWxwwOSKBbTsvxXK4CXrbrxowUOhzrwK0k+bW2z+2KO46uP
E8h9lEux/hgRkYQRhj3n/vVpfU74t/4b4ad8JsnI7aS2IpP1vbOycTTAJ+ivAMvl
If1HBaH7Wv7ksr/f1HBtFp9IzDDwBItRuH/R4vJFlv1yr4tdKcxAhnzdZ4+hBVG6
AjtWGiLXUmeBIMh99i6GCg==
--pragma protect end_data_block
--pragma protect digest_block
PhX0whUHmarT3JNdO6DVz8VdQYs=
--pragma protect end_digest_block
--pragma protect end_protected
