-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Jt9Pe6zO5G/KmICbmrWuL2L9WqOYEFTnYIHtWedEm2TZicfxRMlLaY2P5QFWoBp4
GjwQEDakQ6PA+IqKICofLdmMCGIJ8WFHJBRP903pbrgL8XbbUceG8MKfFha1qx4y
he/VzB6GQQAw+ZLvjzgyQm3P2Qf1vlUErFkW0LPyw1PJ4SseUmKA1A==
--pragma protect end_key_block
--pragma protect digest_block
j0XJ3uJvZL43kPmFYlgP6Thug+E=
--pragma protect end_digest_block
--pragma protect data_block
18j35sSdwo9vRum6ARHbImyqaMz97qakFfIMVXxDPgmJPqzEALBGnSLYnicqgvJa
NI8Iq84u7PNYPe8iVU2tMSKa1bJXCghRbe15nKDaJLNv7h1pb8wC45nBCnoJsw91
rYdx3b68W8UCDvhVBldYI7Rw2UzQJv+WkdfGZqRYK+69RGy6aQlBjfwTkUftQAZv
VUjqf5046tisZs2jeWhLGJQM/61512Xv865Rxq6EUXPFVAG3XIYNka2vfkydsxPa
WnNbAkanNBHzQ9dldmGZQnTLiUyfMLPl5Vm3CyhlVsKiy5oREDNjDXfqI6Gm9Zn1
5BD1AeEOJqq5Ns9094zk7A9RONcIYso/BNTIpk3Ic2Sjt2VgcyjMdk1Fzm9Sb7z4
8cuVGocwbQEv/zLOlMZhW6wqn1J7ZEBm7in4lSRCjiwLWjIPgAASI6C2Lyzb0kO9
cMv6vNwQdJ2oXfjtkEOc+q0+SxXp0KF6DsJO9eZaRxigSBltT8LUxWKMDW05vR7E
3nz2cp+DgVY1DmMTn+EgAzGa0RuQjAy+gR4bhBtk9fc1rG04cF/wHBPGqkBkiKY3
YoZuBeZFA4GOb7pAlG0Fpovm0On1CIhEwSqQIdR0YGNRLWPgZMpymF/8N/hhuPSO
8R3leV6ymsAtCeNG23fBeg+cISWHEW7e+k8E2KcvCtHpEASqZ14yhEch7pHCalOT
JiTxweYz/aLvWU+rWYjaM7dSSmfwU8MN2aQIFT4Qinhw7ZUzTzKFlO6v5P74yQOX
wke3E5+ozTSs+rY03mfrAifZtW2qja0xoh6m5GUZwJ250TDQ+G1O2rnVAUoB4FbC
3u3ltsr/8Mp9RvzM6p0z5CPjoMr68o75Xw4EQwZJgVt9mT/IlSIyPKYuT0UiZYmu
d7LXzfY2/wbmK9mv0x28ZSbxsTc03TZtzDwcI/UAan3xn0jOOxfX2JtMRrE7DLZp
T0ME3JQhYTXq5kwQkdomNd4aAeFHWZoTBEqA/UVHnAS8qaECXOOVWG1hIdgsZXBJ
nLW1j/rgsdT41fLUAzIrSFxEThZmF6raufBi3iam/nq356ZcU9n6+UtQcFSaNbsZ
TDMILvy3RyW/6v/jILlDwltlmzledOLBNi/M9Hse46oPMnZ+qyr5w2w20C+9DhHW
xG27TDK9rkJ+cVBo6R/8WjUlfPX03gvuKQENAHvTLgZ9I4sFt/XXGCPYamFb/eRp
xtdxMlM2eJci1FGl3n7gnH3hoP2o8SgwwV/T8Mnb1eBz6mYu3UaO58/cbbmT5jFa
9mOG0dPgeDopvhL4Xs34HRTMj1Qbblze+YeGPqyynJkLLLQEMZxXk/fEZezB7nYs
ezVZb7+U9zO3MfWeataaDYvSkpd0HnX6FfvMcgRfiyKjXjsEQepe+u+k5S1jRN79
eXjT57WSHElg6E8hQZud2NAJ0+yyK4CyVfmCDx9RERoaXM4W3rgH42kCrAhoiA6c
jzLuAFt1siBPjYdyksQbSfVnB02mlLuQXUL14gS3DnPvPdJmuxM5uYjbrYOUYI2y
UruDzGKVYl+10rL93RHZzWOvLtw32IljaM7fgFRU5mXM/ufFfr+LYoDAocdBCkiU
ybcUTDeD/oeH0Qj1gBaVRXG1bTSa+GBm7kKUwojOgk4JZ1YOQ1HTDLxonM2rQrz/
0uF006QmY3PIZthZsBR1XwQAKs5NfXT9HBDZhePFmqXRTSUq2LCl0GsGGt28P50+
ATYFqvWYcj42hYlaGwHP5mM++A44KO4I7rF5h1Dd7VvrdigLVB6u7thKCPn7SrAF
x9GAQMrMLv0P4FSaUWBn1O0Sj7sVyommcsLhYGXXaBTGBl+qX905Y+QOcWtv7jxE
6No1s9DuGtEPXyz6FfJTCUoNqR0eQq97+PHhg32NeMN2PhpLjQ+TQZWmXtfgnRiv
YWcuqJX4UwOzkHnrFVN955M4jytRhYtR4wPqRlztNpraktjovxhe9QTU3y4skbkH
ZMfLt4FyNG/qzovmWzi34SbyMie/hbDJBUpN1gbjvfFWOD3ItcyIFuWxFgkS5ZVu
V7aTk5+0/550arPrUhEctuAGNpWxDFFPcsKhrLO+AjXw9jlMA9pt8xMu7wewqQEc
3TpxdGMpD7seOxR7EgHNvPqj24NJikO0iSHvDrUk0EzNceoa3iDT0TW1/Qpjv+UR
gnGLtBTkFeR3Rn9krO5G6P3liQEJBygO+usv7iAuKjNGg5w5BU4sBl+tUXq7jv39
AIHNMo481nY/kcOIKD//szxAEmwZB1URV7kdEtebhiAL/nM6QvWDqoX18tYzfIh8
acbphiip4R5JAy8WFVTeRRnvpkizbb309PwQxhmQfRy6+WtBTGkSGtiaD11cmFQF
MHTkC6GnIMTxjt3CTlw0y2u4bm173w79J9oowW6IUAu31yas3ifMdEH4oHzwpJpO
PDJWIXQofSAzSre/T87W7fkLHAAJNGafiYjEF0zvTMk8FAqDUv5Z4VSKri6IF+ox
NJwAhug9gBVRLpmmp25DtE+94gUgrZCiglV1WhFRViyRUg5xfPkVUcjzOAOclVeK
hgRL5M2SaYiaCOz4uTlzNRhdk+W557wu5mJioEwKgeLaIAVPJP32L9I0ipX+A0x3
UXHawlvPokfRp/wSJZMIPf0EqPi6INWoC0tN/fKp9Ho4wm04WcSn09n/q02pmhhE
Xo4lq1Jd6aQtBB5j2t3NlIOwxbi4NyrCbXETWOMu+E5czDFQReieZLYq8drC3iuP
T3KMwHZd6ywJgnWiFJYG4JVAyzct8gYowdFFRiJWtqhTAT0daqcYxMDUTcRniLnJ
89ho0G0wHD71d4bah58zqkNB08o/2elMGWPIMKC2KXOEy4r6mBxNDeIuvejV1QfG
gkrxQZjHAthvWyz1tBLwhdr69IcGLat7ECXQournBgdoe3J3C2OlJZj5hZeG7jka
159E0aH++6wAkUvPGH+65Pb5cOge/TYngBaLx4KmirfZ4W3GoJ4P+BzthegjcOF3
pgp8CV6h5KRE89BgjWnH50X4uGU/ptRoRgFa54V+h0vsu3AaxKDWNN6YjycwsM/T
QrKNsU4i97zP6b0NmDhNNAPtQrT2ipQj6lx1KTlNF9toJRxuSzFj+PzG/vQVp13I
PsZrvFAyttYWZsbDMHpNeSsqMHE8kajAhdBDc+obnJh+5XZHAdwvPTw8tZvb5BH3
HAFtX0aFpPiWDurTtnpd4lMXnaVm9otrAcQ0KCe1J/cq5vZcjp3EuXQDZMC4CaAC
LVv/S+kmA+yv/DFBexLF9qTSwNFKIdnUMdeHhp1phAZol6TDIxTtFP/w0HaPppTC
MQi89IKoxoCmEb7azRBXRrxb5RfBYrNyXXA61z8fA3n5uB5QU0dTfdAb7Z/rupfa
yLAxx6HliX1BGyYri6DrGooFPY+v/7D7Z0U/cnp8x8VkCrzBkvufhMDVHOvvhW5K
zj3kCev9l/m+L5wQoXvKHgTZefoEWezbVHrQsToblroQK/UE8cXmN7efqwTeINys
ZnOpo8mMCsV0NHWAHnnRjRg42Hrh6iEHaBG2Kz8w4w6zE0axJow8/Z/8h5d1/Vyd
V+LFS/KCV7/1hXmcZ+y18NHSqK+pyWSINlm8ddzQSX6zh+m9PENs5WBiV0LBGMLF
ZBj/OLR8EDOU1fkhheJkjTFmd39P64bLhIG0zwkGRsPdg0bnLDKCKZ1N6Tf1Boqc
K5e0ko5wiH8J8U2vVLQwLMZBeN4Vp7g2tDlXJXSw+nPGagK8GvCUioUbx/K3xJfe
agXqQCQF1HOq0ky6MrF8p4Cvztrrr4eZKOLCqe1rwFTqe1w0u3JrGwPcwsQ9B9cD
oyPxaQRPrQst+SdELM8FecOdcVkRnMUwYExrrebU9RUmEE4AsaIFA+G3eNdZYS53
NPICcYBxW60hGdMRxAI5JJYlIQLYXiO3pGySdaIqe7Ts7uK3+gM/2nv7j8E5Wy4U
hnd17Dzj7Vli4yKbiCFvt1pqsXOFUNnkjY61ESK2dYyzMgRksy2TgQlqHCdM+uPL
gJu6/G2jbNh0zzv9am0VkrP33jyYjQsc+NHShfVrpafmKCpT4vbaVIy66pdpiyJT
bjNmcvtOxoSVHppozfY3FdnaXndAy7c3jZa0I7PYU5jIkC8kQH+ZkDG4POEffYAQ
0jx1X/GneTiL4luAlLTeg8GGZw4D4F+MNwE/SzVCOAp+Dpj6K3r3i+UULzMK2Vc/
5wwTxclfAgljkWPW4zsgW6roiFmtH6dlBTIhOYnmkOriR6801AgSs2fFr2sXfZL1
E09xH11LbVIwiO4uyn0tsLGfPd4EutCcyEc8Xz/bAJQ21AVHTTvkMXXQ1Ivh6pzZ
J/Cu+qeaEmgPlZV8mQvovmnxxWwCqiesr5QvqFKdap4dhk5vKKQsvIwBmZSZU1Mn
0zG2h9hMPA/0l2eACZ+XVylZVff5tWQbZEAZqi7BtDt1goQY4GSVKmyHvQgtYa9W
vXZq8ZTv1i6nGsPZw14N4t9at42xzOnd1fSNMba6IBWcEry35II+WwYRBR9AUIGi
HfMMYlyvp88U1pLV/lxwni/bA7udNLvnRrD8vm9yqt9K5aM7EMYC7poUsa/fp1NA
PNx6mUJGmX7OLTdB0wTDQhZFu8EIQWxgx1zTcqvDJUtdQGPxkINM2NdgP2HTPKk0
qFJTu/IEUhTXfzQwrrcXiC9Gif8/51IyRnXMtlA+R0EbLFRKMpU9NqR7Mojwgfak
LPobqE8YOOUAqGMPsEhUjooaQQS9zQEUmfR2pYeNExqJqj1dxD88ZbzmfhFwkMyv
6FEAMtTUruqxz2hEJeK0C/L3HQfuvvrRQ9221AMGBwxHpSWTRymejVlyc6W8ufqS
y9U7oER1FY4AD0WcKF3eFD9whVot/+l42yUPxix5lZYQ8nXj3/pUTCPdgUvU5Zp2
lDWzFCztT9zwaVIkqtx+xn2PDLpoBmcRfSdU1PVksC6VxLDLxk9dp4uaKrN2ET8G
mc5rSIyqNuaw9zgnkQDsznd9r/uN/cZ1Pm+xV5tibwO+yEDAYTEzVvmEXcs7InVQ
HNQfADR3Ouu76tyPaFrgDpQDg/BOt69/z/n9uPxQJ2nDNIR3cZcfFWRf0fEAoQS2
MpD/b8VkBM35E8DY6sHzzaVqRVfMnAOuRalpxPEkDYQT7VWQxOJa3DtghSu98hWI
rL+oQSPz67YIJOefHw1dzVVsztAtAPybIJE8lUbQf24ggbpmI+uZnlSuFZs4HyhB
fb+J9fr0YsK3mgBAX24laZEaXL+bCgXxUcoViGYc3XsOfZNxhGnxALwBpIPVVqx+
vdY91adwFyoKhv4QBxXwZyiimTNKJeWGfg67ffXuzl8ulzLE92NWuio7v2hQ8Yd5
vBEuGtuBa12PoVxrARyw1yCyem/iOYphz1aueArYnoAvgsQycMX3n4ZQ583+thox
GEPng/LM/9EoMiahBZkepq5tZHTluZdvgCmWZe+eDw4Q9FLmgWADqJSGOrmWDExk
jS9EGJvt0mdv1uKxdddliiUUN9zt2qMiZuFrk2Yw8Z4du36DwezE/pITS8A0Q4xk
CFgx5buSelIeB1CdCquaUgiAe+r6BbuiFsFnfPXieAEiV3RwpqDqqRgudCtWEeIU
VxpQgY9btWpzWj8qvuhWGvnXMA9BtkOa/9NX87KE70vSw31I26pG+ZX763hJsHD2
r3VijLwW6C4cASQu9Urv/uQxx8Z9H9HOQkLiQo5qPpKWpb3r7RjT18ELmmxDkeZk
GLBnqPrhjArTntJzOEuHJDg2va400CvOZU3rxnNjRCLYrS4Pkb8v5Obfyhja9GC7
BL+PhkdAd5MObmQsPs3mrwW9Oa90WAYznqGVnmdli3rPIA6XGxXiDcIrPhCKdIz0
ecFlPn2g/WSoLufd0KM9oS9IOHhNeKmnkWbqXJhQLALfMfZ9vWXNO3WOpzaAQ/bC
qsqAXuj0q00hPcstu7+5OuJmZMGWoCTV4wZNrLYtgu+lfPOjICSPUf+UUr9S+wDo
guMjehIOnYkiYl3rUWm9sEyt8BoEyVEFe2dTtkNd3EKP+a9cX6g8BmN86I9NY5Jx
gmDpA248Q9ztq1C75i3ND+bMOiC+HVuW6Wketm3o1h9aLVhZI+qptN1YSBrH5LoC
nXiepkq8v7clqm3vgo2YH1PVpyXe2kBuhQ/MH8/WEKwTzZy3uNCwZegMOJz8b6Cr
NXWgsB1VCKVfa6ZD6GgX89+4L6+/65bzjesxjJtJzqLgNN7mLMEitnIX3+vgKgxT
zIrVq42WOiot5TxMvm+FKdJwTJ7rZiYmDvYz0a4EDdQc9tlIqRo+WeGbu1r1p7gL
PPJEVlDqOgrCgcRthBgdEai+zegTrGdSSv/w97XOM83l0XhFu9f0xxykblzQ7iXW
7mcGhQv+3Oez4hkRQCkX/1a8bUSzgtqw0xfQ3gJWndN6WCZeYYx57AZK5S0PHocY
lYv5P921d0bSxR9+zSkLpAyTfcZqA9CysPghn9n+F75+tTS0XZyMg4tDKX2Hi0vP
g/jJD1Q7x/37xNUSeAFUBpTMCrbewXAq+H3ukaKaZASlzRoaORvPpBq3WCKdiaLk
F34bPJ79XsPUSELxCr6m3ig5IWKRJMuH/1GByCgSqQOXA+KmIFHkVChi0x9sakQZ
ctXhpIhLtQcL+iyIiue1XNoCsGmsQ3Wd4UgO6pVEWFBPXhKFrkvQk+9Aco3uB3aN
W+t8HYhCR0CRZR3/1qVCGXXSniTEoGVdDajj97pFHf1JEXPdTv5NUxczaflEeh7h
t8gzrzAB3myTttFjEyxO2aLd6CMCIS3whNkwEDZNWv2LSeON7GTihRbr1Yt8hk1t
ddefoY1ufP0UsXoTrGcV3j/s/ywTDr7ekJU8KjglE813tq2avS6vJsJSFyznyR3W
U3BpkUgVKJVhxgz3Q1zltJwWO7LkxB5LoB8oyRcK/xuSP829qUvsQpi1raLxryfs
mZDcuhLPCfqw7Bjj0SW81TkQdU0hcMw35pw1fsNrfmcjLWw/vcXyowo0PLejLoia
87xYLPB39J0tyD7QKut+Cl2MlGXx3AyQeaWP6nbC2MFcsJoZFM2I710BicCDL/DR
7Q/UhqkzOndDeyCHebUGj91x6MAn4nMv++I2doANy/w0w8khnNrvZbKhB7K7mqn8
r84C9yMfJEkR+TUhm1fDMkxM+LrJ9/fZNhSZD6yUrPuaLqbyHwgiCjWbwFwoWHd/
N0FMp6zjWobStYwYyxRxNSZyKKzO6gxymhtnQBbRZK58fzHy6mox2louK05f0cU7
GImT7Eh7OkiPeiscWJBUMbcHMc+Xsb/S9r+geeAlEFmgJhNjgfp0+mKjDCwEncDm
JLnnx38vxqUcvnB27qQVHloH1R12s1aUZKJCNfWdkIXCITLLRJb0+WsTFs/GGPhH
bHhSZE6HemiJgSWBD7NZN6XJrR1LRGTOh89uVEB5I4Fe8Ha9uTt3n4UO2ZzRvB00
fqs6gHiOw8wuIotvLE/wgCSQgb4bhOonBOfF7QaGqXmFa4EKzGq36A6+ZIFwEpNf
W0yd5Kx3KY8KZWBnPW+eDjbPw4odOet4j2pQMC7CRqLiywDabVkVJQil7v7KhMAu
EXI4UuF5ehGg/vjvZHzdQGWo87uFJgCuv98QkdNPiyaA0OQ8VNHun2zuqdUlg+ld
HdYBFhoWWOt6YvFbio8mbfn0sQ5Kawd0wR+ZbvIgzQz3Pu3v7zax4ufZHXa3FUJI
JifCLNq7TvHAKrwhwzBNNSdp1NH9EUh3F8tyvmakgSl57jUE4IhNgQbGY6q6jgqm
lfG5ucun0Rf82M+/cjQx4rKzsjZGNFOmyFzsORHyAPULlTiSi3S98A2vDSjdmjI0
MpckhFGiuuKruyDIi1a+wSupG/LzYkN44HmjCEhbxLyK5EToTxXUCDa1mbUG8EP8
9m4xsnUaYT+iVqC0xIj+BCEdMSNfibVAosqbJle1bpHQKDunPoLv8Fa6ukPrCbBM
kw0t1eBxXp+5j8tOWhH8FF++VE0ryq65VIERYrlbq/gps8ncAlne2W/iTbRI1hMX
khsocqED33YXzhyRUzQt/mnEjZPug+tyXNKPiUGFnaFtSLb+VCX3lUbv+r4rcqvI
wQCqDl2BPZuY8tql49TJ345DGnFAigbwhgv1N28jFDmVYTmSxPejtdzAzZdOWt4b
X8EIsvOgZ5vYll3TovETBk2FoBzVvuAshU1s1C4sPzuXx5nn+vjI6h3hfjX7b/b+
mquROVUQkNJCHuahdyJ+4+equhsjwdDr9lBmRqKvY57wLgNRh5T1T4J2YHXichje
HiCtOW3UYFp3E3bN8OdEsOdVBjz0LK9kcOIKFjex3+xsOcR8mhJxreVlvY3QapUP
/OxEice+QZWfBinFy3CBjW2vCQVsSIIowG+7PH8KHIaJJMOo0vMIAqHfk02Da6ny
I9bfaOk9WlQ1U21M6VCf190RW0acJw4J2AAvCNsGsYziZspsMV+bDJzFjx8wceA0
YeBXFjxuhZW0RgXlULTO3KPrNR0e7yXtcmSftO5SlC/on0+DN6Vs43NCGN91SUt2
cP4Pzj2zz8S6tzW7u+0o01GK0wKUZfMS1Yc4zpoAeL7jRAgQMn3YpDRP7BQPNtDC
oOfyXhsMGBK6fz3WXFYYA03fuXQmEehby5M6cTsP0lpDSVNKAaiva3BFQKS+kJ6N
FrrHBzicq5AE4XfNVkkiPTcEXX8M+19xDRozKKbu1okkypgzs4guWQJEWzIhGrnK
IswA1+LAe5hpWzN/2WGoxxs7feiv0PPxDGAQzxL5MktrVrfM1PRvjks1B7MR99+V
8OoUPmLt/chQL4dnos+UGV9XwZKRERukV91RrnFj5Cuq5aREgqHnsOYDzdv++9rI
VjvcmdzLfX3Gmlaw49k0oUTP7aaX0Vgen8A1N/MUvfjnL+B4GFCD60Hhplfk6gBj
Es9M/4TU8wF7qZA1nXLxEJuod7K6CaCfE3AL/4xHI0iw1FbuflIycN09edOE+Hf5
YJFxpEYSiQQDHd9VE06SneJ0Xidx3DGO5yO8LfwA830qJ8CkiCJ3WcKc8OsKCw7g
4haq1NLkIixVC2HmbsPUVum1qG/t8PZbstn4JZiMyO2+ayqKSs2WnvEE2ZBtAUlt
Qm9e9HKEhsNywFEvxrLQ5DbeqrcRqUPPonTq85rwI40WoWM5FLTbOfPwbHPkcZnh
qDhMP0bPBcQNBV7BHz5vFtpQ1fcp87WVkHfOWmAGY37Vf20/ayoAi+bN3bKKoCIm
4DkVZSoUrtNRNkUMUX937D/vEnv2M/xRLpCYImNvWdkooIxC4v59vX2n3eSAnhNJ
ojQbd3QXjarqYiNEq+gpq0lWJ2gbM4DCbb+oeplPPzoKNcvFPnlMLfgFgXRoszj3
DJD45jGoSwciLiYESkUEXtYyPCZtdDlZ4Qz5xfObzsW3sDpzyLeDvNt/LgvPlPAX
pG8VdhEa3q6EURFJmQxDhTcV5nh8oukd8x1gXS6Yj5pi5Kp7FhWkVgzHhdOlL21a
W0MxFqW2VD7iFHBfMmJXlZGtBXUreX/zth+4p9Ia48U8hZcb97QkTc37MpW8wmaB
lwbRsalrcYH72hUM9B8irN+ihtwYn10+gXTsJjDf/uhdO1obh25XWFPnxbY+mWXO
OA2dzFM1YGG3vD8jIPBSuQz7mmbcHEISb4YBbcgj+EUamsghyaJBvZamLaeQ93s4
kbQUSNHu8IpkzlAma9on5pfZY4+CR6tvy5U/vDlVy4+VLrCGghlT6qBHBiQiHfV5
A2zSUCKfV6L4L7X/cMXXRS4j+kN3qcLH5W21ELd+z7Rn2H/zZtO7aAKB/jtPv+yX
yxJRpITqbxKqCtGfjq2mvabH1VV8fbAuHpKxmC9x8VMxYtE3LuCbf146fMkzB4EE
FFKvBNdlKbWU3IqzZ0rceqpivQ6F153tFO4+CWc0Kug8uqd+UP1ocpMzgwtvFhHP
7S6e2jFDvPr4Q1DsYsEdpRTFd5hu0O/WNR4cHsMZP8ck0PAX+al1mA94czPjm6Dq
s7g64XP0F4wI3qSvi7ACGbDL1HZ9fN5u9Ht0Mp8JQMoipxZ1PKT8Ft5wDUeHo/lD
8GEa13DeVO8TLNenPRx2hqVzcq1q6Ptl4um+ezDo5z1BoFIu16VduLlr+cPsuKl3
ZovX3yrnMhFhoICGpZRQ+aBupVbKGet9woI53/DqCWiOvwUL9EdvD1SE0LhLRciu
U3kbCI9StA7Vf6gy99gx3xp//YgoGf1iGLBQTQDxEgjuGsVD5PsiIW6XC5W6KRY+
JAtsqhztTn7WwcG27mHtnn0fT5ty/YYfORoXyCo8cLTMHpiQZXT3XdCYxAjLLrp/
+9+Wdz1+pp6DfbGIsyJSXknF2JF8kU8hwVqhG8QY8z46+DpD/fDX2ir+QOUC9LKU
hXyItrh/riPmOyjtsZ3J4OAdtj5Ja9/0hR1vn7H0YgWwl+t9tsACfcFjyjdqluyb
Ik2I6j3hQNbU1JexGcEaw69I8NqPFzqOIjoneDJfc2md9bY5s/bwi6p5WqTxxS4T
Jkhoyg51ahP/7xq3IkHSicgxS4me+KazVEnIVLjjkcN8tM48Ja03Y/6YUmWTrhg/
N5rhUIn8bGH6oozx3xiNIktSh2CvJjjKK39eTKc2DrAFm9H/+noVhaxevnODC8XS
Mi7bLrVUnfnOmBt/lu3hXAz5QFuV1uERbyNV1TwkiITK34riNfEICCxrISyXHmOf
i7Ieqt74ay2BNELpXe3ZajOUL7w8qxFdO5as3kCxwTXAjFsHJSkK6Fpqi76relJN
5ARi/QIhSsrzhuocGXZuByNt3LpTTg6A7Z13F+03m6dWM8wPiZjlbErz6y8f1ksD
P9JdUs4NwWw2xKP29YS2FNmXCsHAe/zreDVffltHiU23RYNwle9ZA0WGijJUmI5l
5HDKiDbNg+KwK6y9S+qDBAEKDxHDelx04oiZhnTa4yCGoSxQ0DoVLmBtU0HjmuLX
oVMjBHg6Auwxlsb/54dTk3ac3mYEpfM0cKvqcpMDjIfGWrrfmU6glnw+wf06IiuQ
F9Arc2ogjBuk09lPPti+U0Jyi+JlO5sD1IHcSkBlDolbWnCOj/4LEKKoBm/3WtgP
noC+/+dvsjA+qkvxn8uxFUMUCh7XmT9U6GdByuqt39aNwCtkvFYMlItJaGD8BqxI
oPVtiBUhPeOZz8uyor04C2bDQFp+Uf0JZEDBj7WLTYsiMGwgTrG2MoesU9SeY3aX
61G7vERBY3wqxtolQWnLEfGCWfsUKG6C6l5Y8sr2V8PWbj2EUlfIis8ztHruyK8n
M2FpDJ5O8zCIQpGRbj6aa4CRNgh9rXI+x+CV3HQl6sHf8AbPs/GYhjlvAQw59y2x
aj4otcBR4AJxj6ilFvKmwdVYIbQbXlfIv3roNbzGL7JMsS+wW3QtzPTCsYjQQGw3
8oMEFxGkyQ6gm35w+QTdiQBWg12wdJO92rsldd3bCFXj2Barg7CQba2YdnaBNymJ
5NwWkQgIm6tMnSP5Goqbi/Hv8pjqXqSObjzv3/7mRomoW/Fx95ua3k49WeQRRLnx
HzCrBi6J7iZwil90T/k1C6D7uebDedPkfwvGr7V7LtPDmlKwvFBkKAwkRbIVRs5M
AakQV29rA0Rp73ru3ZuFNbMrm60lmHAx7lH0LpGgFwlZUELnhJs0MIFVAk0B3gyR
YAvB6ujJamGgIxZxSWjTW+tuW+l4XnW/AI+sX23yDigQdSgXx7e8TKHjBbHC4PFJ
NbjJGOtftEOvuccN1lFHP6lVk9hXgTLaOnMijuOGs6y4WIFE+aMc7BomRzE9H2WK
B8c8PCN0M68Kcjb9yjtliUNBDtRP3IGniFx0Q3Y3yDTkyVk2GkNoL7IJrBouUVfw
uBpoHO9hrMPOCKjcU+XqtRXUDKnGxfpEo+Z97mIkYV+hquPm/hlsRKg7kcqCd1lY
/EwQBGDPeMQcCLeMMU9N9m6sBUJNciJ+LyXI3Ud+sFiOa4m1bbMlZfTy+SKpIZx+
KabNZiJ7cfSstvCxX+EgY3FFUCsWzJ9ZOoZ9nR/AQNSOEnjsCW0+n7A9QVsPFFsv
sudLU+d2r/QDZwkDW4DPJTrFk2iTKo9W0hCAs3/ckdnyGxDAu/jBRaeH7DAoLxW5
ZPBXGRh++QkC2rTrXX699i+oZh7gmXH3cgc9DLbWarRGeXNTMaVwycejFBlr51vw
DY6Jxc5cap1knPXTF4ThMUgQdFKJx9jp/1CXbLhGDYOHRBky/TCZTJFq31b9uiA9
X8sT6hsp5qdWgO14dUGT9Mkq4uZbNwFRdeaFUdfExepnbq71JaJLaDOiaKU3uRqX
dVfB9HvYhXlmqmvRM4OluYzilQazYiNgTyxATvTaM8LNPxgywxp92FzEECbZCnWv
rbnfY43B+ExVVohnwxC1qMhvGNVXB1OOlRQynkDyJuDdFYCNjDh1/x4facFDvlNW
fRo4ZPXm4LLjOUDieL5GQU7pc4/1g5FkpSafHqxVJO5w8uehax3YOMXI790R0cFd
b/Z15YeybKSb7U875GhEGypFZEsBppr6ttbjSEF5zhcTdCnfGgH8qKevbOERr6wq
zY+945P9Oop5QcbXvecP5Sw79E3dEPXDwg2J1vlYkfLKsUEBaV4kLzBRUeOzYlkB
l0U8dNLtQ5IzVosgTtuJh1tb0+yi+OulLf8s+04cfxrv0qhm9arPmm0P/bYZOz+l
Jbz5Q9juRQewawi6nQ+OZUZYUkc+YDoN+5PNuPq56KISy7hRdb1gblI216esw7El
2toyc6neN67/z0wSn8C1SEbF7lv4snDS1y/rH9xV3iFbGs27/snIO7pr0ZTRA4cw
yap88QQTuXLGQ/jDKSM9ejtBH/Xirch2vXHrquzR6fZZX1dJHALXESTEtskCrbG2
D/KraNnB3KJUTQ6+op2BtlfNzXvHagZqwFa0HX0iYFBnpdPRXJOCtDZuDYz2NQec
nbYXsw3rPLDVazW887AhyNYKAcfoAkpQ4pZEVpjp5m6e2J3rVob0vq93aKqYEjei
s4mCGhZgKqWCs0b0OPUird0lS9/ken1i2vQr4RIQrBKUw9R/vigvXvrZ9XA98VLq
NEmcXNMOo9vLzJ6cLPbutRJgppNISSwaCSgm1+mNZBDZakWy28x9HxoBB93n2pu8
ghOC2KyAzSEVJ8iDg4iOlgg8D6acJar3KES1qeUDYS8K6ewBVxNV4X3hmNFqKIAS
ZtKWmxVeqJw9m0dmOPqsj6/Ilh4qhifyJyBKUA6lNdRn0pS1porNn6ozmbR0NsFW
+5ucQKLAwufD7iSikLC3z6TwiLxTxgvkGkFMi76UiJwaJ0CdyG1phAcPsaMVT2Lm
TFiVQijNmREbZGshjQyREDOoeNvLmggDkrTgUhpUbgNlzZcVzXgNmEO5aKJlAdWq
lZs0AzsgNmX5iJ64XKmACL1GWOTo/9VlwUNkAgZOBBRNWjnIH3XolHfiZc5yTKWk
CcRdKYi0c2ly9odffRvgw3gmlgaH90wthV19tjaUkh/ypCRX4RfgpeLVhAS3r4Xk
YKAm+P6UUpdnbAl+argv2DhI3GanV5AWBdcYWTnk1QSyZQko8GVhRv1ENCsa0l5h
GMcGWyzLSagXpbqpdaU64S/FWYmkF0LiQpOXhKsQvIiwxNmWxBdieHjB/KsqoLCh
xkPA3kmY2I0nAE66uqjqpMWtIRryRYQlgwFdCUo6tE4/PFpUEMAShoIjn27I5FJv
eR2aMHc5ijcS6q0a8a4quSs+Iu3DFdv0OPphr/rcYJUZQXMZ3MXUjPHBO4qaB9xj
b6vxmfdDTVBDXcYLLcuiXK46ZS1lXUyL2SELvnPTjix0K0jDjIpmaLFQ5DONHT0n
Xr2MGrPdb9tkKsWQmStZJAG9qHLIJW7z17fxLQVhYVG7uLoCcL5FENuSgLQ1QGXG
qx/7TfjW0nYViA/chUBUgcvvOYX/Jfr1Spms+Ur7DY0Gb/yTi/JGSXu9DWAhXpGG
42c9Lo11V6lysEbyKHmq1O7dC+kTZWu2WlPNgxRMYyjlUF6D7dcnKJcfPLERZDvx
DytB3BVnlfHnWmNMmhglEUrK6uj8bA9pFgIkzeLerrMr432qqd8vPTLsdZOG8XMl
gkSwxGSoW0Kd4NSrfGUbxLz7wveLiKqoHxRmXVz4zyIzQFjBrX8hwKy159ySYTxt
RQSGi0uuYj2EyynltVqGzb5OdCuKbof6wm9i5bd9gi7LoItrGZalJ92K4OMee/a2
sB3VLSWPDkzkukTxqiXjrCM8rB8csbz6yAmTEU52J/7fa1/3AYIhP/dBNXSBFjEQ
vO+j9zYFAr0w6BJVMELURQgTThO7UR76Lgz/F7QAQmUN9jPqPsh4mwIz0+QzOvDt
sWhC4Y4DMMEOKzpQPmQUXCwP93l0dgDC8T0d9yN7RMUx2Hcloroyiy3LLJY64+nZ
uPuk5aZzTOiATnqc8NhCQuaelAMRfa9K2aywNnD+YYg7k4FO1x0rYPxpIlDVMRI+
zuOlQUYbSmDeOFXK/kxrYZNeIzEfLjGgC+sDsNxDww8KVSlc8COEn8wbv+4KfaYv
Ml2NlNA9pNpEr88dSTeHccTOmbAgECVFP4jZP9ALWCyUn8a74rKZRagH2RUf0yo2
opKttrCVhejFAwdpEgo6G2Ms4ScwbY2SdgX7GcmA4kEGjjVpR0kO7eR3UoXxkRR+
Nld5SUUykXduHW9aqm0TT0NttVo4etHXiYYqsgjv22xakL527BT2oB810wmncV1R
cKXSzHUZVZYw57TuI4b4Hq/DLMv4lv24ouMeqMf9uolrXz8vE3QJploZm+Jr1T8J
VtVJHjV0quvz43aptysUOj+8irPSIpor0kFdVMlLbdE0lHmKw0vfhmWav8/lS/wD
RGFBpSSYlEpx3CvVl2LR9K4tKaYIuChGtePtxCnTJcus9v2c71lyie4awOg58fVn
ihjIrXmDl+LslaGV6ltGqAFPg3Etxdd/p/bkPKwHgqK+PFvAjW8ziMQeV6VxA9t8
WpoNMi8meNYXWJTG7Uav4pvqQFvzleoANMiEOPKY7rP4gbJg+why4nHgI9TYfQGb
Zf/sC6aecZ6JuqRNhsNx6Cko7+j956A5YueK7t0PnofRqKhB16w/Abmjk4C7CeZ6
aI37ENnW61oyz3TkQHOHiQM7HKxbQ3EKoxej9mzjWFZTWJdg73zNleZAkWElUwZH
g3SUoS0zNC/1+xD0aRrhyziPOmhK43jvJXIG6Q3FkDSmVrE4weSeGoA9gCJ4amQ/
zL2I3dqR8mOhEx4k50D5JATsj71f+cQPPnOTb/9pbcJ1zNoWRmh3PFR3zj+vmjiH
ZtkaR2+wXGEIwIptrDeo11M2eppPpdtkNb+ojBs7KImVCtGz1F7C83KeDybyf6aA
AD+cb2sgy9xwM1Fh9RFV8MlcJbPZQV1s1UX9LNLL1ySo0k5p6fmVnT1ChfPNHJwI
02tmAnsrI3bM+DHrC79dbb+99l0aoEY6ey4ww6kZVlAP2SvSPHypctPHx74il9tu
o0uspSXTNl4SxHHKKfZnEEnZcxjIpleXkmz+6VjC3tSNzVRh/MYnp/+qr/er/bFF
Nu8qp2PIw5KYrIbEekpMJyspJTD7nqdYVKPLGer1NOD0a7eqR69ZcaquPLh1wl+2
G9ykC0EVlkKSJHsMw6bt+fEE7/bnoKLZqnNVobRIFILwJk5wd0UhG0hJmEtxIxUi
naBvpJtYRXxvGdTeEjnDg6FXdcUhBHhYGzyfWbD2KtQEHHDzng0J0+DZlxZoRX1Q
ENw9yGc8D+EeEzzjZqFLiRqPvKPdcr7YXdk9kRZeK1phVUiVDS3vjO4Ey/4Pwg6m
JviBnEEE4vWizYy7hIMC/oxeyDVDxpn/6E1Z/joKYx1uas3Rc8pI6hxbAWxLamo8
SW73cOHatN4EHuES6ujkl7ORCJM0E0nXm7DwlAeBQrqAbrynnpN8TA2yojS5lP2V
Lh+tq4C9UFncssq5r0r35cI9iefP+TDngdzBae7shWRE5Cb/yXSyWBe9bDssqtnp
GCJbvxzmhrmUhqeBTIRn6Uw776ntHW4KNdwRmazuO6G0HVHKkGc7gSL14cDcZv0f
0MCJkrYRd1lOw5LFQTXJysqDjWoetx3rNy8QUWuRO1iJBD+Hyub5+lQ17iKucScG
AFJ1ZHqvox89mZptI4ilyqTh0XnZcsAbHhxN9szxbtbk184dSktgEig3Ymkk4e33
Xt0vMLyGTkvEYsucRKmnfYjnCau76TyYIHiGNZ8Jz8E2IrB/eLB/jjppAlALY7iH
fc/JoPLCv+wM9QES9ZP5rzytujLbKMMZvf4zTShTRg2Kgk8F/kLoYpXSSXuvJqQW
qdqU48DIomx0DobpFuke3mQkyHIAYeLMirWKtEFl3zOad9ojL1TVv3m2mpliWsV7
Su3MthCXbHI0Osdq1okX77adxMBgDsXVSR9VgfvBUl5pKWj5518u6CqX9zAqCT9+
P0CmucvKBDECGVYz5ysZ2vAaXWCUPbarlMBAuHMeC4B8wVqUpHhSdZ1cS2kVAwC8
tPDlm5D2s85HaZxfyCg3jjkQyFqIWdrD2sflsUWxyDdx8nPJ9/jtZMvnIVCgD6I1
wOC3ZqL3OhUBgfvvkf1ScJk/txGr+43tDQOOzdIkrjovupQ+lsV3PMDXxMtYi8r9
pd9cyvJN8pNeSsKUWXsKK5m6MGJHCkwuW7jX/7aQROsVa9CqzmGulLaclg8Dh/J5
3MIed9ngS0yGA+1N7P4TINhNwVQRGi8UdI1LCww4SmcbbrBlhxDm1g8zRq0DrkcP
FYhgJNP3K34ChmRsDojwQrR7zJTxV5TmGsp5ryknQ09GzwP9UFnGdqkrFDIR88vR
vz+RaH+jT5qjLTnA+VUP8uMoqTQ3wiPTkYMGXMZEur7Ic/e2XgJZsi2tVYw7WaWg
fRDFnbzSc+J6csALUhAgg6AawuFT81DvEF+nONpTWDcTfKCQtdrCzjqho+Dlvvcq
5BCrcMDxVP7NBC/GyeK4pja897WJaeZftGhUHd3Zq/r6vGnpqrWzPLf9Y5Btl5XS
A6y9M44WL8VmG56DDNapVZpiaYu+DhvyqtQF8yghCivIwrRfsuFlxq7ph8KIKwGt
1nln15YLskWCKJllGpUFCrn02tkH4VmwSbxkRK/ixNP06fQ9YOkcbreaqd4g6+Lw
M6dRdxH7JwG5cgSCSBJZm5r8RDBctLu6shUkzcBVb9QBzfKpriKY2crhC48reD0X
o9QeTk9qTlmEks7tzXBa6u67XjmprgQfqzya31qZbZd0nXeObYkNSk0JiCQVYemG
i3j6tNTMNdecVN/QWrMtbiMBuajkRyQ6alxUx+O2l8iWxmJ/2bghebp/h1pQie+P
wCPZNVuPn+MKaA0AcYzs4hr9kuCERTRQzGPQw+DjObLMtZMv+7NoLiWKYSieuYR2
58TGKixVphI6OLh3BmO34EECDvKtBlj7jrwiX2kx/ZrmIq1aVQj97YxqfR9MmDRj
b2U3vsE49HWtEC+b52EYPz9kvpOs3k2+ZEC5y7Op6iuq1wTX48YQ41RbMQdqbN6O
F0T/N4yos3lE4OwZ/7p9cgspsaOhcKTLu0BFTtsF7W8hrmjR5F304ehagegnsy+k
cMhIK7F2OURCSvHiPDcxPFXi0CHiM6AX2SSYylyuRxjKlvCUccCOEMqctQqtnXf/
9YlLDjwO7tP8P7xCE0Rf8zPWDOXvVsG6LZgXCytbBNRxSvhH+7MclUcfryfLHwf2
1mngmqcJsweNQM0Qlw2LvlJXoVrHv6/ZV206LUfyJT0H09rJsQQPH/DOiTHiQPVK
DVx+8mXP7ju8oUUv2Ei4Umwb1JaD3uIPy/Dw0HS/35/aKjVG0zX5dyo3qnpthMI4
mOwZhi3aE2BlIqLPzutEcr2kuPXPznORzgRE9x7NEJM4UDU/hNDqz5uxxf1bCqUy
fKR1LIzxJ3noXl12GjGwbv89EPapbxVU8egNCj6MB863URiDpTFZvqtsqc96CuFF
QvMbKVM7ziDFrBDyTtomqFKnhwJZdgEtdBw8qmcpMAqpe8/HdVEGA7YvjC5vSPi+
/UgynhDZsB1utIG1l52hdV/11Stywz29tv43E71JdIXL6cm9lRL/uBp6snE/kkax
xo4DOh2viai2+DAPz6ryT1qS1k7ONh1DmnymASyf+aq4dD+IAbqUZvvT62j6VJsp
5uQQBpmdNZ/KR1kdYrhbg01njzZKB4OFj34ucA9xqjEyESZiDlcTjlBcQkzF2mWg
4NVOVYSeKfQDqiPFmjaUFzqFhWbTyxpWHJqvWGvFYTFDAAvPB3qN5kMebr8Q0MTD
3ru+YT/r2sovVh+NsnaSVzfw6LhwotjQ6O0V0QfwTjySb8dOjqJ3/KCuZN4G6eXY
5PDZrigPK5m1YeIZCazDU1G1ey3hftCSA5qivc2YrNBnRuCCIRDOmOibCwI6T9/5
m2OeFueAoeice//4CxogSzN6622CJ26dVM+wgCtbMibLv29akECViNbGTaTjuc3+
Eic/HGNCvWD8foH9DGnGtRDfwjUwy0IvM7gOgGYb879WX1VOGatEREz9wOpSyFQ5
E+wsPhbUpUZ7NPX2nACYRr8DYMhUfPFokhGpDz22m49Jl4dLRL6GS9+/6ktsiHZ4
/U/8xApG+gMnjya0PXsVz8IfB71NDX+vLvGMetpHkAQ8778fgsSzMHh07QOZXCr4
C2teSbdNmxeiGU5P9+SdA6ubXr8VtbysmSMt5YIBaYHZHY/rXKJvfbzYeuqUQO8V
cQdu0N13EQ4esVH3W2F28hqs64RLJ5aazbSDopkqjAvRmQ4Csl+5KHsVbokEvY/8
2vyf7WX6j36UWmUjl1xyO8M2WmIi14RMpLAiZAEY+M3OFpUpvmEbPtWqLbDVqKcz
NElLn/bFOHroIckyT77ZQO1A/BTDab8R6xTY+KU4emloxA3PbhI5zV/zAondMmvA
/b03YWzliG2yU/Priy2K6fNvU+XsCtBE5nPM5zSpc4cjpEr6VwAFD5hPK9q2qpk8
CbTY3f5znDK6UMzTOV/WqSFzQ/r3IlJjpQ5Zs4ufONbmteqr1ZXHyOdThXv88Ain
1wsZnox5QOZ68m4ssSImLrlz+qhqkHs4HXtN+E7mn9eco635PIk0QV4NYG7/I71b
GPPtVxHPEw/1ROe4G5Y+WiA/ikNlAJNwpxBCYK+u3XOSQspUWTNWutPS3JlZAbBq
xik2fP7sOmqk+ZEOamYzL53FD3WY2mlmOBCs/GTSub+2yKwvXRM2eQw9RPsfRV8k
oi8EZajQDLWws3aU8qRPtEJ1/rqqpo0XfsOB4MbcIzk2GhtiznYd3SgsxSuInbyd
KaXZWyDkPahVTcPoA5o2EKlsMm/XKyiY+u7UuP7HFEDNsCD1RhH1TCzpvG58cQYf
76Z7vSBT/68U/htyZszV400EM2QwJM8321cGvRhE1HFg/khHWn/3TgIKbH6PTG+i
S8UBeYp07oaXQ9ArX0wzx1LnrgiEbe37hugMb+C8K2j00F+hfQDssoADDmu8bT6T
XeESBScYlJ7hK6MYLB8ot/HPmotsK9x8ZHby7jGaalvX3Tz3KgsnBetNa2p7+3hW
Shz/R1PgaTim0y37/lh+Uwfg4cVFmuJn0bfMAcHluSBzw2YCZOkUa+vwIXY1iVaU
2+EUt5N/VMPHnuMvBC2qkIZkgOSJPl/nnNRQBUmZn6yy+M5WcoUh9Hfgx/0qwb75
v+/PmZsJ8rQyO7j7w5V0p3EIHnE+xs3JlCHGZt1LFugPthrwaiqJcabCVs9nKQmz
nLExJ+qCs37HOq6ErdKtwi1cLpZ3kdx+g2khGHekFuf6MUZDvjPGPlgxnBRLJtzf
alpbunoAEBpKjuePnHmWYD98WbrZxvH2LOI4Ao44NXB+QKY2KfRRoNIOX1C1u1B9
2rNeFrQ6gfWKYuDdqTtMBvfegG4B2j6GTxcghKhtPaXHiwD3hvFZ2W16TN+CNmcL
VsY9CaekQiP/VCg2qQ9SU9/8IFYxCRX7pYeamDEV2sTqu8gQh8OxhRz2VNFs9UKE
5mpr6sBVp0Kb41ZLZ3a4uiFR8Sr4j32mpgUgyGDbP9FU7wNzvte8Ph8uOd0nOO6/
9qZKrJETQaTIkOGNMJQ2WFDclkaoaTgp89WcD/s7syMmWowDcMX1qCKltxSpycRD
SsHyfqTV5z57OwW1qLMwGiRXcKfIUzedOyxlu8LKpc4pch4Q2Bw95G/B3gZaRIF1
UgaWaPlsVcXLcFKmIJtnhm6cKyQNdriW3CdaGA/0kiuFuL/geL7GI7+dX4PUWVC0
fq/GG7mD8rumgh+6AeMnkl4F5gDaHfnJYvyVcnAu7W/RBRLzfI1Q164CQFDB93AY
Noz6OPjDO8aeeYcQl5EYWSitHEPiszMtOFHnkRDgH0d1LfvAWdZ074V4Dq5Rm9k7
3w9B7IOaAqjqqPtICJ2/L7mkFW2ozFAenV1i/yaFTa88oyZNC/PoFJmJZDyWiXvC
WD+rBJ0Zv7SEO2LJRGENj/RMRlKt4Ko2utz4qlRtjYE+odeLHoSbfnhFAtoKz4yj
l0U27cPTJo0FBN1R4ZJ9CFsBCtSBnmzs3atdk7PbpTfeRdbXZQmYDRUDAsacsfEJ
MkwLbl5IIzkemTAFOKFJJ1sBplDow6FC8bQp7zgp45FdtbWizAtdy/RYOLNVu290
7l5WE9RnLS6U3+RKM7rlCg/CBMIqpT/SAGt+rjWfQNA5bKf0rsDhpoReqP5HhHy+
kC7aNq8QUJo32Vb8wQ27xUdibkYgdiETzDo49GBxbIT8aevcuVo9mFZAy+Cztdye
ssonLkaJlClJFL73Av6yMQoPcVpbl3gYqibwGO0z+StMKEN+/y/beIvw1QGfOeoa
jrl2F+qpFcp3reTlxZEf4ovQfMsHy5tVXCQjPQfkAOZUGgKEGAUrQzUOXtTQXokv
lIzgyz7NVMgBG6IDYKb9uK55ZdP8j0+E8BJhaJ5DANu6rk26tb+x2mUIwV5PgMNB
jGJThPPYJ0SYn/ehtuYWwMRmlvojm3okwNYrB2eO8XNXHJzjQvWYSEbDbzeUzOi+
KZGauoie9be1D9jn/VRhLkz8JQ+L1Ufet8w0QktwbeIf8J1/+NcuuTyIbnZ1WZ3d
MScA5oTqp56zm97g2mnuO9iHnKwGgSryZlgv8K0E0mmLmuoj86bbFw9B99suKWrI
2ebT5LujWm+lSKoZZM+KPlgNh8dBc4nzRYRiK8E2yDet8JwNy0f3s+lEteVCPdl3
lx/fQWFOEHN6V1oONXkrm510eSgmr6gXDMIzuqAfPHNkYPXSPXd63JOMBM8u1Ndb
I8motXRSTfSI5iZEH7IKDB7RrRHfP7yTxD1PScS1HRK7qkk2Uf+wnNs7gkPgfKdz
cM5n1cL5gLimQOU7+hq2NYUlbg1xInvuvYs+z/N+hLiNsCuJjpkk0e/Qhgxqxm/+
lVE9eDSmr8adUhkm+2ktZsCKGfENmThKgMz9vgZszfq2SHMgOnwtz4nQyJX5guea
EuXl9y3cKk/okZC8X3qk+UWpDWNt+DGXae/YsnE3x0X1Ke8onKLL9SMgFWH2SFYt
koRy//IhpPNStZdjiGyXy6XLzsKlIjcSjn2NpOXC351aWUjTR5RqKvWUzrBY52AH
RjY25+Mit7xcCxzNQlRTqjUt5f+sW3dqFyzJM0r+PzGp9HU4uw9rOwJKoEvPOdt+
ytWTi1tPxz1AyQjc2kSkHiG2yHFYT2XAUFZtucZt/qg+OGOZgqQrM0fb7Uh35+KD
2gihIaOYMdfnAqrCVzngQ9xzuQI0/zhIoFPW3NUzMIBmsb73tDnRF3DgtB9wfCwo
rfNyohoMss13MAFGb21wXrloriY/tS8QlrPllE6Y96LUr5slhEtP0xMd5YUgcmcB
8VXoaHwCBio52ofrM7jbcOmjt9z5ACDOw9rwBlGP4n3Fk5Vrt2ZcxZB5s6WxiPs1
emHZpulk16iFj32klc8JfQ/fCA50iOvht6zgZYjnJXneezWMMPDDbiGhzG4dt02j
Dp9TrJLY6gJqHK0irt03RchfuNrLUWymkq0RJ590qmpYi3jwk9Um0xiNLEbqrh/C
/uWhiHt9NiRnPov8xTyUpyxbhJQ5eIKZf4OqEYy2H9rIZiriLo9c4bRRkLBBdDFx
EZfZrLfxQRKmhn92x+Dqjk1LTMEQUVFQ1Jv5WKqTjd9gxetnF87q1fMyofBwZTao
iIB8vs79Uk4aWajVoCSDlU2c2v4ASMH/4czNTSHEDlAW5zhuLLPf/jWR9KwIM7Sh
BoCGZbZmp+jqRT9d3iAos76O92/zFQiKFQOkv4K2mfPyFDNS5N2CgGjp3ve1p7WQ
RYzPkm+H40k8c/uozrLKuwwIAj7XUAWPlwTnEh1X605mu3CEB0pgcSGUouPIES6n
xoQ49VhAwAme+kZA72gAl01LawKVEtaagiJ2DTIxPG7iJI4owLPCrWvU23sfI5aQ
0WVWtArrgqzC4z5PquydkgBoeatko0XKwo+fCsQSKsVMKPwVAswPh3Ozyv+sdLrb
2jip0TFHhcGerJkGaDB3RkAPRe/S0l9kHQLS69VSH8UQQ8Tx500nGy3Nz5AoJJNb
Mf5ZdJ//RHJznAjE3v/LEK28GB5MuK7FEwzuFuUZsqvZUFr+m8pmtoQEP3fNN6kp
Zg2/RDVePgrMBF4XbkB6MaJP17UplsTqF9B3h3dEwDg6rcaE+kupKr/gNHUpTMCm
dJ/W9ivHRAL6PvDnRTYNlBpIagLBLVG8VjB1rRNo1DVZEYsqTQhfhFtBDqcvSF5S
tXSSK7Fj40+dNnXFbNBO2qEPHnA3Cjb2M3TiE5dRLg/H1GGQf6hKX4b/qkbNLHjg
er54kY0PzIAprne1dtYR6ZTvIMbvEBujh7W2rgHBXcT8H42SzTOxwq+0cQaYL1MG
MBg3Sjgxznr73sIcS1sfLx/IfWOx3iJ/Ipnaz5dtenr8mz1DGToNlsCLtD8kIe3T
qWj1YSuC0ZhWHBz/0BRYX6qBZFLYNLjSUn/fkVFtTE6thlnnGrrLHV6sH5K++hGZ
RCk4CJureO1snBgSUiNDl/HZPJBC8teIn02OxsekmDz+g+U0ZmoJmfxXPgnl23EG
6w3BR9HPBJOBzHRhiqc/6tLMZ/WfF5Rb18hXbnqi6JcOH+TlrF9D66YgFFEMxV5W
Cgr+5kP0N0qAhAgqW7rpZrxtPNmacHFDKsm30QlWfYA4zVp6oY4BBjmWDmp1tapr
0dyBKLwTif8XcnFDWJTpE90maqH0xAT7nSipKzlhOCehbkT9oyBeSrd5M+IM3nBS
Ut0SSkxwXdgTjq4oEG9jAmeIALHY4mMD6Q3iLJ2IQRRRxVS4RTDU7mID4A5Zjzkv
cas2ZrAd21r7lwGYvYDv/8g14pmfcuz2yM2sci0Cv+of87uGmjPRU9/OqsELX7fK
/HL+2PFJkTUKvZXJfRG1i6kfcooacizO/GXbPpW2qPIHD1sflbX6judLevTqwYyi
cdV3jc8VCZFSqk00QEQ43+LeHb9zzdjpb8eAENLVJOtO5s1cwWUho0jSWTvxSxc+
Kw9VeaVYFJUg9qH3QdGTTSmRZIy3bJF9R44rVQDA5e/km1gVId+0Y1CXBxlbiRRW
5Os+JPutDzZDtt+A81oTuAcT/PiAoxiUIlqbIpCYI05PVLAqTS6koA09gDa/5WlW
vI6I45PBfECA+0WufvHeyljJGtUjQKoDgrE4j4c2NTI+Zey9uOiRzgrffzSY1mrh
rVfcpHVuYq6ylc4FXXN1CFfcbS0VhnTEEuuLhuq8VE31rPtswfAs376WPdJXXt6M
zflAeB0mC8LK5Jac6kBGKXXp+Ck5xrNAdnDvpfe0ePHAEmDTIIlaIJfhLvzK+ZKK
CGD5peKjHII59iBEfot1L7bknlzamgGM8TQ9+U8sRxI4jyssPWV5+q+0pUFLGpoR
m2UFllRKTkt8sxCIn3y9weupxHhkyo2UKTWOm22r9hLnaC/i57ywi2T0opjlpvvW
ffT9PbxYJNCc/49sASaNYfs9hBhvZ5WmBAwzIInavROtyhHsWRKcBRkR0nwKRaMf
s2No6xv6iudhIoY8YoEGtYE6+9avfWouLmSjFQMboajGb0orMfroFiHmB9ixfHxK
xQ+ItAzL0y03CwZQK2BPrFye5wtlLdLS7M4B7t+Z4Ghr4FCETICOpzeofeYNqFy3
hbS4/+BNECXQHnMn2GOd8y86vau48TmTMK59UMKqAneEm4X8w7gBk5xC+xqTxHn6
5CEKv7JRBlz4F327poSZxuNI6G3lEGqp41a90WnKKI8bIELVSsvnaySoo5mVABiu
3UT0MQxvjkcU28p6UEbgcOSVu6B/tB2bmc5/gXzOcyKAV2W1ylmo9IHmB/PaZt+/
Yk88jJj8JqJjceBqwQ62sl9m/LRLHbYHBewfdJGWptgkTJ8xUxHDhi57bIoCj5uQ
eJQmUT1y8CDLJ3/fn8w8/W4fsqdFbvne8FiWzYrjDB7DJ6GXVVw/bScn0imsr8ZU
/LCh6nieSWzipOyxNm77fISKsn3WFxyY7kyfB7lTI2ZyG42MNe+XqJzChaMjS5M2
oCrDy0qarqZ8i/MKtUY2zEkjTU9uXCnTIhfG+/bsGfjuk+ifsEPJo+wzPoEX6AFB
iY25NElhHuXpqwXeHbpucWw4jM9kOtq2Q6ez9ui7mLMaWEk5sSKvs3EQAwqt+HW6
5d3zDEbkmqWleWHlBhRdT4gUKnT9DwAok+5AXOKqm36uGxDqQud/Qro5/dexSMiw
xcxN1kTjvSa8MvNMJVIKetxO8GpcFTd8SJeV+QA4T/c4ozxs2fymz/uuycPxJW51
Iv9H2k1libYhF5AE78tTwPDwTDq1k+OsSSnhumOO0pLfCB7AG6ZD2x/9XJAkwMyC
NvFfPhDlhGYyUSvBOxPd/Tj7DmQkdQTttWB1mbF35N/juwlg3EGyjsCQMVKdIee2
LcGfypHGepO8LW8yCkmQ4/dkCZhcml90kW87Pyinjx6rXtKZXylWaV7wEyFOTE0N
ozFev22IaNVjjeKBgns6tuYRY6Za224XnvQTfO7beJ2QNkSwb3N/svK+lFem2PhI
FQgn+RAhKGH8XLIaOMPWAXuXjL3HLYqfmBGPOnWALnGKr4CG5t9vCrdY1ptxaD5p
Hbez5KgRh6M3otGoYMkYzSfiFxtVRoxGdjIKdw8pz9Awhuls7dqcnZPx/gnwspjp
0ok8SiZ8BkyLQnQhUEDux/qXEVWC7hiOr6mli4zkOFSIOVLeZG4XRNLw4FTF81Jg
gn6g190eAij2LgxqR2KcSufcTrfKG+GmlBW2PwkHJm+HvTVoySlbBKm5AYgYQj6U
QZVcZyq5rinKLxXqpbG5CpWi7Gu9D/Z98o2sg1tkCW+Iyzn7ePD5tU4sjGLu4VnO
ZGHKsLaVw/uCfCAmqmnm0l/Ms6tzb92iH2muQ98k5vb9VWNgdnz4XVYYkD0zhabi
zv0ZUfQluuk8pEmzF6QkortWIS8s/sU4E0z7sxXCq8ky2jAhvfIc4A094xydMXhb
MZO33vobf/bMHt33AosUzxquUuY8rGfhJvCN5TirA1VniFe4G6HuVNwpCVkEqDW9
60Xvi4CR0gyPVM8Qo87Hx/tV6JhEJfk8jUeXWunSOK96Fyo1wEVwqMIBkP5XzBoI
GyoN+ZVbn+tkXxYZDZlWlrPfsh6QjlFfwWoxyuhHjPQ0JZqNvMvWSgpqJmIDnr/q
oMisPIWnoNx7rom3/zjWrBUA9irwPLYInr17NwPYwDwos+/fgl9gTlvlG4r660p2
HNtG/JWuo77T1Fnddrz2UU5x/dsgk1esigFaIm7m1PFDx9QBt/hkP4MQ0RfC3t43
BYeie4LZZhznPIrncY98MebG4gFPfJ7XWQruVkDp+wyvZ6a13jCTm+sI5QyHvsfp
7EEz4Bium2czJZ2YhYRXvQ9TD4QMVoMg4aNahGy1ezfbL3DaJPD1Bsp40+pRXBt2
GlxVcS/PwDfdf6tHZKkAkfmaf7X8+4rPrEsyWyF9cvgyWQCmgNpd4OGMLKy8W0ib
YPa/+CehWoxvQ0cdgwrXzCPTOCbzRkKj8l1P5Kuf4HrlTU8VOS8fWv7JB7RtUh6Q
PxTYDvL0s93p9t9W/+z58Sa2qIe1gqNAWIhQeKxsPgcurmBb7UBo63wH+8+5YhBj
4QOhMNzbMo0t048ZbkYxhEPYNlUa9uDFRDQSfCBr/fY3tBBUdv5JuBR3+0RY2uLR
++U2JePl7zezgD14HvtgdeSJYAUf9hJ300ggbISIL4mRGZBisyqt9FJGYnEKg6EX
VzHC8Wm30yEmS7xiZEzy5QVSBhX8yERgXh5YLoY7MUFWoWJiQurHcVYNn4qbENwa
Wln7T6cyiRakJJnj81sGmw0ffbltprmqsfjXXJ9w6ypLUPmArMCvgX1/OKWk1JMx
e+GiZQi93NyxqFLWmPyieZbYvOt/LE1e21FivTiMJ96qhRcyUeWymKVbIt+Eg9yg
fQ4QtOuADN1Df8Gz7dEItgusgWh4TQiehOcHKNM+lNy6tdp1ww6ttN410pK1StWU
kCIJCuD1q+W5CHPiwRQlOoff+6TrH1tX7rmAo95oDtRPHSIvvkn8OjSo5yxl1Igd
sulj6yTm6mA3KtMAuI5TcvxXdynPb+sI5SvoT83/4mb9IKse/Pc8gftsDkhbTNz5
N2Wq9Ryq+oQETOJO91KDQoI0hSFNT6mp4D6Fc25lwJzr6N4wjcdYjd7GlJlgnHOH
KxYqnJSnzzv4VSuk1AssT8OliXnmrZ973r/GW1iq/fH4kJA6cH3uTMY9qE1MIXfJ
+wn2PSaPsbHl+VsfryQwEQzRX5Hho90EKFaj30xx4v+R/MgdjZcrhFY6IsOFhoDX
MXefft3DNPk3mjveySt+Tc+qpVZgiu6+6jdTzqP4153ay0ICJDB0YdG7UyzvFzVz
hGDG9LqXkB2Wj4RUILB4qAr33e8CyycZrdQaUtetazOArvv2zlJ6s7SsFwp7LbWM
Rd8ExlbLfHazAKABBJtmUeuPfTBKoRTf29djv+2uNv5LW0VUiDEFZqYWbqPehwpt
kfFf75dWW1DwJsD55NSsZECMBIExKuZBHbHeqKBTWDXK5+CBAilBEo4vh3pLdPK1
DW0rDvP9UpvvRdS+l4jZVcFvJBsMuWMRcNC2GOjqR4w9En8wC7wsZJwf+kvGZ4dn
h1JDVkxfI9joOGhRoN1FpYugLmbIYQrGzMAn9dbTnb9Uy3/H1idgahOsALKhlF/l
JROBGUZ+WWOqhRSpAs1P/I6uaA8tgbfPyyJ4j9bm/EyC5jrLqKMsLiJ0EAdF+kDw
6+QQMmi0M0Q3e4ItIIj5y14dat/iooteoXtFrOcR775RUoX3jaHzsuCk23NH65VB
pPb6xegapCRBoHroZ8xDSCkcMcU/VZm6lXZHwLNGyYkf5tOAzLicotf2O9h4nZsU
3r/s2tla3E+7bQDz8LA6hMqfgElROX1XcOs41yS73a3CleZpbDjgU2UV4HH3Kb/9
XY5QfkIQjXSmoAERrd/YA053P0GTpx69x4Drvj9BzTCL5Tl+N2J9DOIqSu/VFxEa
v12DfeV+zytIQbXPG1QYTzMJW7kqm6OT9LvBiC7iVA2cdYSi2aQoxZXAFHOnENet
2/2YamHkDjikHGGiri0JkMivlY9zF6K3YlZYnAzLYuDylNSOCRiBjIDJGRGi0hO1
XP/X0Poz+1hpKBwnC236BKWGJg1s1nbOdTbTANzxi257Un8ODBS4BwA7iY8Mf5xA
0CTFrqOqG7EDevdZqIx+4+GlHHDxLHXYblnX8WOYZ9/dA0ZHzJhQGXafvC8M55tp
wnaRC5rRtk4A5wzUpNedc9ACjEwrWmg51WW5+YymdF1iTuMEx+FzPh978SRwiWY9
sbGAhcsdxxd/uAJH3JHQ9AmonQA0kDKNWdRP/cPTd+CjrKRVp1moVuvkAn7RoL3s
1lmz5nYP2xZQvovf6xW3gIm80F56KBzo/HlTVxDDX7gHYSakENt/TRy5S+wgRX2n
Dqtl1+dONojS8WM8Oa7ETDKjjPi6/OWGJNkOD8jaKcdG/CAv2cIhEWLoYDSI01xB
rVcU3NQbTVG2+L1hzN0k4Z934rwjuIaCDb8bNrgmO9ghNIMmdBv4Y9GjEQ72DfAA
tdcRAV8isyQgDtCQu9bu5KN8BqssUOFpD0NSQLCoReq/APygbDAxdCHkh7o0jNhe
0DVLwdNGVocA/G8UggjGYrYBbVlqoEn/BWAiLCrhF5uoQP0g0BoCmVzx9+SsTbJr
5W3tqdTyURu9LHWVERERaEsl+ITXtB1Pro3kpkioZYppSXKJboOwwZZELYoblQaM
pK/K/eAXMa1YCMQX5LUUMiOAypzCYrqdYjGzVtA9DNit38KjM8lvIGlwQsBVbGn9
euREmezw0miXNttOxTzRsb+qzP5XrN5iwtB21K0RDnk5fwF0QlqWEJO3wO0g9R0D
WjbHC/cANY4tiXo6jDQhsb48fXXvAU0CGs4RhcE+i7ydvtDhK/fz82dYKTgU6T2w
gB57fcBppSdIizUwFbG9tMVgITewS6EVxv0RjF1iaaggZ/ZOxGLqtrq9Pm8cbi9T
ZLU1hsPgoOOHv+p3GNtVucYjIrEHUa3wz9pzbTC5rneCw764Uwg6N6lGRJ2DIkSB
Vmcq8m1ggEPcoFI7ek+4+Hgn+DDwMLy8qFi4LXMTFV5JAHFd1hdqUKiCV+rriPuw
zjnj81TZVj+UGB0CGaKZRPNjlCtOdDjhfF1x7CiK7MN9eSq+kQObe+oHyql1r3WS
h3LQgzZbOg3AZgEaxSJ0Qik783722DB6vRVBIf3fmbt7GvC6c4fkV6bttZv7DDw4
0l9SLyC9F5L2Mo3rWgeV3tgn6JoEyw8hZColtAVeDG/wWtwVXmni9HJgRapWHB3t
ld4mnJ8LvOFK+eQiOX9zYBKaxT0COzBYfzBlLqNn6zJUJpovAaknWmLN5v9lqQ9f
9pA34Zbs8lSf0JTCH3iK4GttehfnNV/EnFOpE+pXDNf6BT99EhHGy9SMSZQEo2wy
BrCH2lsZuiZB/ZW+3qbZqgQ0AY3WpfvhPHuYDGVTEo59yI73ypMiU7EWtsNjbA+H
cgiEiJM/ItuUxjBqE9EzXifBy5h5Kvacd1MJu6y61cSxVsDJhxbjNQAXNKD7DZ03
WBwauaU69qmQ2vAQQfTZordKU6muabRltDnrDh1Md+zghDnnCdbVy7JoONL/qadX
zqT/EUUlVumsOhqjNCdn8dY3sJODQ07iwykOymoNgxpSPV7i7YR6WSFgBNQWHnZA
5yhtvx0P2o0RF2XVGuVsWx96eexZPzxnGDVw7JqeDOuJnFZSICL3JnhCHGAw1zt6
1toAxiW+S0bRk/8zvqhxQhiYFuBEhhyyTEJtJklWm2y3WNlgVGroyAGRu10ujCOQ
9BxweIPsVwCjytHB5B883kO1J4iAyJZdJMV4L8sCSC7Kjn2Y2Lv42qYvWxNVzlEk
N+DaF0tUTs/t8W5x4iJc1dpzSc9YUH1Rz8ZgP8VKPevc5gtvAmcVoHRwJND95s2i
rKmtPAMbamLwe9WltOjyNxQhom32y1S11O7SAGhvSU7VnPpaK9zDRfpTf8hpqAiR
9HaIYrSB9BUvCp+bsFyeMf47EPV54MnBYJ9g3q9Jb/CrP4jsKP/HSVCiqiI4eCYr
NrNbp3U48T7bfh/ptwdCM2l1hr1tSOm2Biyqhmw14jvHY3f74Sq/8dKziEx5Xvol
C2+gCZY2aJGiHeorxCS+gvwyGCx9x/2rJFMHsch9SZP88GW6iuUCaGssFctJ0035
V9sXRyLhHdJhbv7prgKEuPd2nllXZ1WqozmeAtm5ZsENGgEzg6fYOelgCdrvcBwN
OX3q2B8jxvIPGz92Iu+DaNPPL2PEUcfi5LrAKJjKCHkQZoGCHIpwp2xyfWgmes30
qDbY296UZAMW+dC0E1KR1qC8YSYfiHMriRk1zGEeeKOj4wK1oL8asa9egUKBCVJt
zEx+9GLt+EvSb9elf2g3VtneAFjiqnClczeVow94HidVkfL3t3nwSfXZ6vmvpPnY
yTaVyyWdHqlTdu76Y33bsEx8V3QN4h6+BIeYzXsD7fO16oFqriP+82uHYuIxgmla
d53cJnzfFbCickKgEh4JsKkMUa7PDtaONbXBAx/G+aMp6yYLHwK+1+u0B0nde/Yy
7eTSbXXQNHNO0/TV9aJu13ncf3qIcqQiI+R0l4eiYE5qyVgp36QokzdJVFCMTSoa
+lvgXKWrsR+pYxNFgNtIkSct3gNxll1MB0Slw+SHlkybyRdj1YbdAIW76TxDnYxr
QYAuRpz4NkNigkCfPFRT/MixVDBOKLLlHJbnI3LdPQCclBJYAUgZTZdJw1v12Zm3
0/fhnwu+otd3hoGNPkkjRzRi4Cd2ZF3SGYgVDd7VkoA+48vka6mrEixeeBOv+UBA
lRPgjvN9X5HeE7aW1Wz4U8Oye0EmdZPuD5vDAObFfASF/hW5p1/kc3OHmZy9I5S1
4H783ENwos+6h6n1LJDF3tKc9Jnl1baIGp2ZvW0LbnuO9o+22YLWuZHysXREkpu4
chWpk4PWeoGbrXHcc03E359xCd6V0c4/fjnI27zTyYWSGFDdZu72wLpB2IGqlrWC
w+Hq9fEV2etFwqxbFdcy9pDWKHnYtbJHJ9Rf2cXviXYRIe9bfPPBf/hsE/iQwaue
UVKv/XXCK2vSRyOV92b/CYvYSi1B/MjpyPeANZP7LBlicx2yE8OQwLCfC0dF/VFT
SpRmq4Ku8F8hRRXa+9xQKXqxW1t6pjRdTKZZo2tJ7WAX8jtdtxd5RnQ/DZXvaZYJ
EVO6hAnXD4QjoDfKxrtghHdVKMZp4T+LsmAPtH6bOqhSXwPpDZXwqJ85jcCCHUsq
ZIRWeSwSN+75zWgw89GHmR9k/TOLes2JpMDLblIiN1GvSvHIaGpZydxUWqgVw52z
EKO8TAO+pgWZYh0GH10iabDnkrOuVT5cvSV1U2+TYKfhgvMbGOF9hcbU2hqk/71K
GzdnsX2a1xBmQWDXRp/2xnyZkNbXQCUtjg1rcj5co2ziUqt4hBgd+5F3npJhOWYf
sHRDyHKYLORdhBrH3RoyuQfaYc3EuN7dHPAbBnbDdl/QjCn442weJOrSHehD3tBE
DooJ0UUHatAYZTojT3NtvodBsdFU6VRKgOAwDkksHOI6jVSeXvtbL7R+5p1CpT3R
meblMPOhf7js+D2aCUlJfoLS+MRxHTq2P3b5njLvpB9nABI9grJCE9jUFfIKh94+
X71Q9yJbJlKqJBLqWStU7NRHTCCIEehmVSIA2r+Jm5J+eN093j1x7CgqtQOoVny9
GbLUBqWHNLfxC0HH4gA6i7gwwy6NF+kBC4pljAaDeUErhfmd0boaoePTalzzELqk
RSegtnLT1r7L0/xo0gzcKw==
--pragma protect end_data_block
--pragma protect digest_block
VFfmbKeGUWN1tGE6zsRUYuiQwBs=
--pragma protect end_digest_block
--pragma protect end_protected
