��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�������B���8���"���FE�Ҧ�@�Q\_������C]���5��1)2���� hڻu1ǯ�C�ƾ���kT��_W�p.=�@�0�2A-��JSk:�2~VE{+�������b3%r��ӿs4�j���3�}TEN�/�Z�6A��q��P%�Q-Y?��n��wbu���<<{�&8�o���h�D��:��0�ބKG�Z��R�h���W5��$��k|�'ɘj]+�]���Nb��EM2��`W6]GD����׭�{w���K��G'A�ySd�䩸gݘ�ي�kIֽc�j�^�\��<mf��"J�E��﫩_�㋗}2*Yה���GBl��H�������AD1xM��2HmĹU+�K/#���C�|���ΏY�x��y�hHu���
z�k2�&�K�%6�����+�E6�%��w��6ת*y����/���&]��V����]:����zIt���܈�uwÀ�s����0-������ٍ>y���܈^?�pޖnĤІ����ܗ{�E��U�5o_P��<�_�2( �ٖ�U�����'-]  W�K�����7r��[��7����3Z�\��uSq�%����H����VH�xpJ���t���׃��+_��`���;xB�q����+�ֲ��O��g�\��DI�E'�r�\�{K3�Э�!G1�6�Nf��"?�8P=_����fG)&i�K3�EIk�~P�rUq���t6�XY�yy)�N�N/γ���h�<Mi:�Uׇ�H�@n0%�����#]}D6A(�S@"S���7u	�$�=�ؾoQDl��޸�Z᫤���`�B�:�h���ك�@����S@�I�Ѡ����jm�x�f� �<t�_y0�MӎT�-�[��deE
`��s?�L�3���/�Zs#Ub�'��׻����ߙj�G�\�U���s>�mх<�FZC�"L�:_:�1% �c��0��S{��(�*"��|),E}�bJۍ%����!��*wÒ��nvõ��]��39��<�E� ��d��}f�����P��xѫ�n=!��"oF�����~#|,�g"�x������t� +Ѝ�ė**��eSh�5���_&��='�Q_�n���W���Bii3p��*�Ϛ��-Q?N"͍�=818��J�/��3�uRհ3��Σ���_)�X�u��/yց"`_ҳ�we� Q�����N�%:�F�0��E��)*GlWW$U�� %?�_1�ğ;�Mt1��4h�������c�ܥ(-���v�;\�<{?'͘'u��H��)A���ꠚ��g�;�KV�%C��,�՛���<��7j�7&~�Y�Q�z�D���� �����<O�j}b����۫%�nmB��8��D���&�o8�v� }�	�0C<[!��d��Wqx�Hy.[�M���m�|�F�����6Z��6)~5U��Ue��\��g�>F̝=�Ir�}>
��8�V�DN'~H���Rp &�V<���Y �2�`�	�xX7 �Қ�%:���C����O31�8kV�g�����/���΃�/Kj���D���o�/��~s���K����L+B��p2l6W�M=7�ۤH�sK6q�$2�L�$%a�S�:ߺ��x͟s��u����O��gR�8����b"H]~�ݱl`�3ʑ��<I���	��c��;��1���� ��}/~U��]���ayxy��ëЁ�	�޻�Y]�Cޡ�����{��c�=Q��/*�)�9^E&�C�p˕��5��F��lx���j7�ݵ}��3��4��%��l��]X ���9.zC�;���s���G(�ֆ�D
[ՀQv='��7�Y��>M4��U��ih��EK�)Q�^j绻&KYKi�������]wM B�8=Ē�o���=J��6w��ǑC �5>Z�,�߬:U���j__�����x�siΧ�9�_�LX�JQ!��m�Գ��,{,v��ON��V��K�ۉLN'������tN3l�n��v�=U�p��P.�`&s��'����Әc��
*�,��D��nԃ�h�a+�]Ct�Ӭ�_;�~T�-�ʿ�u˽�/� �U�rS�!*zh	�f�vRo�B�q�Mxp�lϝ��s��#�w����b�(���@Th�K ���V^��{}�l[$���1TmɆ����蔥7w�c7�,�.��66I݄�&$Q��h�P����]& e�д���=M�wձO���͉�T M��ڣ@���[�q�aA="�:<ΐ�b���D�︑��y4ݚ!�!�� �9���'�G�]Z��^v9� ��e����ti �^�����%�j�2`Iş��L�2���H1,��e&����f�2(nqv�JY�_���SP �w�K\RR��C�{V����u��̄/�4� �c��7�Ȓ��U�
A����Ĭ˳/�O2S�o���f�A%7̱>�E������q��¯�c[N	��� ���Ǵ�8-���u�o"X���>+���n�o	���
_{6tF��L~9 �;��U�s��o,tC�Ey�{ָ=2�Z��-$37x�)y��L&�]�QBe���mMV���^Z��j��<F	��m���`u�F�қ��06�+�zKJi��s^��j٩`��
�&2�� �u�m�u���L�GNP��w"I��Μ��e��WR
��CQ��1�[�K[�/��8Ѳ�� !����M8�bSn.�J�6c-njo��M�RP��_9.�����o�6h�J������)��9r�U���W�Ŗ*~aQූ�~;T��ֻ��z|?Ә'9�LN�Ӷ�&󪁈x�Z�,�%������H��,f\�<���#H������c���^v�}:K��?�뗮ݖљ�/���E!�D��h���)y��"9d����Q�����P�<{�q�,k$���h~�Y�{���/��(Őw��ɤp����r6�q��x?@�v�y�[�ԕ�F'6��(���G��OB�7�nG�)�J��ǽ"��>�˔Y�y��o�5Z��w�\o�]Y�i����˞%��J���P�B�z��p��>�:?R�S���0ɻ�e�CW�&�z�2� L����Z��U(t�P�n�~0A~'�ɴ�h^[^OҔ���ZAB�Q�B虿:EjD�1&�����r	�E`���;���"����k��7�l& ��^`A-�Aso�GY>��b�UAj����X*I^�A5D��O����s�69bvS�ٌ6C0 ٷ�`cs?t��6)�`�k�1��w�c������%E�ŕ�E_@ƕ;a�@��Q{�[��ڭc��O(�~-z��&�A��˪�Kg�p���{wz>.B��y7��»��;+�d�SůE���|ɧG7�F�T!{�kfj��Gl�h�M�MbJ��T	a�U@�Z��$�Ԣ")ÿ���j{�A˸%� T��X�8�3ѣ��,3Z�\A¦u�F��=גBOz��p���G�R�Ƹ8�蘛����-=��Q���1=��y��i�9��ѹz�4�A����b��s&"L1Z���0�R�xZE�k`�Sw�����}~�@���rQZ��)����,Ii*S8�������+��l/�Z� "k����^�1s�|�+��	���=@�G\��B][�N�n�۟g'�ZƦ�Ҫ��-|"���a�zR�B�*ʩÃ�+p8A*�IN)�l��J�9Tn�,��F�9웘�`3w�ABa����m�f*lZQ�h��V@+۬�W9?��Jv�v���Rz7¬��"XʨB��o��0���W��Rᅳ�"J�K��Xv�='D(mBe�Ԑ@_�s;�D�t ��-ހ�%���]���%1쏘����>򊔢<2Ձ�G�o�8rC��kk�,c��^��Ar��bՐ�]+K+3��T��	}���b���x©܊�_�ƘZfa��8��e#ҧ0q���s�\{�, �p��ق��jD؈�E�@�rk��%2
�s�PĤ�X�^�j7{R��Z�t�G�l���vT��9.~�͢���06��Z��x�1�%sQ�OG[[>/)�7��5��k�N�	D�dG����p����9�e�N�#��0�:���
8N>M�u�,?f�b.`3iQm����U�Q�m8"�V��"�8�Q*^���0�W�D��(��q�J���+��i���9�s��B?r�s��J�a�c�s�����R(�k���cԂ���7�g���&q�2&c��c�!����@�xnY��O.���;�ވ���x��Ӿx�s�"ϚD❌�����)cÜh˹��C���%cNE8Z�j�@EXa�|v�K����Ibbֲ�:ZK�>VzݵGX*]s�/_�ܑ���6O��n�H'�[�,s(�Ǩ��A����|�-0�F�b]r*��R��;�w�^'v��w�es�_l�
�5�df���K���5m�u4��g�$I~+v�DH�:�I��:$I���Fׯ�<R��cS=) �=��J��� O,��7ǵUi�;����gDuS���)�W���Y�G��	�j��<xN���ZQk�y2΂����I�����.�����q+R�,�7�:bn'�Q�M�`n�i0h�B��jE�?�r
O���%�����6L�8�oW�}M��%���a,y��6*��Yj'������"!7G���*&�j��;�2&���*�[�kSS�򶕔xAq�����}CDLV8���F�0OCd{��	��Y5?��{�!�^�2���4`�I~�(Iǽ4�}mJ�1�����	��;M-q2(r���ʘ��`K�Ή�j�-g�����fw�Em�4���\=x_!MK9TB
8�"z�X��*.��pm�è����
�Gj�-�#�����c�࢈��5�w���弴��k>A���Y�m,�Y2�A3�i���!��8f(y?±DG�F�̳\2�^SDʡ�)5i�w$���,%�%n��˥_���ߞ>�?H(m�}5�i#X[6Ew����(z�h&G�3�[�h��`��z��<�g|����2H ��fCU�E�4�_�)��e�]1��
xc�������^'�����eE+3��Ӝ�ϱ���N��������#jL<��_�b�C#B,�)�F�𘓝�H�"�b4�+>xͭ�PS�T����r5�&'Թ�Q�&u�3@��.NÏ2t�nF��*�^�>�E��B�1���f�F&Ӏn�!��3�[3]����Ϩ�}^�@vR]�~�"!��-�#nE~�/�f��r��J�}��ůÑx�?g�V���oZ$��nkR�W9�D�ߗº�O��(�`+�U�5�I��@�p�`w�?����)�ӑ%��ią��͘sO0���
��#X	-�ې���5��=蚛F��%=K��>B��Iw��z���=�}�K�^2�U=KׅԶe<�u���ZT��(�7EV_�cp����
2������&��W�|hΧ�.q�9����Gr`���������Ʌ�!泎Wӛ����N��|ʍϪ܄�gD&şڅ�A[���RXh�Z�;�%N#U_�\N�ny?D$����+� ~N�G��c�9J�� �����E�?�<u�:�g8�ei�i��Tޒ��68���V�	+g@�X��)�w��?����J�����<D��}B"��࢒_�iX����y)G�"�F*��ɐ^	W���2(���}�O�Cx릃��X�d%���lƇ�~>�qn�2�sb+@��)��e<��^��H��&�յ/��춳��h�ٻ����+��|��w����n�g�d�x43���@C�5��$2�l�>�����Y��}#���}���v�`Sp��I��D��h�L�~]o�6+�*���V�9N,d��؎RM�n^s6�9	��Fep�'5�'i�7� �u�֞�''T�G�UdO�Y��Ծl\m��Ur���y]�Ltit���0���eL�sHV�����(����!��Lm����P�����u��N��4���+ si������ȕ���[Q�c67��iG�X��te�`A�������-k���k��#,Vi�W<�3�w��8�6S(�+֪MC�T[&��2�w^���	�Scx�3��=�%̝�Ʃ�i<��G�*2CoA����]^X�JQ5���kA�qw1K��U�Ljג�Bi�3+a�%L���ɹئ�&��u�fߺ���2n���>�m�F�M��Փ��v�$�(��a$����	��^A�ޡl
To��U$'�:۰�U~"+Tu ��xU���p��K�7�Q�tH �#��p=��������Ȅ4f{c�S��"��R�P�mrٳ�� ��AQ=dد���- (�i�M���u�IP���%��Nؑ��Q�6��*"�MӞT��c�W5�����9*��OC����аy�g[c|ωkbw	<�mO �D�3�!0�����Ą9�?�b-~�]��d�m7u�Ĺm���M��ё�� ����5��=Q�ް٢��~��fɶ���������w6!��������nS��fj/!�aWe���'K�Ω�<T�fN4C�WA"�׻k���y.CLq�f6\��Rb��@�`�+?Ø*	ۂ�����"�|�J�]X�r�S�U+�G]�\"�dhx$c�BW���e:S'%&
��mnDS���41���������ڄ�>��q���Y'|��D�S�XC�NLb�����r��&6ܝ�V�Mnfq�#��Y��_�j)�z'�����hg�8���p��k&��i,�<ް�&�2"�����a[�e!?�ŜI�%p*��̱̬�+�H��$Cq
�m�Ջ�e	�G2�=g
p����u}W1/���Sq�����+��%~Y������Kx]�"ܤ/����'� �χ��T���s�x��"�THQ� ���_&mmp���(�����Ѐv��`2�Թ��6��U=ɚ���w dy8���4�<q��C��VF������=���\��/�<�d�\��;���d|@�+5|�����i2����g���ř���wp� =�Mma�ƭG]^u�HT�J!Y7�0���b|����1(F��1�:m����$���(wuP�B^�G5�^(�K�q�ͫ��=�J|6��­#�b)A�����dq��D���_�
�E�* �"D�����N�?a��(;��e6��1�VЦ��9�kH~��#Ԥ��=�3���Ew�2���{�|�n,F�Q��������j�O�,�S:L=p�rC�99%�/��΍���V�*8ÀA�[U��zIܙ���;�v��~�I�k�Y�꯺	�FB�g)}'��)=�=F�b�J�Et�tݎ�8��:uI��1�R�u�87��)Y_]XQ�"�00%BXt�;ط`E2�0%���DGڑ}0ɖ�_����mhj���j�xv�@X��x>�?�K��vb�����~N8Vfǆ��/�=OtPIg���j}I�4�V �K���{;�F�lW��o~<A;	��2QhY[��Y%�=?Z�3�3i!�{���Qw��r�{��2g��-J�nm|L:�׉�w)�lSA�큉
M	,��.�AxX��ٲ��%PE �����T��
~s�!�P�]#W�l�%���xуǭ��W��PBܘo�Si0�/�+��tI��螹��;�.�{zL��_s�w��T�1%Us��pR.Gh�r���Ҧf�����A�^.�3�9%ic�i#�Ͽ3va��"�a�rPo�A_ ���m^�6v���tqĀ�V��X�{Z��>���.��>�}�a���r��6#fZ���v��O �1Jh�f]�ߍXB�j�XKƤ	�&B�#e��c���B�t��Q�L-��i�\����z�!�,�Q�z^��e}o%8�o���=�>�|�����>'L(.N�#63� ?�ǣuY#/4�
�,9��[ ��Rۇ��:m7�S�I� �}�7H)�����aRȵB��L�hjų1�z�˥�P���E��"�L)�����3;h��
�Pm���7�8�Xd�ѠR�ů)T�K��?���x��2Y%���� d�*�9�b3f�X��/�����AQ����Έ*6� �nM�"���5[:�v�gԦ?���q�A[y�#Gi?�u)���gj<Z�}���z�C��^��y�z��]�1�G.�,���`��[��xԖ V��/�j�bO�����f�s=�|���%����b&B *<�&{�v:����
�Z��2���G	R�>�-H&S��E,�)ڄ7�w^k�&�vZ�Ь/��1xD���kH2~��]�1�qo�	���b�����^C�<�3�j���{c���'�'��ϧмK����K�ju#6j+��8H1K8E2�@D�V:�<��T��u�F���>��E�k��*_��0�
�x�������5v��
���(�ۢn�c�g�S�֢��t��8�j+o�Zx��x��O<�g��wΫ!k@�����F�E�^f���Z��_��ӕ�	 �*"OJ�['`Äݥ�S��ۋI�y�3������w:E/m/�g؊��g�&L�y3�������2��:��r>ux�����J������Y���UC����Ҳ٣��	�� ��q�)����=?��_I���\��JْK$��t(
;f���i����߃��y���rnX8�`^W_Ə�Κ�(ۥ��TD��T�~8�����f��f��&@�n��{dc�"�A�F�5�vX�]ؖP��ùb{�U�q��_�3)�NAL�.�N��^�@�$ޟ$ݸ�T��Pj�i2r����b��V���U��3�[_<�3g����L����F��Ӿ�^_��ƞ�ܰTQ�H~���i�r�ɍ���r^	��-�6�h�
�H��=�27Kg��b"zW���C�A!S�5�b%E��0�Ƣ¯��5�Whi5��z��xŉ��o�5���	�����Y�:|��u����&u���F��BśR	�n��]ہ�Y7��w(/^���T�|l~�x(�����a,o�qxu�x�6_nK�++)��j���
V�K$?A���%A��D�r���	;q��#q�F2��BrH��)���,�mG���WM0_-�"��͡��s���ކ�)>u��,`p���;S�P	[G��)��Px�Gcx�R�(���/.�њ����C���1x�Krp�����Wl����2O�H����O�PG�V.Own��Q���I�dԕ.��,\1-�����H?�r
��O�6m�;�fҿ�6��mx���t�67u��
(�aۍI����z6�4���+J��\�%��jk�Z�p��XZe���P��^���c�G0/������`�|�s7�8���0Gr}`-܏�{G��A�x;#6/*g5��ɆJ#�'��	mN�c�s��q���,��h)��e�%�`y)zR~E��Cqj,�����oӄ��=_1��ص�y}�h�T$d�-Q���xZ��,���c�{��y��z㹋[g;ʕ��恬w�c�W]�+����?�^�%F%Y���D��B:w����yV	6�-�7�~�o���������}Mf�[
:����w�a��e�=�=�W��W��\x.u0K]n����o���
�!r_p�v`�<�ddn���^�t&�����=�m���{N������ӡ�iS��?�V%�gm�2N4Y7���ݍ.snʏ1�d(%،��WT�X'�>q&�����9�7�2��DSM���V�`?%C6Sh�G#�?������(�1��1s���.�kI$h`YzݎI�É��h��}Ճ��A�)�#�3�Ԫ�~�,�1�=����o*�ʐ'� �,�rwX >�>���9���ԓw	���'���_�Qye��4������O�Q6�O���3��.�L1�;U��l�$��ѬX�D�J����a���ә�V3�d���`lX��z6�Y����{�*��;d��b��	��@�iM�J���*��^�o�/ڵ�������c.%Kx�@��T�1�iB�~�j'�}
�������׹|E�#�D�
�� �^�&�����$��w՗��23�r�mi�����&	�s��D�.��c�S�M��2S2_�G�kQ�F6��)B��
�m�H̄(�������A���Psa�5z����%�[�s���H���������Cz��z@�5��޿�b���\�~O�l;��[��Q���\�p��F���i�s���;ݱ�ʐѡ�g���)8t�(a���� *5d�v�]���d��tҼk�I��) ;5�uiΰ�� �����K��`!�(�������������	+y?7�1�3��z
W!Ӹ�#��1o������d���^�i��v8ڊ�Y�O�lA�] 8�8$�6]�
�:�qP���F�-��[������2p
��� =����ɢ��:�4cV|��$�($�<��z�m=j�l[t���EY�!�l�4����:y�vL���A-:�<ǹ�͂��)��ئ���1E�<�����He�q��Կ���ԸT4Ɖ��n�Q���NK����2_[R٣�MK��EB�6�J\�]��䐖1�A��`��s���/R�R��Ep�k|��5��� bI��E��e�8�HZ��~����N�=��.r��˩�Fk�op������Y��Iۘ���mF���l՗+��A���fsO�@������k�Q�[Ƨ���TUR�+�4t,��O������v�b�X��@��E�χk&����z�������|��K{$P0�!��wod�������#�F�}K�:����w�c�}�q�f��=Q��@.	�`?�H�y�%�s��� xs�iacoY��dz̽�KG��!����N24�0�딈���S�'��u'��a28�N���C<��hMB�U����h�z���6خ݊8بKb�Z�d��|�HNl�2YWZB��)!|gDxI��1�Q�O�r�"1F���d�vC��P+_��ϴ��G��oׂu���(�g��0g���jc�����N0�sa��~P��N$���˟Il�+�A��I���?�&�/ �9�����Z��n3Y`��9<ft�쉐"^Dm��������ec��~�[Cxmi+��#�&0l�{�������B��hO;�����?�i{`q Q�e�6m���]����,A�� I�"�c#�C�B��'����ϓ�;DQ��'��g���G�S�H��-�g�jJ�֌�$YU ����%�$� ��&��A���9�Ns��t��HHµ�\$�`�tBG��Z3��_�����la�?a��Oo(<��^��v���%��P%��k�r*�����%rG�m�� G�bc��t}N���W˫jf��I���.> U�ϽM8x�M�`4���\�k��Tq�-�
i����� p�����w]��wt��\)'�S�V/�C!�I^A��#�7�TG��'t�8&��vɽ�{R�4*W��)\*m����}O~��g�_[�h�����]���}�P����QQ3���0�ˇ�t�xi.��ka�ap5.c��z�4q��""�:��Yh6fZ-��=V@n�4�	Vp�-����g�r���k��;�ywQn]��tZa�]��bn��Q��	:�_'��D*�8�y��*������Q��"\]�x�����O�d��I�l[�~
�2I�3���~*�hdnz�&�Ӆ)�Y���Q�����[ �����i���l�z������ �=��uO9�@
z��t�"� ��2�z-=����.�j!v@��+Z�:��F�q��̑�g�)�AQ�/C�m��Ԯ�a������Um���j|b(ge�L�k�� �yC�©&έ���L���oN:�:,y�i�hlQ�(v(�D�E�d_��G{�B�i(��A�\�(��.N�g�AC�rJ�O �*ڬ�N��BR&���I#�����+r�
�4B����dI��<\�:'pP�[�~��K��]4�&