-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
BF0yNaq6qCor/UDeMbQno8jMD514ecTVirtTZQzh1b6YXR1o1cJOnbqPb9/kM2fr
QbCBZensDk5FKOY2Yewa3G8dupPujYYmZUdcTM/+PMzfY3M5GITyDltX8en2TURy
nMRHYUiH+EvSr2cvuAke/UVl3c+jYHXaLsDJJ9M9D+siUPskf/1ZpA==
--pragma protect end_key_block
--pragma protect digest_block
OS+UfkGqtePVqrEy30eD9yfM78k=
--pragma protect end_digest_block
--pragma protect data_block
Y/7zki07GcKToEnn+e6IZIsSxDkf5gdRWeFSi0roJRHNh22Tj6RffZ067rrn40DS
mgfX9E1jnIYy3nWt+qCJBDgTUke09GX9abaO485U3e4CcevjJxzhWhpOv225rY3C
DdwmAVbfLPcAAnU82iHU9w1BZFVbM8Wsyl+hqVJo7B4BlTaA/JqzHF6ddj0bpr8W
EjNhA/f4zyTiHSC+koq9GUFmxAxy/oYuKsS+h6eUDq3gp5LO06JPKvWbvbndSCMB
Az4WZOxMeMSea88Uir7Sw2RjLKJPAf0NCSMaUWYaDXQc2eHzHdkarfqmDSrAYntI
tR4yjgtBXYNCCFFQ8dPfkgYMYJBBzJ7rjDMYBGQ1z5flGQ+Alpmbr44dTk84yXW7
OQCq/Fuf8g4melWk1JhzH7X+PkvpJWF5dVqHk8jAhHN4qrTBh1CeRR9kZ4ZxQs/J
bBWXWVlVIKszhxe2nXIloy1x3tPSXtEX0mNjfUOP7Rb6tqAEO6HjUOxvtm9T6DeD
E7NgVjgx/FkDTKVZfgokf2xVnY7SJjSTnKolfZ7EsH7eyBmU22eUnXY20wVRylyh
qbtSm8myrFx8B2XRXwJu+JlhJ3o1zbfeRMvTUleWNdhx40d7UtFc5xHSXCBLH3Ni
ca9Yrmad0NJmw2pJxJjiO28v77xXZz2ZHhKhaL5mup741qHtoujQokyd6/the1FL
jN+9ZgeNlIzEw0RCIXmtoq4uIy0hMfvdhi9ldMwC+SpGlT0ZbTu4RbPIdN/YU95i
R9PMNBu5M3cEXEv/HOtIWPnNfLTmjnWGsQkZyG2ox3MnHYMWRlEuzPCd2i9tBfjb
Gil4AjVSFStqH4fRgkbzWiZQsnU6GXMxY2t31A+NfK7QDGhsWne5MwuI3Un7xTwi
YhX3phVu2QOdJIupYCnfFi7u8qa8ofH4x9Ym14/hkl6N9wACkRl3InKF7LsXC6e2
utc8R6yNvCLGzDrUpabO5IjmacYNOzyUtmKFdttuqcg9y+QQmDWcoyNDAPxshNTu
7elO8WjX+BD87UUqY9SHIEhnmCKvROzftnCpzra4LeBsVa946nuaLZBo4IVRWI7S
xj1CzjxALUUWcfwhJFPalj6BCBbjfWMsyXeEBichYNCQWmbU1NIMstua/shS+GwL
zqv6SDGOow/DxYeOqDNlmZ/goQ9U3NuIe0Ff7b07eDWyv1p0eVuz6Thr54hNws8z
Xycc0BnaMlcmWgSJE9ooq2sIZ2sX9kwS0v5Yr/WY76SF0Uu8R2KA1Mrpkzk5Yc9h
erRB4F7uYcAzJzWjmzg/Fwes9bvKwxUQC5GL0vMpv1Y+A99BjtpCn5+hvYdvqwBH
FMd8xN1KC5JeiTTPAboexlayWze/dJ+AwGujSd6mVlx7Epe587PruKwWki+njKuA
wP9UkWWC/UIL9o8/KBe+G9kY6y6fciwY3HZvsxD4i0xrc/RXi2W7gVKhbS1BKBsZ
njqXPK5JE6HQh7afqhfRivSFBzfh/1vQo/cLhUlyCBgXWVNgqC5F0FOPt4EMXzqi
sT/Cz42jbHqcEumXLhG1YdhsxrJCXOacscJQin0yLBVrdfX8poK/Mu9gDWICU3Ma
FETGADVuobdHaN5PYBHr80f0OlnzTe4GhIWpzwgY2WYS63PsGJRZJCw7On8iOzcV
Z8YdQ3PLnbaHRZk56YtTALJlxbtRfl8trKOxGKe80QYRjKCUY5jajQEM+JS3bOQE
d3EjrOLGQlQkac/ZJpzSyBrqPrdJbIzBVCcZX/MiVM1cCPNI7mh6mhpuIUxgYVho
DNNRLCfC1I9C5WJiDwUWe284C1M/nzJJ6vgfPdU3duwiJapLRvIMyOz9KOVesgPk
YAiGakkMuK6GRw8LwGxmv/PEKviFkYyBxZpDU32lfnFs3POQ9qaVL1lQN5UgrnQX
pIDqFCP7upzujBciyaTi/Z05rw4+G60HwIoYak1FouNiMfATOqT1kbONNOBvUCFQ
Gl19VPP1LDHGqGymb2heVD/ZuYjeZLxXJ/lmD9zZLibO0D6+3oqPpRnUUe8gadRc
496OBt6Ta5ARprVFWeC5UMG2HOqgwImmWKV85vuoK1SNc0te1xQ/jZHOJIRgOgC3
Ondt64MgCg/o3hTwOJQeYEuyMd+QKlYuca4nyXCXc3UA/wvqmK+59EyWsoS0ssI7
Jw3QnFHJJvaeIK1jrmZ7+bo0w/MbR/g0gUY31UutEFe/ZvOrjJ8WzIudFiOckPz1
M7WymXIM8fBcAwyye09tOt5et4n/mNL3RON4QcWjRb1Vr7yHTXk5RcHgaNzMY4UO
LBkZodGG1ICgDWfR0b2vGtyYdfx2pBBB2a8QLl/PlTs7vc8FgieAcAj/abie1m2z
h86+k7PqWuDfzi3jl6J3fa06ofRPRzcgRSjptVw8yWAFFL9A+lkMKWEBymHOiCFX
TXc3/x+FWxyUEmtrqxjxrZBsbhBMgL4pPWOj4j3XsBEBmCCxd1wqYQg2cjYBUTO2
lOLfPEjhbdr3yomtdFqQ4PTJrTSIXE53UiQXjbvyCviyw9PuyJNKUgbzj2eUllzf
Z6w8UnE3G32cFgpdiITfbG1HvYN8CfVPilAM8TOKxuIZ9SLmVle/abYJ6xkd0cvb
uejnoeDeiungnFQ0V4G3wumx+w2SWdYG3985U76rm1Npoizll+hKJDfsiE1gjeMT
K4CGiUHw3VzGf9aYdy6GadhkRsnuDf8Q4ypVVejxVluewfkRavFIZgaWRrmB4k92
gmMreQNlMrY8RVq/WSQkbLDeQQBiwelRSXjxwzjmuE/FUWo9VjQm8whlsKOKOzkN
ofqmtb0h0Ggsr7GdLlz5/oUnmiRBM4KbJuVhNIv46ePEIoUyqwsFTdJcdcTFiyse
E+DhPvgNHQEdGAI0CDgNX9a1dN8R2hH4cGpg4FFum2JDnEHEixQMrZvKVKzAhpER
dxDSX6MsQYnaHEqEvdPKnbUxaek1XnV3mp6xhneMW0EhaRqrDuwc6r0DDqswXrWm
OLYIsLYKcectSzzTivY0KMXovosOnLxBs2kiQzMH2ph7WZeEkSU/m6VQwyris22o
kIECJYKXjV2rjGlTCFGJ7S1OA/SRcSUoes6PbXXwXFPx04/dZrQdMCRIr0FAcOlI
hAz8sg0TMnCjMNGz7sU0GE0hS57WRr5fVKE6aSVi38JhfryagisdIruz0jedUB5p
Jj5/ZBRzyHYcTZw7WFwIQ34yOzl4AypdNPaFbMpoWAVqosiWh5zZL7Q1HZ9Sy2+k
Ra/hHE6RRYl0Xf7ryPUGLVMny0jos75L5b3dJMPfn31WFhMm13CjKkry3DC7W11K
4fVNM7bssBvoimIVaDaZvwCd+MI9PlPVVs2/dXY49tBDoNCHQcHD55KxhihsQG1n
pkBDoOr4gAzP4txht5qqAuVHHv9ePklFyvQKpxAtEGRVz1EiUI6NmzhE6/Cz+DHS
piGV56f0eeg4SPNeE8b/VQFuym/mJ4dFWORxZtPRVYmTzb1IaqccbeE2PyIkWvZz
W8iiStYVPmoAT9i3pnSvxDmmDwuvZe8coxzV8FlI35FSGPZE77ButCtlfCVtxGgf
zIrW69lO5RbH22zJpD8xTTJBXSf3HjCwyNHXegV/AI5M7mFMwF0psNoxTIN6lR3L
goQBBz9LL71jwZ1Vit+YBrVCEM1gTo1gSKi60YOVCMCioQajXKqrYzMmHHi5TP9S
9CT01iKAncSAxFr5+gP1NrF4JsUZl7QdnxyPF8/35CU2gfYf0Nv/TKMnakSTZI+n
9QnpjDkAKtR+m/9b9mavI+Lz8GptfME4jMeWUOy6qVJpeBT1+OjxIZtmBsbq2BKI
SDUoIN63aKsHYXp8EUoNu7Yybf/mW2C2xvYNJp19siGiOV4LPRzHIwB8lOWlO7/j
TaeqeiihNJEZCJeQtpHzqSujgsAl5vI0P/MAT0jsaUxR/e3x8Hz+4eUMipryxg44
73uNETGV+FU3DUPb2RXKedOGfcANELKG9ggljLRz81KQsBHOQ4P4skuyIMil9f8f
NF109VmaUxKp6UtRLv1p+85LYik6Xdj/oUZP6ff0AFoHsaNDl5hBrU69lnNKqulF
J9AKHtH/Q1mnYmPnx11gGPNJ2sRr7wACwbUrfi9elRYabvTLQKL97SJ7TDC2/vCt
dGwENga6LuwT1Yid/yhB3YB2dD2t5yCqdBReV7BmjvTe662oQgTH4bIDvYYHfO1m
onh+RaCNN9St2KYuyEou5D7JW2O6bp381K/xF6KZrtXPJKGWISWc+Ock+BedAHmf
DcMb4gQ2REjmZgbgKQZbn+ZBTxKY2yG9g53Bjw8KMVVyd470jVDXnfds3BfGbUkI
yH7T6qLpErSIqmJqO/kabxYf/6i1jPqCaG7PXl58ZMmMTvLVM3YUKCQJGiMboxU3
uELwgtydFqpU7QU9rRVpum3yKF956Z5q8JLUa38Nms/IQACGQMpbq9R/fjLe5Mrc
ZBhb561QJhoVPVnyPidg81wgXEUDST1RHsS/PdXpdDw3L6EQiICyEq9IbPMFivFR
CeT0qIA0CxunwpLTS0fMRfQ76L277CjstqACCkfJ9N314/qQUHVlIRRi2KHzqcoj
XbdfZLY7P/uLCPyJqVzK0cuO84bnVCIUUZdL/uT7Xi1aXkU9AHyqqj+O7ijSXq8Y
KiB+EMApqdpkf/i4/oHVtLwuDilyBlKlBWHPVqgI/ElFwmoAC7NbVukneAp/cboz
73EhMMOqDmk8mSjs379wq4YPuR6uSXtbClMasGaLkubaIqFP71dCAuiYoI5eIn3e
uBbTmERRcfTDklgNp0MUN7yl3Dd4f4NNIC5KtWk4XHuLaerZaP9ti3tCl5RBfpks
YteAbCRenL6HKHI+A4+am763p9OXZDnT18M7CoyccMAlQ+jM0qlDoIubYlV1Z8BW
+mn0U3/wFQqzoMVBmZetJqILVdLAZrd2+roMgaJqyodvBBs3tSKIa3RtHei54lpf
HhYZG30uukqWaqO323iOrgSTm5OgIjmcJR417Ecx7hcQVIXCWc0i+oybsFlywBSi
4uMlSQNHURTqBnVjtmsiSq1qDHoi327iPooGF1LrF9/ejvbEGxNtr6SwZ8YIt8Qi
4p7bUOcQMBZQ7DEuVVdgvPhpPMjWO4RICcJwHDZiUmlGeWFljnWiO1g+t5qyYIO2
3+e6PI1POq43PpF0dlkewKAKgSJImyI/LwOsL0iF9uKpTSr7gWAI+qCFhLVeBuPI
+QLJKb1mTF9BEi/TUuIe2sdS5q25mAo0uD0+xs269QcMk7p6k2zx1TObxvNxWW/c
MwtLqCStyy7tdaqg8n+3uLWlKB0pKjfAzvEbhLyMg9QzDs9RO8UYvzqbLAM60ExC
CpBbK6aAIHjILSkm8PJIoHRUcdh9yFFpIw1GMq4sjpeeKQTPsRpRn5t4VuPsR+nX
VY3P4f+F4EX2mSJ2NjSK8pDQIre0LTT3iOIDP0XkbsK1MUh3GnOWnDz1OurArEZk
X9DRhf9NkcOCUZ1GnaQGm8i1FYUD0GdXb858PBtVhVqXOZwov7uNqThmlnLYF43P
JKwLYMWqsQSUUQdEELGqCFL6Uz2geBM81HCf9VcwZYmacrhNBjcS3g9noePMVCq9
cL56xBIjWXTWf5Y59I4JnvokhtpHZpWNLFxdsgs9p3H/fdEM2HjdcBp1FyPm9XSI
GQRn7f/LdMLp38wRtAY6T2Ca5txKmQKMQcSG7ZTLMMXuPM4dN5sm4eMLWRStqxmC
uLV6Il+kybkQqmLwg587CPY7Ih4MqPHmF333Ue/NlzAMn8grtWXBrYjpnThzRjJO
2BK3QXsFxfNKl6Z54N3jvKWFZus5/Ndi9PLWN4dcxGe8/+nl0sAPiCT0OCWw4P/h
BlCBxi01ZW061599arOSCLJ97e3Arz2luUxrk4gikbcTr3id9X4ZT4cLs+X0hqLn
8MCkpaNZbL9FG8vkjNM/BlUSQl7KPl2UGw8CxKAw8yI9rta9PkUscdvLSb8xC0cS
xKSKUjGo563bQCJJU7RB0NDbgFXsAeaZ6jCcxjJx8oBBH8EqPn8ZfJd4QBXfC6cs
/y5sOdz1lFmUqvBq9MRCxXDKNvucO7m1QeAnMZZzr7XciH2r8rn+5LP+7s6/5N79
haGG+Vg83PvWTaktCW5EYM2m1z26pCkXx2hHCIdXgPb2k9nCge/MPLmaiBSYqtGd
WTdkQ0nv4+XmLVxaa60DwDc+LMOOCwLhFEbbV3W2u/v/vJEqcRo+hFLfjt4ROz41
GsRvU4aY4B85Ce8KVSThdjbueR7D3J5nvK+A/3xfDCC8q9/vvZeoWNcSoeN3zbSJ
3pka7vZ2VsFK30LaxF8q+Wbs+kPOHLM42YaYdf4crs3wXcIbXajpu2zxf6M3aN5y
lHOSqO5TssSF+/y/yjqSjZLIvB/i036UxYJL/KYhAlgX2l20CRWXwUyQLdsJxMiK
K4DuEfCcaXtkLgJls/YDJ3Bd8r6DPUnOr/ZVVBUBa3JXEo8llD84wcz38p1lHsKa
UD5Lz6HNto8WUM4ixEQxRR59l1ZVd96BvkBviU+W6/eDBchRHTiS72uko2/WCYzM
Y9mmDljSVS2/U7aJOGRoKGqr1k0rm1vk6AJzIPUoAwWFw7Iiv+c/+PeaGW2z6uBn
zKVqMS5dFSakKVjYCm8IrONSy2/C0XkRS9tWlZCHN64ENOD0YW3E/1S52GVCThG0
55I6L9kuTSdOGfapcikVJ/bUrymu8yDYfNVPwEL4Uh9KoGFmNPaEtgJeQl+qnuy9
P8gnNr5pwq2LVy3rR8zlTrI0r5uywY8gsKuzg4ewFEKX+skeZTJSB+gnHQZEkfpQ
7J/4RdZrD4MvYPiyJW9jsSCHK+JtOK55QxTDwzXR1UaLR0GtM2YpM6lTf+LIXxHP
PREpBKDb7mkH90zHMMp0/lDZOmNPvyASh9287N2lx0COfJKEF53PaqXopq4tq1dr
9k6iHVBipHyJEPArt4KPPAGCXLaC6Yl4NU19I1H+6fj57R/2Et/SmQEtFCORXeJf
vSdz9UJzNBQNWqtLVItudsYCpCdvExmV/QnB2XR4ENQt6MUvOIekbAtHW+0Gf3Mw
chZnn7Ut6unMCgs1pLvw+dH7rE2xIU4DqQGd83sye8LnQQ+Zm4Wmfx8hT6xiT4UV
C1TSh0Xrvj4lp8WRWQ4mOD0ZrHSYWLvBdOWG3/FX3Wj57+1fm2B/g/un/xhXSXEJ
UiQyv5BrGtPI+woWjWuRhVQPNeiqOUwUn6M6Ytd/XaoJmRbv7qVBmI0rIZHy04OW
Ry/VsHoVAgCmFfCv/gI6jYSUwb1Jpb9HYfWA9rHR5rAkq6twsbLdRz+qvGzw9+9i
Sh0Od9NCQ6b4leoI8NYV/JBRNDghyhwvn3psovipFCLWxGxfczhDiHsM7JMsqIEJ
5aqNsLg7Kc8JsiluAOg75fP3kXNS2t7vKO33FXb+QZGQBg58hsSdlMETbx3RxB1g
6CDjQjA22UfeW1Jj1sdaf2KorJ6wDBRAd6XH8t+a3QlEtPHjdauVC8jy1t/hfUCm
C4Km4MZZRyE73yOeY8xHDB2GMBjWJr4y3N4mtv4GgDya/SerctW9I7/8y8LExoSm
I1ejhCMfYjC4w2WzZKtsy/ZcGVO11B0gHNL0yu/sdFjXQQ87/6KF+7P396T4TBzt
RPK0+kXu2jb0LP1Jbcz/+ob4Jv9qm1gixWNFeU+2r9KQUaGl63nkR9l27yAlT1J9
ld2Zb9SMBVVfgYw3nmXjmkzFTEBWv/TaldXTWDOOdcvvtKl2bEJqHVGI6Jnvl5n5
pWUFbP7vLE4Gpl0Q0vAvoEBPqzt5vTDLCTdmHLmP6jqMthV5IPa/Nv01VlDh5W7S
mltUMDf9KW3cGy8l33swtzkQEJ3a0nuaHWFnIdMS4ATlaAJrDuKWh/XN7OHm4YFn
dYogRs9FVOU++/Wl8rfRutAIu7PuT82n5HcE/r/bGBYwEcGY4kmKM/pbjm90iidc
VYtLJ9aBUayiw5DTKrcAzirtCtA8bT2xWzpO7Hj1gDLWVaq739SL28wnnX6aV5m5
rX8h/s4NnFqcbBdJ40Oaj3s+p1Y0tWZ5hEg0xDYoF9UYJ3UTiOZcyQSMY3GEwB+1
SjthrGlA2EYOEyXeyqxpB+9hCH7N6XuwehhcJuDluYivDDisfRXzAbdbITJtjAs+
w0K0EXpYpIoQ8dE7sGFfFC0vkLStrMvI9PMHqyZyXkchCHepEUWeNBTEyn8aYprk
z9gOvH5X7uEZqkcaBwBjm1vjqe84GbCuQTEgGrnHKkKmsWJNyiFMx7rV64zluQn7
EAhFlKCX5GMQNZMCxq51BZZB8vHvLocaV6bnETSz0++9MWglGtZ90ywKNgJ+w8Zg
SBlBomb+Bu9ggua0pHdECDdd6ashrOxEZUWHgbDhxE+lho1pf0Os09muszKtBc3P
6mlpgW83vUoLDNBwlN0SF/P+ahKSzk9uUSFomFP04h0DA1qAoDg5Ii5hP/KaNsRU
T3WpJpblXaIfqFVeE+sqx9n1knDBerATThWQPEGLjghqC7vQ9V0+RZ46xGC9c2hh
1hIBcXRI4SvMy+2f9Cj9NAeEKlYHr97JHs7D5nISadcLgmZIehh7hHj/h60C+Z94
NzYPnlHF4EYMSZ2/w25u/UnmohAE0WcJpFppFAJCqWJxbNEh+FXYdyLmCSwvekRh
iAmNS3SlXPzBe8wzfYGu0wx3awpVml+V9qd7eL5Z/avbJJgprhYJi5XP5uP6hEhy
UTikSbfIcs7M5JRU+mTJmGeHuMdl31QbqAXcxBaax3Sixpqj4Z5eaqZv5l3rHkoS
kNpfkukCmtkjM9HLAGv8uY2Ci+D5CxRUtajlu8dwWq8+kYd7so8+b1OvzedmPHJA
6t7oN3ri066nq2MN+0k3chaQrIlhfBdSFmIIg0yTpvUygpHX0iUtD2tEck2zO9O6
hKbSJGPV3Wz9n/fIU0/Rv5uniAiOP1rK2+fpVexNcyKJt6dUA4bDQn0kmyvyy2y0
Ij0uyY7lz5Rp75LWfjtpmlR2DXJ0KbLVrlY3zPEVVRmDXk65By1LT+q6sjJCS9Uk
DDUKs/P/Gkbr7OyTM4QOc3GZ+J6LS7TA/dpvSKoSAhgUbOxHhncVvjN+jbNRVyRA
wpaq0W1gxHM/f1kYzLYivAAyYJlGj5zJ66FvmpZzprCl+4TIFB28HGsmpGhG0wAj
FX5XSZ88lO1Rq6FUPR0XcPb+Kz0e3fQQZPhxQiD2TTNw3TqPqVBYs7VIB1zEatF6
iZoDBjvEYxgDDJwR3eRvTwi61D6hMmGrFieQDPxnJMHRM4k71WbzBpNEn6Q8HXRd
XMyRrKEzUzbO0oODlEM4SoseCsXxPqxBFTSMTRo/lhgq2XOoLq0PeuR2BC4yQIeS
33TAa3Nqwmi9H8ITmII4z2QiAp3DaZNw5mV2owlFwjRKP4KAIHjnN8ozQ9vqOVEp
nyWQamDsYRwZ388UnoWL9doOGOIOSB6gymtvNuk0QrI8TteotBQelxPMu0TIYNsS
S7j6HwKbqSUHrCi/24Na7g3uEJxg9bCIsDQdz08pK3DDLgs8QvC1Nu0A2XYekUtZ
56uoSlHXD8JeZqi0Tj69GaF5mDPeqTLAAEhSeXFvqgLFotZuDt9GJreuZaT+Llxy
APhE/9+DQkVeIVmLw5OBb05WBzWl9z3cjeE45UMx+lgkG/QKxAq4ciipZLSTFO0c
U5WEI4guf/k/zddj/yER88zxejDaNRnQoBXgTdSTG9qjrv6AqfzMT49zxsCMJzyn
wK+myg5FvjBrM7O6o/DN6zhVgPsj30r+fVOwzEbi29A6plsIAcj9QYghrBrqdciC
BKLdb/ayj/LD6ubng+o8FmOVRpC048UrG4VwIoh8RZwT2zbWil6iPjevBCeeKw1Q
xwX/8ElDJWRLp/YH3npDgJBkpqinNjrIYz/jWvzxskdN4yxIdFbrYgOTXGuLo6Hq
/F1/pohUwSUMdat+O48wvI7gnKcE/ET0MoHISnJ3j+S/8SGnTCqFRgxA4X6O8bR+
I5Hq88+fKQl4QiCKtRgRFmqWd5CtxPSmChJlJL1g3KB4rHMeCA7sbhlmjRuM8wTO
jt62/2XkEQcL893um6FGc9zo950D7Yzg+jQTGah/Qdqkc0xKQTthq+2tBA0ayCsZ
lopkFgHKiYbHdw+61Bqiy0p3KbK681WVY6FbTqjEr01H12UfQXx0vtHL7JLBaxdg
2tbgLorcg2OchdBoA9OM4fzHRUo/+ntPxwe+XMf7IbuLH8hLNLmLICY2CpTxiabp
SE8RQL5CvVaw5kTIDQBf0dmKxE4wQ5I2Hl6/OfVWtObXHkyxLXQzyzvC+j17lWFb
8hzmqMyuMbgF0rD9tL6zcYeec7FEkw2Azc41JDyluKbkMDg5Lo8Xh6F1bTCU/uV9
pG9dblqYgUe5inguni4LJAazZTSzk0otYQq3IrKR+op/tX+qzM13nqQGqDWTBEyq
UQeCzHVb21Yjpgy6UidybPl8zhcWC66YfNqBy/iUHJI8ZapMafUDsLj8gHD2pwt2
IfkBOvQzUhcIJyvrcJ9VDVFwqPcTupkTa7An9Dylw1rj9zEyPJnwmuqGiqi7zCjn
/WYokBuo4cc2ZgNygaq9vii8UwMNn4CyNHaz/OjCOMeo3r+cscYEc7CnSfkbLtNd
S69TsHACddd+BxGcFyA73yJVB2RlKbXUPnsNcsvNfzKDaL0+IOfl8rYUq8JmBe9d
hU9yNWZ7IVAYO6iedbxLlxyBmD9l2Dqqzg6h/gq14S8oa4qQPZQMYjQORiagnqWw
hGlNHME3tXvNRncNP/zrbxcX6xMJL02ZiMmYYxyjBxBqwGJLajftH8Omt0QeO8ih
Khm65U7sC1zRxiGos/sagHxU3tOA2319tvnXmWY7EEWkW26iSM2Zqmbo7tB6ACzg
c9Q3VoCzh+ppzErrirGHvYYXUSG3+1cBVwVxQ4Hzvy3IDxiOJHiLsgFnxkQL095b
DVfGHintyL8jTkaEAX4FEZEunh3US2BvUl5jw/PSe1E0xlDKjoeAySvwK/eRrk3o
pYIl811yj8IP96kmwIqJ72p7R7eBrIlxx9we676a4Ntoll8OBnDFP5SaZ2LGOIe6
oMQ+vzbDa811TuhQpw1wYgM7PKsSnl9wRYbCjf/N724rOgYZhHUnSKFc/ZjeE2Ld
arm1mWRhoKW2qy15D+NHkZdSYXixrcUW/6vlxSgRmP5+hfWIdSnJM/6bfSBCLeJV
tXfyO4C96cGpDvVPpB8mNipl6UuoBjWcF6UR4cVLMxIEZvhKK7NXu7gfJ2cTJo4O
AiKUScNfT/MZt25bFp3hnIZG6lVeRbSpQZBVWEkRjPWptyVEnr3Jh8P84W3zS4/M
acuSFkJGkvs1XG+U2L+A975/ZLD1BLFdkp36xiMuHDJP3VFFu8IjgvlVeKv5n1VF
OBHtCMT5Ou8ZA2sF98WsWq9ciTpJ+l6f8N+0zZYIJpHkhiiNegpUP3gEhz1LrLaE
M78MhGw8xMNf5Hze0dev9yGJzzS/xia/5Gzb5jB+LJnd0JzyoAOCPW1mHvKnrT31
YRDiYyjO9b2b3KJYZK8LqnP1XPf3BwjtO2nK1q3rLHh2ujDVVmOdGREsA+qxYtHS
Gysh0UmhylPChQ4GupzejqbwijYBPq5O9kwu00w+rahBe/03TBFZK/RCaL1Rna+2
8RWscomneABvc00/aMyUYC0zMNhmPLfQjQwPklY3gDewhZORp2XAKXLNASjzGf02
FqSDlIjYs/ZWV8yqpY9/+Pb7J0sz66FCFAQaC7ry8dfAJzWixbvabcIEqCzYZC86
3oghmNoboMpGP+xeZmp/FWBkIOMbBka9WQRL+xO9y5bIklZvaGcJkgJfQ/S6tJIw
79pauAdRlxh8YqGzc2gP+qpSg2fd2inhyUpPTiUHvH/pexxovZ39gdmBwl/2nhSS
yPat4HM5UVNd0Zfr3O15M/7DYIRbJGxbHYC3+DW7J+bJ4sfGWmdMOAZFJ2QygYs+
FyLgflUZ7BKkTVWbRCckteV0bK4qrmX4kKPbYsrIlZZrpJFVAGzcfuy12KEUaId+
rfl7Xxky+h3PDnfXFA2yIK5yJ9T5o5Jk+XtyvuR+vdLS6bpwl7FEeezPzS/ZSWro
z9xJRVf4MvUevJNd975/poMWmJlyYL6PYO44OnvutBLGdpXM6LmR1EEGKz7V3PL3
6s53hwPZxQFtCIaesYqHCl5CZVXtu4R0T02lD54vD3PiJm1Hnshw+YzltqsacljO
UDvXuvR2zwf8OdC/L0restATxTPc2DVPhHy5nS7SzKrMoXIvNxWUAGXYsVZd4Top
hS1H5JD6I02Kl5ueUk/oUg97tpZxD5rsBVRxo56Jb1HApC4e81yskTKVUa6MBj27
FFWkKCpQ5YsUWdgqOeLzusranQ0lqO7hML2IKxlf79DNgD7F9F8i21ObGQSSu5Oj
GfjLBEtgjRBvnR/vjndwb47wCPbTf1jRIjGi/9fyvAKvAGeWlRRy7rP54UcHha5c
RrMrVIH3y/5BJ8zr/Ocx356Rx/tgFI1Dx9fOQV/Lfi5bJyLO80e2FLMDrvP7RcY/
FxL+wGUw+6BV3YOynGDP5GUjwFNd7aTRN09aCnpoWgiq8hPYlN7ghPMnO+ha5e8K
K7HyqHKRwdiIwDL/i3at0bmataqUKbgBEDn4CjZA3+taF8Om20jTySbWQwhsGFbu
ntNxkyUlJxfjVeB/fnxKGwBA1uBXy0KdcRF6Jf8/x9ngFjrK0FKbmCZjDWM8dXIr
C4ZNPpufXR7StmMSVX6vfl/QHQ8W4lZ1fuvNRji8CeiMLoL9Rtl6f6El7/Wd8985
FiLDIE6yJzWrEXRGh4NFgbuLENqwDVQ2v9+wsQ+RM/QriH1m76amsK3loVqjWpC7
tM+ylgyCGMBRraa8/M7vG8Ms3p+Rk7Ol2RrEK5Sq8XnvEzYgZys9ts1t9pFhcXvR
7bsytJDPYE7LIEvP16lQquAR0Rht9vPtGYma69lCTeuSCQuRYma8EF3whfQ6A/rJ
dzwtIrSIDcWD3atL/Bk0OVKb7tECrLQeypKJYRw6gb+p/u89EdSg7CZqiDf/MZgA
w/Hxlnky7+fswqSE/gc7SM2kqVuuA56E7dcOir96uBpia/jKgLUY/3khmje5AHOh
f3lXrWmzWrkGkOCTqxDn+PrGE5/CTgu8m4rW4x0XHu2URN1Y2qrz05x4zV/rYyhM
o6HTm4IM7LqsRw/Txcj4hMJnxYYlHsZ9yJSmvsA9h5fB+DqSTYLWzbvflRpVCMk1
RDQzswYyUL9Ues2lvXyeW7tZW2I7BQ8c5X35tXPZbNhyHqT7nhAN71nTGHEUrQHn
NxHDNGJd2PeOESyA9MUujw5JteIxGjGvsZrIX4HaN3zqb0QlSUPseJUFAKQCV3jj
/bY6/OSjAfXhXmDRS8vZtDWk3xy3GZqFUq3SZ3BU9FC3VYyZ/BoUmWhFU0dYoS77
XEOOjQksO6ym9YYpplxQr9z/kDBiEr2IZl6/HDN1RPqvROqvkHPzRrxbOzKQiKl6
FxmO3tiB2HTda7PFxvx3skS0Wme+IQIbXu5wQGb1hSHxi3ebjrRbFN5QFnbaxa8R
qmb/cVrsZyDAWFM4lP2cXnlm5y/elYAe+0KFZkW+bTCFYRnOGUn9GiLp2sH2hST6
0m3X8yg2iENEwtp32xib4aqz80dTOPQz0PiOkhERiQ0AIkvIfPwsyMkBFkmxIplz
X8xZEY3OFiHWzY8cV1kUQetiSUgQbOGPE3Lbvbc3lZFDeK0HChzGzhXer2TL9949
EpTft54aBbP5/0ai4RZcEE/3qQHazaNZy6+QT0ZeT2iagZeog3H5KQzIMKJt43pu
7P0xfIFCVsS5ScrAwgkDRalgVQd3IvitmgBr4VT6tmPN66L/4osTHkYJKIlqcHzM
ytLeWY6QWX3tuRu93x2CzK9p+1xRGqFGE/bgMsbKALV7UFFDOvdS3KRZar0I9j5B
xgNcz0kiGlV6R6E1+mhxHFqbwxXgJHV8WpK4RBjz+B4R+9Z23GBOZhCDaWjNSrhV
NGmaqRZXY7LfGL6BZNO0nimiXhHSKlhiXVP3U6zUqgiT5wBpU1pb3zS812qaburi
mGs0oZtYCZl03367XuUqT+o3mtYOF7zMrcIljk35760h907TObRU9kiv7PlQMiYR
gq2tYsJAHi9e7GsvnEoaMoAn89DZCVD7yY5fyrqBgg6FqiwLswlPdVwAl/e9H0Cz
h5i1bBAAldBNXVV4xezCji220PQrMo+GseTg7su8oVI7TprxRnP5IrI4rJaFAZBl
iWPHR2rgaJb6Lcpfp2GoFqQoNYm8CMuufyvTE/L98b9PgRwL257k6G33eDEFeMui
Ncnpxz2jP/1UFM8QGeGV134A1LNcW0+ZbrypAedrgXNN6jbRPMSVhKrOkGaNhqB0
k/P1Km0ipQiGbiA9vCAf6p/pBGJMg/4mGFh7VkaV+loh+P3hcHdJtC/a53sxfO+y
5A21SHUuFKDFKCfgdHQL3D2WtIypRHpubVsvM60uLfRmwv5w4EB6IXuQ613g4MaB
Bg9QIMWcjLEjks2ecxgxY5kE5Q1AOaTrG9oFZcMrXDadUKIZqoPLYQkofGpRz5/h
UI1V7C1oGQRaYhhbEOvR9DnP2MnReYnJRzkMuRTCfOAr/g9oYo9VF1UZLwMFMGS8
HhFEjphBsra8IPE6r7ZEETLSo3iDDyMiLn4yrNbn0Pp8vdL9ygPGXubHVFW+1Mch
U3tT268m/0Gokj6F2/PgZr8RdJqXRw5pHhYJYHQRnEl56Ox7U3GbQjia4PUblW6B
pmvPEWnzKrFRYqbcVNB0YYaUa2DNHniulGAhD/J3SNNCynzI2mNjLoqkdC2tIewG
CR1MJmB7v6X1z52DOE/Om1cuJYjTTzm6tJvqHeJrmLEEV7G8nERJ+QSRlCr1BGP2
fSzPVN9HNtEA9UcQeGOCvnSFxAkyslA9J0C2wHQ4VxQPow6lWtlghM3pRxbg6dgc
5/rGEuoVEpUrqU2M1sbMAsMVWpAbDa08F45IDSDOI0TtakWI1fWauZJt78uNSBet
1mEDl/zHCP70p0futZ9pOKiMWM6gl7a+dJKc2fdKYzMuLB8FNK3QINXrM1yY7cMd
XD/coUeqhh/YWYmquclcs+zYAL/MDrnqe1wJwLYgy6CKtL5ac+ILxa1T9j+46Obv
ZNDEKtw2gkuldvlz53rLIBifByO2/w3gJRKxrXGADGSH1sT+eqdeJGXJbGjs9xmW
VKZkrtrSQyvwh2LQZgNwNZc3S6mEZaibH9mPTi3ZjJ1eIH2EYj/svNgczh1vkoJR
ZdcE27vGdO8KWkUPqjrnLtz5P4aWrNg0fkrCRN+C5kTfe7KY3qkDQGNsx6m3aHIF
PNbm33ys7lLZo663JYA1RkdZZznzH3HVGAi5q27Pp+QpoYkl21E2CNSbfzo8pT1c
8pBXD0vjZ3s54teeRtkERe+jPwcIVcn/xSIYNRJqJ887Dp5OzNTt4R0T6ZkhUpGv
fStjTbchU40cF5/sWHL1vU4TBkIv0J+WMRu2QK2BvIBN3pmek1p6oQishIG+C1ug
VDEBEYfarmhqDWn08SptaPvVmkWCeabTIe6HgpXWs7rSCZ/Y70fGWYX/ExaHmyCN
i3416cc6qHEoJCZ2XWiSLzkUJ1eSZc5DmyZnBXcJ0G2d/ThUnboSZLcN2qxPfrfN
hRR5kx0qdnXUXVS5f6oZkdiT5VdY0xW7x4IFwinmRG9JArBfS9Uy/wQC4wo5cbTI
a+5Yx9kgND6A+c7Mb3SrO4mwfe86X31kTioyOVNFDQZpjkuWiY3cDxMN3uAgUWbr
1fai+TRvHSz2RVzOjhgZgTC6gB4zqFv2exlhJSQ4Z+qPI6pQV1eDvDCr7H1/zKky
xNrqWLxghop/aUkGV69XhjEB0wg/OFwRXTlahT99Iz+85j7NDp1VzL0WfFLWdI1i
WyFGCpekzQE6ieYh3q4Zue440R7K2p4LngHo6SmG0hBnCHiCtdmPqtkk9Iw9RPDO
jAd3die386X+7oj5l73wDNIG/78myDo07HNui9xUOhNj7XK1WCiCAdev3S3eHHZ6
lcdMMLn5LtHf+kkOm8rRYkOA5hVpGS53PJw8Ym7hiRprw7bn1zXbiRXS7NIRke1M
L1OUtBdzA+JVH8XdRD1Ek7Is7AcSm1gzFWwE0URZ6Cdu3hCOvpqF0nMbrigS4eOk
MDEkFHNa35Hk6vtWk4cA0llveqpAIfkretR28BGBsOr/6DAa3aTLtFSAuiNTuSN4
gAlIJRayXoMyx+0YLmQMIapJ2BCXSLy6rsN+HORwyRSA6DQaduVfxY/8JTmi93lJ
GOYRm9KNXdlfDhByrk5f/12GnFIWlOMrjw7zUattAem+msYPHqbclEREG8w1FnnD
7IYU9Je/HupN0r72pK1aMw9+WNgWy3Y+ccT8WorxjlTbMQbEdBnGI7yP9esrfE9V
TpC/HGeGpuDhJvV26ep9q4rayKtnNqEIKwk7X1ubMWjok/KNBLMYg2ycRANArXqy
ybqIJmeOk4Js03N/VsYhC60m6aDxD7rGgKwzMd4jMn72nFVuGs3H17vrfGyp/Bik
YiCEOvZ5nIM7jeT/H/Du404g2FfjX26v5SKYyWNnCngw+PCtRinpTRSxUiB+6tXE
118ap9Z1qMn10yKF7T9bq+m3qM5YYJjG7uYwoLbzu4a79FbZtP52CeX2NwMCp/AJ
cPyM4GYgLLr9z4o5KUnJ7ogudTyjmkJcZqe8TWb7QbyxbYOOO/CMETAcAYbV60wS
in/pLMisTLPanC4a1+14oK/MNGBekr5pJGusrWswNSNS61+483RRoGwH+y32mxxw
x3YIYpRiELpQyRigx9Xu2QaFKPxUTU7L1+dzIViqnnG/vlZPsk/qljBWJd17eiM2
lxPbASPQmKgl802jm3M5sEfh2EZRXpc/Y+rbGx4LkP01/6baa9pK0sLFHOSdwVCa
ulZtHpAF6yp4wdG9UC/x1g+NpJ2JGZjcUf5tAE/YPykrXv/nV8x2PwagMDnMLlI+
tfhhm/6kVLP1EdYi+6znxVKzKluf62NPV6/DwCaZHsRsvWpDCUFBxF2Rne4y9hEf
fNrGzSmp/r55VEMS2JVyj/Z6X/PbybcvCnZ+j1UGjZiyqOLYuLygGGe4mvw3rbSQ
gwuv1Aw4IkEMFbq3/dfNEbgsmcaujSE3dMRSYhoc2u/sbufouXSWGKzilmFz3waU
/sgEd7pw2eqoRPQ0m4oM0cM8+AO541ly/TdUxBHp/rE66ShlTRSTCLLT2p1QHtPY
9yWuR9bnJcPBRAWxz9IJc2vuuT+fyjN1ET0CkadZkp0rXF2BYV1PUYb5FRUGETNK
PHMW/ZDP0CVcskxp4h8Y6RCuC2pJIlEfIARcyY0/XTvekmzYLWMKzItiQtrlv6Z5
o8HjHZE4QJz0SqJAJMo7vJ1/AOgSyw7c13xDhbQKjzyfh+LN6+oOqpZIO5ou5BF/
MAaZsz8YXQ+jzPKyEJvIWLDT1G2d0+7qBIeX+trWd2YztK56pYx15yyzeupjDnjl
LGzDoTwVPAqxbaj1azpKIHfWbwSoPld6S8lpwc9T1gtTNdnz+CjdVCwJ/LREVqwI
gFgVjkG+XzjoSPQyeE4VReswFv1wSBs5No/WuG9za2v76E3dIQYMfdYEUSr6b7JM
AdFqB08fJORtXpzkjLAjl+Hiys/A5aR4YqSVxsgPuxDMfqSYgO1Ro2cxEPm+ajQh
E0Q7s9AY4z8Cod1T7gexnU4pNFCJP5/NpHRstKO9+1jic1rGQxZkhSfRuXJu8Jfa
ph7Y2XKvNPm5ShZF/kbqrf5+o2pj5rZGG4C0BURWhfyu65FrI+YJAd5dAdEk+l6E
L3N8Y6X4FJxVWpib0sFFFo9YQK3QEhdkUimwHfodfaZEgxrRpsHrSIRp/PSjt14L
8lLxh6lSzvRRnqbg+QlUZAkjzEUfeme4CPOh+CWQxgUHAeoIPOc1Os/Hqrk1XJAW
pGLb3Ezi7342dRYZq9ISzuOVWfDAOfCTZD9Dh0NMsKlzOGKJKhteGwidWR7DOeGu
OiiLazwVu8pMgKCUwNlZKEpAEEblm76auWkb77ZxVlU7l1qf2+jpoJ5EZSdFCdyl
PfqfVjSJ9/ZqxztDLa8ON/83q6Hx4tFut+tbSk4/Gps7WjyIQr7YZmVx9OfjNu/k
MeTV+KzgSAL9rCfMl7/qADB9uD2pHwf2HtnC8M0EVNR83ppKojnJvBtWIjKRUc0U
nidnBrKZMIZQttiTfSVvkQx7opS8EQhGTeVIyAF4d54Kl4jFnljwePIMXAISyLCm
qLsyitLxmvt1AbXod2ufpYyXVVOPGaEM9nucWP6snica/AtJqczgbkO/LDM5J3G6
5p8ztYlXm2JKZigrhutqrHTxiZkjj0GzebJG+9PQ2JSJGdoFdbPljhQu0cNioCT/
FssyZg6j6NRS4IH7DZWzM7nZdVku/fIRVGHZPuXg1JK6BqLkuUJuLBLS+oJQTMEr
FGVWOakwnRbad0xFvh1KriI6om703LvVpRMYvOC7J8vj77ajdh2zRW8rbeWpwCcc
4QklbT6SS2Do1OMgDqupJwRM1bqY1fhtWRYRXcM9G4yf/JAs+DMQbjzq1dyTN/Xp
wBWtdUrtQ3L5ahkzJu0DBrsC/jfzh+7p9HuUcAupy6Hmivy62L0llK51q6NqNwYD
CTP0D1+eTKB/nz1lrQLw5ce81SvaztQL/ES3Qsp5db7rA+MKq3gPKVQ3ltzVTazk
gPUCsG2+XTyy519bc2lQS9ml6KpbcDlqS3KZrToRWKQ8FFlcS/Mz6rgWxh74Om3K
6uEMZqJHTkzXdatZij7ihEnB6obpdXpg6jLGUJul9YgLsYFL2PELu5R6xyZNuqEb
ID2HoaDSOauHRvZHzDQ+JTC4Z0Q4Ew42eF1TjBq9I8b9uCYFwY6Rzc76FAn+0whQ
7npt8/6ltSsC3gKaBIQCLPnYPO22gWUkb4i8nhN4xtdTUQ6xGTi4zaVQ9pQLIIgY
9ldHHD4bsB9O9tp/rspMPzeuLb3yzvRD+Fzugh0eMIHaomevSbQXrkeGNKV9BaSv
A7SceKkOgxDE4ubaJlBnxWiGV4378Vb2mqglk1rceTZ1G+wqOSNHHX+RFamZ+TTa
ysIoTqYccawuyCk9jD2OFFOSiLfEpWxVCkANBnXkdSTNjLMcm+xk54A7BYyxsjTX
m9TMWksmJOAqndrz4CqBoYfbXTce4Uc8mSHBAClF6UykKhLzU/uybhv2qWL5lf+p
1HaEk6umLKCCCh6ZhPZHVCMfUHpU1H7K3h2kOeENK5VZ/K2CJHsdlEnlOQ9nRNOW
P19PoKUlJLmM8OEDMEXj5+t2gw74NMx3FMKMRM0JPOanm+2lwayo1NXNozELR6/X
xBzy3AYZQY93fxzbDf5qr62wFVaNP3/lnihQUiANndxT4d7s3scNcoyO5cBZhiMR
kXYZv4hURSqVsu6MTBpPHoH01+Sime5uKamiNwoIVnJBy6l2EO55MryE02WgignG
RyXADhfynD36RYrQpS8t/3jmuxSo7Dj7CdARk9lzcVCc/IpwoPipZsbKmtsL9uz6
tEeBOclF9Rv+rAGrXM7GlMjT7amohAvCrwkW/Ubpwcd5QuPWMZkXxbtts7L6MShU
zQKthKvQ0TeQgDd2ufBmiuekWWUSKYnAm9Sq966YkRnwDDZqFF2MPuUNWa9U1VIH
HYv4SHzuGLH+t8FyGyOD/f7ADxdQdjQwPi0ekBsOEPg+HqPZcVjBHZBybJzyEs/W
auR3mU902mMeMYJDn3RdtJ2o82iTsvFF7xNOdDLqZyDNcRf3pI7DfVKBifPowDnf
VOnTssRg7Pr+iRYnxXOeLByfvwxgTYtHynUQhhFGsAoCnJVKonFwWqZpPoAWBWa7
52Wva7hZedhaKVAYQ4uZ8H1/aqNOMsOmWuj/6Nva8WOZf+kkxN3iuCeVi3eZ/Ic1
j80jJUPUwbN0FOdHz/2TgRgpyF95SNeAWtoLcC1qjBturXDkoN/pL3d7CtDL7VE9
QPXh2jsyn2FrYLEugScoaVDXOankR1qyKcx9+/L+ihdlwl0o9vYHtMC9UShbGa77
cNWUaf86y1kC7/itxgkf3IxOyTTN5VOvOok1/RjZgBS4JzTqXOibXNpJrHyR3aWo
TqFbu2Fj4RBt7yaaKsZwVJxqsoIfmC5fbFvafsa5vy9izWiu54EFjg4k/ljb2eOc
n/jjfkKFDGJPM00WmP0F8SQN9mPJGH5DmUy8lhp1JBVgSt0CbEOSvPkBwp4AE7ue
HW8GTB2DABx2hvFHy99o1vNiWQ5EEi+Bmj4JNOrAZEi95/M6SC7QAwxIFJiQRWsJ
xUmreKY2peOle6a69YXZCtcXh8gyk0rug7az1A/u/Iy34SjoJVxP05Qz4MI/N/yp
NlnzRpXs1Q2XxAg++OHfaEICMHKDL/eFhylzyBjNO18CcKwkKCap91/e0gRGphAd
iqhII26LfeQhdvBc17Xb20HwUhanf/N97U+zjkellUrf3yW5NK2GbKN3quymv9r9
DUq8AHdoAtRhoK7P2k8+iFMNpmXuc3VVYrIdsk16PVmzlmx0cDlxryYcg4EZhKuU
o1tfJ59Nu8rBTR2NjC86/Q7iiYJqhQU5MIrUFMRjsMgVAjPXoyHTmmGUKW4jYi+D
01vyv2XFDMSsur6XSUT5giG2Zd6q4+rjlZ5jSEO83diPir/sT4ewqhzmrx42WNed
T3+Orz7Z5+1olEn01k1indeGnSScpIYtaTkdRt1antbUiE3q0cc9XinOGrPbP2Pt
IpqgZx7JzkE6LjCK7fe32xOt7bSA6j5PB9m/LNmU5Biyl7DNj5CPASCqY3mX2fML
Fjxkncdi9l+aSk2YTC4Wx6YPw3jXt/aGtvKRERgvbthHhtIwx994qOlwQDbWq/GF
+e5XKtKrrPFivRgITyhXrGKo2SrkvTCWPs2rk92y8gmwsxXdsmOvc7fV4Pi3wCJg
zjzCDFDyuEX/qVirPnE5K1Cx7jtvNecalw2d8pp19cwHuYltK28BCgsCuqmZQ4tz
SHLnQ9PEAA/wFUp+p5dtfj3L3TajyWO84ZOMxyhXZTrJ4KxHhyxf2cb2EBrP+uFM
CrKr78fy0LIOY81N4VGwVnNeJq0oWG+IuqLPi5Ykd/Di3sQ0SFp8DvRu6WWGXYYq
gmQJ9zMndRRHpifT1zHuhBLpiGIQgeTegGeVQDXYM/apEtd90WIoDdqs0q0R51MB
vIHcw7f11eIsFJk22SxdHwmMl9SyHobgFMk8saoxSB0HjWcf9VM4SXbR6VECT0BU
TM/to2gC8qT0HAgBvYDA+vZ9158cDrgMzsn8uFz5Ac8PJd2xxvjO3S/swvySZV5k
bnegqFZ+nkrmDiyeyf6UTIXj3ljWD+XTB2tLj4Ky2Y9uNrTN/TwpocgWJjAt4mk9
ncB7xmRm0uxASSxetS3OuKs7yY/CzkPxYXh5z96uuYV6LzLeu5W64qjpLA+ocRVl
BobS3sKv6Fa1XZv634M1wfbMy5bA5idNc/DVXzhNf3n+wIkqkfZCjbcVSy4y44r5
C3e03ppxeip53HrTIxGGRl5PtCV+CQrN/piS+zvSBIekXWQsy5mqwXF3GkWvukZ3
tfZs5E2+Ftexva7UBg/KQTvhVcDb+mwpFogVvZUba3t8/aZsdqqaEI0oih9co35I
boB6fOPzH2LPMwzPC2KdDnCtIVGAECykeb+jFVGccyrvmCiaphqZ0n1GCTS426uM
N2maYrhtV9A0TqMtVfnTs1qN0A0fm40R3Q4/EB6k4PaZRT9m2cB9zUVZKtDocghj
RubAcMAknB0sCQDpQv/H7RQSVfIEaqwoLwZOuarHRZ4vG0zRqYqSN74GuwZgkogm
40r45CcpDlEnGM+d9b3ZG6WkXguKPfoVWi21G6L9XW0AWlNk5OfbnNbqGM6AlOMS
A66QNSJ5DT3KHR3bBAQzlJPlLBsbgVfjqz/rO8ARSSs4mJANb5K1YrxW1GcXR21b
zyO3QcwaW1c2YqtBSaGFh/lYcOWE02RWtyjSwxbrpdd0xBam8A6Fh+bgy3fcZqWU
k4jn0pHgg7Umu/w26Zq2cAlqu/DkOHNpExuRNG78y3TB4tIERxNCQnqyY3XuyUv+
HJTG2IXEqDHRS0JH/MVDYlNWYnN3gCxElUXVaxGk2PNtmWZhZGc5XX6lE36iBabn
moNyQ/DikVEM5wKmX1mxTIEUQhaGW3kaeK2AAxNnJmQ4QRYCq5mKq8KWa40//7rE
WaiQ93y3CYHq/q8jJXh/dwsvJ2jpPteVqBWUDQeI2EVfW06+HfxX1md8dY5Mpe5d
89b2ruITVpgST7t+3hZLACu6zQIX4RMzIkUsc1+5G76eNxZaPZQ/8ZvjmToowzkk
geFd3SfcAnb3kaV6D1qEhJZbGv8F9JKCYrba2JAmTrdLXltNQQtepFBuzB2t73ny
xLoHrtn6uIb3qA0aNXLSFMV7D52tgT79l7o0/fTWDtHaeS0lIWwAPZA9CPIs7aRj
jMZ3BzKGAOgSOiaWxJ5PGUzLniCtzsPs6o+KGLm4UxoPWCuPzMzAo7aOtiwbTnMU
6P1brD5WmkjVtQtPWYepE9hC3YWG05Okovq3fvQmhaUeV9xyRlfFEfeVqJgmn+WR
UoGcEL9oobWEVdavSdjqNxS+cZ98qffpbZrSOh790X38bQh3eQcdN6oZVOplUV41
cK1ks/Gt8/NJjsD5SvRLNQsZP8Hk84vVi7nFZ69lOV1WEluyEEgw8dtcs0+aH/Pk
ONdFKrsdns2lX/2bGtOBRc09D3GIgwaWdNLA3H9C25SD/Qhx+5xQiFuQ3XprhH76
MaBmkZu+h+apgwrTwMXpPeij/hqJAcPBTQqu+FyjWqSfGtzAaynCWDL1SJ401f9w
tfM3JsVumaf0kDUuhtk0BvlOkvp3sY/a92Z8oC0yYErgLxtJbR6Z5Qmd0Ejmt+C0
dl8tTwZMXaZlXZitF/AfwCU+lTm1cNOBCFpM1hg0HTDXbIykEEP26MwXFL8VH0Wo
RynKgKjkuy+JRgSunX/CZSwu3i5BjrBgaM8dZyzMXUBCLWFE8VwgydPjUss3v1P4
uJ+bIIanB9G0EtAjt15FTqdpW4rMxAIwqxZIccsXhHvBlv3f7YMh6MCxBGJfBBSD
5YaxchmLGBbbRwh6YvJqPDvAdhOu9iw91ydKhQ7g5LwC+cv2dWZ+cKJUUXVvEGv2
Hn2bjTad/Sxj5zTQwLiPZ7s26hvV5s1xXEf12/rHarbWJ2JZ0aKUja1E0oPiOMQW
M+D2uXzOz9G2DiaODS1rOTimM3dgztnXt0iM03TkKru6LifBR6vXN1rMlh0VnIAc
wupv0/1Mc17TqTzsvpQEKI1rhSTjl08P8+sFRF6PMLIF5FhxlaT7LfUHcE9PxdLi
OTWKmbfrYHdaiJK0g1gUd706uJOaN89SP/zxcd9mj5jzLWqAHEI/QaRKqNMPikAn
pe3Cze3YZ1fgwZBVxzA7gfExTzNkuPq+GnDjrgvLdaZWpIKWgD7tj+5H52nTqFle
dSeAk+EW30mnaEcdccFiG0eMMlGfVdTOsMZ9pHbSbmywCP8utcnWIbdCQgthVYba
JS+e917lqe3MqB9zj6KBFPuYM9bRByjpP7x77C5KmLyBYubIU2QRwIetnAg3Szi8
5Fc2i1rBNS5v2nRMfbLLw4iC1PJG/JlDL+JbFgPZILc0sBbT4iogBbC5Qb3O5wld
2busxnh63dkuH4bvSrEMG4b2VdUiUmIzwdeBn8CZ5/CYRlGKlDVHd9sbpVSofFT2
P1RXqxauYi1YayOuBMLIWLOwZVpNVXvYAenvvMxhERgd2QaXVU+1IV1k6N6GfKDS
nhSDGza8+jeFrtEnQLy7Q79uomsafPsuwcZyefUEV92lIBmz1J8RB6/4dixcSJtU
ZnGsj1Z+augnbRcd/4u6M9OiOJAv9lNXPE2GvLn1If18Qh7VP/5kz0ySvrPg0L+u
AB4wgUyyZCazJNH+4xEz+sb8O2/acSchLd9Dzal0GcKyxjRT5C/ASEXud+VJQ92+
IVtP/Ej4EIifur1Q1YDJAG/J4eHTdQ73ZIWZuLghtFfBnvwNH6Z5uJw41kWr+MF8
7jyjrgC++MAaN0zVivId/85DEUYOfeX76Tv/Zgl3xaoXufjVxhAmcf7yUHjXzA7c
Yp5QytpiXBTCW2EMYMWNMf8Yog99qr2SH89NHy3aOZNz3DGLUBW2G6xT/XHtPPi7
rOdeKN797Ec5SILbD1jg3Ruyz0JzHcqkgsB8pNvpUeq4LAWyO2OcjXUoD/WZKCLg
6yqZqVLNsj3eT4/AxLv5SMinBQiFD+AlLYc1S7RRxWJ6wFcHFcbgM7VoAAaANYC6
ErRYcRNVDv1zwgStz2p3nShmOQ+WENDLX2CYQoWZ/89FFQ/okqS/opb5Isz6cSXE
+TPE4+wHd4YTp/MvjlI+Q4DmgQ16aVtD7DITV77LbdHBr+kgoxTZiEfkg3Gqkqri
I0VUZ5QlCsycRARWINCM1rUulLK0QBx+P6t/9epamDRutFAUVDFlv40eL9HB85XJ
4gg0sinuhMVk7F6luuT2X0f2SlsLsjz8ldDRbcJxejzLidqaJqvqrUd5Md9t2IJl
MkXF7OnkhA3NFuoKhmrOjScigqRR8lsqLdeOyUaHFC4T1PPlTSxYpKgGVqMHfrns
3fucMekvMcfXpg/cC3EjJf9o0mM18pduCE5IERPTF/FEdWyAL4316orAxukPtCSG
DPyWjvRQ5jxFVExe/Re/XOTDE75Qx385j1tmjqpyngiVLOBvZ4yVvobSasZT6clA
uTmLf71ZyD1TBIuuYR7ZTBtPmoF4M2vZ9Szywr0pDwJplIoqgjzY4+gWWxuSnql4
hCL7YRPcYAX7R4cVAw97DvOrr/K8/u6GGz8YPQxqo/DTJOKgz/2LFiupgVtnRIz4
LVARoQgDxXA19P8EPvwSo153u4wueUqe55jPoZf8GTJVu0evL2oEEzUAFB6czlkV
qqzcP41TwCkOryJKW/QGzdfEorOyeAj+wBxs115/NQH+CRW3YykLbLs9vjv1P6wl
LQwydytVS94swa+KtD6gXoagwiBUMFq1l6b/VTdXAgATg3AgSS8BRipb7Y+oTCpW
+D3RY+fyold3FcKP0W90ggyieLyeXcVDgj61zUwDcT+JonAMhaeuKgk/swuu9L2/
0xw8Mn+txsd5zt/R46ITAGnzEJm/Ndvj+et9EosfzfKEKWnS+cjBly+sy4jRpuLU
ulgywEyhIdoHvipYJsYXaE7Vycr6RpkkwGwOPBcfoPhIPM8NxpAOC0m4xQuBhkeP
VU2K8RmyBHY6KxsLR+dG2KkCwaMIelrX8qEozl+9nQdNTqL37Jk1sIg25cI07Toj
Fm7YYIM3+ZUZl1u94KwwxjiscL5SIH1iWg1/CqqPQZB5tbUyAuOEr3sXKvvlrAiS
hTpnWLa6PC3DUo39k4PZwUVf682l9ufRfD2FzizGNC4eDulaVQ5w/BS/ClAhVm5B
dMxcAdgxoJRVsdvNoNHZVRrTxWconmvjE+sJXrT7Hj9zM1KRZFRNu9wMNIHc3ESy
HrCtiCLy3BtTU9XDqcqsXY+DOqdk7jRzTLWffGVSUDV8r/8nloLIKk95JWrsKDP7
N20AGWcxq/0jTEuKOQbazyktJEBGaRrQTxGuLFQTqKwxuge2U0AqAq6HBE/P1/y/
OgTcL6ItjAwa19Mgk7f80DDa5JsG4d35ie0ZlZ8wJUf6xLFDJUFi16u0ZQ99wJ4Z
K+NvCH+vWazlQP8N9pIeFGhkqM2TQMCi+LKcIOw2UNfRraY1diHMvZs+/KYkFDYJ
eTbhtjRH0w4fx66MFmfzOY5kuDu4M4ib8uVtsTsZBrPVl1he7UImcr1GSq9nqCLZ
M6WrzBHvil2KYUNERBD1bcklrDGlrZH+mL2tuv4XQbowNyZ79hp6L5dgicPEUshT
2bASuuukZXvtT1u2PCsTwIdlaoKR3wExqzafCHlG0eSoy3QaOvKuQvtBARAJ99sK
rQGFKfkPE1eDFMpvFhfLOTl3N0ALkJyD1J1LvxDkl5uG3J4CcStCmE1h+Nykx5+t
ncFcDy4loLn7EJ5r76OdrXaNwwMxDPXBmuyNhsbOkRx9W/rs/vdXmRRkOOuBOcrT
TqQrLdyTUvJ8ArkSpTwyTfYII85RRn5BFh2tkFE+UsEY852mzdQTiaUJWeGuv3uA
74cQrDJgrnE1c1qie4hSgu/rvG6T1HmO0jD/qJZsPwnufET+jbIeT0L8HXO7wkU9
smesZTNT3pqHezV7/GmMSgP6FgPgxQ4qy6shoMaMrn5JAcM8/BNX5M9MNyOGmt4m
VKMebhYNRPCt64cFjRGGzwrhNImP/KOBx+ALDihQuMVb6FTgNjkQBQ5A238LL5e5
FjbSvCths9IHhoREec0Jz2yWu8ODG+e4p+/vwZ27Zmg9l0pDQNfpPS00ss7JIi+G
a/Lwws9WrLREMQ/++TQa1ztfCJNE99R2qka4NrpZJRQthIMrBEammfRLgeHGdhGp
fj4l86Yi5rP1/cn2RG89QS7NskO3U8znr+YZjnGFm6SyHLxjGNjN33COM+wtGFV1
U8rfbRL5dnWz8uUU1p0X1dLZLLjUmEU5KpIxXIywZtpSxsgeeKG6pmugGfi7wtFp
yAVctZy21P975VqK3ZAVw7hVvUNHRd5YV33uenKNPy2k39sdLzumN1Ce66srtlus
K7+hRcnAQNadsBEve51Gvclp5mfZcGEguOw610zjSljegjFT5Ac2Gr1S5XmXzxQn
aUT4aiME2AeiXGQv35i29HLZd93VOwNnbaYRd4kN+GI7QkzqPb2pP9dD/fTC7RSO
mXNcikUrex+y/rS/22o7GyLNf1BZPqfFiKtaEV8jVNoKMTN8I55bR1/G3eFbJZHv
SIoGEDnM5OPoEvrxb+WQWE6T9ReLJnyue3PFw2N9jM4YCKNpkngupa5ErMN4En+T
NTmwc3wWhqyIqzcGrLM4E8LVWxqGEIPIYiOVb3cPkp5sesa2dzduE3Slc+3ytvwN
R4fLs1U+TyHZ8gNe6iZg5q8lOY3aALtj80jOWNR12nHo8FyLTouJx1YqHoMGJjoR
xuc0/I48wfBbgAOJNVlYTA9qb865Xgq82hkWjBzgYtNsY9+Gjr0WZpFKVudLZhPR
wZtFSQmc089h6l63wwVCmsXfE1lND/RPaLJPAvd1Q/BjV+jvqJs6wmKNI3mfcDr2
zrwtvTOpRvfcJ/JIy8SDKW2eubyl69gGgIFN38RLZiRL0Duwf5+vt7WKP0jKMdpc
2Eflt06RlO4nMSTzqguRBYLhX5EpsfaWezuLFf//fPoRcZ3eLkNbIDcClyzzuhRb
0+ENl+3pNw/A2ebphtaMbaHdrKQIJkXWcFBuZkd/AyqQeVJqCZ7gtrTRT7gQ0baH
gcaWjP2IqCnm4oT5IzG/pH/4ghSa2bLIdbbgU2qXbAJezhh8tpeTKT+BIsKMS0YV
7X/BYszpOaUkkDmkI38XkCDUzNSSeWY6cpcBSt3npaDuxq/rvNrEagRrP1zHo/+4
JRdHFUGNix+qkkNBEWO8azLX+BL5kKLx4YUKuyiWH+jyrmbG6CvHyDmLJsbEkDrI
3A0RTAh+8CZRb9qsN7hQPH7Oo2qnu38WKKZP8adTDJsZJMkd89nJGb67Hw00GhKz
GLtfCrSNCwplfS1pLrxUX04lEHONcHlRWPZ4LyxB3+9vkPg5rdlvNDAtXoYfpOCF
qAfMJBYktzvCXVNEqAYSJ3q2PHLKbBA9zHvi0Y7Ot8x0ZV7wprJarL7/rXCvff9p
hwBs7rJss9YI/Fbgsm/h/qipMcRil2/DaQrOB9usZ/bOK/DeH7IXWxhJa/nul+OZ
B3zflT0y6S8UI++6X6gTYrslR8NsTw5azZrvmFRyArbvpZ3sWCxU2QUN9bjzDTVn
jV15PAZ1W1TjW1GoqJL0dXivMrh4h1X6ROI8y0/7hdltdGzvRIeQ3H8SD1rZNAWk
gZCnCBqIcPOf9J9DbjkYcsrsAO98lCTxrI71eyV1V/PqZJfdtMd67BfqNVlPGhxD
RHtSlxBTHsOwqpchYwdkh7asTQ4N5LL70dVyXvsQmkTX87RBaqKLoBNlAac907fC
jgADncfMkZq3h9DNan/OkrE05ut/Mk48dY0ItHmsHMXDFDVBSSKEpxTRDzFEi82/
VgXYGxDsUeAJRB2p7YX0uMqScgrr8X/1QDgJglfmFSrRVhnLzwJ0FFd4B2CBXJRf
qTVNl8nLT74RHvyC/NO/EOvGbNJs+rrjBHnKVvIyT3SQvSTHkEnRSZeCdV1d+A9e
HMtMbyqQQkyAMj6TXB3pwSDs7YvjGTenldVH1R8SL7Awy6l3wWn6/LhhpDXt0kZA
qkVqERz329kvwrEM5BwhEJZbCwebSMSZyxZpso5hZVoOAEdJSFCwGeRC8QXy79NI
MXfYLdkPI3XWeHr0C6oLg2iuVW7C8etX/y7lkNPxyRewbB8hamePPjbgONWJf8XW
nvguODuPhZKgaw0sgFfUlnyxto51qNGeyPuGRk+REtwwSwzEGLf9qHKTmzbsgiip
QI8O5uYe08KKR0/86g45XdfptJC1QedxZM/MfDFehlZ2X3L4FHlUf5mZzCXHXfjR
IJ+W24mA04YgyTYD7xa0oD3ePPEUY5JRJORdY5+wNxMbrw5Mv5fNTwzvIm6YHkjo
yuyGDt0ZaiCZJOKbZ6nNlsJH03bHrYCRXhD8+9vKWe8Plrb7due6yAjyALNUB/HR
L4nZYk8C+0CHiKd5tySeR+IaT7dQ1k39RbSxOdkPEDDBHWIdI4pOMi5fcQPb5SH4
YrjyLqR0TT7ixtTqo/4J+9xwCG7aNiS2rl3sRu9KeUSuU9zgnuPePlHhSR6UoFfk
DlswmUkzba0AX2ziopfAWEoruUPDHYtzn1iNOREQcICDppMEQcwyJUsb1pbWShyU
5bAbnY3Ks9QQSlaY5BnATcpAaf5SQMv0ujBWFFPxLD+Q/x/m1vPmpLqTYEDLAqT1
VJBLPTegStrTQdR6dTU4Drj9URCY0M1ItS7DGB3GcXpSP17P5NoAy4TqXjK5H2d+
Q2AdV7Ju+uFM89GDNKDARYx4+q+YU3b02TSbUoeWiAZEAv0DFovWYqLmlFna/OMB
Z1SAroRn1HjF+HVE3pmmOxwe9MKZufBXrBOlSunweOT9mh6FXcEkWvl9SFruekkl
pxyLJdc1/v65p7plnDRqvt4AUvL3iEJmJLwyBGPjg4evq5jv0A5OBAdYo2DgC8CC
8W8QnWtdlRZMtK/fK5dIRGuQ8kKuSVaV6v6j3o+lpOuMGuXnXSF60c28TS7iI9/b
CNCcRVCjHRCtkhdiJFF1lAgR5IzLT+fOXylWHxpOY6Cif2iWdZsF5iqTCwECT1AT
/MeJCXnNKR3XDRFuQA26RqeunBUn1ugpBmr/ezr5RhZPa+QnUvCqzE+UgLPOfeYf
ltL0eauKHgsLR+VUTLg4vxPfAVR1tRVIf1d94OvVuj5XWwa0xgDUV0CYUACSkDEQ
uipORjSi1tCLFrWwuURMdJ8erQrBAmdJlndYEZHwmvgtj6uEsnzmb96aDY5lWyUb
HpyXuXbmUsiew4/UvfX7SK0Q0iGzIzQuhMVp1IFrBOwUWLGXT7I11ENa8glV+DZf
6scQirMUfxU/qESpmNy2qsP6nNmBkfTiTqOUqHsNEs8y+7Ed1t8P4Uz7w4l5mVB2
C8Fx3zudtI8ueeoWvRfKs5uKH/YcWQKZA7YsbCEQuYSqG+JFCPN8RxsPSAnFXM6X
G463iGamXxqxQ+b+I2d+6cBfGvwLcE92RMpSNM1LDJWmN4YN1uPdEcWDcc0U1IIU
Mtsc87nu26LbHCsbD8m+qO8iyhv4MYBB6cdljvl7YJ9WMD8WcsEniqo+aBNwHbMq
RjHvJaqOMYptVhh+JZ8NIUbg1DTuFiNCp16w9dTSWoNwOevLZPQyhLrcUPNiTk+p
o2tkJk6I7kXE25m6rIK1clrTCAeYEM+S8O/KSI7mmLJwxrYLUyYThTi10+3NQp2l
K880fpQC+u75LEg39wiDlSexLh5RsJSm82cdEoTHhGqq0xOvq5Oe4H5YaBhn7kwX
si5EquTUadPbjUmODhyif01fu8/iGYSc/dUNgQdJdskrh2/Lps/JrlD10OzWuRU5
ZJ29BMyc7ku7vLOw/EvjV2inZHDkwYei47G3WcNURSoxzeQ36Fmbhrnd2YYsWpKk
yrWRGbDuBSlNeJEeasqEZrR2m6Cq/kEqjlVGiA6NX5hkhhwj1FgmDe0YFuZgq7SV
CWpZj/IA4lIV0p4TzfbX8uFvnhcsH0qESzVui0wu3S6n+tNfdD5tINiQ/5aTdxws
HO/f9C5PnbYxD0w+xBwk8qLeWjlO5Y9bF3PcoszLlSc=
--pragma protect end_data_block
--pragma protect digest_block
8C3vNQffGW8pfunLs5tTDCeIf9c=
--pragma protect end_digest_block
--pragma protect end_protected
