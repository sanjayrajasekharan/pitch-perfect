-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
iaEIOoVqU1VTzoq0wHbeYCHgHGL9fwLNR+hei34Lce2FO2cNvV735yPrVKmszk8w
+6lJU6RmmdLzAtPkbXUFMFvNE/qT5EES92cnnseK+L+3zuVQVky3rgrOVhHIqIhk
lmxPrIxrPoeLsJ6oVknBMcsAlDrrseqQqLol2B5d5As=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7685)

`protect DATA_BLOCK
XEKYCEQywDNnWJzt+k64GxkDuRwkeyqIHGb6h4s6N+2J/olB6VyPRbdPNFqrf9WZ
FoHHcrlVepFrGYI0ww6jJRXmryNqrWkNUkkBQWnzFeoj5Imsgnt6PxgGES/D7E7b
l5ZMIilVQslcxIigpbqrMArk5j+CRgp9p9TzzmkAaEoWaJkofkKjU3qkRNOCTJDz
juZzHtYH06+DvIUdx+ZTcwXP/EpdJBZUiWskchJDZIegOnCkMJ90o5DaO65Qxrux
cEN0EDauTgdkLo7KZMHQC35aDQ1JPUSqegXB0WCsgBQDBgi0UDJ5k1mXx6TRB2uK
aNOIl9U7s7msCke6e6vbLrg8SSMO0oKDq4BGf57ONjZq/P2JQB27A5R5Kg/nIPjB
pP3cU6yXFafvEvJPjoK+p1voNPe8p6g6KGD2ZPlVtkZlsuAQK457HIKBP8hwTqpr
5lFPeg/HZ7TEE0hnWz3yEN1toEKhMgtqMjCRxyaKNkswXh44v0gBMr8VAe35Tam2
8oI5hJktkWi9FqKWLvTyFZ9NfXcXwcI5FdelznWAYgp8xR0XtEUcSO6r0C/4UiLX
e8WYgP5bcpD2bPumnQfonG/LdsK4bUUjDRbUvsmX6FcWvTDiRakKj9WWxlOqNPq4
BV96FMMXCpGteLtb6LQWatkZHMJFS9KPZX0qLYLURnvHC1HA/nYBH36+RpEFuAto
EVqijQU3PlaKVgTiu61/oWtXt9bQqBb+sBFWpT70btlcKwHvlNiXNP98lGb0iyQ4
WPhV7/ZBCtOvBxtsYz+zl7OroCuHdcO/f8zhwa9JWdJ0l9DUHcpncXALBZppwg+F
8SBaKVfE4ycUtElXJDZzt7A8NMeSbvgWstr7XlpdZSOm98kEfNifVDXsUg0XD35A
MBUuRnra9663EdVy1p/Dr49dgr9PY240U7uGeji+RMkEIZNYu7soIUtr/RM9JFoM
twGnr2uUE9ZsuxC7Lj+BCbQpqB1GJTX8F8uXh9qSqzh7M4uBzWdBuxz7SJ/+5H3K
HLpR1dST87RBTqAXoWHL+W66bbxPVEXPIzVZy131h6KURAbssknv+8NEsFqJaL0a
GX4llnXFirxcsnNVpGuh/e40b6zdEQRjfoAXl0LaF9lre3HuCruyCaEzkm2paiUo
FEecBWuK4LwYXePSKeqC0j+NtAQ+Nvfjrw2HQvOdicpJr9WkfjPZPPbGlH1ShTHm
7dc4EFWnzcpuDhaZgeeKSAwRWBtGbKLL+XHZJN+hGxHRrSe0OLIz/OSMo1b4Qpgj
/ZNbF1XYlpVF4NznQ+Fqcrr7X0U+EHTvtfXPknKbZhTItrtTujxjWwpLfS+PdSgp
suplz1xpgzb4NyGm44MnXny/RWYDsXEUz4pDQ+8hEyppIisB8j1wlxZArBOvNHEE
rpR8B/nAuxF3ricGA2UyUU0nRdTX9sfx11qLieGvojWtMpqoZJds7/IxKuVbCRxH
UDxRX6i0rxhP9eFt+yMkG0lhWL5qsGXjc7yjDoIszPlX6FpmarLjdLDNhJPCyX+E
vy0yUwnG9NfjCj6MsKfuH8T5snUmYzAgGJjKE4R9LXBtqeK+nDI30p/bKIsJWSqQ
hkfdtDOgZYDT2kfbg9SJ2gbfkSpBGDxRJQ5y7eTpl95rZl69+cgSFS8E4ElfWH/P
lJ8+TN2xaJunk60fohU8UkYFE1nFyFIMHCeL5vZvYsLO30B4ekU+BReU3frhv08J
NJiAvFVGfXTNQnzBoimFkVeMosHYQIfFjxfdmY5OxqiMz790EUC/gB49qXtp/WpS
o33upAda+5D6mmhlPDLhz+PFur+tOPs0QsP00GR5bd2cp+q20GpEAsBUQUT5SHvN
4Xj1l4lN4XJOLeo76qKScW2l7CrV0cTjdq3YT8V/K7hfG9oI4kzaQm0NgTqYR7YH
2GbGzO0sDFMo2DR3zbrNKTTJLXWbX6ixMZjYJfJRwcKLMKuRM6vnFkVlnMZ5AOQo
oIZLK5dEPBruwng4nf6mh0t7NyATwD8plSpxDZjHZEMzrCe3g0cT+R3XYiLW5lu4
PkNKBvSNSLRrh3C6ATRtJh4bjuV157K2SzjOKGrMl3GreLL9sdxfkvqh9tgXCgr3
E4sAMBgjUsqmsg0LnhrujehmQYTFeFyquOUcxcF2rbhJ7ODF7cXLbmNlqu7/F2Xi
Zi0hlkoAwhIKq/i1qjujfu2OcRkABR/nunhSwczO/bKR5iUF8QKUTXDqJzSPX4Er
zXN91yyWOD46oigpRZDEmVGLN0uvnYXZoVrqAaE61HVgabo+IpWWSngYWFSxOJCx
P/eUaovuLPYigUkpEGHLAuablqvFmhLkWPOkY53t6xJCjKDfkkHvnVfX0CY6BPbY
zg9xyClosGugQyRuoFaKFd0hzqOZxKHQ6pQGBWfs1/Qh3+shuit/H2Z3O4Wz9thd
Bn3pW/EPBhBD4mjtFDqFPINDXINCxvYqtl0nZnYPCdZp1+ZQDMGCZgkxMQOEZ7e5
8Cb6R66Lir5FwEwSX1s63JWQiGu/vUPEVbY4/jyjOwTar+W+OttxWAwwyDGPc4aZ
IrOJD8gEK+qHjgAJ6S72UD5oPsSIZLdS/LJHt/mprlaXnRl4GKzbifHgfD/o2kkv
3WJ+bKB1mZ8S/+/8Y4BXYhcXdJKV8XsNuKDx2rEuOtOJqiW9ONg8c2oVbRWuzq5h
ZPoq74UDdkBgxrYA+w/WGL+vSfZ8BNIaR9BHR6v6pSoBoYyumOuvwkwKmwFb7cxG
+GLB2s7al4On4YIwIW+EOzY01MTcN9sysru1ZaCxCOD+lMY2pprq86ViWH8TsiKW
xw94rqRBFqB554YrV73AmmWISX719DQQUo9nPFWJCSlmR+BRz7jeSi2M73Xw0SiX
iOVhxHmkPe2+OILMP4PetI7/u9kLt/EzbWWOVyQygiGPDEPus4r5XeMVu/iurjPi
yskqvee4eVpiWXOWnUljb+K9Px6XnWrl8T/DR3FnYHU6T2Ew50fib2Af13kOJWRN
1Zlh+u0lYGBh2/0E+V6ZbHTt+J7PsSAKjZyPMPNFuDnZc0JVsxbqC3fu2RPeWMfl
nSl95yOtyD/cWXDTjCrOTdwADNQeocWmXh2TGIQQRgvzn0jTMvfP5ZsbIJ4JZM18
0UWKDnefNrQNGFga09EJkxS0VW3hQIu7CNKBl30gCjCu7zcpor93qqpQOm2vGQuP
QR/hUJtCBHY3AAyFWjUP7dosBpCgM16dKh9Y2zztKJ5l4TXJ/Q0vocEe+7uZARPp
Iotv1mW/13T2Qf4lqS6IPwQzcw4ykK3PaV3cyQlgFSio+cCnQzgnI24TC25/eNTN
g5U5uND0ZeHVP6Onb0Wdrszri+91J7StI4xLqluQSBA1twZX7/pMmn7Hyu/7GTfw
l50ZOFyqLS3RmId5ka1Q2yO6uMns0IAUI1i4nnCmqOvhowM/85O4TDrf5sRv9lSI
bp9njGUcKSy3c+0uwjik8npTD9ETpenXwbS/MQmVyCwyYMYO+EBC4QTHS4B2iMGo
7KrfRhu9b2cpCnMXXAUNOy3kD7TrT1Q2rUZMP4TVOk2lQjge1gVIutxe5WcZChpI
uUTFgbIDCbF46xIixV602mbXqULhN/IqAkUp2t1oQ0XsrGopKFdRLcsXboJFo9fo
nyRPDVp4DXT+bs1PIlURitmonUAYxAy8BiaNxopeSI0oJBCcCSBwOWcIVCAL/KAY
aKykVEHUA17ZQ3df84kjzq/EEIs9AksCdrDi4v+0ll3BNRaBLDQhtJzLMxnNFi89
FxdXNPe32kTWnEMbtXJL99xVaghjT/EN+/VKQjQyo/hJRHT0VgPy2sxSBXYLwJWZ
souTULEJcJ35xlsijJq7/yC1/PmdTIT5cdyDJCGyW71y+uTpiUq9TxmMcu4xNHFh
9xP3BlMWIo9tTsBGdYRkfn9GTjjzs5K20olyAbyQpcebKNgcpmhX/YDit6t4yv3H
OM2Bac5ELpfW/5hAIeESavAjXuWGGOljXgMcOl6HcO+kP04wi9JRS3MrpKoiJdex
C7m6lqGwzjBEUAW9DRQGrKo4Nbjq7vkukIb1w+vGcB+28A0fSCbj6TlSl8qGwh63
x+r2+VWmq0DpWB0WXj7rDoqYUQ5GiFOLZbU7Mtv2FkE1wD4cKrTG7ouu/17ZRhtQ
zn2LCPFFn/Hv7cc5m3Pt7wGVEBFFOD/eJQejuYk1OKZXvcxaMZK+cOJOtVm42et6
jlOXICOQp6Ha/yAn1y/Pcc9UBmX9v27o9lBzDbPsfqSl/vLlRXFbTvAzptXlO7Lo
D5Ch/9S3JPJOJPw/0CETprKeJyMRW+guExLDycQuUm9j2oKjYiSFbIRU2nA1DTOW
JDq3qDrIqXUjFhPgWBbe26aVt5JljhZXxO1hblttUKCtyyJeah8GVjYyJWsSXLK8
vo7VTa+7pp5tlxBZDYHJ7QmOYSfyuKLsfOorrfbgRdQu4o5YgRZFidPTA9vSra0O
WZ5hxrMFamgHBqMYLZLoBtJ623BGTR/Gnc3VIOIJ7nxhNTeeTeDvvpwibhHhPpE8
5YIpcezWvqKq08bhixgAcPfFzKiLR05AQ4xXbdtQQ45+5En11e8RErg58xaZ+dNw
yGw1CG14DnlyONCSpaDpFw0J2S0Pdkt3/yicGuazZyWCK1mLi46RIdpzGmmA0evU
46xraA3udwxUOUK2NAnEfs+SfxkcXnWVYcfrpkm8Ika7NlFIoN1K3WmWE9DbkxnD
WElJFLTs11A6OEYq4lro4GFuhNPPzB2QbC/5NPTCL6Ois5obV0/ZL8GchI+GQksw
cuAXTWiWGh8kk4KLLfDGzcBvJcBfi965tOuxkHjq5DRMKupIUKTQB/hw9S1Jh9lJ
yBZtw47voydnP25ZKegUExuMpz8T3s7wXoq+5fCH081+EJEzJHuqsQ3E7LxWs20B
DIzIMun99Dnzy46UVDcUHEyewBY+fOBUd96fOcwYE5NodPNvCQqGhajPr7yu7h/u
W+9xCUQWTDnquqRL+FKU66T4iUvisIc5Yo9foj2507P61nsFi8eeiCfmPhsbZzsi
RfxoQDWEe9xU46f6OpcDXTAZgObIAia/31gU5Ol+arCEYcxMwIvPHbfgHv+CiyYy
ovPdL0TXTRlj30DLJE6ZbVMPVD3jZuH3e8DwljZs5afJv2GKd/UT3afH3S5kc0Qu
3vD9AnQ1UCIaDhQtJ0rHJxFirMMSIlNbwU4MVzESwxOF4OO7bLm4z7M652k5g0AE
Lbx1n/QpqY/iXKaemTmibcHyvH5xBqHp3ae8mUnjGli6hZwtZ5Xcy2vcoGuKUAmD
1Ui+xUSpNRqwOFZwp21iKdFT1Df+xXjTNO0Wzco2/vIf60Zv3eXM8xA1omAtc36C
Jxe1NMpjHoGmOoBt0n7vlbx/xr2ZlcHEQ4ZACg+MAAthYj+HzumNnAZxh4J6mB37
XmSrKBP71v2MxZuXXWS9rkx0j7pLHQY2V0duVU9s7ThuzeFuPh9EKS1f7zLOzQNU
9zWo+6Kn7x6lUwFB81KhQ9txbVFkUZHoJTeDTNxuu+LANSByybzivRjO1f6KJq4v
kawQ6GlOVWpVHsuvqc5X3waiLyUat2jMiKJfuri4gBBqxmW5cEcM3VbK9+OvjkYG
u/f+U1iDCnS79XHZwtjOKTxnQ8/YgXbbasGizNEuWxESxTt5lvX4AbEMf/N69jAc
RHu6p0YFd9F+9i1H3+xvPqNa/kFmUQ+3Iz5DbPzARh1CFGI8HYpwJxkNH1FpoVlh
RtN8dQpgORmOCHlRQ690dII8WpDyJuKRXKcMSoeVVCRrasTd9FJ5MGgdzrYTTqU+
zzH2cuGeanuFrLDluwIiW81S53TzoqmJk+SOWteEHvKSAB1hAW9grznI3gFYiwzF
W4wo0xpHCW7+dMykzFfa/xIn8AsRtENfX4aSa0T8THe8PFuCdbjCEETSW25N2z2T
uT98ka2puzCsnKEOr5axQjLcSELpafS7LbrS7ApNCX23CZZld4YdOcQE8QdFKXgL
S8m62EDWO4I48Xr2Ul4QuoMTMMx87Zrxv21abu5f3Fh4DbWJZWFhykky/JoiOds/
F1z6wbJAhrDZ3thzz0zl24yf4TGY394mqg4OVWjZ7XC4PL2VMEDDdM4yLnX22QrO
rPBGaETzPmXa6uWB2yBGsbkyondF/u6aZQ9bIvYA2ye/Mij8GQZNOaOpMldKL9KA
8lDGuVogEccmkeHi2tIfGLNbsxGhrGiHR4sb11O+Pcc1iKkZZ/7VQd9OTyrd2Jm7
AFNhd5rZr1WZBkr9beI8A0E9ZoD4Oc99+lgItTHqEvhgDeeI6JZIsmq4aWxVcEUj
5Z+lOpNknen039S5a2I3l754zA7doqMdQPSXwQWRSKbAYYM+WqaxPYJINeQyEONg
XJvZMgZcOCY4042TbYmBfVHPtbUwsldByW+t0BdOI6c/VuSzHaiZuWCTjqsyMQsC
sJ8jQoS+rafctnqwC2v9W9nMYG7qZnm3h8zgGvAP2ugjs6pB6mRwEklF42Z+X8M7
cptePElPRV/lohtMoEWxuZwDRhAp4vgBcI1NTrmhGE8wedIbB9wL+AoZofSUsQDK
F7nUXH4edqOdPCRJnARKVA7EAEdWHNWA4SZHnCqBHXb+ED3D8SkgA2VDzhb9Jq2V
lfXWZlUdSLl0UMJpIQni8hCcQqOe6EWg8G/bLSAL+RF+fOEZBGdPXB/WQ7m0rrly
zwynRBPdB28NSAUHUMP96eIgmiGwhvkRkbmGFNhdUphQPdzB7/s9fr1x0GIiUmfS
RwxOOBXLGvWoQouCgCRyAN57kZupZoBTmCPuU1c12huCghS6vOGNaT5zG6Yz58BC
TfiWdKmlpsYVLMYZNX0n1lkg1j83MjFXKnxG6dDi32n4gn1715ozMARft/TEHqFy
A1MGfrsngZQuU8RLqo88c4GE9Y7gEl8rKeu3aOP6MYzLSxQ+PuYRFRpyaa4knIQm
urOTXSWWgJqE1UeGeJ1FDr34ZcRCGKQ+35H3zFddisGt1OqL9fbxzUp42Omf3ygv
/kTkUu+BAB9+ZftY7DpvABJp4OaA/toQAxP9lIfMOzUs0eaKf3SGaLLqDD/FtrJI
s0vgtJT2BYUQxLEb2eQquodIxTHa2hFcwayxUEI3VZzWUPQnyRlsdcEWWQuL31Rk
8HwmS812dR9LlhjT5C9P0MEpJN7Q0QEVKmcXWjgMIc+BUI95FqHlesVUaTsH3oVY
3u/ycHu6tvH0PEHhQCdFAdKvOPVfZvlDULpRZpGu2P+o6cRUthba84UcEexfn0HC
6bq4wlLFgF1OnWTGHYW7Im3SUgT+H0dboD2aFkyIUAT1EDzzxVA9whWy5aGe6D9p
dJTS+J8yKPP14p8z4bEXUJTZu14pOR6g7qM1kAy+H5skR3o4Ownl5OaVqxfs3o23
w4Djao3kw9T54D6zLqgMGr3swtbKLbCm41PyllSkg1DXpHUXLnyd80/Q/b7s5/3A
bUlyCBOjpCgwVbfGCpg8WMxqXnrHIv4GJTOE49Y2ZqBH/y3LeXY12bgoNn+LYzHn
xr4JxFkTueXMJZJ8NhSFWxushXNL93hGzHZ1qdqHb7YP4fHFnyyurkUfecfQC267
+bOaJpwP67UYkNTfWlSQ3YKtp/RCTtvZkDq3FjJQ/AdpVBG673dMunuF+amd9dgV
kUZDQfsVnYDgVhIZ3RwsA/j9vHM7NWuRJnfb7yTpGTmiPL9q4VnXXgwNJUrvv2s4
DHDD+Itfjbg/dr/cP41cE6JfVO7yfuct6FznqeR/QdpJpEaKxY7MhlmhvrgN5Tp3
N6iso45nM5LMb81crk0MBE1sP+CKzkRewzx2i6Q6u4P8E3Uqbhc7wzc5mubCd3iG
Ny8bafyJh2dWvdboaya5EbiUpl5TIUgvKNeXlJNx4OQJoGvZyjjV0zour63yE5jZ
M5+y6fX6UREr3JgGxMx08/kXG+yYRy9FulvgitdCk5sCPXm7mITJeZPuSLB1zOiK
DS9P2kDsVzFyXowjJV1ZBiPCffg4Kn1GOOY/Mz2AZuDUh6mUKFS9MRuSqu7KIp3T
GQVsQ4nj5lQHXHI8bXr3h9wOD3T0PIEOh87QSm4BX7xX9Cs40x/cyyFENSe/zacl
3uaasyr12xtxUnfeowH5xvFikLz9v9tVfHWZwsbEVVnIkvqw4JmyXG1lVb7UAg8H
8q5ZrkBTkMFFNFV4Z2oFkyxRJB57wv/yStXajCAQsIQVaNkuTjE8sD0huMCPXH9p
qgApSI+kYgCLJUFMtGJjC+Z6AhfjyHXyRsPd0Xk0ApwKCU31UK+tADgvjZEnGQy+
cJfhd48pf3A17CANQuNMjKrYFwZpU5sTxtWU8IS7E1IMZeuNoFyzMNUEo8Vt6bMg
yGYtgql1ddx4pzUehgU7ixyU60WxkxzI5Uscyi05uxrqet1wAde+qGmFpddgn2mL
GKdQJif7vjCG56s+YKZnNbBYQnocFNmSeuclIUCcVpODhM1myVEquNBpFvUQEC7U
dMlJ7hMYMvtEaG9Wv10vTqiT3wY5qW4J4oBqhzZhBZ+ii1NlU2TLLNAD+IMp4VKe
CPVUrOVt8geyRjd+G36tiXKRvbd5ln2GVhkKLsU9IJFfiaUTe2owVtdUOX1GMNxA
AfE4hHYTu0p6hq3+FHxLQBBnfFg4XUW1F/Ajl0txY4ThC5QtuZdDJpf1qVxik3IN
xPlRYWFaZmFC/dXxLKoabSJajrpYDjlCSXCUPjwFpGAqUmRw+ThwnZBG/dIhufhz
co1ooycaRBS5+1j1P9Zi4SWP7gX/DVZBcj9U1Dq2mALKjZBDX1GoMSG30X72SCnK
A+KqtolTQEeZw9d1huMQ3mOrh8y0P7LSilxvKq1vjMWtK7bnVdZFRiTdGAhAD5Yk
DebvHrq0UNT/27E7oucT37YPFiYVzphkDryc8p6HquynmTUg4m1UCU5BqZfhy7T8
wScIELRR1RG6XI6cX05KQ4+HltgvseJEb7miVJJEEMTCjE2e4kgfGfjCP45FqvNR
K7CZAZwJ+YaU70f9y1vx1V8Qo2w1YSfdpEoFinM6EwjGHX4vfM2IwlRLqcen7SDT
YUSx1okO39F4gzM/H83XI6DAyEzBV51JXCEHcmLFW7DvMyara4ww3jsVZxKw5mbf
v9x/6dclqsBWOYPkS41WKyt12W8sBJzpQ6w4vNBY88omgZ2jeDH1GuAzNL2x2XbE
eI6Q/x10sqkcSVFpM0l7l4Dc2H1PYHo5h9f9wr8PkuApZ6qE8aYKvu7v6UaXnTNu
Ox6knWPXUjbPxBbuQMGAul+xFQPPtdhlrwiyudLYY0a+15I/0UUUFxuQjMlJuSOb
UY0PpqbhK4sjYeOUo668OPGwycjlrziPMc3Fwm3pW1gKhmecpkEk6Bz7blf5Y98r
wPlRVF5x3NpocVX9omNB6dHxFUJV+ohiAk8B6X6xkaBNu7GQ/io3EmNeUj3fzonk
loXNy2EuNyPo6chdu5fWrXrE9zWKhJJSIJjkSZtl1BgCMQBSoYqcXFLLCqv4VpKB
mV/4hb6iyezcSRvL2ujVJb6uEEN7/g1iWEkXxbjkKTnnRFg35+CgBhyNjySZEg7M
Y1nQqNbCBSom8evYfuKjjFRZ8eUP6rdtkgnmtrfQTd1yV+9oS6vBingoT72ertQF
YXoMTjxfqc0/iiBB75GzBAYDUTx5yACslUXsv2y1G/l474eF4dEizZ5PHB7qcXdu
n+S/Ji/6ykkaMf10kXVkLjl/D1nkqyWmY6E5/gu04VFAoNhJkWs+belEjxNfsr3b
qEaHZW9sC26c4tnf5au2UosxghD6Vfl9nA/snAWa3CosoGu0dH1HyV+0mmzCI/LE
ySVECqaKklRQeaFlEOpwPjaV6bik5ATV/GWf2A58w44whe54k4REus2EgcVWc/iC
lTh6LqVP7xaq9DM6UIZkj/fb99KZz9zj9vHYby6TZqSieuTDtqccCob6aePCpQn9
S9U+3rb7tpSL6s+TJ/wqhApXv0IDC5G2IOY2PxQVlhRjEYNCxo++C49hvFsJJvG3
tekZf6NjajD4BGk82DEmum0gj2KHIU3SHU626R195agy+x0+Vp+dlKljdETSngIt
V/F7Cxo5LoVQBsc7345FGzhIlaV6L6+Jl4L7UewwbPeELJKq6BVFEIxxQ7oSBgyT
zASu6TfGB2VuMTftIzvv8taHvKTj2B0bKFKxuQBPpYSq83mTv7oC1BfFYm22IKlP
OBn+fxxke5t8ETH+1kpr2RFoG6ki27tRJvukTeE47Vg=
`protect END_PROTECTED