-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
IG+Fm8gbenz2hJdSPFfmrWDrYXfg6VPYB9VYG0v9VGX88EnP4F3LmhLfEzkAjScS
GAjSP6Kaax0+sAzHc8vPbxnyn0yy5AMeNSTTWZfHxNBta8M9EhuwYv2b8c1x86gM
HuV1tnj8IjjZG4vJB/QarVuQCvviP2wuA4Ue3dkIq3bkSF+x3pmGpg==
--pragma protect end_key_block
--pragma protect digest_block
SMw1n8VssxwRnBc9Z1LvoSZ6dm4=
--pragma protect end_digest_block
--pragma protect data_block
D6SxuT0sDvam3GZXIP3kLMuxwcxAdhH2/kt3FAA+YdB+GYXbc9UaVbk/YF2gAl3Y
FveC/So1B4zjiRTO6WsglRICWHJY1+UsQJNgjq9hkDzpLizdZGmKb6LJpli9TQrA
HK9uw4DmEToSoXA8X6Av/94p1LWLHePrAzoMfMVuFPsFO+ggRM0/IopfbvTn5p5M
zC94zmMI1aw5rS+M6F4PbIpa2tr7BNdjG1otjUwrUBM9ZiCZYp72qDLb9jPdui2x
a0pDGI7DjbKrAQhmhOitTSNQqwEUkrq8+M2idh1YtVhTcViKd3nv7bXomJgRSQIX
8LRIaLAeuaNsGfHhh5fDGLrrrJrpsj5aheGclRAdGFi6uGCbHVjBnvbE8yz1jMWz
nW0wgB5C+CnWCGrrInlaVR8tLKv+JzAh440e4Xjr53iJS8TIoWwHHnOh1Zq4JDBY
zyr4cwoK441RNXOirqsLlzel4377gIt/hcxpjlGpmHXSrZARbIiIi2cSaPoXPe9x
qYQyGo5MWmWr+XWzUweZ1EXyuuKjpqstC3h3cSsRSTm9agq31bevqXEQba/ImASi
d4M4Q7KSp6OgpkqQximUMPHv5ifdScsYTe6i9Kge2BQWdl1y6YPoOvAjc+SrVwC5
0d/OG3Vuj027mNkM1KlH50AF6PVxKmNXV0m6g3hHGpLSiyyjiIn4of6dn8+hsB7D
jWzqn0OIhFP45r/8Xmb/Vi5j6pQRdcr24ZahURIYCRIu68tH2LgNBsFCIZLvx23O
gJtB3EIsDTd6v0DQ5oZpYH19Giv0v9qT71dY/l3A+EnfoKxz/z/GqPC/MrhXNXJm
sZ8MrcqQ1Tvp2FXe+rNs9maoEo5FlTGrj9gYxMHSfcQIf9tG7UCQNKKwBIbEl9Lp
TMo1wLWDA4cRXeRB9LDLlm+/F0enQsBIJmsEvZaQyHbK6qH7yGEpo4WqD/ae9k2n
A4lDTKCAMy1bDqQ/jQkTMtltcAlB/jg51ds3IABHfHr8VK5LXgswWyQ3C5IfiYdY
MUTwvgtFuRpo6oCysMyivBaP+zqlFhlC3vSKEjHciPGrF9GUAbEpjqry8w7ou3Hq
Sm6dxZu7dP/T7iXpgFUrcU8NhNeh2qFCuXcAiCKbxmCMNZjkfvmRD1y2LqCZ6Qi5
FHYVghoB7C9BOLLQenA1YzShM9GI9LmTLw1EMg8rDh+dQwOhvBfViKjmSpETBGWs
PRYolBgZWHZKiCkyWFASi8lUqyfEdXIXJydi8TkjDFz0rR0k2bPL8q0ckr80uzO8
0cCFMU6pQHGtn/gk9DmwWj9tJp2i59YBXSUxMKNNNjKI2ZV+CKiz/y9CBIQhEh65
8LY9oAyaVk3pfuivUC7K4LkGofzbewk5W/odYCA52KluUFxMXCktv8cEanweg3Jk
SPwABb5xA90RoK9LfvOfsC6o9Vpp7ZvL9KwADbDkrQY1o9KIwZJmQMO/F6GbzD49
JOOkvUBp6n7drDWrr0Sij0qw0qMqHYiqx/rhCCo1s4iwFWXjYeqhLNfGrKaoqgsY
O6wgqfW7w/qfA9lFTK7ber1h81Q53rwtjjIu37WvyWksV5FbuvIVAADRRkZ6ZIAy
gvMAwxG0c0L5BQl+KN11FoDXGs8NVmR2v73mCDrI/HdSk9tjwXuYTqPJaZWTAilk
g5JfkS1ZgYRI2fPJfT/dZ9MCkEUnoebFmRNozRa3L38U9U5x1B++iwZ8RmQcmU1r
tHivWttkpM+0UvUO3++LGSHi0tLdyd0UPUfSRO9vFCEsCKwwuD0cufb3maif8q7t
3+a6RcVDbGQFy0V4mOD9nVOpi2DiZW4HaBdtkeW53BIwvxwtTkHHDITRW+GTezUV
V6nKNRsIvRywcu8gfOMZBpDFH+h2nVoQt3XqjupZJGd5ECCHBhr8VZ0RdA6EfqdQ
+T4kAECNyLF1wliNAOW/i1rqfAnlctoX75HmwA6RXkTKd947qmJtidAQEdPYvRpj
et1/iSLD1eVMSfTwUvwQ1XSn02K48v5t4dCDeFq0uHfFUMYa5AsHl0dwrmveP1CJ
QTWW280D2NLS9Oc+1o+urfPoZsF/0FTMC/XX8gnfTF7sawq7KseHUuQOP/8XOKDH
PGlUXmIrfzIz6Ugh77Zd6k2kPP+mbkknMZ4oi9hbv19T1ImB0hy9yzPM1OP95D1K
S4v6xYWq+ijj4YdupV81bE0pZeEE0r23CnYMBDyxVxsFSHREwOTUA08Txo04HNBk
aKI6/iHQ2dQxUlZFV4hik9wTM9lJOHo6IGT9LD6royNH8aVz5TGELN8Oh4L7rTwu
R7gRnDBE+BeqxG0sXgI6LVcYUzpQsz1v+52SijRZl1AkbJW7I8/O0O65Vo0dntjJ
2bRu2BY0qxTPVGgrB71Aqb6naBe+4jDRSPG0+MeD+H8qTsf1VDA3oZd42PdAlSSA
ncgL6hucA+iuMSwyEqGQxO/lvCWIxaiGVDYM5HjgWbNNJ5O2WcqZlLHgPenE5Z9p
ZwKdsWNjcfCUg3927IZ26l1yCHSpm4kkZ0Mc18Ro6mD3HSlCzPYZuFdqRq3g2D+R
mfFRPT4n70wLtwNifNrfZnsouvyzjSNtSrB3o/GBr8wUjn7IINZxGN+Fw+I2lkfn
ciIe3i/Xk/0btNy8dmWWgZKgPX1U4hoACAMsQYVVA22Bq9YBtQkzZTlbjXHpowF4
XKewRL9BESeoAbnCNTS/n3wtWW0E68sW/FNVyOfymwGXjy1OfpUPuzbN1qwi70Hd
BtQKWHWoyGIPOag7PsTqakq67Z5duOH0o1KUfxwyUQwfjEndDuAPIqSXYBBjig8P
7SefgJ8Swi3NJXXdNLbzFsqLMeCL4VezPUFOEYWNq8YP+9jyMtL/mSFrXJhY+Ljy
duehS3K92lN+svQbwP1F3ZrPRlaE78S/X2R/AqWqJVRHEwdMmaGxxp9YWmnZhnkc
J2KpIghABaiYDAsSh6fNZTYnbI82AC0x4+cTlYdsytUrtEogSE/RDrKbIlIAc52Q
N2DkloHy8Ypn4gGGWVBA8EkTILYA0Tdt4dVKYDBfW1wCSkgCgmRCAEkC1nhysP9A
ft8QELUvQT4jCq2mQPsvbf47huek/j0Tu0nUmkWrKIfkAL5/I2Faa9SWIyLVQAZq
CFS+6X5HWVX91BHNoZFBne+4x9B/BqVEQyAqzy4mRIiFxrFzEVNBW7ULX0dWiM7E
lW3wjFKtuD8LJh21srpliNG/gR6SPGEo0wTIn8d9sG3MSg8PKfs1Cx4dQunSzjqP
OCq3rHKQTHhJeO8FH3M07Hjjpqi82D2cPPY2aa3NiZWmzLW3nuB6WO4kNmPHI9hj
MOKf7+qcDlpjwA5XosHVmrYzKs9fh1jR9VrcCNIeIdLFp3EtbDFoJl3CnrGm94NF
5eLdwLbPXGr/h1AzNe0QDoD1zpbw9KNKviOfN+o0WlN0T7W0ZP2HZ12rFWvj5oYS
Meh3uIDLvawxy2LkqrNTtLpmrhSdzeATsKZU3J7ZU36Yl4NqJev81Lbd1luqJXSo
qvBSaU9YPJlyloUINpO7JPh5b74tjgU7P5LOs627IuNwrdaRoRbx3rU0QXXwNCOL
IHiBZ6Qvt49vm3plbGSgXLoFiBU5jsayOyKnZrXn7i+bA8AYJ4dLp4/+pW6fZTzH
tWa35Rp+4OQVHB7b+KXJUWS5LNmFtj1Zhr+PgU70BfPWiftKVh199yEWIT0up5qp
qUxeOh/wKlFLw7+EybjIYml52es68MOj566zx/Cm8C5xlskgNjGdIiEfK/7Wmeni
qe2JrsQzpgBYbM3kFTbFl8JmOznwuJ9smng69bzKNPeZ9kY3numnn5rGvEZbewfU
p6bVLGWRc7U9MXxG3Oi39rca0Xe5t8RG2bxOdI6P+q2z/qvKfMVwnxCEtQ6bim7+
4DWk3lKYx14ud4WgjZhBRWeEz7SpSLmFj7JZo9MqExps7lhzUhmNwCbo+0E3TkbH
aeixWOggTOTRtdskVtKq9uI4XLNL+TWm0tncn8uJGeppvr16YBvdZ7ENdKqPRf2y
KK1/0adlX/scaMPISMnJq3/AAqzVgTTqznk/pf/kXYkxDCcy7wb9fGB+DmEo9fIK
fAl/s1qSgGH0raTovDsMhAksOZuZ/wzEu1kEJ7bJtTMM1Ho7eoqo+nM6Uu4mTFDe
9bPePPTftASuy2bfwUQpHwyZ2iAyN/+ic4kDQIS0ddYnoo9aZott7WB2QjMxYMqQ
mEa/YNvpJXcxRs1j2OY3UEkmDugRWLPlWLnMK8ChQajzXZOx3Tm3C975NK0BkKzE
I63Jf8SCtYtlzi3130N+VMPz6FVzLw55+zUfANkeLWvqIpyhaRCn5snC+z+hj9QO
3tcuFnCnzQ0Btoz0LjUnQeat2bbo6U4ZTtY/ky+61avA3ewWB72BX9dexGadK2UY
l4fCj8w4K3O8dKtB/TVxy1Ng8YS70isZG1GDEzs/5r6/yLGc0u4zT/RiFSZfvBaQ
FSe+ZPqWt3o1zieTnbgEiO/W+rLXlJO4nlEJmATKxPJdnITlReJuhLz4z9uagpTn
mrKhgrjg5sVzrahiWFunXyqMjrMTZOzQnhzo9MfZVrsK7GXGtTmSFSM7GWSPeUjh
kkLN0sd/wIMSYsmZldvqntBPnQNNPVkcqe8ntIW5AppWKJuic7L1NaQ+rup0r+Z7
pDO61+nnCT+MTnhPy2YP3lWazRwc9N3mIqa4kAIRS0td2AQ42SiB2pzMU77iv8p+
zzxmyPWh4vnvgCClvEJl/cad+UKDYOW2/lczcdFy8D3mRbHEGpFiJ4MLmMWevuvD
HN1Rrs1DjT2rC0RBofRd4d0E7H4HZdPerSv5K0EX9ghoTaikrPx/lepneQ/gHe59
fBX8SMMzolf6XFAtl2DQ8zQG3v4DGA+RbyFze74LooXdh2IUrNLLsTYBsbk/YGB7
JEsw2TIrbA9IU/Im1umWc8Z1/4rvurS1qxhsySj8Sq+WQaDrQ2IazX8+ggjOoaNE
Oo8uVW2c6gMzWFPgqdXsOagfPZZa/ymowtRO9EDqsBki3ynMITyv2IENoi8MvSXs
1n0oYUhpNPZL0cVFSQUUQOWRKc3n5e+O2Cwr30gR8MBEoimUvLz3ccofP4ye/EJy
YeP+PY9hR35TUSSzLmwHO2EfiD3IXS8p+FrfRZglM/1t5krKLZAQzdlA2k65wQ8W
rUvPPccMzMtwvatqYNijHk4CkoZw3dtn2FTTQKxkuh1BoPAHNXWsJESpQXsCWoFK
2FaciV+Omgzqoz6c3Z09N/+oIsrNQfN+zfaToRDoLnwqHPryXgU/AMSX5v3XlTd+
Fxms+rgC7iSPs3Zq6L0uPWoFWttv+pOgCcF9p5K6kOZOQpv/ijFt5d5SpBq4a9LG
F2lgIw7l6p3EZNk/wnTA/GVlsR3yzyrRdCUyFjbTxq2R7+cDWh+zHFZRrpJfV18k
+y40SykmGM7QpqYP8r0TUA6ASN+MYntwd/5+KIPMCqduQya+cDb5OfZRTVh/iUmU
xEZ00FiSMnnVLBxhcwRsu1Dny4/Vs7aCTrj3RSqrjw1Z8PAu4p9DKDbPktu3NliW
ktaa1YUDQwyHRvn81kgGGd+78sS2ROqdAjqcSNyJSdNIVXX/ZehqlJAVMyiVTNKk
ezpgN8ESS5eNx0+Ccw//Zs5O3fjBvdtTAkfpU6omatkAKXkFra8sCDJrs6QuZgz3
8KhPqIxl33q1Gje6YPEvqr+qAQgzY9qYlFaOGXUdw+PaoyTQ+SECO2Mz6LCpirN/
7GfGj31ZVjZz5lKLbcck4hOJ45NPYYNM67mVqZ3WUv1hYlhrUXIDcakb5zt5T1Wq
08UoYlHU/ILD4zTbsduahbltqUcqug6pL4BZ1kbGi6d1uRJmmHyYS1LdUG2lczen
Clnrck6aJdPZcDkrtFMHkkcW9Mj3mMjMjvaFH1BcYPmIS6QF9GxndzrO7ZLHXoTE
K4qzuXG77pKdTmruxedI1A3hN2QkfZ7WINBvN2eUzzyoA0JF6xZSNs2ZVcpJ0cNI
RRqlw51F4XAL4vWCHvo5ZAYPPi11FCINJ++EuREeerPxekYcDHnDYsdHuIrm+5ed
dRer2ZCuouetKo1wvmjiVpd66XiMaPqqrCCXW5oTt3Kx/btuUx0697XVFEkOHHjN
Inj9iELwYpMBhsSNe+NjIuDgnPpvJovkLWrsITuGp0NAmJHCXM/7lgu+R37+VuST
3tU3F6dTRg5BFJNdN51HyVcfNyKYjLZG2QEdNI2Lizq5a7rB1uW3QuVYAKGCUEnP
Ld1ifUpcYR8t3H/L+JpKGN6TuMN0wVBgWBIA+McfQeLk/xMZoigv/o7uGMWpwiMl
zIPzCu6oRfdtjH6cK52p4EOMUv844Vp2J7OQfjfDIJICQQ33Kp7WCqJ2xFRmb+j4
KI2Vm1dLEs5v2bJtYbiT/8OaYzfsuZHkCvvV4syTSZp5qeaQ64BWzI7Y3L3Uw3t6
4RvHQ6tVN09BbuZAHGaSyQBo7BkeNrtkBmZqffXyqWdUdBUIOj8YU6BH7aqlv1V3
fzKiofT3w0svE72PcXX+r8mQwZHS3H7g4UwdJAhrJuQGQMBaBgi3P2jG+Njc3Uxc
rVfF+YLefdxDqZhOV/MNGuYBYJxxsyn3LRXUEHWO8rjYfUYNek5IEg8rzeXhIAwa
5mcm8lOspUweH6ItbjHpIKzkibMRPv3eWpfOo6cs3QTF3c0pFnQqvzgKKth0r/11
qpo3PHyMSd7Vb0oUFq+G80LE13Ij7RZR2DSyBsfYmxp/ZUCMu51VOmJu+gaEZkce
KzgjltqmL17/YfzV8C9sOU2RGGUgKn5xuVtvP7aTUAHThgIbEUGSWbGijSzz2lyo
LOzLTpvPomjm4b3rxujItgJxtZQRwqelGh7X7IIlqdh+KtJ32kwOU49Dwj0HfF8k
j+iSDFZghDGiv8lC6kFeQ1iHDSXKG3oUuz0YroiFHwXLUmrNGLBv/4w++BdAdTgp
Zt1oXJ85gnbMmiy796D+1ABEXcxPaRE6Zv5sJZwwq0xUPEgkic/sOe4HlJyWXXyZ
NQ4TQ52sNS5aaMwn0e/4sswdV0kHYaPDJXUz61ynCnP/ompg2XPvvySb6ZAUZ+Z+
EwkdxT94J/aThHVqhVY/MJgCGfWk6MWryOIRvahXSMk/593DPBPbV/iK3myKAcbA
SiEBZ1+zzv38H8Pwkq1hi5iAAKA497iSE8UKS/I2Fxe3TKJUFmoihhwpSIDBeSpZ
ljKocP+Crvw4r0Z3pjJJE0+elyvvFi5H5eQKuy0QceVac27R/saBsNSWin2iyd/U
xHOdNfYsDJ7hl4URE2s6xy8AA7alqGW7DRaKIm6FUhe8l6GC0L0WTbHObImYHAMI
UlDPppp/edd74RQqZ812LnbZ4PKpSacDH23vPaUKK2a2C/MV/HVB9Og4liybkugQ
h6B4sEYQ+uOCCUCM2LX0k08Qq/5j9fl8Y7HICEqQtQz5Vw/IN1nxAnjURkGmEBgE
z3oWTi6IK/aoPnde9GTnpXP0qVwKf2cVssLpS6NarjX0/CPF17kChdRZOPCTcQer
7y+WOdCC/L+25g0r97G4oG4tntAU6lu/FczxnDRWj4+uIh4EnSJwNGXeeLnRbui/
FMZKjtdxRgbsyzly4eq+q0NNI/H+r/mhQM0ppmTi1fgAT2r+l6fVhIIvoH9BsHvz
VHk7M1KT1vOh0S7KRFu0Q/DiG8UYD+hcr26GK+RarCy4x8O/elNvjEDAsekJEjBX
PpLLCzTyDtdJxpyZfxlQqse6Q/VgJM4kilWc4eKdNdlQzzjF4Me71Kf37k5/WLj/
OquOusp5C0OTE3HOiOYT4veYYDSdbYI/nuT5RcFBSKujZn4j9crS61JfW8neYJra
JY61h6k1cgifU5uo95naz8bzKbFkDS/+nCbObSqWJKz5K/PJj6Z90ffo3JQddmA5
4GBrNvZMfIR2cZ2U6zPkd0SQFMf4a62hqi6kjGR3ab+n6wVXOkVtGlWnl5vkMdrh
DVyTx/OiPaRwYf6+0KyzDwHrmvHot9hhsl6/48+1yULC1KrVGXz6EKDPWWeFAMXW
g3i15Eq/hU6tibavb7owMNUq7O8GsrtmZG8JA25yXe8+0lHEIhQxWavXKtG38sM2
7t3adzeVeGxEqePq+UaXEfN+GgVdaYb3T+hRGb/2kgJBYYp63qJaEYwx0CVK+62P
Bf2146x/Q2nkypACw6nUsFlDGjBb3jGxuWR0BbrjNa2PL+o0Q3HKiPGQw3dXPvp1
XsRZ+MELEiWzh4YTayQL2tI73X1kGQKRzW49gxUZmnpWX6G18hSL42J4IVocxNja
UqgzPuU6q9oSDdBYD6UQEPfcxEw5F7xKg1GbI5aVcgcOh/fNbIH1mK4TjbWgSn9z
XIOA7nEiEmFbgwru7OL+VKXoAYmjHBVJ/MOys0cV6ZAHdOZFyOJ1e21CxrFyDmP1
1c8lwfa9ZyFdQfYwJ/mfHaaVNMax2eh595KzF3yXOUnZLDhGI5qLOmkZCjGS+2TT
MrEdDn6z70ZSSRShe2BDLjqIzW3QC4h8uPgvTQVbh+1jrEE7gtH89pEBqXEj+osn
yljuiuRiRuiP3Jdg6dNgfO8pHwxaTW5wahBs49anj7b6OD4qQtxpe4Osk0Duu8u5
v0oe49PW7Z6TOF4CyabB10LtowfnGEGXYn7M1OBRKScJGvhiDOdJtt8EbJ/592yD
Su7BUb3y/LYnf9ncE40pfhpbs5m/j+4pKCS+PNjBP0FN+woduZoyINfh4oB80Fbg
K6GM+lZXDl8mJ3M1vGxAp8mKleLvEU++k8JLSzp9DmBvXnSgcMj7q6TTrdU6LT4i
WpAbOAxdpjadz/nTVOr6bGb7b77FOIYSqDdGMGHbPBs/BRwzAdICK2qd0u37JvD2
yudDhPtyvgWzfGrLPLQgnrKDYcgLh4v5MmWCPwxaYSu23WdIVo87gJ5be4sQaV6A
uAF6C6JVk1FbnV4mnNb7Z4CZl92ulpE5KrsTkWqBep58Tx1+oycpzNVn8xiBcb9e
H3/MNgaNc4mVh9n4nOuYvuiBAWP9D5O8UfRxcbkTuc2lGGRJo1yD71SKUD6ysywB
hSWyK8ZJftgNR6OYPXZpCXjCwt9XqtUSLacnc07yu/tVkE2QWbb4e4OYtQqXv/bk
98QDAoI4gRu1/6sNpIaJQMYFB6iLg2Su4DESERVnf6AxhfQ+T9q0jrj9RhTgDtj0
jTi2vF2K/7EWU3LxqhiJ6DC4hVPMwNedX1u9mrwqlcfjHQYkl6hr2tAe0//PXbZ7
SbxobY2iiNqrHUxTtF7Pg+7z90VAEM1wf3K8ANPWv8pzjgS3+k7ixJw6mwW0CWS9
CqogjiPlVB5hfWbIBO2jsukwQitkYAe3zWVb8jZC1Sg1588ZjCfaWxPcXzAmsUKT
5PBo2H97wG4lFxLVRE/DJ7DCzj7An5jRElVfwoRzZEDbR3LEc1Iqiot2cZk7mHlA
1H+/OK3duDaMw58H2ckeIksJDmlnTKgMjryltwKlQpWngo6K0yX0n2qSzQAZXg/X
xXund6ikcKApgRZwjW8nvyc21XYurj3q+VOqaoNkCNvk6gFYZIsbFZf4vs2W0Jjb
euYIkcKaBZULULJzCDIY18Xns9/lGm1Jdiha7Lq1Joxk/zjtmW6PDTUODNWeHVoM
NLQ/QFzlTo1LJ86IdqMYmI9JZQCwVAqgCnhq6MWnD7iaMCUQMuktFhHQfzVE8iaw
WJUO5uGWTmaA+3l11RbapptAmRl8CJlpKLfFFm3XDcpoqW3YqljsoxyO4W1UqZ9R
OulDn6EySLwrfhLMytdv+C06LycLPS5oDEoULXLtryWPapBxkXeWT2AVXYXmBAj2
AptqzXvf3LY1+gltSVmpur+F8VJtk1KO3hdGsz1nGH0+w+dkiTbTz2DLpblrLB05
/sB9eS8ivLhQDbGNMMHlT02rIFRsS3G8QXVZgj5/q4NudzohxiyEQhXxkx3xXO1h
ixG1uWD6fTq7OYU2W9Q9pH8KrovEn3d6171QLUMC8n79Nq+mtmwuFPDRBwKRqFqc
DcS8om/lM/NbbETXFnBGplskP9hjwLqZmW/a8bnO8jG9/EKzHpeI8w+kh24sBvvC
7NMdO2GQgkv2IkItVscj3kg7Y8I3HdVWpsijaSouenUaJwmmS18hFXP/kCylxg4u
FkFaPBXRmcjPj46lwlyn7yEhgMxmvb6FHpQFdX2dVMJ0yZ+oO89zdiSAjzpPx68T
CieSwCmtPKcAe9Y++IEBgIyMeRqcP0em4fEkkRpMbTrfR5UrUFjQBLw+f2aliuGk
1Q1Fpf78j5HbVOOlAuM0K6PxyBmHeyRT9GZ4i+3z5MXTcGWTddYLr+H2ZDxUMXaY
KbJTL3e/76hQ5JqCOmWBE01z4ifm+Q86YfghJG/mMXkUxVp3YqqzTQtEqRFPdnFc
Bkq7eJ4OaXvl0zj9n0ts9v5x0cLvMVKKYr49+jCkU6j6MULYLvqjuC40TIS7yCyI
IZPRWb+sRRsdhGpDTsa/qQ9WewC1M8jZvnVAUa/HDS2TaJZ908tb30yU6Ca3cspC
qQJBg6CCij9CMC5LkTCjsEVAOd9R+ZwoQmKkB7mrw2hCwL0na7xhy/WRZRi2JIZJ
EFG/zGwmWXPcM3br/UEPJAxqThJbNGndU93hqFCPAkp4HsgFJGyHRNSCQIsebRU0
AtlIVLD33RKab3ypFUeD8MnX/6XDxCMM4Op2JnpwvpGfwLYLfEVmD6lSZAgGVR92
3SUVNRsE2gzef3lACo1ES4XnVyfqx9N/Vw+Nu/Fj3D7Y4JBjFw61vGG4NO3C7qbE
rG2I+kTwlB/056AYWR3Lshsw4BRPTcSETtqlOF3Aapex4U89T+ip/z9GdnQwdyKA
BUkJM5ayKSwFR9YwR34SNN05nR4Wp6LfVnwbfr1p3J3GEkwexJ1FfU4MYnLJWdsC
ZUEo0oVAQw0IkpsJzkhpT0Ct46Yq/xoftNFgAleKcidGIk/qcDbGy3chGPZMjsHI
EgZo/dphy5JOyrwfA/pYO4Lk/5iYQNCKkPzJoDtdkt0Hxu8lel45ygwVZhwyaJse
jy+5V7RNqSM9myfamZqzB5Qyf4niTs04WGQiRmqkG8vPdmTwwTTylWIBvFZgBUSG
Q6eXfZg6kVKvE7nzfNx6M4Oh1bNwCX/Qcxh7WAdVhCDPuJc0aYnGJmBiIR8V2toA
trFz+ciC5UIwSJZXC5CCdj5fPgE2+bN4v4VHamMUndLgW0UyuHiSSwdozEQBh8Aq
M/jINOPsFrt+ccJ7NPEjOpRP9ntBYHzuSLcGfFDm5bnCbS+1/skPe4GDpn6ommuD
d5BmUJ+M/cZOghK01uFy46qZzXKbBtx5mnhMaFOzgrCl7yxfD0HKmNISb9uB67zF
Lq5S1CKTbwJOG9BuCJ+bQpDu3TByuef5VNMu2HGanrX3UsEktPw+dsh0EzLZgEIu
+mR2B9yXWMdtmR9VCc6pwKBzXv+C0xFRYXMJbik/RYuTdh+X9gJwA6vNkpS2I2SJ
tlrl+0tyTebPmre4mv/H1+LSg3nMkItEwMkX/A+dW6/xyh2GcQTsbj2/blDZ2HoM
fXZfybbLrmH1r3gt/Abs7++kkl9nA0ZLMNUrvQ60mKdcJtqD0ivk1XUCWYBWBTav
DIdQWydQdWtkolgfuszraqev48rqLvS9hIa0ili3JMTmj7hFnEOW/r/X1oJ8nNfw
b4aGmEiuSLp3eJZb+xgQB9NMcaFFJQ6IJuNrpBzyZI9P3C58dG9vF6K4YgnO2Pdi
Cc02gMXzeigRgKNxcb2O+hD/PMphR5iJgHqlZnZtxsY4YwrwENnn1QPLyEuikGo7
xaMhifhVYkU3knDdpMfysUZbppNHjgj/rFqa1kRCYJ50ZAW6kj/CqeG6DiiB416s
7jNQJDm0Q49u8NuakkM2FvvfQYb8uNV8Gjj406w0wir81kqPyhWX0cJa/FSZzUiz
gGX/08xEcZ40dWWSH/yq36DZO5WiECKY3GiCZkBnU2QFOhzh9ofi9Yg0IzE1g4ci
+QNFgRxCqMaN29YT6mog19OjPT6EDAxJ7+4XfG6dSt6JKQ3C0UUE+P0Xcj45SPOM
korcIRT+qjQZJsS9Xr3BbfFTIwX9pK1LI+6HFwQVpLPeE0aZi8ikoYrLTBku+1it
iSjTeByP4t7LUpKNTXrlYPzue3zGqAZEwu68tYJrd7JOIBG2rj2HVf/gJzlKjVfq
pJ638m4J1gss+g9aqwWguHD9fWTIos7LPVZauz2L0zn5v2fOaKHGHg+cJ//Tq7i0
ZhXhY6fwORNlE8i43OtQnh9gaxj4j4zOMA7IT7FPjrMh/s6hECHf/JLDHa5nvD3z
JHvAKoBH+8TA++LVNhUUgEWpmkWyB1ubcs/aAaVzVEuXbMPBR/CIHjGvIFwpnpx8
3CZSXdzbJk57ig1zn6gg0gc8V/4k99ybNV61rWurbQvgG11PtjImYRnSZfAN05Az
7iv2FUkz94vCsPRwVkjk8rnAL+rVG6HQ9URCVMbzdMZajR/snx2XjuDy/njn3moB
lvV8JPQ2sT/GHZnNN8iJll0K+P5c+BFjV1Ue0Fm1rKPNdaBQ+JOfHHP7he69JydH
BhVBvf/RC71h2XZZFvuqeyuISfiYyoZ7nCblxwV2hGsQVFEjG2yDfB8PaJ0vgD2n
aryToagI5M/FF2tVMTI97T72RgVjCqCj6kV4v6vLzLGD6PL60dgDU5C9JQkNVQtG
kiuN3FKpl3NWTK1lf6liwSo6oC3eLjX0WXsEF4swNkeSo+zUsXyE/8KAX97If/X1
ur7x74TrGpEc/nJTpOYAPpLgIR5fGbjzBJLCo/0o2gqinlCmsgf9e5yido/dKkGU
9Q9yLzI03V9uCG6yMxgrcqOOgymydTgIFFVri6G0EPTfCZRBEQvyNw3jVvWpiTaq
A3DttIEVvumNPffTRCdXGImy5KNMiMhipatDMFJiE3H3/bF/rkNcztQVlEFSJf6V
tVA4qrkg2BL4j/KRPoyhIIqBazsmEIfLzaV+/9VldhMKGDI4L/+62Nxh8HUTU6Zs
lrtbs2RsStBrNVx5za475yrkrSZwWtRcBaWSH/BnNLaL53utSn7uF+MI0im5Jha1
E31KkrhrYmO7S4orlFH5su8emYyCXB3ip5Td6LUUPvEiXwfGj7Lrv9NLYGnJ9v2+
mgVAtQYHwcz5acfEuyUkRcBsRHzffzv70GIONPIFLe5au+G+zEsPjyFF7CJg74dp
TQ0ZWwsJAmyGbf32Lfz2aY9osUawVyUFq4KsmUn4MrfncjmHMV3t1UPW1OniG/jg
nCgxStiyu5JfGBxHMYXPRVnH28KJ3+5XM9Jk+jh7/WG/gv9nZyqz23dcgehi9TDt
5irIWJRQXz1s1nJR6zGF/MyNsuZTfqzcBfD2hf5+9VSKEV+ZWQairiClkqa/exII
QFswHwoJF5SSLumWqX5EcNCxByNzSIqnA/npOXa3WTk6BsobCrLgnnb3EEePgse7
yFCaQwamy7Pa4P+XIOYPHBbhQOG757NEe6/T/TiZ/2sC1ZuJPldICxXbAsLiyYju
+pDtMxYCuOHVdgMgo9ofpF9LAJmNY7QDwYE69sthAXPbvv6jAHhyqH+QMk/kBH11
XRq0m/VOJVuprvZYsL8+CF6EWLLd2GepfyJIpv0Ck20TEhhcvTBwQ+wRWcistiua
yGY5zngqR9MUKErRc/N6fIjIBn0QXavAz97q+ngxm+BAmW11g8/G71s31TP2km7w
/h6OEtLDnH/Xmzn0uA9gTFRCrCMN9LnjjIV1l1pBzeDkSeNVmZ6gTLfWlUHBlHm4
Ub7vWOwGR+XWQbPyCIsXqjJAhIEtcDWgLg6swGQWp4cok8eRuCuqwPSprWKs334r
RisNAoJHTIyI47qlRHyCzPqpdhwUNdD5SCFxifIyc5fIT1u7mvgrnTO+RBqSNTkM
BJcYYMEl7a6kDxDghzZLnBgweHGhfgJuQ24hlnZY/8kZk+YffUy1FE0abMv9nQP6
DEEQJVV14hprY7ESba9ftnzgHN7M188/azkUWf2zIxDnympLzncZmTtAXqmQyz/k
foy7u7VAjEpDuC9VVnC/XSOVh60soR0cVf6qhV6zQ/DfLvkOp9QnETIbP9claAab
Z+0dlh14areF7OrcBkFZt09GzBwxFCL1iKYwlczsI6QSZByD8vg2apbbQv0OlAAR
Q3BK0Hbjew6Ovjsx8/rPFSOZCYbUaR/ldc75yual0AUjQ74mcvKufIqs4kONM7/o
STn+VfQ6VXnghXbZiYCNQCHurSFirqd4gXAuz9I6ftiTJIWit7myaQw69U8+6HZV
7viasXNuPvmDD3DaIxOGW2BCv32allBuWoJ8NjxjfuvrwGDrYREk167c2ZS4G80H
O8J8pijQrluQy1ON/9O8mb943KFCoDPx0/wYieWzxI570xnKK1xmky2JRRH7N7ma
eJ/Aip8kXisw6Jh/8L2s8I361Jm3jDCUdSeffBfYnXmMAuc5wPtPPnoTj2f8qCP7
Rb6by33mxA+WoQ/RjeaAKEbMGCf1UWBzlt+L5oBu5TpNRIe8BVSc3mEbRM7daJ+h
2sVzzG8XIeKgWP8/jtx4wNU5KRN4p4Vlvt+zL6b0krEU6zXNiX85pW5riLIYEpns
+LzUmk/pSkD4hAyCrOg2G0eslwVK5BbKY3rlV6c0IBgApSOpy8TwHZvQ50FEoD8b
/vP3CBjjPU05ujfUFw0o6yGVEEM19V186U5xIp9jWzf8C1MR2LlUmp602wh65Mrq
Iiza/XAqqNft8iyEX9v3Pwjl7t5e6gu8zWBcmOcdgHbcSbzJpUfx0mpj478H5miF
FLzc6zSWFfDcUVR9cf8XSA1kGx7HcJXLij4FuihV3ZO0gyhRFiHJXsrIRYJ+NeeV
sdKD41MKjVdGFesoiAQSz8vshh6OHxUI11PRWQCzY3TFyoAz6wWjV6ZSpRkiMCfh
rrRMxUj9DCR9OLTUmTfj1wwb4aRWdqPFd6g8gKZNq/vny65PBVE8QNLgiMMJ51Mi
DcKc16IXIrJA358SihcurSpKyLPn2xpeTB4iDlCGMARQPWA01hIuRIZmO3wDWpeg
EnXKisrUHWYADDRdGQZyeUmFa5gKndnc4ewbN2yEjbFwj1R2HJ6SFmF3S8EmKGUI
UHRToE+SBjoq7mE9IoZjlIi0M1Arial41R9fFaUQ29kUnViFW0SOrPiAAEF7AwbY
tG0FL7+oHUNvTidJWqixc23PrpqdjPGdLMqheoONZiysmBnlyYKlhII7Wf2mSznT
YDw+m8Z8Cd7rNolHrVIfgxyfzCXLzNvxnqk5TBC9DBKR1mrFvU+5UTiSCqEKMSLc
OVF/B44J68z1grWAb3gkX1wChDXKQST/9+pNoxo4AeJfHRfeTrrK5WIVo/2Isn7n
Y6OoeHo+zpu0Q9fLwWH+y2vjpgB4SVcgAJ72uxvwePUTHXh1mx6Xg2bJwVnE3P54
ZWlVdHv5awz4X17F1NelWO3U8quaeJfliFmrpkQ+SY/Dq0wpM025yHbrEfj6h8fn
Fs9dmkFMlNnmoOQKCQ+6ocSfh7v40hi3vR0t84Lrn2h+uPxTlUBU2uWmfiqr8gtc
iayttPlfkIDpmeLAuzuVh1YwKjZtHjlG511wONiqMrHKp5IgceXkxD+2L3RCRvU6
shK/U4nWcMP58iMK5WWWyZnX9N7kd4p11Ag9jEto1j0yiJp4NBg5j9r/4M0fE8+U
f5ZH3y/xYdWV+kviFfgd5+f22UArQal1vUAZHDRn7mYoN43ElWb+SS7t7a+YGSkO
1CsyhoC3udbWDMaHengAufs/lJnUrdb471G/nOIwmZAW3mTBsxZJO6c3vI8rvwpN
yhYxUwOB7S0x+zt1eWJFuq60kC63MckqZl4m5rHCq/lirNcFzCpYbXd7In9H7F+K
eNqEvWS8xNbq1znQOBB8l87HIqrQ3jlnDRR8YX96Zgd8M3C//rJA/CU1L+Rg0PL6
5qUdfBK4sXIm+QV+KV7uUBO65qRkKfu0q96FuipQOeigcC2y88CPDF5pUcGe0A39
Gex6luvNb3//9bgwWyvR8nqOV6m6KiiG+TOQW01optkjyeJpjguQW4tJ3mIS4APB
PmVlVNv6oudPds7499tkac0wg1wWYTsv6bhL0DVRH5Eut+JIitC1894QKQuCdhH7
4U8kAH0ZYJm+ngGaHAnpRqksjfTW0MSIEwjdgjsLL56LBDHk6GRaYXjJFHtQMLD5
H23TFAIrWqvTCNRy48IbueelmyNpbhA+zZDqdO+G1vHNDdwSNBg7ANk6BsZr4S4I
V3N0wgR7yiK8h+nLJSWA4mPPPjpcRefPmdIY/VJ8ibFFNnYNZMLqS3CmWminqZxJ
f7CUpgm3C/BV4X6vgaiXZILFVbhJadImbfXDGi0ceDOIa/07MYC9lfu6zU0fqEWH
lW6+wrP54BCTUUNllUppf9aWa0APzxoLxZNttRr/WltEqZTzF0iwTgn+idy2NW3e
FuJZSP3av6ZL1fC8KgBShUe093Crfor8dtllVGeHMuiSHM756mSZ0lxfE8p5wdgD
pCPB9CJmRr+FOeyoMh+pSNquZVpBFUCIgIDS4e4SHA+VEpG2eaIMF37Lo1QRLsv3
7uoQBv6g6yKNC8jpXwRC5HbN4ojw8+SygeoPlS3khUT+OG3H0XwDtubXdpLpmdtr
10AshJ9EPG5S2rjItGQuAVMM1w7gGKRE2mkNc/JIgtpgv2ToRTK8IJe8YQIVObcW
ezHlo6auJGj2jQSon/9VPTgvhk6ePFlcv/UUDhiLY5QpI1mJPEIrxd2ZFdKZyJod
Wvbhua4SSF8krZyKfpOh5KjBxQkrWZW+7CEwS2rJz/GZZ3AR14iIHzNTjRTEKjvD
1a454ZSG4uaoD19PeQChH02rvEim7D0QDRFXvMWJMctAaPs9h0wOkhg3SjACMviM
CirAaDEDi1ZEUWX+Sb6g5vnr1S3hyfP5og6VuvSbNHsvaiBYGrctZJOlamVEs2tK
QBSDZOwJwWgiwjO2oOC+aMq2rc2iskb4tHdDadcRSY4rCpJaXBSt/VLkB+R48hBc
nV52U6xTWTeO/JKYWQQIjdJeTXdgBhpXTMYOZKu9k9IvsP+02VQedgykhOe0Tw/z
TekYaqWAguVBQPNGgdlQsDbLmIyQyfJY03a4JC8NBSvBWfxfE1qOW6NEAy6Qa8mb
nKoVBe1WqGFC2ODUhClQASw5bE6DsJOj7s/IPq0xeoTSSPXb8bzwrtB+Ybyb+bzf
bdv2GoVM3IcumfT0mR+0ykEKMVQkGy7/QjAIHghspSaQu7q2w+xo9J6caE5MbDMf
ogwhJDQ/hzppAIX/OocyxuppofHj9FlrwlD3rO7d7+WDmSGNVAwgvfO9JoJsHMzj
aSPvJ8MYKsgPtjYDCdxIBkmi81ufRgJr8tiREWOLHL9OXFopS2a58DpHiDCN5rkz
jhx8S88hAw8IeJOoeZemxrT4yBRolJDH220bWKPfzkLdeQbTNpLI1K7rgVuh/5KF
xsF8CQ2kBd7VgHme2L1DB+VpOaDuIy5vHpfGZt90rg+JE4V8Bz4xSunpqtnaoJR+
oxaIlyovuCGyocan8HrcFYeZyhB2ZnDOikjteSlurkf7LQ23xge6MzA9PMaCjQjK
yAXriqG/SU1I8JI2KhO3mlV83GZLnVmwJwM9dnIsvx+yuqTbpqf86Wmsa1hSmXni

--pragma protect end_data_block
--pragma protect digest_block
XS43/WnTiRkGGr1GiEyoY/rNiIo=
--pragma protect end_digest_block
--pragma protect end_protected
