-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dJjgVH+NwZoF+J0xRoSL0k99ta+Ra3CStqC99um1qp20DzGnPWJQQIR+CnISJKqVZyAIbUgyFWHb
f7+D9pCEti3WWKSk4+/IBD0G5P8+37hH6uNyCj1o33VHBAlX7nQ307ZHvRJkmAmLjNHSDd8xg05O
nidyqK16mpkCw58iH9+/tVENZB22Vw0g9BPadCV3bFVYYvgm7vV+trLn3u8GTSYcYvLi6gGbOqUm
4zpj2sQ8XBf3lyOrLhyq/7ZwKkqmnbYCXlD6cc2b31fWTpp030PpmHksD9f9J5MYYNrStv4X9gsC
XxtJ3tV6nAoYdzpKin6TvpBV39WSLRARH7EITA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 16528)
`protect data_block
AUtx9RlXqLFYfrwZjQNlAOH+U3OOt6QkJFcFg9rONgaaeJYBmDUFrlchn/TT/aqidJqx1K60+Aa+
g+VBoBnI821bbZ1URUMkfWFygB0uYASebPnGpN2HFsomX3pWATHR5JFlSWrExcGyR35av2CpA86u
AuFsKy65vg7B8Nb2y+Dr+fayIkDXGFdtS4imBYiH8jzYv71o773cqHaCk6iG/25Xa7YCEIHkhQst
4AGHHbxAe9wvw2g9oASC1TJRwDKuWwWT6oWQD2ex3XfBE7X+uKMjRp84ybyYvMCFIKMrSpjNJnZq
+4/Z5GDNTzt2/TcRZsW85Nqz48/4FNk9bfikQFFdWoBYF/Xw4ffVEc3SKOg3k08Js5NIDaR4ipH3
Ejtu5CfVB+gxTAn3yoC8bnYBvXR9TWGa4JYMS/itxSLojPJGxSWb1SV1WgIWAroSSTKB/N52EA8n
eHh8ZDqdzhpWTn81pfd31ICkXkLISE0espkME886/vrOpL3gecSrc/vT6hw68mjbqJhrLeBchW1F
cmT3AJTtw9iRuHwZf1F+c3TaJsXgbLxTCJsuOoDa6hNt4O99F3efSF8ErdgegJ0f41/5yLu3ltLH
fZ+gQgI1yKwTpTCSTkx5XR9y6MlP7gqPTd2bg13girsrUm/e4eR53YCpEsfv9409D2+ISLnqpXWL
9q/3koKNP3GofKqQ2S7O0UQTzWlavA2jOeMLHGWg8g7R4/f+ZDh8Um6Ky+Zcu4WIArDOwru97cSc
fxJj0SM7tx7reGvXH/AB1DgTqhn9iDoVxE8JARVAXYoNqdtSjb81OtzN38OkUEwdcI+ivX1SvDic
/pS1VXZ2G92moQTadESvC5kqCI1JdTWveBredZCRqZcEm6JXTw1/j7OZ9ckP1zHu+I+3MAEU+HGA
p1GAeKeE6Pdkb/X7RJxlnh+peqajy98v6QiDnWUnHLJ6LFRk3geJ7BnLIrzLiKCKxEjf4UKO7/3A
xbCEhMsJobK5ZH+fjKwCt2MlCGtgG8dyyYWqbK2DP/o6okUb4FXH/pLI+GGH2q8X+L3ul/rmFu6V
wMbKTtI41NPoSWi1Y56A2gPsupsRpjgp9+7gv+bIROcxBg+w4JrsODbj1Be47gdJU5fd+F3Km3x0
Wtt1SckYuDKaKSKJCJ/CHBkf8dqJ9GzROTId0nvUngSc/pTE7exUJ232OcELNDOwtQMlQHqq1ehf
pY/A4qad9BbOvad9Fxw/U3ngoLOe5MAES2MB78242SlUBXSADQAEH3NA+lh27U7RAGRkKd6Xgluv
Hvii4X8bW0OIq5SQJI6eD7IiiWZonHJNjIAE0nn1kYt8H4giKYwjFmPds/GrruBrR9oTmLpLqQdg
DfP9q9wSbDXbBSryP6btHBj8AcW5KQI/tzk2KBXQ916lipcpL1jIFudOvdZCBZu/N0OeQO3oHp1M
kZ+XMDd8d44b3atakzypj95OttEOCXApFDfkzZTc2I+OZ+ZtzzB5dJttTUIyhDyEsXA4mTviRhCs
XZNQkYmplMtllSfEvcdz+t0EwhL8s5aYQrkqX4ZOXyVJ+KqseVNOlH0jq3Q9TnW2Cyc3dI7jDU+1
esRns7KOoXc2E2xYQRuZtq6qkGi32Km4o9Xn2qUGUoFt5KxcDWiQukLuWymRBPWj2pU3hbfpDXXn
WwGOCYMF/08NrYVnOQTda6saYapDFQ7YbaspPifmNke3/WjxjmrOeIHCUcMxXMR+yHnobuLWwiCT
BvlW/J7E/FjORHXb1kjy1dLTD5M8IbhrY0IRkp2FCkvveOTKwHh6VuKxn1LvpPwa84nW6iBIWRcM
+WfLhOcMR6cTumETNhtBT+iJex3OU7nMyMjXBIT9TmCnU16igZT2P7RHUHLxIsrMKORF0v/yokpo
HCs6OTM+D9X1dGf+5hPDCUlipjBjskU4stR5nyY97RcVBWSbYWmcOer5S7ssxDY4dZ4d8+Tkkfw4
nHqv2AoBhTX/B2Y5NgNTuGhiqiD0MWLUKPpHp9lPrNwnYEFX4LUm2pRDrfAVI0LRPhetoLLsLsdR
KRjSZycbeo48uM5U7JmRINLXYyF8qL1D8Wc2vNLddgUsngv9udTgJ+x3/9hfWcBo6y+W1KNlkyC9
Gb9ANmao6tUc+ZZ43S9a87WPcehOZfWcwWydVbzQhMunTXvT/gLFtR93H9PEgL1W7BwQyLWHVB3S
pK6Vzy2p9YtiX6g+ampqeI30j9SgyjnH3od2NgTkzqdh9ORBVsGkC7t7Bbls/Byt7EMNqLTHE+g+
aqDMO3zTaIC6lRZUL1AmhufGJt6MZCsNh3qGpgVNaSgsrawqiH3YBlHcn7mQdtDKEJ8hOYCvv12x
G4Zty00nzbh5yTnFwydhedff+61n0nIg2yvOg4oSO+QuLsTdXLjDcss2ardZOLZtw5wmRBEQavvr
vzOwJmtMMTfBXLIxpwD2daYGltHpiwvLs8UZEbQL0FniJeEpa3TrGU2iHUXptLgSq0lqMJO+uJHK
OADO9FZdqDJ2DNZOuyQJW8jzf9TWbTh6lE0kACacLdWILozEtCtR2lFVQMDBIGeCq3AD5DUjLFJE
7PgU282GGbhNhuHtc4Gmr8SDmPpBdsOE11MHRElqQ1iiT7FEbhg9KW3f/LELL6Wtgfh2r8Nm1TYT
Y0sDeHXiMk7RO/hRY3byzKh8pQK/BxUdQ6noX0Y7Br7sANZS4tjIx1uTtmIwgpEzkL7AZq7wmKhz
6i2Jugx2PmTQ5EBjEJFwIiMw+7LBaoU4SuIHG6SIwIoa2X7hHbYYt+Pkaof6ZYzyCNGP7gTmPKXI
8vCCqoReLlwYliIxq3GWRVY0xbH8VgXAceCwzOVDqX92WaHZTGCuDAGnDAQ97bAee4e8AkafVigl
aKjh07ICWAKMu6N4eJHWWKKvlya9hhGRePdNJ8qvy1AobPNw3i1U0KcBhfUzv3aYEOXcG94vJqi6
DUCJL+Ti0TP+M27n4TuLLiPBtdzPUnAAWTXWcR196Nnxk/weuzsK8NRtJu4jzrf3b9zRXnLwrIxc
3xjgeGi7lVGoxF/RAMutxR1EWT8Rx5qby9Mhebq/JSQqcHH871yZR7ISy7e4SfpQxY8vXEspdfkw
4pg8A/DfaFJbEnCTlbI7o2s2PlhU4WB9aoJPJfMRM4EweNK4EbZ7eSM5fLN7QgfUqIlGjWqeItfX
H4Kn5BTBa7LhUkwTk7x1ao7aF+pNFUQXsqFTTN92DU48s49gEY7stSLjK5VDUMNGnR9wsMHBCrD/
sNS5NlG0414uu1ZD6UBkyY/yG8VGcZMX59OZ0MNOsFXU+cE4NEHqaLnBFhU6jmSV9T6/UKdk8O8x
y/GluDNzv3fyesjrQ0g0zNfE4jjD03Os4wyrzkiJuf7MRHGHgMaTPG6eYOcg8t0UCDduEw9d9fLl
Jgpc45KaW+bs1t1PycalwnCT7W3g5XHoCZb8E4s9ImUp2sOhk2KlchW7ktsVgGIefxMJ52l9o0aX
I8WV6jHkPPX1WHibpz1EW4lQwof8oo0oP3MSuQIyVhtgpjC76TgaptM6vFibxmxyCVAc91Mvggf8
yJs9+E51imHxXPxeZS9mgkJypECSLcZYn7CAO4MvNempiHgJxEYLv29tbOieolMADBtiTHqnyupz
HhF7ckh2/zv6x2sfBhHIDICywyAKzrF1kro6GhEUMZWYP7bhpaq9zNAF2l106x3wICe9a1AJ1fcm
xvqPQ6FiutMiM6h+4a4WRFWngAPaG98szSM7DE7Wcs3lnh13Nr172TAAWfBjoTozsP/+hjQXNCTR
VYx51ZK6Pqqy1xOFvNeg3NeGLwViIA1NrrOlECYX0OvYeCAtiUfKeqpjkBnCOQvXm92SiRGWoXc0
FzPLBa3Fm1gEQTboM+agvrx08RXyMoxOXk2eGVJfsOKIli1QzcSWsIEnGaXzCAA/hm5JifqXt8aH
jRKYWZZl960J8kOmEy46uX/NMua8i0+t302bWVNNCuZqBy47mcSyxwYiS2fvvs19GH2LrTBMne0I
mlMIwn9BjFdjlW5CtJ2xX9KmkR6XgIyqWbNE8sf7xIklEhAeZjP6EOwRk41nUcM/O8Z/J12A+xWF
M5lXKrqfKdYaQpO2lOiBdYZ0Umo72GcXcLGyj28YOuZuD2wWyFg9wVey2roRafXarsI2WhTVSs+B
ViQPx8sXH0olxq0nYWyP7MRsvitGPlNy1ul3ePlnDl/gY5bvtcV85TzQDX5btH9Tkly7CTmEei7i
AKEBXvOHbuDu70ztZz5OycEDuY7SIMTgQrg8S1oH7G6E15hY2fiaSUp8GPqC9z6ESw///3ZoS52c
sXcrrippwM2uYlXCBuMP5SxebstT7h44Ic5dSS19qsraBF5n21byUUTvTzHbXkjTsYdaEl7Drc1p
jir23jn6wep2Neg4g2iWQs3jWSycuy0yBsZrtPSc/bg0ujj15Mrunvi1a0ZsP99X8Ez+VwyipVXD
+2/C11R53eGZgQyjTo5qVqog5Hbjq7F6Zteg0MJkLhlAkxQUiSoKxUwkkgZH1YfIkBfZzjDZTUXu
p/7i35WG/qbk4kXEs0KzZYcYTWsygoH4TesKmWKz31hDmEEPYdqPmUnqqPIoewvq4WnTnwIm16tZ
L3LLion4BWS0H2BlMOxXW9HfQGD2dnRmI7XpfTXIEEI0y4CByMMExCAKP5o3qTSF1C15uXn3pe2/
/nLLmPQ6R9oM7LifnZltMyp/sHfbSAn1mdTQysXIikRcZafilp7TRKaxQaMl2T18Mly9V4HtcuCX
xEaRVtOW/IGjQruiNSHfbmOPdjx2TXtjbaCYE7Q4p5qOvjHaYY2uCk1/SAayTghI8MRWCxpmcaib
iNgFgRZFxFqOmphab2eOizp7N0OsVCeWYGMA7l92sLgOm+unlprtVdnmtjfTDZ9vnzQ+gXVO5+Yo
8D5wujBPzArwDRrGrPCSpOby/ILCPYl76DUC/djRwIVtxHShWVCp/2zWrIr7OdWHADwmzLDgiqr9
oVMJhHUsFlWdwFL7IPp19f5WewfgK6j9xGyrNVNLYXKvqvYRtTvaQRVmQgTwaeDHksOBPBJx0k+Q
215bVIG+x5ZZ42SdkmPaewiZvOdotTtAddCY0RD1Fg+c7IICRc9xuR1toOUyqG6aViD7wVQjog43
gySbzpsNVZSS8rmzoAaeChJDHtvHRC31vdcpzryZen5GRxLaY7PzweGnzcme5+TNApYfLhVoHeXu
dd2qia/jAhBl0X4J055LeW21BGoLCTDp+3LjbRDiUgJniKpTX7rYieDgY883+AROlMAp6vbI3NOx
Pjb/HHKOHi5FCYGjav1FTgXPOZhl6z9DCNCDlzIT7tSDh6WqBHpPtmOzWqbtk9AEaofm6lErX9wQ
I6t/WYKLP9m5mq5BBn+DjCjD4AGyjSnE3tBhJ0GJ4Pqqw/U0sr68izXNU8Jyz5n08NUbO+sXimLv
vPH7od6Pxmqaa/gl2pLPtt3hhQWx992AAG2LOAnPr7/oBZX0yKK5IKdQFj1FD+fVGWWlBP7ZBWLs
d7kIVJCkO3muGtT8V67n6e0u0QWIVzCOHaaRQSOz4SmjY2Dy/qgBwboLtsd6LDLwKxIIkuDqsrYk
bvSLgiJe9yVmthV6GtfQIX8T8UB6CahmdFRF1EAyUIPmm4PJhVZzzJ9n2NMi/ct16Q/1u/sJC28w
/z11hTR26VU22qQcUkswFtW4selba/JoTLhr0BBPglAXyadvDfa/fAiRv8WDMMfjVJqXNF2R24SE
qE61NPhus+ekpcTHFIUkQ9t5zr7b4dPXQHDqYKAfTryZKRF0tB4pTSovNCoef9EkHpyzIi26HIMd
HFPeCQRFnEHAuePZWtwEyNW4vCVnz8NcdeUIM+n2UCbTuWGrBNxcPCTUX7naIMzil9Grkn38j/1h
00t7I7sYfQTd1o76GL6dVmbrCi/wdZJ5PSrMtRGqHmhHm9rGAf3Da4pMDQoZD9p172vw9A0ebxT4
cw+JNfK5pkwbcZMEvMDmFMAIBZg0f6BnZzmR6KAZK7gy0/dczqo2iEblXk/q3jkO6uCW7m2TVwZj
YSMWHzVEZLOi29znaLvkV572jrp41CiYxv4UPlJo6vaCUDU3On4HqvXt22uRyejGnx8O4Kyf8m9I
Ef0srVPIobNlMnn4f+vQE6x46UIqDxyRZ6LrcYqqo1TBRgIow5rK5piQCFTMsoE4Y9d3DIZGtyGQ
XB4zU/uE25xpyXkClAK7o80vSKAKsXFqyqUqyEGkv+KDfa91Qw9VHwwfrZMn5QIiNfyLGevjuFZD
0G7qF4GitqHgGWYnu96n3fCi9lYwMlyBccUTlzgFhHUWpk5GPz0b0ZigCNgolHhw4Vh6XkAnt+dB
ehva6xXyxZYtcIuXuW5i72E5VqIKmK8YVEBYT1lEeyC9rKMLErbn9+d/5gJ1cH5CwTkDUrROLlqa
PROL+bwn7q/88C7calss6aBPlpdxq10LnytuiZADcD34Hyb8ygBf7bHjavQ4TlE3aFMLm0WnwevN
XkQVFWjpC8yBenvfKWH+utwFERvAqCeKGPsHznlq1daiqUNdonPO9+MT0JXGQzzZjajFhPokcxxy
j5Y6mZSAkbqAQ4owDfN5WqzTO6d1bmxsFuRuX+3pQNCuygHe32HeatRz2OxhFPOtN7RXc4J6PQ2c
Wg4BpcMMX8xgKWRbtml4jCjdZVNzWnsqoZ6XtfKZM8WMfgfi0Zz46ezMrADEpYwUnlfUqn73Y2rp
PS4Rsj60CSzfmrEnaaRy2ZXbDTAvUb0RdNeD5PbNZIqRSYleEnCOLH2kB8v2b5bcD4U/bB7WUEjc
XJ764OoiH6FN7WZCzsN5vWuNRoqTfc1BrnN8+0qTvgDbkv3NTJdgz4zFSXMysDsCB5FrFJDW7ovd
aJhwm/VWJlktocqpCpM2gFce5koGtQQwfCTSjQj5o4inO8LTlCWqPz6Q4/Z6Blfv8Ya9HxLuFf8E
YY6F9jDWpuyCuOmKhJ1T4mH1gRbyGRzvAu5DedZhgLmW6JwlETf/HLXg6EVnCTC4TRo1qRXfDD54
uzNOrwhvFieUt2JKoF3Y/SIxWxyZc8Bzvp0ljKsOO9cI2lLFl+dbLWk6WQO61Qj9nxlQ9ufVX0hr
+NBFEqI7pWvnhnF9DpSL5DeH4h2ZneUYsnqVHIMjKk7EJ4/1v6nNXAjk+cNG9MrY3ESh0zBeOE9M
aubHPSYkNATi60Z4ee/B9kykx67SHp9mNt0zmVbRY/B3CGqKj6HvaFVXlFhqy5Gn30W+AlfjQRH8
p00oMbheK4clwwbeCtPJ86esIlSJqHv/N/yxG2Z1ysVLZw13DhX6Z5YXgWc7XbrQ2nv82FjcXzT8
iVM4qC4f0/9Nn1LOLMvg37KrMfm43Fu/tzt+MbPG1rzc2F21llCPdGyKskS0DplLOy6Q7AahtKLD
k+Oj8aWZgEBXjNQp8eDJ95abygpybM2148aDIzvpN9tYMRYaVOSRtqXUAQnk+kmdcQVp4mSelPDU
/tsk7+9rw6lQYCeZG5juVQvcaJrRRprW+HqEK41wpNPXFOdyTKNiXSV6vhlsCKam1/yn0DVJzoOB
4Vxqf+3tl0X1xCmQlGnDfnN+rYXW4UwcOHBDmCPl0fTcQ8HfWCIGBKhtO6WkaQAVcn+yKPYRW2Pa
awYcO7t2n/OR1s8V0OTMSnuorSn7e/37LvyWItkzx7In5k3jHITzpmOG8YsYtXG3qpGXPdiTicew
GMJHOCmqNOWKnbpkyILfOXXqhDgvMbKy/paD8MTjpmfsK5CtqOI4jNj0S778Tiahy3CJwqlspBIN
M+BNzzVwIDJu2iv/1ShfKvWLrlF+XEUShMihSWfRrzcqXogik2Ye/fsAItKLZiJtDS6cupqW24X5
ZMI2Wx4M+cYubGiZxi8T59z36zidfnvX2fe0AjO1w5vmcj9cHEtpcE4/X0yESIKDBYiEbdv6E80m
ZLeg9Ynveh7B/8nxNMDTV5FMjV/xPj3S2U5z/YVM6HgC/4AZ9dILeOEC0/DXlwZENMUgexm2IKsZ
Nj/1Fo2e6pqiKm8m7FK8s1eMJWCppMXb2ccWC51O0qtiValduAfzNgJqv4A8roHMjOE+OtLJFXnk
JjQ1KDwrtrae4RDd2CTJLokLtkGYdsI+GF4FGhfcImiFL7mGFFlJQUkL/mnXEXCBXHEM3bnNm7q4
84Ozy0dP7RWLTV3JfFf1GLBO2o518Tzpdx+F0yxyfNfx5R35tQOA2V54ZtTYYkpdZH8P+FkKWXfI
kUkjqq5ADFJyKgjYcasT89a5r13BiwnDEjCldcDM3zI1S+aElZHRHqZ3WI8bkHCHug8txCBRAQ2r
1qmVctvA2MoOLxNwR46S736OnOwZ2nN+UGxx28pPH7sS28+FVfiuo9ChK+pAAhncOqzJ4p12CKo9
+mOcZmQjK4AdEniXRi8p2vkizseKzwEk6kOb/7P42amBagtN/iRzfmICyKk7rOTetb7De17VexFL
/gRC6oTYdZLcvdZhAgBXuyAAf+wBTU3ip2A78qftaHmmpzGIuGu7T/mi1gTLS6yJGqyeCz925Nc5
28iRLT7jWz/CfAS7LWHExNCDpv0aWSIiRtAzzH0HhUBP1MgtrDAhp58909ea10UkLmDT70zGjePu
UO36P+4cFcgLw4UP64GsSXKws5s+0iEh/wRpxnbh3SduIjZB9m/uLrfDsT6phAdWSTy6FUzLpxf0
m0fI1hiCaKns52a2FHIxQfNOPiQ5DGnvtNnE2INTjZZpaqh9Vi87DhZnA9KHLOAiXFx2SoIcn02z
AEg6++FFQBzNgsxq4aUPWhPb/a9kDPOGz0+b2UQi8977yCROZO6/v7A6EYiT3tx5jzil57Z8jVsO
wtQmHcPTcaph6RJSVWkD1hI1+aUKq3LRiDTdzYA/b0IjiF9Cdr7BAhEjsrgiA7KadDgcT86Cde5f
MdUajLOFS64tV9GAaSKW10vJfyc5PIUse1LDsS1i009XasvRefdgtB1H8qqHmAhPCwJe5AfZj1Qe
nFdq52bdU0XuzsotKeCo+HzVcAYImbemnVlxfPcoKGHjILGbSmGzQul3vpjA/Qzc3pJhjBYPVTJu
1JOoQP4BMjaF8H4WSIjO2z/333C/SAoP2QscVp3IUBj4I2vlVqyUw6Udztqfm3NV1TeoK7wW09FL
PgGDbfnbeWFuxH0AVvypg+fXOW+XJM8G0/HAFLvne6SOOVcxsOJwR6IRztI7DaIA1Ks39dLhQ5Ud
Ep3R3Hw+Y5cBkESQFmVmRYvhl3xB4rpa0tOeiOKvrviqnvP0NI6nM06Ct9sOeHocZmNEsPg2gnFC
sLicHaxuG81nyn6Oi0S4eEP+878lPuL0vfjhNncIA+RyCgHO16/D+qiEHYgJlADhaL1iet178MdK
2BhUwnJqCmUV60xgvJDFxauhdTfg4so+6Tqwh1xstJR3AS4tFAKRoH/+7CrQ2elN2/fh+X9x8e+d
j/ZfZZH0fxYTE5exTHE8iTUhWAfdpQahb+GrK85887xthQ9A4ccaxbK7SZLlaGNiUHBzo5sv1DoW
6s2iNrR8HM0vLU2QMm7J0wpMR229+Sj5Eo39izEE/+7lIl3OhNlFzhqm53tMxAFV7Cd480CKDus8
yiNy3mCid3bp3Ko8MWWjxQj11lH6BPLokb2KRAfHVd4nxe3pCUPyMUROeojnX/WKWG5H8TzhYo7J
FRiQvwYfq32Mkr6MhAy/BNH9ecLeq6amIZbD7b36WzAU//QqHQHyaRQV5cHEc/ioNNu2eoDFz3MU
JbxcyrazqMfBujGQaCfL4s7kwrONm68CEIGq81nfBIjXm5nfayiF+0nF69cFSY4DU++uIggPFRcc
TUoGZSrGTvtz6pUQcpnnuj7h0QjEYfrVSWczRG8h0cmt8OIig9/P8IWrDEgHCuiPf9M3Ks7kx8UY
rt2wnPRPk+QePhfLeHQypTN8NCwRjqZ6pm0OMQMbcwtIMCiqY5zN97zzHXWbh4bUNl5KwCErWnxW
RrgbQdg+Qlftg7olDvVRX0Pe1o9rLqbXl5PbzKVqEnnROU2Uh962f7ZlUGLVKy1LMNzhi5/MGAha
9J1WYDBGa8vE92dtuGs14lo0d4DaT4LGMeAMjfFzQ/EnuHNPXWiT7Nmr8IcncGWWxXAY8DYmHeVv
asQSEhq99Jkw6fvS5IfvrM7fgzpWhiW3X2cg9Poqj79uzOpmRwyc1Q1tE+HS1BmLohe4h9aTgp3f
QXe6dzm/td86NHAUBgEcEHOoE/i4/T3yJvk4LnKBLc+XMvZ+Re+GNrI6oQcZOSNrl4Td38J26QG2
R2r2Ec4KxtKYHthIstzySwodRR8q6IhmcheURg5c/zq+NXYXfouY8tRUQOf1irODHbgYDgP/AsKB
xrMk7kCWunpIsO2CkuWmlyRJATb974AsChAmRU0d3ZrFC+i8i5lL7CRsLG/zopvIeSn7i6pOzuI7
uB/HRm/5KVWdZWS7GhNIetWlntn+z6/aiQhg0AwC+OFWxMlSUOralhnrOAQtzO/qxaOXY79WCBgw
sHfuTHO9AxRrFME51+XIgMwG7b/Og8+oY+Cao5pv/3Pmr8sBbfafycZAUIc0yoxMp1E6KOVAeUki
hbL1S2BAaUVkcNDkMBTGKDyS9iys1wOiswykN5aDwYOQcxBObEA9VItLmiT8toT5sDb/xQoZnNER
r+cImyiB1FHDixBSMYmMwjTjbgG9EGIFaXDB1cenaUmdDLBHfvworUuNZwtNl+yEJ8sDRbb8TDlf
m4xBjjuAu89uUPC0KLLR/qi+0RnepUMlhEb2i4mN0Svi4ikFCYkx64N8PEqn9FNz0V7EriNrXZFf
v5rLBRtpOHxzDTAej2Yv1+OTcIH7Gt1M6ZQ4hnohuL+N7opoEgGr67mcBU+iM2vs25QA+/ozf9KR
Yl3DUvZeskmmL6hQe+JRTcDRG6ds/8C8FNhnWEqB+7JxcS9N1sXDS75bEKoaqeI+MCU5GeR/jsDw
d58pN/QYLK4ap+/T8cz6k2q+StsH1Zqzl+IzPuBxLTIDoZNSBvUuY1aAvNVzggKSzOEchCahKQ/Y
aWz45i9DYGeFG9Gshjxq0kustjGKCbgoZc2tW/9q8aaVUbajG1y7gtsogLUtQc4XB88CJ3h26iww
ICX+4vAYeaGvNpnhhBQhxp6m73kkO5Hc3uzHOiF/xAvH2AIiBfeIYnTI195RIqVJ9YjufYIpQ0AK
Z/zYFMxQM0t9Dq1p4gYA+HACeUVn5qxnj1K9HNoCICnYcG8aSCjafOFgt0UfaE6+5RDO2HnsYzZt
QhjFgpBmZaeTlYWIWxaE7Ga8naIc8ftDEfGb+06ZhotOLjX0ovJUJmP1pyrOpy/h3HE0A3VKxTc0
iRKwHtUF+ujurz/yHkXbw96+saGTCM2PIE8Rvxxuk/raHhC/ZaKJZ7ln0hldNI9YSwDTlX/+DjsR
p2S2arxWXeGVT2sX14zPjsmBy80zSvshbZM+NQh3fdUMMu3FdRo6VKzEJeFVKCOlnSDtDNlp3gbT
OA8iXiTxMQY6Pas+MGhuFO4BI3eIL8v6dJ0eOa5acKMU6D1Rib6q/ChywIplX6GuysRMa5WH6j6K
yNHViY8kQWmaQ4Fzlg2kfXHdzReibuA4p7Fg1KUcr9nt11JeVIHhbVTssSjY6Rcs4zxqchx7UTmC
jWM4l9yq7SfzhJxuNo448MBpztRjIRUPXLLS15b7jytnQj1wCA/sYBiKx+Vl6LrO6IYMpDJkm0Kg
Mx2h412QlCVAb18eoSN3+/pk/925LsIWtdmQFV/GipkiyzIWi/rK6zwFuEMbQRGrmIW/2v/HaIX4
iCMNMKAJAxoNrxKQGf8/L/fMS3wjyfNa1U1a7Lnn3L2XAQau4/e63BesCWaLacnhrGIJZScftR8H
1a1Ayt0uOb92UNisL61nJjVdIwasHsg/F4LPcwCEnEsEnb6t8DWp4bB74Cr4guhcTeiBmj7eOz6f
N00U62cO23XKMeZKQx/8/wZIVDSwNr9KnYzz1qrN/GuxAU3YZoGvf9WaPvX3EYYoNgzkuUKLqyRq
NQZKKlbRpUiP50Eysm1Ney3b4h9v8mxg/Uud8NhA24mo4iiMrpVYEok+xGQH1dk1tl7cOxeUlStN
tezAovMpQf1JnwIE02i+TM/WMkui2Waj74elBZfaAAua7d+ujZb7ujos8vluca7LQX2ECpfE38Xf
4PmjxHShbXa9LEoKEAd3JOzXXfo4094GQZwBSH0hSfRYcsLdkBzHt02wyT4KrHk0hjNQd5W7fvIG
c4w4hLzLVrNEWP4AjlsBTHnrm+B1LMrLVUNFX//d6aUbePN2338gZMCyzYOGgRWc3LqAer8WRaOx
tTPIDJB4Us4RPdOPACEc0t+fCNtACQfJ337LXaQW2Vu9z2Rt0qMVlhgtKz5AdHBxhYKFiFo/7Ybq
is4DlJehogWOqLKcdnoJFPseaavZzbGhBu0RJzCydxZCMsjHYrfDLx7uvWX/PfjJVG1R1UnJo4yv
7zCZTK9zJhqXUageAgts/FpOyYbGcCELk218wA4G8Ma9Mg29rhPcEKf82Cmg1d9Vr0cwMEBDTtwP
uTbluMzd9GFjVvb+TRZaNqRKqLm7nlk3CqMqAyYPgW35xWMFMxEo7C9lo3f2v65aze76wpL/XXM9
+wsNfW6okr2mvSpyxxp0uoYmwmAaTMMA7aWER+E67+EDvW3wy6iEsiQLSV9dsaLT754RsXGNIXcG
Il74/nFDkSk5e1vY/wSNiLpuvcRqd7FhqKuMJa6s30M+96usA1KuKiVXPNhjyJVIk1Kl3nOC/aST
F3uJbQ6wv8oeNuI2k2EEQm6BsInGogdWNrl7wngDKXJq2yIbG+HEVPicxlDnQxZN6URh5sI0wKZW
3rvIVWTwa5ow834tERQiMeNGrqld4lSOGBsrLxm4vJI/FhTtNKosz3QhbepH00MYp28jAePtGe0q
LUqNBMNCZ8lGjMyN207jUAl4bBNPpqczOlBH8GhvXbrl5zT6v0Qhp3Dr3SY6oW5GLvMxr5ks7jHe
srpDqm4Tr6npcBgZB9AdOHcBqHBE5peqEoUU4spvhmTloRsePgQ5t+SzGBjaB8E5vyTGAIN8V4Z+
5ELbGTFha6M58TwqV0f2PJCEda6vtu25fqi5tkz5i1qkGE3IE+Iu/6bFYMe+vrTkNpTz5Di0Bd0X
ER/Crgxh+bUApmdN+tRcT7yxbNT47e3VSm2tdShPEFWyDmaSi+vYXIVdUTyWxGlP0i4VnT4FOvSl
WKh/MEcPa58Zylp9KuaP4M/1AVoKgrvKuXiIZhHr6MG+8akyjWg8Y9S/k7ymOYMBP9cr8jxP8avR
3jxFlcvb3+JfJO8K0jSG6k6LIrUKv6I3bs77JpLAtxMDKp/Ym4Zg2xxwQnMjkZxAod6i8b6P92TJ
Lu4CDdTmahQEpcbnR/kQl84HmDR91wxclgvTIEpHibXZvNz851hV5+g1+s9BAjIPjBKe2IdSPOZJ
TMtcQ5gEwrX8fvU/vqQ6T+zl9SXAfbKrxC2Gh2lRiBmCZg5a+UXLsN56FArskhMa2OCUJh+P8Dzr
h4EDx+UkWFOIHiEA9gFR+tzWfOOyMVoCFRYgEdfZbGSlbfr4lSlisLHw6vc06sMA6UXaEWESNMP+
V4OxpUmFt5vMzvV8AEQXGl1ag2hEZN23KsXeTuzjgpPIjrlhrnkbinrG0USrf6s93LZV8hNG9wJB
GsS3hUibbI/6Jz5T+qCzcBWnWlnswZQYAveXiY6LBs7NkITI+rmmfsV1YpGMZQ6adMFm9w2hdPJw
hMvJA7qKrfQENYzEFzaOzuLMmn7i5Du66xFZG2zoRaUfJLHwDpgEMIwlY70rRmNFtNmZjfmX/Se9
9rT8zoct/+yTSFYWpy2RyKN3B/GWqeB1WLwJth3DxY+fgvID0fT5uTwq5YXlKgym6Y2mCFi38DLJ
MsPxR11fu+KFNZuAB2VdWMWuwitB2tv25y+1WL+Ua2RQ5K2k5jJ/BpXcb1G49ZT+jhjYnHlQWoYM
2NxVXmbGcsk6w8k1YXxlldOi8bKCSJlCh5Ck+oTSU+A+ol3+LdMRVTT/48Z0qllIk9UlBB8gQxB9
riSXMzmy5Oa85kSgwt5y6FH1i18MFxCbQVyYFArdUo3eifzf41jl+Ujva5n3X/YxbNryln0FP9YC
Os56LNey9L44bf7DwVzYaBT/Op820x9iTHeT1lgja3pdZqUQLkPrBTWnLvlF6Nzzu94KUqAgtp5G
pFPI1HOFS+rU5MjeRfLDf+EaGyWAWN9+75Lm4+/7ut0Q+N2gLDAWXZYWXl0MU183wxGCfuqAzquh
wHGZKP0dqN4T/RfgpwZkxo/kDLbufvo1F5wai6FG2ncBf3/RfDQZAlRJYdit51yxC4iXTU8Wy36x
UiCES1JCDAOFMHJ/P7BO77DdiGmyKGMaQ9Jwn/E0gpqzeJANhrLj/rqIYFUrA71NYOo1AZ8kamM2
Ga/s0yqM4jfWdgRBe0AjkPe04rkLjo9COdWeATp9l0Wu1kvZh9IfBhxykRa1VtWFguM9JcSgxyI9
uj8jkGsf/Ei88nlF2rTStTVdgYX3xBc4UGZ/at0OvdlffFk+P6PQtxaBPqSHSyNwwsD/pxf+TfUQ
5N646fsDu/ZV/siTMabD+t8gCLARhsXvz3BE+lSnnj21bSZm69lwXQIVM0JuscQFcgT/jaoDxRg0
EWd+rzWlhsFwNw3gWjnMPvaow3B+MObv8aS12zeAxVNOC2awwz5r2PhFoHpOB2iOK3Ore6mfTiM5
3SnHrXpguFK5ZeAB76CctYXU8U+ZS/7bI0Qwd5Tz+t6+b/+9UrGlQ3Rnr/ooj92t52jErh/ebhcc
aB6F7T+L1stG2jEPsGk2Jf2haiqaBtJGVBoXJffrYlUIsM+neYmUNLgbOyCma8NUSZs6D5VDGyFz
ndKuQFK5ycIcjcPnS7A0BGKzuwaqzSVrJvWZLCU1e63uaTfkDTfTM58bJg6f2ssFMN4BeMu9qJTF
GHpNAX3Kil7nBuoGD1e8vcL0SJ674CSim5GDgDrQ3Idsyx/Qf0CxEihY5ozYOCPtx3s7rF5qnnVs
SLD6+2YkxFD/Anw3OJ3z1/Z9egRQOArqKgisnfXsEpn5wIJ/3YF/wVAoa3QsPvloVrcnKbocZiZS
152heNn80EMHW5oq22zn0pyFCV77qnKDf0PWKyKPrT6weVAe0oVpJ1YvL4qojqU47D9M04rIO2yL
ajBOpfXXBdjtiirR+niMpSvMtQWJEwp3cqcCZq8JkUO6drH+S3HwlO1/fgdwQc/MTs1uY3/0TQDG
tbdwrxO1izzfuBFwkWfgr/7kpKj2KnudqifadvndEi9GN16EsGBL2b5eeLugnUgIZBghM0uZRGPw
MFYNHGArEwbVCWa9ieUqu9WNad4tlCj6yQCPkWDF6OWUyv4oxurv2UN1rTnCHYgs5/e9krHTUNAR
Ty0mcXgRHXlZ5pf9fZ10dh+x6ElKsBgSASU9+AkDCV6M9SEO09jgZtpGgZpVnmTsdjwJP7Bih00C
Yp8n8AGefS99u24sH0yof246x5jME3G7R3bBchlwZorPBxtpwkdqWOV+lgD94ROTw/H8FQkczN6P
f3uCEsBIoEN+j1j9OCLWFUHqbJJdVA8UEOXjvt5tEdJLg6fCl9RoEAxucGjmJnsoQhKtfx+Zv0Jc
aJ35780qhUmTk0GnqwiUV4MjlMfuOd0vowrmwY9i7YtjHSoddgjwClyH+A5TPAIh2k3IaJmGoz0c
mCDnyQfaBrPejJza6BA9KsKJjk+66lhqmKWgf58d185S8bMSrpAueUMUeOZxINuQeBP685ZyK1qq
cFUaSqdgl9uoQ7lhTNKXiG27J+swSmjtge8aDi/q/nh6f5ZBdfJEGZFuDW3UFVT2eOn6WNqjiuQB
RknYC3W0fjs8IZD9ojVjLHU/MvN5C7NY7jpZtQxDJf4X+XNk4F6+g7/+eEgT7296mWBZSUAQZY0Z
4EUmj9s9TsJ61N7VLjsr7QCJUga4Y9odqxCnUS94gugRNd6j7Z5UiOuD57yQCnKw+DXNwfI47D9b
WUkpRX+IDr84uWNO1IDYLGICHLV/3OZ1uiI1efLekDbtPDf4XLQg2OXFSlMWodO7uy7fSGe4FvFM
/fCDf1xYyTMZFXgHfxxQJOvTYsS/sxnd7O9fp2FIw7eiBk7UjwmbofuFaOb48sZX2T0F4MlIDiim
ks6F2ytyY84TrbvCmoXMYKhqHIjETu4K33lfYY26CF0fsfy4zSQqn0P+P4h+YJqEoFKxVilw97k3
g2Nl7WHj+UV+BNP93MOAGYDslnpUvdKyk1rmQl+8mizkcbt6cky7/XjkbVUHVhc75t6m9ErtFgQH
YhqKQjh+qBPeLDGpxsXpJPFYIE3cXxGI7vEI8a7YvA1H7dmEhG/RCU+LJE1IwbI+GE/lB6QkjSMK
7p9PWq4/eWn04ujT3sWMi+fBlh8ZBjH/ptic/SHtlb69LhPcDKH4IiQNZ/Zzp6pqgVhga8p/s4MZ
Z77nVsC8PHOmteoWj/It3dYYyIxFZUx3rDBGf6HEfs1EcZzlf6d+Z7sisg0y+fz18I4iAoa5ZQ2F
iJLKIXNQzYOjF23WfBWmDj4zWerEg01GemWuYu75DqKtLwkGbUw2wnLCPZ48LNg9SccS59xU5Gm0
kWucgNMWkpjG7Vrfs9yBJ8dKyE+6qEEc0E39UYAFxdl6AaMIe0pcaupmDxDIXnVD232bRw9RCk2S
AHAubParoZlW59feZ1ybZDIW2VPqKDN8jX6DLydV8tR10as3q/cXc29WCSf8yEpWEvkvMKsJXU7r
8QzLHFZEUThcl3he7fewPWf+RykE4qkpljoNVwFy4MacDPDCGN3edBftL+bwLktJWRDF7fR7CK0F
endMwS6DHQsHw82ccRoTjPe7/+EjV1f63S+w+jIOSbIQ567t2VIKtUwu+vGwbF99cxNjPvZtXq2/
DX3OXBDSgBDJ6LTXJcu5x7HhzXXZe17PJnauxfypxbPQb2iVZHLY/Y4JlhDd1Gyrl2x78cpwmUuQ
sZTprRaYv+/Vbkm9cmoT72bnx+DTUcGwwCZFP5aImkUMiQP7R/7/oGhGSW5cPSZTSLhps5MYEH0N
UlOxSAbUtGQ19jIrJEqmHN3WYilZH/G+JAPPqW67o2dGBDcgfhjnyXNgMyrTpjTZEwqEWXo2iqS2
NifAWR1D5SwndeNiNyuwcK7yln+kpUidlmfzsypMyiRg0+3wdornDRgswrWKStx1DMhUMX09L0bL
GRDrl3YJsnx1HVG2WKA4y0xDWSax7lQCxmDKqX6mnqKi/6xHOaKDBQgJP15JA1QTV8r+Wp08N1Cv
xU/KgNRlFstNsrz+OwyvrGyaVMp3U+GuimWryhwJS00pc24mdxRwnuMtfZqXbHdsl8xXY5L4pabM
VPtmXnxlJT5696o3NWPfV/Ly/Q3+jj0NLE+btB7KK60H97LPh4TSTwPTdiXxOmbAkV5CQtMOo3Hh
piAcinS70qu7HJ1ig+fmzKofohvev1nQGaeIbLMRew3ChrurkaCEyVXFpJzHSE9wy6K5+KwUKPt+
h3fY8NBeo03jdJFASFTVpEgyInQfJJYTldsu2/VvElk0QD8UfsHzbHTF1I06d+VHLowvcu4Ir0Hr
V+yXolcgHaSnVbdJ/UZb7tBMg0b5ujAdSaxPemPkwrDgVQNZ7yDIRZdrFauCoxSr/g1jyObBAWXk
Lb/NpvEAzR7tP7NzQRdczJEjkkiHbOw9lWEzkrRmu/2mf6mohCbUB4sGm5muPJxMfLb7SanlCT2o
om6QozzMDxA6bHfS8vUWh/NyW9Q/2JuCKAKhXMVQjxmHeaq3eCkjFAuo+bv2XTJhlluNGrj9LdWo
R9lBBX0eKOwPyYCeAN5nVhN8+QNkx6Cqr550m0LUz2ca1zcnA0VeBfxPOqq1FuqHb9vjERrYH+Ea
JaDeJoF1VCh1D9Jutelj0YJYm6GYkXERSSaGCzxiSO1wjMEsDw6U+juoTITYQn1c0hEc659Whgwv
5xzZT/5FplgaOc8KZ/BQ13dzZ4ojW5W1erXaJ6ib1vFviWimJ8SOwyWXkuXC3gY3C6VCHqCc5OIk
huFVCCu5YTAB1B8+NsW36zv3aGqLYSs27Ag3mD15Fm72AEaHTTScjUoQnmp9m4Fmj8M6TrBgLOMX
UWml67smJAz9bqvr5pk9gCIOWyEp82q+Je1eOsasW47t/rt1eAVChIqBsCRMLFahTKQsfxlR4Q+3
uj/sxEhpbwZIYFHp4MYntWTPncKOKg4VibDwCyOfG9tnv22ifEXXCXnf7LyZ0m4hutJczn5kr5Tw
7DOvL33xDjepfRIrUf3UHmBTr+ZlqZXuRZaFdC2Z2ui4OjYW/p7TqZ4uTQrZjXMBxKVBWLSpA5dJ
ToSTBjB5OgKZrTZEivVcLMl71uMBAehRVJxznkuErQxjK/RqmLxMUfqNDudGOubM95EMqmtaXSd5
WPb7JLqdIO013nFJ+ePv6b6hK+ZV+VMJcBQ9j7/lRiVsHW0zslv1P+L+99Po5H+FdGjFStmSFY0r
7Hjk8cq0FC10swsFCDae4LgY67pscY4tROrNRN25l9RMD74arULi4Rwv20xCoHNCbgLsyAhLOJUb
VaZ1TGXrLCQgvsEZIvDoP/wKoGKgwETomYs/Wch+LLM4P7ZX8dFcEtuDXfVgkgPLhakwv/c49a3R
8Dh0VtPznJNbJpjjyGy1+4iMEXGQLO/E88A+mlFZNSo1yTenHcloGz+ZotvKPoGDddqr0XwgAR98
xgv2IraCkmynakEv3L3n5f7JYCEi+u3NuuLBtgyk7q+QobnjQSFDOOcWKrHvz2EzI2PI5uOF68w9
/Py6cZNxaBOXbnc4lv0SJP8X33NasOxcNfVQmyQFmylJ2JurUW8JXXmhkS+IxiIwWdEplfi1s6/Q
0IE3aSIDkeQk1HxT/F+pDAHp/tVnW5+sQqyBiE13DFgTTi4f/2wymtS9Qoezedqn+cVRXTtyYRQV
yXGfxOyxjIOxc5UlZoVaM6uaF8vD0+XIC/qSbvAgJhkqTkLmXo45RoMHxU4ONeqtTjfzbLvn/Wao
8RLn0PDcWaofHii7bF0dQeV/LiIdsFeh9SpdXwAGIbO/eBWtP7JH0fdxLAzcO80n2Osn6SzkytaZ
INgx6plyXRggKic/yMi86Wsid0oYJJszst3JYiHdLWbpGh9RU/bV7blRv74BcmNlFbFVK4SFY+V5
rapZ0Fkl7X2wktT1q9FUlR3JKU82xesyUrcx0mZHNJROZlAkRK8EYEAuorl/pimxnCp3iFRsIt+2
jQ/pjbAPIefKcry1oPYwod6XXKKn4gkrEwJ2nEC2BDvHnuD6HlOy/by4sKCAesWJBdXgLtj4jdDT
WB53qbYSsqh1GECE7tO445jmsUpQ1Mko8Q4WXdNnutOXIgmcrPcJSmTTzqFkarU3hfzBQ+t66hMb
a8RV6PNYd0bASuAKvWZ/jtQEzUyoKAlQFmnr8ah3lBwWoP3d9Whjj3XRTtBLy6XHcKWoRYkgLN0d
AUuRxeIjEf8rapGISsrPh7f3dvpHNEP3Qy9XcGxYvfUWo6fcehE8yHCs0N/jlhasr/FIXTzcA1qE
aHfAPS1fTzrRj+B/IJQ5wB6l0X0R7Dl8jKRr4ghIxtSais3Qk4oHdcBee04kX/MbeLW75i+OnT4Q
yh2WKMypPZj56XtsshPA/H8PrKlIllNBQPE8LEWoSAgS1NamKHjnVXtqU4YebjoCK8OvMraVh6Ok
BwDuVduXypyE2C21bUGXHoftndOpFthE6yWQ9CRmh2unt+HUR0YxbRYm54aFoBAe+cuWcEXqhemu
dTZGXvPgKz+I9kaMy24rXcqkNl3bl9wJR2JYtlVZH2JC2q0tKr/uX0a8WX477DMVHSoZYYmwbcb9
M+5/vqKbCLaomzB/Q4p70EE4OgOANiAQUK0mHdLJUFC2x/hl9O1bR3c9rFhALNa2xGeltvM2Oo4q
JgPnyn2qKLgdfm0t3NXUYsxeImCjA1qel0huxuOSu/ZbRj5jVI68qFgGfFmO3Pgy8BWKXCom1DZt
L+I7jKcsJya9Ax3afC7OtERUQW1lUQSwsxvNEpH9zPTTw8lQtVLKFlVv0aQb04xXS/N7CcxM98dS
7U2bAnsQeWDpy1K4xhLeh5r/s5pBAmega+e8x5gnjnicCxfDx0g0D/Ow4Sh2GSj+ja+oYppow0s9
PNuSsCHZDOYaxV/yTMhCEA11pOUTvDd10Pu5VkX1hMPwhlnGr53jIaro+GT0+vCSRVZWiQdXemsI
mAzoYaOIxtnjI863Bf7uvWh+4zVP5WLTnw6Q5DuAe92+84fKcIFeyMM4bF34h6NgOQq1YDe8j6t8
LOhaWsSOb98w3c+socKqzErYKVQ1wLa7DYW9Hm/nP/IUpOGbDGeFJsx6bgZF7vIukc1AfOxaF5xS
WZjiau2l4E81e205p/eWG6meJ0gBcfVQ2f/z5Tr3xaIB1IY/c7zcrRlHQkA8R8yDNiVvajWpjjVf
hK59f7koHCs88lNuuMJlh2+MOaPZjQAj5cVgRoizhM/LAwKBRUsUiWkd2Pp9Q0lim2olu+3bvA4T
ncuUbYxzuHoA9d4ZjhLNHj95tyJ3VZGili5DV8S5VJiYq7fy3slOeqd2LSC9Vdj+X9+ZVqMgSCKS
FtUbDIGSa+F8fpADFayhLWfl87nwG5+QJLyc43fvhP5anahVWMwX+pNRTiXShIbZmoMRGalSEC1T
CodwR84eRer6I/qEMMyQ2J2uM17GYvNzf4AIbAoFiJbKzrQTb6qEWFUXHnShxtwZWzPk3G9JnsmX
WeaigKxdKdbj59neefpHrjqVZ1S3TVFz+xYiLrx7JaWY7n7ZV5z+a03b4ZN7WfzLbcgnQbbrcCnB
yFTGwduUe/02dZG8nnaakfOftCQWcMoKMypPZpzC8W4M1By0Ov6I9tjN76744pGygoT7rsoWEXoe
2eMu6FQg2CiayLvbBeztHMFVIv1tDbAvHMuchquBFq6PaBFwwe2d/5fjRcK6V+daKA7ccmhAjBVy
REePQ2VYxDcvaVVbZO3qf+LVcpxmu7RMb/YbS2rW8i22gVRearwmZ3ko6TT2fAxUlcHIFXV+mZ/z
giAsZVP8J4odleerZKOJKy48QpkD58nYzM82Ep4RoFTe+w/X8ekYqqIJbKQ4pAWxhUsC2DshTtkE
9lN8HSsOlAqfDWSKc/BsaJ/XuLKAN9wGCbgsShPUfqoc1OxrULhfSTMyRHJBF7Gft/xXbjbyEooE
D5NdO3amuOn45Sx7TDy+dyX9mPzPFxQvN9Lpn5g04y7fmagzVPYV+upVk9AZdOt6vHT5c6Cgl/uC
sp3m2MwAXMYZVnwT9YH+54xg3Xc6oinckWTwHX5xLBIkBgshXcydMtR1xbOEgGJKSuO8OLIJtOn7
26JwSgVbjyg4bLAh9jgRtX9XlYaFGHza8Xsf4pm0PAK35JjDahYjWfuhdy//Zze6OSRkNUV9lISf
XXvU+O/4TRIzpcjESSTGSD3aNQ2rDC9UUwRbVXlrRFuA2DoXlFe+gHlRtchSebwv2HFy/CFN29pc
GmeOcE5ShqIoAV6ai7XgDZLtAYwFA/DeAd1GzYDuiSXqVsXGHZVDPSVKCgIVPgb8KuHqgO4oWeJZ
UeMjhTjzU6fDwzqgEgsUsSgoNnMoVGr5E8eEJJ1FC/aeSZDJ7lrZJ2+Eoh0NTbwJr+DIGqVmH4CY
EqrQKnKKqXM849XxA9/0Q/qc2ff3hTlfe2Xgy05WPyfpJzYTJgpk2/OJtYaRNycbSM7EZRTbPkKe
ZHsnuFbJ9IV3vMzrRpLZwIbi3pxVEiPbIppPdpCIAKR8OE1+VW2+mziNv69DmwulZtn4q8kkA0r6
gU4zaobz0BpYS9Mqi4uyjCTgD2LdDMK6XBIYM1flSi8AL2LQJf/WEKKQmmwLjcv0rVN13h/K9g==
`protect end_protected
