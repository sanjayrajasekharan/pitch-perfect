-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rVwsMz9X/oTM5XWE2iac6S0UBAttBE4maG97DClK2RabG6OaP8SOsrqX5Z9Re5fxbtP9ubMObjrh
MXuZtYF8uPRs4WnZiyaA3z9tNI1r5jCOKI9tgWjqJn7ksmiCx4Imy5XHSICijO+vQQAm9y73YD0H
1UPbcpyQ3gB8hLGSM5J/oq2gGyP97vQBwi4CveWNDKb/uHrbFXyAJvHfhe+vOM3Rj4DT3AzeoovS
yjyeX/vcPXWHDeCoiI6eWqQnon+ULCbBGkYRtaKCD0wBZu/AwgfpLP4ucNxyz8IXY1FRa+rrsg1n
qtQIB/FHwi9QelfokBnmhx8ud/jFvZiktSezQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
9R5xOL0h2diQ3A0FKTC49AoukGoMi7e6fHH0Cd6gqOJR3jFMYX/ybH4pFJamFWE1f821dv1hQEIg
JSOE6vDebPzjCYQsLCeQb6QhBKHeSMkTzqauNHVghOMQ02lf/vtIgGi8ylNpVOWgMaepJjrSUCIV
YzQmGHp4UH2z6yd4769+jz8aYygVvOIERancpetBe3BsbUGqgd1VV3VUGOzCzGet9/ncCAZDYpWn
op4y+S1AplRJffXgF8NzX2meBobyreDPs69i1FKT5jPUa2I+f7O2VJX5tH2imLNkkDTTxbbEQuEr
o4HibyOHJTStlUIN8MgpzIjdlDZlijPfOk5AyPus3++19ZSzt2YdP2PySFzmcdJGZPe8BuYmC7We
8ZXtq4HN3vgYAS5ctx3VAELCg/eyQRQoej9lBsQ165NdUJiiYoOzSAbL49iDdpZVcJ8udJntucQv
j1rDItk7N+il66tVFFpq63mvJlaoxPrPCovlZWUnZFGN90OuUtjZ0KEMgBgTQW3zv0Wqs46iV7tP
T/KTBSbs5V/ENJnwt5tsBil06Y+YGoYykmRDK9t0/PupxXdyyCn9NXh8pjkntDOdteI/X/kfRwIQ
jIb08QhmhlJv1M4dOHddD4onsqPJUcsL5sZM3CXlSAW/pNMXREKnbeyZ0e/jhDc4qlz+EjPQmRjN
wGeaoEqZAFWIRwcNMeEbRVcNniXenbwJyVupQ2QtaLjzeCsGp/p++70Hy1WodRA2B8oOdKhU33SS
zGIhfZS9HHZQIhAiMblbFVQ7wJE0FkGgQy4xqAIPp5qDEHQ59HS6I5BkjQ9dMIWTCNjSFYcfa7sj
RmCUOP4mxUZX9+eVn2HOveAtZt95mLnNp6Lysz4PMUbVKuCik1GKgbjGNfd8ZwlKdHLKGcFFgK78
27blYtyN4cTpuslDaXbVBPiQrzKuc4clHUtWN8zKf3u81XWpBDxVLm+trLkPZTS00kMZUZI8nf5R
lByVjGyZ0n4pTTkwdtQHN2jxa4lOqa574m+Oa+PrikXiSS3F4xjst5DwwgFhwLr+GrPHe0UU5WgZ
qMVSq90nN39M80oOxJSgrUMEh6oHcOPXUoSlRJm+BDitMlBE7m5yakczvBlMcCa+CR7sZ+vdBhbn
WLUy5Nr0XNqBSX1+SHdVhjBAlGImbpfv2V9hsB3Qxj9JsEK2qqaz2eoAllqRHn51W+kykTy4904C
jVYUwuhbCct4YmYR4ycZgccKbget94oBZl65arSz5wjucYmDmCycKaa4v3jLXqArvrRMaeYhEc9T
Y/+B3B1HY7okAFqSpfpipG6fmq5HeLJpovqNoWXD5MYsfAf4NfmNYj9dfjy6Ng1Y6QMqJE9TM3B5
zOGmzRJTDkfuG8zVM933Hg3IeCc7X9LsVPYq56YIa5SoIwn9CECnqKFzsK2U2s4VeeaZMfy3hh8P
Aoe+heEL/frzSIZ2E0WBXUYzXryuZbKK5Idd6+wNbGzPOWCJSwEUfKPtA89LiUyevq4lBk7Aj+Wa
QnXQ2c9TJ3CEVqzysg8w2yNHo7O0gGdDNfZ0WBcc+OJKalcHQ9jzrh3XeEt70f2ZoTZz3yzOsPu3
2LBEOTEr5k6CLFan8TcSt7dqhpZqghmcth1SgSszX+FVjfeOtffh5VjvcbEfgY7Z2ZyFuGizOMRH
Jfwg/XFMvEvdBjxVmHfjmJdJ/HYjKE2vU5u4cjRdyPRmG3bXxSoPlycqo9qFVV8tFGpoQ4Ghv7OX
dONm1WZy1czD+Ox6hYWmCqO0cGFZFA7U/Vfz6wDsbWIY4GAm8UvzAD30S3JPRIKdqYDepanmXxdm
Hh+UoYzfaL80SXVBTXIfFDkBN14slhL2Bix84pNuG7ABunDq4YAejJi/YZw5+h/PdX0b8fxDsqyZ
PIHQL5lorzMdySE+k6ll6ArsPkjfYOj54d2ZnH44Wh5a7rmHsdra8GbD2rOaX5axFoMzt1uZ5d5T
kItnwFU+aqpBpysIEi74Rdryb5EJwyP0KSwNBF7Crys6Z8byokTj+c7DqQgerFzJfAO4/3IWBUCt
Bn8mkJHtpzfJzI01G/N3Uy4OBKuk5g/+XE035NUFd4iPJyAVGCajvM04v7e9q08JfGUXz+N8Toxg
kU0ykcQ4x+RhEovK9RgIjz9mRvjBImi90zKZ/+doDrBN+dj/+1ok2IshaoPRIDClePqPtr4hV2Uo
TLtHIYNDZD4tr9P2StGLdktKhCNHObIBLazUPccnLKisCvFVcQEm8T+K5fPDMosaPQziL1+/z5u1
0ysKnAtBTM1aLBfMq1BnkNxXvCDBTzfBY9oK9zCleCNejoN0RVMPu2LWY/s1VUhv0/NkcJ6yVHzx
44rmH5GTwfQmjgsB2r/cD9ZmsVVh4/O8j4zmbbqx8F6hMlsS5wqzkOPQQKHpJWiGdcnjY5UA5hOq
7vfPzq6995JqcBKJ5ryKHtvZVujnOGdSNWYotoqyQSARuQDytOCuQyvHg1EUefXR+n4NZQYEREdJ
wbA5+W3ZVNtiTgcrg5pOzXxevBr8YFZ3v0ih9ii5OkySLz7VJlJrEK0FzZfwlg3Z4eodH4bkExB4
mP762VFeWeA5+kZdjxhuLo/4d7zCWHNbe7m+dyfbXY6QJfzc0r+wUI5CsiU88REeOAbh8Hm/Xe5j
AyYbL8TTWrin/9bS0+H05AK0hV8HJtTK0FUqX16e/khFaq28wWY8G+R2Sj+NxEcqPoJYo8VDy38N
sT3VU+zyDUEkPgFetcx+JhgKyJK5MTK/mVwVb3dWUleQNEEBX8jLbomF+C1DEx53VoQEcYQ1rX9p
1Da2p/sE5WDwKVVUZ+KB9l3CP0uc8xVY+1manJ4yfDZdQOtx4MCdan59r7Ug+9iI5oYgxP3vCMOb
aMGj5WX14UyY9CXE58GcROHpLS0vswd942XwUNyWR4vLi9JrVE7T7c5EmaITPkatFW4I3G0NVEgN
By2NokbsBDb7VPGKMRXq3duhbODLBQevuhLIMj8QOXF2mNaGcBbbP61LQjXFNC8smkI3LdSQepqc
Yca1srAAJ5+jKEt1NbEGWp9/BW7tSUtWB8Wy0V7TD3u13baDLaFFvk/8iQnWv8rn2RYFdY/le6fJ
ZxIwIwoPgzSYpV2agcHN+w1MdL4mZDDu7vjR4AzwBT/YO++nrcd6ZUuJ//75mYjUulRg8EKDr01i
weL4pnlE9Ykgzj/a7X4WLB0zqC01JJKDJ6seqPrGATs8QbeRlsCw11nGBPVZKw+lpJ6yvN3DtCdC
uFJM1mvaw4UQj6MytZdl2x1Ca42ZBme6pGkPNo11X5qHYlzrYcoc73NTQuv/MCjIvQlekfeAEN2v
OTmYT7vHsAfDF3VQAIj+n8Q7BpVA5h3TdagL2Gn0FYUzlcaP5OUz1MwyB3+M7+R/KDDfP5A/gJWd
Vgb6wFDqkkvkF4txJY+DFFauuaSMEU9UznXiZqXLEy6LqUjjZlhOuytWcCiLHyu1Ioe0rT2QqWD3
BKhww2VbzW6I820CuIStY4I2D3tnio4eL+k3Lq1ouCMtq6mwXCdjFrm0H1r9ht6vEKz7r29B3FeQ
GVcjF0/xlANFnndHRqVl6GAyEniIsovno/RTdL+bctSsUd29JMzfccCeES+ZJmjsCkUMxm5nkP/c
3ox91KdYojVXWflXsoBBHW9eTRObHTFGejxM5ti77DClaKruBlMW+Eq0uxxTFrmkbRe/Ngw0R13H
21NM6M3HEXO+7f9R1hNIG6+jPhK0HtWIOHzfQ+8ngt1Ci9bF3lbCRfcvzX+GSnqReuyxpN/Cag6F
g3UR0RDchc+lvn5/b1MFBbVC5kq8myHZrdlNtchTFsm6sEt8QYvuG9IKV51eeYKR0cJmYnshzzrT
ViwnYJHiXq7LMYCSnrpo7woWvB01Jmr740yt5OOQhv+SLQGiGbqKKK9ytlMi5jSfx8wvVIf0kLGj
T0t1LH+weBrdvRWbQy3BrjpAmFnTxMGq3Z/p7fBq1nJ5N87fS7Nz1oAMrdj6PDTqLdVpjVzu5D1y
sF9Uo9dMp2wBdeHCAIArWYkhnNBVv6cqEFgF1izUxTki1XjhyIDIhoztaK5TYzfQI353BCZmaC0/
A8LgUEJHPNEMg8KPYtUrO8NWyJtoAd6nbcKJx48zny/gDgKLQLODMO21rLKQqJnqG5Xt1rLENsKc
qIJOuXftLlqgrJUqcIFYKrB3OGEVWQvCORp6qmuCDx91oYT+vPm2d+1adD0hkJOeiGhH+sTneDU0
KziUvgAm+xQLti+anUejvkLyTFr8kr3rZFdOYqVoBsi8B9gjFYjlRBE6Q8hUE1DJSnIP2QnVG54G
jhsyk9YGobLztGfvixNpWfSLOIWdOCsF1d0Iet0DFFTOwo3FUIx/WcGuYMcN8/rz7Lq3a/hDg22W
h/h/tAUuuj7IZOTYXY9gf7yWk6JeQm5LaIuO109Kpq4f8nONcsQcJJtdumVV4ESZXIaJbBHpUD2Q
ZiBH9BVntVlSOfw6oorGzB6z4XoZohamVtqqGuy+Rac1Khl7jAp4293+pm+ayADXBpG/jAxkQ/Ko
PFjhnzSLI5j7pZgMjfT3h/Qa0OJZv5WvFidXu4MKsJuGQx5YwsMRRAk37Bb7udxtVl6TfGl8k2yK
gHIcbiVVUcOSSwhREXT+xhnD04efCHPRQXxxAMUh38Z5ETotVeXJgXsa7bptG3TweoV8CGcYoGtM
tvo22OI97Isr9vrnKDLxc/W3be6o7Z+3B1iLtPP+lofQL/XKRQbFd4x43fFiaUULQ6UzUJWgG9uK
hCZb5GDFnr0iaMeewwMGbKv/xAk+v46o8DHHb6S6fYgtPvymhw6UBw68e7TW6HkCCkfPM9hQvr0u
75Kohma4bCdUfjBU+vBHCOuUAgkbz9+8VepLe3cSIMQGcEhHOXGyG5EG/n/UUv2xJQeX7gH32I7R
UWzPcALn9VdySXQoyRPqjNLSa8aLpnx2rBdHLYMgofNkU3NO6nPNVSWDnUPT/L6wASgpU+dgg+tT
Iw2i6+sQZEWn2ozjQAn2aHKLUP4oG6mBuxFQRGrxl6j6LZLk5RVPoEIHT9QScAjV6blfLO+sO2wD
LzpTXNWB6/TjELvLcWLhizytNk2c70kgW+gPYf+awTylwsnSwGp/68OMBFjpdI1oro/KksBn/5Ab
PEXBVi/QAZCtzBf9DWMBRdnzb/pQh7FHayayhAAlxCDO7lcQTlBHGr/0sMPlBC4+Bl1dz1pXxNEg
3GCJYp8QDNCK/geoXSKbjiD7b9xGbN41z7wM6ZMSHkjEIfjHYQQC44zCJyEwKCqSTvkqcpNodelI
rhDvuFYPXnbTZhWRvky7U38O0pqd4ODfm7wmxlyt/S1MyImoqHByD8k6pjkEgl6VF67oKh5owGOs
c1cYuRnTcThEG4+X5IOjGGMAlS2NfdNtLEgx6rfg0E01txV0XzuWdXy9ii/QXKma1stf3o79DuMp
YW5rHx8/e69kDebKcbLu6hIl7uMty8d+Yk3mnEBGG5eC8+uFhNOxamqVnYdUmH6LeZtVIzabC+xy
R+23ss7yo2fO12NS2WRwaRUvf7XNWytRrWYNv2iWhTgecUmWYm4/ShmwbckiQ6xjkL+v/wDu7poq
Y7FPP2AOdwTt4NN6Lodv3MzvKi32QkH3uGd0naUTfhsZ2gwkzFUl9FMD+jmRW7BSJE2nFK3jCZYh
ynGFSlGDklg7FLE82bDhQHqhgDb4W14OLNsbClhNgnFwpVmadKG3r1t7OTplgCjv237HonN0bJrW
XjGFrxcgRhCXIavqfN9bjjrZgfmtmwBEyLkgAz+N4zSx2Z78SNUQBJfjUVGbh+7umnwWgnBxwz+/
Yzc8zIu8zHDnpYRzAUi/u/5pha6yctwGQsLY+tKVBxCsoyXMo3RL6YbhDTxXLeIKIgKBdtgNIWH0
adayDbQjmUCkZPvyOnCAN7jna9DUrBXSO8XSRJ/F/gjGzBGdKTaY7TyU2A7s20Lye+ZPxWlmRzk/
Kg0JVKZ7YTaMI6Lu/b55b2gMOnyiUL3glv2roteYGRGAwikfM3d/lPTnNUlwx//EzT77XjqOpskq
m//0xNgL0iBNX5W+C6U034wuq6IBDeFIlNhJujT52GYaw1cLCvggj+o6Jhb/ewUgugaQvHRETBvi
CbdtOhXPBMJtu8mwrtN/BtyvZTx/rgV/7I5IKWzeOtuBlK7eBAUG4NoqjYVLDhYlVIa1iRH0EXMU
X5YEdmSthA5kUqAgaWwdzPqn7rDcI+hyYC3afGR3WJBjJrHhyykxyOz04FD0ysHEv6YKNQeVX35z
8Z3vgnXY7IdtPPjbwqQcFWjK3F1ywwpcgAh2P+ymfkdX0DTg37u0qQjSg7j81L0Aj4HVzTNHQTeE
c6/Rw/tS5l7umRfTMc95Lli6fFQAU1V5UK530RoYXoKPr4lgF5+9so5K1Z92FHwmyd7ZJPZocNmJ
6WXbmoduaRwxLPuyQKEWGfW2qbyOzuW2LdqjWGpqOWFNhMNaBB/vi//uFFNpPbAdoIJ42oAwBlAA
AF96644znohXIHfeu31SMC2zCviHb18HJHlFUMt7JGn3G/v8yrJ/TSMNYsuy+hyjMcBGe3/X7TYs
qzL8XxAlnyM3JLptfeIXxMauGlG+/n7OQIbnpsTSQZdZ7PgKlv4r9hMyQPJTiOfVFNFfVmVnblxm
YLecfva34UFyBMeVvAF5iG7o1yeBbAdtWTmlyOE0ns8Z+FNfhrugKVT+eZGVhwaBQ6vUwHYcWv61
n3ge8iKPjWv+IJ9TPq2pVqOA2FrCTutBj9NjdMK1VBt1iWrk3SDZJYJkQBDTD1Z9ApJwEaPB/0J3
I19mBFvQpb2GUS+QhK5SnLhZv+kiSuT6JN87ciqjpsg9JaQpaZdY4KQBiJRLWSGgJlfvUH3iVef0
5D+VUM+wqbi6ymqx3gcDBOBIHtYPH5+B4wawDrIvhrU5oJGnOO66FCr4Em7mx1VqY8qYjlS1KWaQ
EIgHWVeVnvJ1forTXm+pBsJOZz4LGHtDSkib46lGtQVlSlVe5hfYAYGM6qYpsmY/3BXwx4qVVLNZ
lPpvvlBuRkR8XC6qvdcsyPC3tXmyFEn2x6YBjTp2+6UWXJfionG+bHIxUApHoGNxaWsKmRLh9FOu
OyfXVxSTHeYC9DOXlmFK4o9bmYHOYIn9yRejVK9JitAcPznc7oMIKfoRhAQUIyeN29iEvsha9zDy
vV9CurdzWh3FfNxgs9NgQqmXQs5fifm8Nn//alGYpqX/PT+e81l9NpCE0NUL4f6CC49ejC0peTt5
hD7G0LkKJfO6YvqMmlFbYdWN3GxvHfpDxB2YGMzHCjYSx0kvMMUYDXcVufYoh7s0VQe31ZFKVMVe
HvA1ELzoml6WHuOJoa3KnDKfWU5FwKyYpowWVeG4ltsRbFUM8KtTq/1vGur+yoSYZcLEr92Q4g9k
KUjnfaKX2pscS9AUDdo+3OFMIb8j9kJJuaxZd3W4aCG/DHdLL7sBFwS6heZKFZQvQIcqM9/ZOq5h
bUwv72+VUyvLUgJRAAAZ0eTy68FK02Oju8HNvatTOHEuNsJQtDMwT+pH4h8zM2cXHObR/tC66a6I
TA+nrlBgj8MgWCB5t+aMx1Tf+MmEvQbFTuiZbq0tLYljjl3AgO6oBkwhssE52Mlwrud1HOFH5+ZO
sUp03GwEL4mSx3h0Q7uSIb9f/NCTqQMF/NKDU/OhKp3Qm3zuZiymF36Ize9ovdJ+ecMguvpa/MOd
7F2RPxD7PqFIJJNYIkFkLwGGFd+mellzcgK0SsKw1ef7F+lnsCuQbibAZby8clQ8MIiSbfNRLILu
Di63qlh0rW5/+Xq5tLAnTivoGwuZL9yLbW1up7/dtpYK0p2CnrDW8l0KW7LGz8oGjzM6n+PFhCTp
JOe6R9SW1UvL5njAkJ4tZj0ZQMqdCv3SnUmD6UOm3WjIskCW9l6gkP2TJk2FVQc8JfDUQguMa5jF
GMcNVaL2y3F98k196W8H7Ry+vlTHIs01+X+sq9KxlmvC0IWlOL6/VSAWk4EA5cuzut8ve6giae2G
eL5pWJGrNAT7Aj6Nm21RiZuEtDzRwzXv/jQwrliYTKjs8SMWP9sCOGD+im+EhQQqyyIFX8J/rek/
XAYX9ADvjrGAMI0DYS+siS9KcjqX3i0ei8aEE46yYdvT3Q7evO+pNVtmP7Zc7WkqAVyYsiwC/fAt
aoNAmnTxzPozP9y//KNMqBEE8h67y8Eimj5groAtgOq1ytIpkss5wRY83hvDCit4GkmgQlmCQQHL
TDycfac+kh/ggeg+eUadmFXKQmgm6iHf5ykiKj68ip/J7j/sHRIrAMM2rEl8os6dYiHsuEaDjynJ
SN31GrHbATr39pLeuc4oXQPsxOfyeTu4CQI+Oi3chQcDbyuXGGGRTN39MEpWtW+Tjnz2tYrX5q9J
T2kC5SyIMDi2T6jLdKgC/wyDUkdgPHoM/HOJrD7fGHencnLeZKrNCNU/DNH6CLMhkp9SUPvKXNM+
3d+6mB31pv/zTP2XVzHR0xHz3TGCGZEidixGzhyHcw48MPVQPF/pSmHncxuLESF/4Jc7Jl5g21aC
QLRbASCkxfyq/CUIxc/l1JdiKEe/gvDj2GpbHraMl/TLnPNCsuV5NVRRgiXLrQmkA8r4W7EDqUz3
NDaoU6EZjjJR9w0BV4098OX8CIofJnbOZ9YZKl1FGt8707Vym44sBhM6k6Vx3pdP/BroNAsSHph/
ZJLdeO8b0qAvG9q3WfAVCDaSjSTw288O5fdDJ1KO1PKN41ioyTLaH7lPRskFR3rdtpD9HIDZi3e0
s17kt8Wk3E3hbzXLktQsqqyBD9Cu6XRbRTFiGMwxb7FTNYsQYdVE+j6trjWQwI9L1p2m8197I7vD
0CbUiqA/yNx8ZEgEsPmMdzR5ZsN74tBI8rx/w9mRlEtZUprSn7dj5kEL+EaeAYZRhhsZquuB0B9R
1mUyne1ZJegLD34YoLj0ooihX0sFpag9kOeEyBgcLEhVNMw5GsJNG6WKrcy8GQ6usr09PGQPVhh2
PLyZlfUf3f9JdZebV1miOxVXjDBUSDbs8P2yC1VsqBTw6Iz/fYUyhifKaODT8+dYJMGztQoTPdOH
cbvGvWuSv1EECJ7HEDptqgNW3UFLIIoNgHwWNb/l6tsGbE+rPKFhUjnXbG4+tu0gXCvV+RQXvOhC
bWK2CvpaOHD3plx7i4G/LZejQpKAAsgv69ZXnznyoEzIrCOI0dPIOC7Ab7Vy/xTU2Xi/H7Bxn3Ns
I+4Vm4caJDzmwwodkVrbL2d6Fo5n5xX7081Dk96gshk8Wiq1tnCb7Pwo2tTwWy8N39mfq3ReOh41
blvxa8KzUe6/P5u5k69tCJnCywPdQO4nQWy3F923D84Inkq36SisGi6+5mODxQVwfWF4WBb9bw/T
9zIywMuV7RU4EqmD0r09jAdxl4dqm4ChwikApwpeZ3fRLTRSDf8qqesUU3rSGEOpLdMSEKFnRsZO
itTPMfjRG+ax8vCz1BLGPRDXE8l+SQ08w2oC+pifwr9HQUvIINBoDieQl0Hn97LFRbNF65IpyEbi
+/Lq65cKv+vZ5lXQ+7nKRivEDJNbLbUtlg6scjG7kRJy3ZWBJCGWAkF9IfaOjjyXzRc2sGZWn6HO
85qMpsifCWrfi2BiszoMCrfyVhIymjLindKkcweCO4c5BKzXHBJBgSkdFMIRBR+DHddetZ4olM3G
rgWOjTMbpnOCfrt4jT+fKXy7yEH2Sshj9+oBtuhMdY1IOQfB8VWMuxLhYIC2DliNr9eUZGLIoJoM
xsa2tJaIZWeFD4C411U+/37WddbCLQKH/fgMoDKauhKVPGqZnfm3QsZtycb3V3fJaJ0y80i6yIO9
0adTz1L0jdLWqVdJagx5X//wN/hfQoBpUWwO6KJQMmGk2Ru6xhlS3kr23/t6z9SaB6S9Mxh0PQ+D
U+AueFXkq3j7WvOmPW2HS0FLnutrN2vj4Jak5nVuzXmOuMFDwrH51HNF6ssiNdUxM2lDNOkYBsKt
EXWdyBn97rU1O1GQFWSoHQJRkluwnCXpBcQVtXT5LmSCScYmkGW9gS8wvYOuehBHoF7Xfnj3MZRB
V9r907fqIvQ7+VkfBOmkmxHScdLrK9XntzdxC3EDmfvCQAlBkcehIS4zDT3b9/BWEekz5DnN5tiq
OLab9ndFBSSzyFZaEbRPkg1fI0Bzu2nHPD+umC0KVNoa3Xt9OcNHWOMj+gBB8KB0jZl0ZLV4IS/W
hNwf8YR0OJEbnLNAlJ/KE5s=
`protect end_protected
