-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oo26J7FnJ2Y6Ul+BSySmH2623Onk6L5XVU7Yjbj4skgfncEdXk6WIl/oeZyOkKbp/laescYzC7+A
gdZEiEpMUVzoH5W0BUYYWhRDEPYMQgMALzwoH5QJpjIoWJhoa3uHVXIxwJsNns2u9C+SN0IxuIPM
8fThaun86WwoFaIvLnlyQSiIuW0pYj8mmaLF5s3iUjIa+WHre37FUvEMGj1PrFDRp1iVgM7Si32l
oFSstRj+i2m4UCyXSymDQJykCApZXZi9qVlK+dWBFtB/KXi8iULnu79EXYR9FRaOXcGnTr19vLO8
D2tcH6lXIHW+NJzwrKCM9OtcU81X/AReVyS+oA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9440)
`protect data_block
qBPN43lNF2SMvUL1k/l/pF1iNu0E1Yr0nYghh47fgJ1dG6wvPizLE7heIE81gF87OrUYvblnV7eY
ne6FFE4poalTfr0vwGkxDAZMb2BU+jKASRvPZJKp7CUlgurVmGHOPNspQngMzXXfIjTW66UjsmoR
XOKDuTpirMROxueq+7lKQ0AQF7+MK9RSp8GuN9s6qiEEzdKiBZH0kOn4VJbg0IhsSSEXsseXAkbG
Tm03c8ZacLfwzVov9VmSQW/hFr2uZP0UPZSMtjxsplZxfJc8xiC8Jnuzyw52oEGe6OEPJf3VGFP6
8lA1UV7aA2P6G/f2PLfwDPwy/ICQyYeklIfAgZtYX8Wnymg1yky71cdZiY2Mkkb8/axNapVOTRBS
UMiSVYBl5l+lunKLAUxYTwhH07fBKKbHapFEqH9/fc995449nEG5iP4ibY52z5NXGZtvjAmZHUcs
ckyotm0nvgsrRVuGXOOVhj0xo9UjlEtlkmkKdI3f/1Dt+g699hkXuojq522t1/VESyhJ3GdImWBs
afzxLMr8qzmHNobT158cObyO2AxtnFKEkLBEU64wFwgQIE+2SVDMPWAa9GDogtTQD7tRS6a/vst7
USDQKOH6JVoh/cGdXaomkXVjkwP7qIgAMh4qxrtNoDp08ezLoCu5rSNvsAq1HFvcfJywKJTgXimX
c5OI963QrmKFadjYiRxr2733uAerfhO+HBWGf2jiJcy6JTzJMhJonKxq50cZ/GN+MuQVhT7WUjiP
UrlevKQUY0pVoR4Q45lm8zdWd3LMFV+WLhzCHLIRCCZIhhMHdzyoYwV9oovc3Tj93tur1xI0VC1S
851B8gzSDfp/l7cVSxSTL+LqpCA9dXgGV0SHDUUkgmreDEqBd9UclIp7+UDwAdV28+AbFJ+8pbly
XUHhjp8dhrN24CNdcaR5wMH7NrmJT6oApgHT6ptN2w78VrKIYCStVP8tAlqiyqQ1WndA8gcJS0Md
jr0di5YYHQbW5/vg8zeCcfaDIzF+33nrPpVR02Fk55FlBrBfnUw40kgDeqjuW1B6DwEeK9s4TYJ4
OAPqJT+2wRL1kXB5D1Z6H6oky89F9znogobH0o8lhsm/nfS6vOE22x0EcJ6JhNZCVPaS+oIr9tJP
ewuZ0ZPWiIH5JcIRcAB1rLZImn9oWvM5Cdc/9WzcMOzWyuvRpp/K62j9o9J1ouJCVFBAjNHeIxlU
hA2VGi3+jhL2zc/vkb3KdOxuazNxnMhTLXuKpdjhqEFmjEyR8Qt/8+/kyDKHqljlGn2PS1Id6FdS
YiqxaK8ocDWNJv6zeVKcFd/PlhUu3M8nx01p3hjxy3SwrbdaJoAIxa0SWvoOG9+pDO7NZbcDoRof
hpwTv2xt8RZJoLog5VkwMoQMPlIgZqemBR7d01PuxbZznh8avdEzK/r4yNR1ZriQ24T+bGhVvSjB
iruxih3H+2vwEoR7JnvKRmevHZbbZqZM67ITpKEPhTrqoCxMV0OwWDtdx0VvmGYjd6C5vT5ekAkK
9PKAu1Rf5hEgmJHo753+ifFGdyuZm6lHHrUTKbE0nCkaNMALNxd7lxPzvlWuPe73dhcrDuAnMafH
ycnaA1+0RqZR8YJZrP5A8/K95FKkrtOhhSxqTTsMpkzsur2iXb+VdUXMiLHHvxymtSxnP4RZdTxG
Vx0xZ0qCZiKLNQsPrUDtteBH8b18BCEmyiOBYV9omvdQyvBYZmB+ptTY4gGgNf35QNn3n+6RNiew
Jc4BdRacLc4Rml7rn0BQT87Uh0NjKdJHq1nfbR5inVpjslQYl/yZgL7g82HLUnxulPlFGd9yl6jz
L3Lx9K1sLPxU4XqA+n9oOnatfbOa/49A/LgH7rd4rvaESGdhfoY47BZ9esILy0tcslN++Q2LIJN8
feCMXoVDWTRwhLjdtBMqxiuJoIbracwzH9BsRAHGe/Zp2wvJDjss6Dv/F/c3XBViJ8xZaKpEEpRc
JB4moeIavPONRo4xyzgVGiO4cOBNyCgjqfe8tEb/2ATOVKwNtiCrMrjCgPYAN7aHHubVblo5XMwD
kvkKENFkKewjK6mudX/rHqlvrYlu2+nZ4llQHOgbVU/OxIsXZ8bBILCWscVDVRvTo7NlM91NsHvj
0lo3+JNuhWRWk3dsKKh0GgmYiwczUbsL9JTfsmFGhS93z0oMKQt7vEJD6HmAlQ9XZydmAvcl2Xjd
MV+uee2IrDJzKLPpVfqQBmpl5xOw8Pd8BFBcgiYn8XTKyCOln4mrbpy/1ZLI/Der6VF1jXyvv7J8
Jb7HYKJKg+wsjr66hC1qLeXuazjp59hX1uZHh0jzL030LKCyeozqmOGVop/EFRVwqCD/XadlL7uf
+qvfWBnNVd3sCUivaSh0b6dPO2kxR/ctEZHSlMyamwSGJKSf6O+9Rwzkb549bBl6DcQGpnh+dlyA
TZDlCCp1kJGtpac2o7YkxhUMTPsMwCdoUIVwihr8/H1IX3UtGZ6cb5K9XD8UTaYoLLHPRmt730Qf
zjlJK8BCFhib+PR96L9WySAXeK4GcAUdkeMOiTdJiZwDIoprHGR+dGeqvUdv36d2SfykgE0cIqc+
bb4X5r27K07I2vjqpkdkJDDyjVtY/6BXWVV8+mZ5u7NEVvc30Aa98DaeZw55uuDFwSvXvov3rmZL
5ZzhZRCGjY4oeV2ZlcoKBAX4vzmaJvwyvWjM/cQ2RMtXENUN6ONsBhlC6K0cSQc6v83oJtQDWKKH
ne8IaEMguTpg5aO7ffcmqRbQusUaUs/QsLA4Qfd8ng6H2WGKGqDEG0LxxhzTMuqbOrbdWC0HDs6N
ph2d1ao+H3HxHUaDfDZZTDuDSJsXYQ5XzQw+i4YQRN/aMMXWaja4wDWmARbf3rjRBt2SFXLePEkv
5qfGAwbHWg+1qHrLlq8bPCBJLiz1aqjwY69TLKc7w5cRgKADEFQ9AWNd0GTV07ojxWuv+iVOakP0
H63tKKG3huYUvvrjB0Qx0N3IQvQT/hTK/rROMmQE4gzCYAwyWFsBQrdn5b6RxEjpSuQbii0RXdh9
J0P87rv5abuAJzKjoxkI79JYkzzNecjJo6ctNAQRF16oWwgSZmAKVRjLcgQfXfEoX0g5n8laR9Rm
uZfLmDqQrTsNdcv/sexiMKGUsn12H2ykX8ffkQb9OJcByCyrX+FRPibzFYTXB6igbJGGXNy9OfjR
uuFIQFkyJLQPYVNuhF5+uVQbnMz5hJB6G2UHNNbDEU2+uUMWl7gAZet8+07godtngah2CDscLdNm
+2BaI9DIDoEJWs1VO5MvaIAYGjJRT5NjHkyioeW9Ko9RF/tFJYyE+yuAUUQed6D+za+3wWMW3RAK
kfXmw5O9VGTHdtvMmTDMR+Es7k4HmswGw8PCiJBIlsW8PH3rBtny236lHlSUWRscyKRkjgTfdQ08
m9DD8IkdXPUDrSUOcLorDhL/PcqE8oTzFX2FE6Bt5goPWwikA/zL061Yeb5hoIGlmW4/qCBurZ8A
IUTJ+nFYZ8kVobTMCY4/P70B+JP0KHkNLskv+D+sZeZCQgrZ6qrHaGlM/UozhfrBtfRLrdkAGU/m
RbyR3edI/aMKtYwXBjReIhOmguRDWVoBHh83s+GE+EdOQtM1Qic6cunDGv0bcDou893siT5llX99
qaFRU+JbwN1lXlO4NEHSSm/rKvApr0XpD+tENLAKTGiAhuAFQI4Sw1Q4zhpKWX07hQuTZJXk6cUP
4cbOys97dPg2l9l96Xo/LQTBaEjOfqm9xAM84Khf1I1DRBdpFEU0gLAts7BMcZ5NLjx8A/RGYcu2
KytXsyAUK9NmAG0f7FnARoTIRggUHzSipkuCvj5IU0sKz9Zqb5SobUhuE7jP99kPYvwa33Ra2wDH
rKt7dgGcac5/1y6QQbVF/dRYm5B6I6l4XHtOrp2DQCxknvYkyuyE6PipXa8Ly4UeAvnlujVl/kFB
I2gDCf9rm+of9PAntUaM1/h/VMyU7klOIFw70LiKUkB9aNak8kwKpBp/KOGnmqsWouMqwmS/a5dS
R6Dn1TsCbbESDneishKGkaJy8+6l+uJ7cEgtMEqoMTZww36W9d1fTP1AAJFLT/JJa1L1ofgQVjXF
p4DwRRB8+CI1HLvYGKeW/mlAEBgFzVuQlfmOo4zyNpW7NrVfpUysj1l3Ky5ZVnNjq/oBc8pm6NeT
ARPLUbRcCZjAY7+FAGsXz6xBIdfbhEwu1EL7XTaWYJfZv6vV3m5WvGqrH7gaoNZd0pCs/OPCLTT4
Po/uKHgC68GJa7NF5VrRa6DAtiNhjYbV2MgFRt8rQANXaEpJ6OhCCSoNcSxEG7jmZHZVbDp5Wawh
u3rNj4Nhh2XLcyFh4/NzPTLX4gMXjR6Jqn2ACQD/JxfCGZVKRXEYNQsDRzBNWV/ZVAPpHIkRahRI
6PP1JJvQM6q9yreFacdNYNKJ3rTMGcHXJOWIb6yPjI02bnVxMsLACREisbT/m4cheBYgiVN8erQv
MCzKaYRgYVFmmhXM88z/miIrOSYFpRk8xTY9lAeNCwwcgnjYETWPkSBULIzmBrrg7cfm+0xKRSa+
TIhTq+7QMH/pt0mtSh82uSypiJ5V417/T71Nto1Gj8Ab+u0eoaJitm863JNH0S8Vgo+vWZCRzz7A
EHutGrigz+qyWsxE0zt/lHbNX4EKEv20fJa364NqaHwYUdqdQM++7iOD0Pn8Tw7gAxGt588lWNr/
VhntRURCxIsGe5/MMDByT6yWjnoREZ7YbSTP15FwcOP6NXIajTxHkV3I2nvW33+DT1by8atMPzrw
M4lGCQO8EKzxulTY+0jFKtT8MO57kiDDQ7O9YZ5JrHHzXT1CdS3SYlApSVN/uZZHTggMJP5D6IzL
+EsNRMl85Ezk3S5vYHww5jFlY3mTp1/t/w820CcJiwAn0P/SwAlMAm9Z2us7JYrFIEELiQdHrpPn
OdZxCn6FZi/pt6Ilsy29DEAnYx65Xa7wtnRYRRo17dDgeYo6YnpCx0fTdGKpdZllgGTs4msFCByX
1fqJJOPLiXEofikTtJLJsivvx3OPRM8iLgFbSeHlusXE8ROnxSa6PgLL49i1FRAsgs7LjlOmwry8
KznCdxATj0NFceS5e5GnzIK7YwCKZvHscg1R0cEAeB9qFRyeB59DPot0rQqnkOQGgLarCsT6SaPU
NoipQ+95CjaT2XJD/ynT44PzoffD48BEviICvZbMSNRxtHmiYXPxGKcKE2bpQdjNvQpeBIqDCdCh
+/iTWYbDp0JZxJB1Gtj5UF6TWPjtC2TSvUjYhEacXsKG3ZmaCU0k58aanwlX7GfXSIhtGxEtW4dI
mdtwl+aCXMe8xuHCiqhhq6UeFMbyN6kyeIUqup4XY+qyWod5C6+r7zvHJt2m6049vqGNCS3aauup
SVeH85Aau/gCaDmdyt8c5QYLOnreswCRrZAdkM65YhHr0MOoewvTVsTeMIEJ4VDR5AC9NwcLAen1
MPGSMD5CDi3ZoX5ZSFrgbr/QHL2+dB7K1G5YKVsXoYpAzSAzchUaP9FS9yekjv3Andk08pD7FBjG
MFWIrz9FCll5JJJu3KsyCmy95Pl/YWoosjfjsJIEXMds9etpSBmpg+fK4gFIB3V5QfbHTu6ZiShb
/tHdVqEx0QrDMvcWy2yyf01MHqkM3VDxuHRqxOOVCvq8eadL8/iHzZagEWbnK2KTff1JyTjYR2JU
+uipszMblLTQ4bnBj8DXeHi2JyWlGOHoC5MJlb5Liz0EQhvJtAA/SnGjnRA5q2f2AKyzF5iFhWEp
KglSjWoTEq8LRGekxkAAlePm8b9z2LF+Qtkndpl8nwpIHUfJYpe7xhHbt+Nr+r+s0DHwghuY3ggb
Qj+gsqwEtBdcnEkKk6TmUT3rIGLEjQeuiTDfd3cGvl69BDdWdXstYdg03cOw0srVF3dwSdgjEK4H
19H5YrKc77V57uqGy3tbmkwVikYhSOd3PPAc8zb4bzsy5o54lFNYhQM8FU0Ezj+VsPUJliXedZ2D
HK//A7jUdr3F7QBJsigR1fQ7x/vx+V9A+sQ/zUI1HksVtP7LKt7YepMO4pAjQJOeRKAXIReSSK3m
4ldUNBfY9dhSgZNnqCRW/EXbeMCVFwSObpM9PYLiMBiYLbpEbP+BBtCZMN9YhSY/FDXf5xZGDxNH
GRG61OsuQ3FqKkMVVbFCYmvAnn7dvQXNMEJnGUlh+zlqrwuHBcQAzzuNxplND8+DItu6wcC/fhoX
lHDiH0XyMjFzhoqeeN7/pP01l4I+Dpb3ptlJNV9kS+OyZzXf7NbSmOlHXG0s1RPRRUrrtbjFIY8N
RWN50PUyUlg9BVEUUzGJKZWioSUUcZuH1sfZOuoZKN+j7eXfisVLxtxgzuyN2blZU3E4WAuDoI37
NsYJBIDqs8hxMWL9WUzXbAbPV/alh6Uwg2ae3mA46FmQW1dnDDkNYDMCRm1sSysJt2bF1qEI1eSM
aTQGUpox13NVenzsZmb95Io4d0XhcbVv1+BLZs5WqGfNrwCQz1x/+FcOMQiWJXJKXvC35GQYW8C4
lpH7Q8v50gxSyI4myY7X9XHIy87afmemzYkXYQR0igaVusA8+YCRFl+Ci3EtOE9P413gpdTisecj
7oVR5RAV8iEU5V0rj+yKt6M7U5SJqpcBydvzZMbXOv6wWMAVTSae1R+uEZnSd/EmGclIzWtvCA1L
RvvZ+nX3yvXlWxeN1qR3Xrb73Z0wO1QqB0pp8bDJi/W/bTWYiWCwB2qizAebIJw8yKnM9ltx6KDK
NP7f+GWqAy9WZe9GSRKjJcwikQ13CoeKPmWqhTyq0fZpe47QMJBkvkPdpju4d1jSM9nN4Th9satw
dfuz7dfFRflsJbP5hWQvIuDW4TuYNO7np3wHPC/2k6ZUjam2aZpOxhQ3pZE3eotkubXphidzeV90
a5oFqGPqLtLJSF+Ct1aTLSqvPG5+sKg78msODgdwnwEAcl7Ttcv4lfDW2gj3pucQS61OfLJn82Rr
P7ugzW35Z0MryMk3XzIEXGuvsUQYyTN410ccrUgE+tO9iLfl3bchLZzqE4dBL0bRDzYQR+r3SIea
1q7QNUFGVs47h7SrAg4jO+z06U2xw7ro3StlPjA1HRtTrUEeKt5vZuxbcRGbStqD6b2EkU2ULl3u
cg2nfPJhxltO/6XfgK+MsPfePa/AVzDMsw0YspBsJHEN/xhUNY8NkdIrHGqtfDd3D4WNU/pYa8b+
pO+6TIj6VV5uW360/TDjJ+th5fA065u9Kx++I4nDX8XW4UyWyciQ4WbLcyEFUkGYRVlqmoZnte59
Cm3ZOvNWOoB+EGW6i79jxqoJu8dcYmxGAd6A7xrsmqdskHzX4O3bOgPNPh7EovR7A47tucK2pek4
pZh5jFs4fivy8XaX4e61yAAtZSqvHrvlFADcZs9NQ8U7svfcQ/gU8OYCexJR3lVZucIFsbKnbIob
3Ghr+C5vMWPOW59bi1H7W5kHFmuuHrlk0lHkAagXHsu+f152hwC3nZMKULuze3UZAmFT7nn1XlnB
s5nCN7fYka06CuqRoAV/oXbdJgseaYlybTLs8o9xDpKaUYVf8J16NEyr80I1R8DUAtVadkAzc6Z5
5oiZmMyIR+eEjX55rHE5HlULgaa+haCHFBnKpS3XFPVan2qTxj2/o5pEUtWg4GR0Lg0bbFEzFWq0
/V2ktYr1E/M+yvpEJjnBgXqB+D8WoC1TGBuC4QrJrxbz4bRq1jWtyyfW5f3PhK+Nm/CN4VEuRA0Q
IJLixAWWq1/OmVs8mvaaUPlhlhJy423PCpFTfJYGmm+rKNY2ek0P0XEbEbcdvYC1mbynzhhTnvQH
zPKvQB+H20c49ZvIVLwHF9r1+FP391Kgsqu1XR53l8LdeIdFE+XWqSzW1yCLQL6TjpHcPlpxgeyI
sKpkFSNun1ECquYm/Mm2QAeZUDPS9orzFiq+7LIzIbTzAyp62HHLaNy9ZRzuoE5wVe6TuSBiB5yN
9GG2B2ifm9+1dnt1rt5hi4w+zqFDDbogT2w1WNT0g7JcBn1OJjvnL/zQC32vTyJ49QYupp/HSZ9J
aAmk1Jm5x9I7Bmt26iIT0UgNpVfAQxtfrqy+bzDJlnigEfM933rrhX68BY1mT56FEIXHWU8ep4G+
3Eb+o1z2pE41KfGv5XjXzYrS1vi0voyco8UORT6tpWr4BMiHgFHaLQ6T7u5hWt+PVDR8plJnR2BA
nUyZDECfAQn4ZSGw1my66Zhr+rSc/Mexy9bg1Ccsllj5HR2f2ux0X7s/QT0+ZLky2eIJ26qx0Fy1
Yk12NoulAJjZBxSX1rijxHKr5DwexWTwYiQ8YZ+BUbH1xYVbWosOHbFFVaFmMYlVY+uK7lHx2J4+
5xR7e0OgF6dXa+vO0K/+5p7bGY5V+U4Icl2uP6xHjz5xIhhBwNr+ccdxLIoOSGPHiP9dL6CryZ3p
Bne6MqLszOFxMK9E4h6yhlPvn0vhe9mhnOF8qUncQgclx1Dx3eDEXTxNWdfym10tqv+E2eUW/RU4
8Ri2YoOcZTn+cwDqWtIFImCciG8UahvsAhHQGvyRkjWQzzo5pLCexoezpGdyd/allalNtxra+Y02
Y2QdLIZkEh5n2m8IW6+9gnfcjs99jMpa/Z/kwKcwJFe+rcy3VxWuUDKxFStr0NX8iJnTjXnClisL
3FgUNAqEv/yiutgIJ9C082oIEuo1lk4/8DbCxk+ZRHtzXOkygeXP2R4a9l7y58QPpJ4K2R6fAtWM
FsQLxJJFvMOUT0H737Kbs682Lr5sxvdmL4/+epG2sTWwnEXGqKV5Pe3KF9ujjVcOi4xCRnNNJfkc
bzMouMpNZVcefty1aRLhECWT/FbSJh9d89V+uqHjMdnxO8Zfme3tYe+lrUmV4G0h+JTkgyf1ghfU
Wqe5bhvniVG0eT8FnuqGFJRzj3KifTgd1Cx4zJwrbAMzh1VxTvdShi3qHv+b/vPaLvIYyMpE2wDW
9xBa6KDVvRUCzr7OIP9FoNzREHSWLXenU2tLCIcpfHDRaVsraC2McxUV6wp7gm+rjUOkof/EDiEz
h3JHtgjkEcEn3Scjzza4x1d5DF23rTRfZ9FZrTiHrUOuGZ3c9uItAfS7roTWEXMjHKmVt2vMtHy5
SYGrUkyF1kqDLBaBrZlNRj2uv3fsBxsN653EoUUEpnmQT4tQSwi+ecsbygnpEPgHFj2EyGtEKeCe
1NFRFDX1UJPKd2sY0tABzmOpbkxzDGW/VVxqLCKU361wGpteIlzz+3Wrg23DIccCaTfRAfTXTQHp
2fhC0Z0H8fsPF/UrD5Pp18MYotUQD38uB2TaHFG3rbaUpzluYt5h8sWneyxHO/50DkfN40CXPe6R
C/AN2M4uwKK0HnIY0SxLA+6yDOXIHBKiLDW1/fJKlp46oMqZnQ7LfKzMQROJVXrEQ1TvVYAbA8fn
q/A/6VpA+IYR1lztboTSnF5I12gt8pZH+Y9bptQCvvG5BmQPhIh2qd3KpTUFfedBkV+/U6FFaU3z
l2WpQyG6KBvpoTp6lvJ9zq28uUwUBzSHv+UhxNTXF7rYf165I9jrj/hiqtmrVw6cbwBQ5PPyNQ3Z
9N9vgkybbLgsBe8xQYdhNC0tyXG6s06nIoU4bUp+4g1lMkwgQSmFhqBt2ThjV6jhHMwNrn/or3ed
n6L3zMPMj1xnxOStrCfiraJNbbTzFr18LQA5am8LDBOEzk6djqG0TjzEXlsXlv5rM/KjvR95KZhc
/5ZlXfC9NCqHSj/yJ87UP0vDSK9CqZAdvkoqi3cQL6OPmTBdGbUTiGnz0O1KYn7R12X4BKjiNZTW
idFeyoCaHBtJmJFNitb6R8vCi+5bT6fAlRUrotsfnrJlqghMT95mO97UoZrd+iCPG6HrRPW8EvLB
GsVQMo4pc7RE7xA/BAPM4wM6ZbkQTkTdL1NoBWsVD8oF02dJCs9KAAabOUCVZA+QVwWh2WhgXBHZ
OA7Fy9OOIQ7GPwyQyNJkvxwD9ZhNMKOYkyjMybcpCr6sn7DeuALBN3wkGG7tsIAS8ue2B2SBEAU9
WGIwu9eYNDlGe3JOyDKkXX5qImxdKbBUPlj6iZRsQLKJPcKIsdbYXBy9UN/i1ii0+p2SFMEDzGkF
gI6ZfucEQWscKKGKmj0CzenR+eOfrCjaSM+Zx+fzcuBkV7utDo1Pl6+4tDvIrwxyhEKmsW/Ha8Kl
xN5/IevRPzvS273eHdi61IaoykQ0fzdQmM0F59mQ1BvjZ1UHUl63zMqi9PTXdGYU7I07GA171kNV
jHISUs9/igTvMIUAqprDqwYbAay6mTqlnozCkk5YyJl9eiWGICxdujBeEmuAivXjwnjhCkY9GqQW
iD4mcL/IrsfGLvn5wFKkrkW/Qz16j+rOjCGKWG9dvYCNyyvRIyrOCeR/ZK7w8YMLHwkT5FkH47Qp
eg6c7VP6jPUyL1D0ZkB0fJwHMRG62f7mutZpwHJPHlgSR+qAq4ZLdsJ94Io5Qvln8/NMEYoOb9mq
APROSTTALFUvcL4R4ZqV2kL8SzpwCLUBg04A5eS0XA91Ih+SKGxHUaG7bGxZQr6A5IfYxjYCQSe/
4tgrtrBs71TDBHVMGwdcxwMg70eRrPJSaM81dLsrGVApUMG34Jxyw3ep/kkFOneFk6l9dtUs+jBi
zQG2+YncszDYYP1331iHuUR9T+XbNg7OoqP5Ot7mptCHPd87YyP6XjISq3YjbzSjTNeIBeF0UKkr
vOGf5Jw8IYXMiVORHagrpzge8j7gt8hu7kGq+uCQpkt3CCgEF/1sRppub1EM5dkVNn1b8V4b5Uwm
3zWPishhv6bGWubCNpia55Kk1ZFnBcH4W6h+O32Fu2PVCYVjdiP+qGjip+rITpXx6UIx/dBQvV8w
Ig8a4KquQ1kO+wR/AJh4AWU8KnINFJOmDYr91hM15jyQyECwgZVHk++TB28PxPwy/SoBNVYjLiUJ
gbla6ikaO5zMgSHFQHa0jn+SYni80dIDKySwelhspUTwM93wIPN/zUsZadfsDK7zGR6jg/A0iUal
Cv3ye07Vv6SI74/buWDpi4Hd8cR9oTyyD7+UhGjn4tRzNeXZO+KTLrThVOdHCOrNq+f1iYgYQ7kf
Gu+4GduC4B//lhBOE1Bi/2loPE79l3+8iIuVkbL4w3XqFRzcxdb/AQT7taOrwVtMYcqbr7ZQbsrj
iMxcBCmF7BJ8bL/zZyN+5lJ1WM2ZlmiA1SLeD1P7bC+mck6evosj6btok6Y1xf93HQMbCx9FDSgZ
DiiJHnMIzgHnr/bqWMB7xMYsl3lIGMdTlfxLFczjiF6WsHlg9zP6Y9yB/drTqmrNtTnDBXl9bkuI
PeMVmBxnBh7wfn0m77qSAUJ7SZ+PwsO+Jp1dOJIXTtscPqvbjnyZFCCwcXwTF6EvaCG/PDrB5N3t
2X9QlRM4VS1lqNc80IIpNItuX4ONnH3yKuDs4FX0XDTEcfkrlheNORk4et6VDVXuSuDRLkqBw4NX
PnkKTLJwK4Hf7tZmRpVMuAimGGwdEy/vikNEIeXVBUOxyTMuG+3+f7IhSE2YmiY8W+E2YQQsYAHt
V8ErVLN9g9XHW51Zxek++wH+kUFWQcAWqbmMpe0BfMhK3w5S7MiFL80i6C2pCG0VIEIarwCqNM88
3yyiLjDIwI6paeNNgNteBEgjOGvaa4ETCZ6JxdhT2OlL3oWgcICYRfeynbqRrTIHA8Qffby1XKJp
blEojN3SLYVXFrEHt1PrjECdD/+TO+yCq7EsHm2dwD9DkVjkGuWK9Xcsh6DSbIJosD9xvXOLZ+Ak
1IC5nEci/9YJFGBkwmCL4jMYQNPmWOlfIB7LUjRK9y9c0lgHyHK4KthOMP3LOlbU/WOZjRSWVfZU
l3gdhVvqUVi9Sz/7XIMe+pnH7AOu/cyjSGrZRcQ/EqK74HDEuiwNnygrL7qVTWWlHkWgYApVedPm
7pFRfpDk2RTZiI/I3OfnrXHS+675IxtWv1xRTXMKsbkVv8dml4pUt+i9CahmlgQy0upIvNLrtcsF
3QciVZTVaB2nWZMiIAWtKLWj/073MWYKmidDwRkIPSIutyz8zxrCjIsCvhjMZB0vj5trUFVpWOSz
kH9gFiZ85H12+JZCVASmcoB0JPLNjeu3T8oIyw+h7lGiJW5iES40yM4RclOZMF40x8BwrlgXg4vq
C4tcMaMvsTcB9drMSAS8pcfq4JOZlG0TKhr024EgUxpwcP0mP4FlqrWEfGZUvcFPZxohR6psqevH
ABXzpjoXVxIXiGznuRzHkO/kRR5TF3UaP4KUqIWd2Y+KT6MkkTgexi28P0Fg7LeGUTXmbJ1Dj3rc
20dpirsVx+5pf3I7gx6TzpJS4u3VrRrTOiiNfW1CSUHbQdq8kuxuBYEOg5zOSrqKJ/YE/3B31azs
HlScpLQvOWmZMVLY8tmjQUS6h/F18Sq8OLinOX4pxjkWpIicAv4XEPJ1eatZmWrTgdo9aH6UT3oT
5PkS8kAaCJwgXtWKTDwPRICk9hF991Q6OXSK5H0fRcIImOGiyNT1S24M/mFZO2paYZpz1cJ5I29+
ZHwFjSvaJFD8WgX+Ez04fHUrd3iX4gW/KYFI0OxM+Cup9pU=
`protect end_protected
