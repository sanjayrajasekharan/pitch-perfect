��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����?%�v��:<σ����i&2�P��%u���di
�MT�6p�����)�╬�b���sssC$~ 1��?��d>{
v��؈D�nݶ�X����O{T�G�ZG�l�Y	,��~�X��h����l���_,���us�\�!٭X�#{O��ܮ�4v��M�� �Yt7��/����S�W��}yZၜ�g��������"�-tu�Z���T�zt��x�&4�:���Mv0�7]?~��ؑ�ۨr�	�8�T��>�>�^	�n4��������L�M��d���=j�ѮSʔd��j�D+��D�D�#�06�xpę�Ժv���9��Y�u-�z9em�]ט-�ϵڭ�E\6�����^
@�VKh�2����>��$�v��Ɛ��n.:ID���Q�nB�^@��A��1������܁cP�Z3�j����@���&���a�)Rw���g�ǎ�+V�+��w�k��Ĝv�Ŋ{xY�.Ճt#�`e�@u7���q��T�^l��c_J�.�'�w-ɦ8�.����wO2f���gu�º���t}��S˱���ʁ�I@�-
h�M�$���\(RJ�_ܮ!cg
7��}jH,gd0�)�D�F�~�P��WxOE]�_��b��9��POdt��-��[���9�b@�>!h8��ި�>ٵ4�6_ʨxXLX��-р�B�{&JOy�+�PD/<p�ow�as��b�i�V�6�O�}L1�#~BK��nm$"a���� ��M�@���b}̼}n��=�6ٻi��_��4@��/��<�������1ޮ\߰@����\o�
A!q:?��9�O6i��m�*C�ϲ(Ga}#��r����մ���c�$��1>�r�d�[�,�#!4�8�R�㕔`�;�������:Tz�k���_&,�zn .n�LQ��T�d�|F����d�\�[�_]5H*��>������W�,i�YN^��)�-���D�;傪�)�u�/>�r��0���m�_+�:��D�Rq��_N�ߑ��%x�����vh�����{G�5�܅*Z�7;;�J�rcvكք�1�+ �WfI"���\u��`�J��:�?�T��$S.%{�H����5����q�eV�f���~Q��w�'�G�.R
oX��M��/�aFf�*_f�dB
}�#:��4qS�yd�T��E�!�~9�SW���W�����˞�����mu;�s��V�����5��wY�!�
�Cǒ�v$��b�SY�䰅f4����:b�c��+�c��ֵ������{iK���ҫg��uk����n��:P]����$�.֢�ۿ{h�|Q��3�R��y�a��ied/�уF����ǪzP����� ���:�|�9�G�<�a>Q������db��3Ek�����h/\��!}�-�
U���m����~�c���W7SI�[o�V�z�n]�����a������qI���R��o0���aE^�<}Փ����3��3BWX/�D�茂�*ó8��\�
����fz���Eր���Ynψ(��y#?T�g��w d�.C�>�����U�$m����7�<�D��/�may--m.Pg��5#a��s�գ�s��ـQ�͕��X꺩��[ȑ�uJϨ��GMφv�+Cô#��"I�_o����9_�Al�/@�xT�LK�P,�7�`'\��>]����C*<�f�u��F$(=!�F.a�A�gK�3ɲ�?���$���Gu[�� T��H)m�S巩�3��f�g��}��̺žM�k4���T �G;4A#�+U�/��Bz_W�~�Y$���BlJ�zX�4�tu���͋��q���͉�(���sk�4�_!#WV�H�ͺc"�8֮.�r�Rr��M�~ȏq����iS�Ҙ{�{�@�{�xr988��_�;W�ԟ� LG�#����.�Q�*��;��?���F�,�_�˅�?R��:A�I�ܶ&�ݏ}�#�Tc4����V%��oK¤9�����۳;?b+t�.aO�YP���j��۽x��Hu޶�3�-�FD6�Ӝ�A��
�u��TwI�n��p��;���_�_�k�0�*K�z:�i[�>�惔���N�'�a���l�[��k�	�n=#�:5h��@�px+b�a&:
��5���.E��;H$n%O�'�X�ќ�f����?XZ.�m�D�.�Y��p;�p]�	��O�y�sO�@�T=^)�-�����v��5����{�!w�CvG��yQ�/D0����N�-�}b�(]I~Њ�n�(���'�IN0i�	<�n�SXZfdL��2�Z��\[38�No��|�#��7H���P�)�yN�}Fr��(\�x�γ�=�/ζ����jJ
9?��-f�ò����\��U�!��ܳ�?7�ȯ���({��u9�u���!�D�uS��2e���`���';����i��{�&��Z�x�����)>�2�o�Zy�M^/��k;bT����I����ĥ��
���n�<��޿|�*���\%�N>�齶9��-�x�ԇ\0{�|q�uI����y�HU����n����4~�����3��Z-�����Y*|o���0{zDʼ������؜�.��Ź�_���i���<����꣖��|
C70%p�~��.̸ �.������Nk@�UEx�I��r�l�.|���R ����1W\Ӡ8�	�;{J��*9p�����g���C�; MYh�J�o���U�>��պn���P�L��[9.�jm�k��q8V.�r8��)�~��M�*;�A C/��KgH����k��^�J��ϱ����ǫS9{�l�'�1�#:c�u�Q
&U8BcON�����O�^L �J������;���s�4\������?Gކ��s5���2sf��1�;9s���[����)9���	�S�S,�>T���O�z4��Hg��^��4�v����&J��1f�A��k�{��#e�o �Eh�<�J��&G���Ue`���i�O��؆`��
����o���Z�8�f֬��V|[�(��0)��	�i�@�&��OqM�9�O�2p�؀%5I�*ʖ��>�%+�*�+��j!����2��I�u��	!�W9�?I*��A�Z��ۺ8Ԝ���������ك?ʫ/ͅ/=�d�	�Vx��V�9OJ�R~�V=����~�;1W��b2�)�\�W�>0-�뮣A�젇Z]ÊZ!%�����!U���q�jا���I$)^����+�	��_i��S$�#�W0� 7�QBb�� �z}kU��@5�7i&S?���`��qȸ��B�z�cb�U���\gK>�a=�����bZ�������'��5|��J"�ʲ�RS/�V2ߌ�c�%Q����^�(�/��k{� ��!i#ʖ\���]~�x��=4w�o�C:c����H���np����Q���u�f��_eixk���o>�Wf����ǋe6��~�����Q`�q�|�cLLN�M���j�0�����/�k�Ԋ������
�˸x�C�c�bT��$��b�X�f4j��&�l���~:���2cR��>�	�#�TI�ſ(�|w��=�\����ί�ܡ�eg�U+�KU�Q�M��3Ku	��^�Q�f�4U�˽�#oR�s��b�F�d���]p(�r>5}RiKdT�:��*NK-��#��S��e���.�Ҧ����`���* ��Z����]M���:�����B�W������mZck6�O����w�N�$;�,����S�,�f#@��ǻ�������h�EKdal��S�:h~�֑P���IْA�5��G��#��%�a\����>tǪ����d�u9����C]��9-�x�a{�����n�4�]h$����x>��G�Fz!o�:�M����bA��c�j���I��|	|�Xv�I¿}t���?��˥��l�$��
�i��DL���`3�R�D�0��/�6�A՘%��p�m*��Pd���|�h&�pv���{�� �+�T��B����O�8��co�l����$Q��:�fZ!kM�r{xo����X��S�5!=!��/������ˁva9#@?@$�:N�+���y�V����Cd���T��<&��1̙cZ�ݤ��8l�r:�x��5B�0C���,RBj�&m8�+���@���|�)��\��I^4z#��}����p����@�1����������F[3���I���I`y�����qR7�z/��:d@+�R��1��`|��Q���-�ʏq�J�0���=0�'I��s��Ld> �͠7u�t�Wq~��.>���y�R��6_�l͖�|�X�k�3���J�6������p
ֽw�0�Q���A�V��V�����$z�j��L���e\�ޑ����fnN~�]�0���J�f�l~A����;+�Ǭh~q������,��"�s�H��&Lܧ3���!�Dǀ��Y^��7�x.{ϳ�^�	� Q��'Im_'4p#�6@+�R��آ;-oLT�J�Jè$?/���ZaX���́�"��� Ԍy��5�1q���m�����+�)p_�qVX���V��.A^��4�������4[���{d��Er���}�T}�ZvYF ����_ìy���;\��՛����E����(.�?��&"bdq��&��0�
�B<��7d7*ЬJ->�����B��Ho�#r�^n�]#�����}.l�t���u�x����Ĵ�
���f����6�L�a�Ϗ;$)�~]�l˄��}��P��-�c91?H7�	6�\�� OIC�۟�F�@La�6��x�p���:��m����C���wVK$���0H��A]Aެ8EX\R:7\����-�0\F�ׇ�����U݀�e����'�a�S���!M&敶�x�x�/~�n�]��Q^�y����ѝP��#�
�0�;�Q�wN&��W�d(��Bʹ&>H}��YLR���� ��.�U�=Y(Zn*9}�iL�c��U<�9���Q	��#+ƘY"��������˅�̾dt="��1���(����=�:��V&ē��n��@�^*�'���ͥxUv�mP�6�gn�Ə�V+X�fP��$:~�H2�'s��߭X�#���?���;������0kZZ��oX/��� lե�K�l�vy���Y-�7�Y�z�ᔷ�n6��������x9���t{ �����Z��a���r��4L�Ѱ���f:�al���_(�ªM�PB�����B!�(�]���0Tӟ�,+�c@-�q�Fٲ(�����J�_f�j;a�����%�'���i4�8	Q���TA�9��5�@J��P�!8W&����D�(Z� ��[^vK�(�H����f��@6����=q�h^�p�����2�cx�4
?r�B�R(ԟY�`V�$��)0�����3R�ZѤpа愧�-	,[O �uj%n�x�^Bi���X�`Q	��s���|
ހ<㘯aF���D�5+�i��p�	�?L'�^iك���X�'��\ͣ6}Y������H�:�,�C4��e�C�`�p��毫_�E;&��b�m�vM�	�����Is��7^�q$�&���yb���sJ�ѯ)��w�6�Ot
�P�HeP3�[h䀏	�d���q��,���k��� ���2'���l;|�0�����ĵ��C-��$�:�2���E$H��XB�p��cA ��:u$�
��)Nb3�雋fwש�d�tc����{��P�(VI9���[��e}�3�E�1')�	u��$���*}�9��*�U�d��}�y4j�M�dN��f?]t����Ć��'-(�#��Vav%>e��m��l��=4�.݀�� ph��H�hPs��h�}�O�|��l�s�kX�+�*P^2s�����O��4U�]����О�{�0��u���Cm������]4����&q)a3��t���/}Rkj[�̻ӝ%	AP �y�A׮���G� ��2 ��α#�a�N��Z.k+ᏽ�IN��0�QHW���po���5�֡�1I�q\��Tu��f�$��g�Z���Cx[���b����du.R���C��&ʹ�9�j{mW^܂"d[~�_�4��Ԩ�����lW�L��Z��XĶ_��-6���	۔����e4��T�p�E9v�K�zv�@���2K�BD���v�Ga]�;w��J�h��h%���KՆ�d�l̡����Y�u���&��rz�6F����ж�$mXPM����w!���\:�����Ř�mRD0�����(��2������b:Od� ,���1���{E���Da!M�3�]�w�7��^j6[y���y��8MFy@�F����� �y�v��!�*�#��s��^I�/
�X��zϑ�|G��<z@��8.��qqȚՑs*�),���Ř<�qoU=��Ps�Ԗ$��0�k�R�_��5S�a v��8�$@�'���U�����.����-?�A�ogp��K�im�nf��p
�Kq_s(Q���h6�������U�]��#.3�;�hD&�Ç�]㲘k��I�����]J�b�����V�s���w���{&[D�s�y�c��͋22��P�����ؐ�فlD0�9���!��/�8�a��׍�F����w����c� M� �w҈���_�W��ܓO	'�맳���i��ͺ��-��eu�T\��P7��̩�{�In�{e˱i\�T���@7:�Y�3A<9�gW��"�b�@7�=�\��0���v�9�u��k�早O�xV�����/XM�C�2 �j��[�ۓʀ8���⒯��,��W������4����.2.��r�S�[F�^��ʳ� ���F�-=�g�����CW��yx��-ET4I֤���Ѻ�k���������YxW1���{�7h$!+�MJ���f���-�m�$�)(;T9qQK0���u���%1MC""6iM���W�R��X6އ`���آ$�8h)�f���xVs�V/�����N��Y���.��O������p�@�����I�CxA�� ����*o����S��fNu��˧�����=}� X�nh3�}�����޿�cjfo�w�.M�%\�_
1=�n��W�2�4�+�R���M�V枤rq�w�U�ųĄj�f_��f"6]��<�p��\̘'�x��wIW$Q�\� �-A92����`3�`VF�Mh7�f� v[�(C�.5v����%(L����{�yH��o�϶Aܵ����n���j�O&+�vE���H !�6y4Y�z�x��`Z�z�(g[��^	o(PD,s�dh�c���9�\��(<�+�%=���X^:ˀ�}܆.���qy�1�v���t_mr�Z5�
�ﱇjE��S
~]��.�h{|��z,Iv�QU��S�{6�ԏ -�F�=T�9�����0��Ll��%HeypZm;��C����FZ�C�o^B!F7�GO��r���^�G���|iy��/칄l~�B�]���2O�`������X��Vi��&y���r�+b)?�+���N!�ϟ��Y�q�?M��6�{�V{�씗�F�1͕�|/`��B�C޴�*&0w�}�>i�QC�Jg���l�\��Z��RxJ��hbF����x���p/�Y4�-�n�f������?���.���B��cX�(�s�Ƥ�������L�R��{!�����%���}�:E�p�N��ul�sG����ĩ:}���_�	_������z�N�l�4S�����&ŘZ!���Wp�CM�6��)�<�=�a��Td�?k�������-r�~��@tD&�4x�e��N���;�+L(�����S�	Y��B�hۣ�κG�u�8��>B� yc�霈k0S��O�5��9M�)���|G���ʿ�Q�TA�B- �ZB}M�ag�v��|�!M[۱�i��}��]�$�Z�5*�tr���pA�M<(��g,�������󼼱.�\ho�"������'%�lCb��=���x<	,y8���?�%����\��Ľ�%�1��}Y���d�.�Q.��0@��`���lr^��c�����f�~2�7���%e[#*���ε�ވ�����u��w;'�z�?V��c�s8����>����T�t(�_k���`����+��Е�1�O,����<C�<��s��� ��+?�?�3��K_�+Cz"�GVWb?�[tF���p�#�x��8�4a�$3�2��܁8a�'np�����)�F�¦��$l��9&_��ᗅ�.��A����_���6d�T�da��T����S�����As�zjX&�BL)��0
�3*�SN,�;	��J,9y�C�&������d�
�0�=j�M��c�G)ϻ�SP����4�W��U�틸3='��׊m�"��՞)�yA�a��pH�M��#�	w��`1~��=�ǤX�!"���4<(��)�y���t��ݜ�mE��-��)��B��6�|j��Ӓh����TK"'m�;����^Jd��P��(M,{r@��\,���h�f8=(�;C���d�tYd$�j��<��r�K���-�y�޳�Q�A�H����MGS�諱+����#�A.i�p����_��&@J
pm�۵*����D)m���X���-�������/�,gں���F�@Ƚ},F������¯����� M,�'�F�B���_3���t>[c��;�r9��A�I��/]�e��~����v˭��:�rX���i�/�M�����:���lXג�ܶ}ʡ9���w�;\K��(�>�V�o'B�ZY;���B�u\�\�h��s�6�B���ʶT,�C�vD�ڭ�n[B�3t��z��N��H �S;�?&�ϖ�n�HF�a2�g<�Ҧ�w��P�����nÙ�u�Q�Ώ«��Z.�J'Py�Q-�1^d���\�����!��&A7Q�ٴ��5��d�ͭO��WӾ
K韭�Y�^� LV]y�}dǑM� ��K��w�$�4v��Z���<���P��d��΁b�§�t�Bl���_.��𱽪P�P��6
� ��m	_�G5��b�ܚ��D׈MB1y��j~�b���|��/�{���q��t%�^��NԓZ������H]��?�9��ra�u��`�ˀ{V����&����O��@�Hnt� �B�˭>��!��(ʹ�� 5U�'rl�Z����5�l������Q���`h�>���1�H⩴X�+vnI�s��vh �}V�y����snᾠD��RE �أ`�t�`�o�XRE/�e&�Q�t�{�3�[a�;U�n\�"|��f3a+K5t��P����0.���A�='GKsV�&�bH��Y5�hN��ԡ�������x��zܝ�[n����a�2�Ɲ,��3&ܿ��*&G�7�z���^����grW��
j�̥n���7�"���R��ޘ�Sg�������"�W�\<��yU�n���xg�����zb�b-��{#K��*��{���$����6{(l�kUO�O��; �χԂ��i��M��j���ƥw�go�0|�eTd5�&5�QJ��O�W��%zaBSf�C���U��~"*=��f�������c���C[J-X��ߣNW���s�!�?��Lߥ������m����Ԏ��/���2]G�I�� 	Ɉ��/E|טV?�5�v9N��!ːR�����neg\٭t���f�WO1L+��
�x_��V�����P������ɦ�1I����td��Cg����Ǯܚ}a��/��[��~�FV�O�m�x����O�|�9|�;��HĤ� Y|o�DE>C"|��;��k�ivP>������F� �,{�j����V>��+D�0e�)��Jl�3� �8j��h�ݦG#�d���&L}9�v͍�b�Y$ N�A�w�@^���<���sT%��v�!Ȼ!"6�S�{�ot�}��9����^C<�@t,$h�f@��tۜ%�pʂ�ζ8�Q�bgg��M޷�ig�x�BI�O�P>�3+7�0
�X06]
6�Z���{���N��3,��%��Ԁ&ڗ�3���P�iS�Qwg�V���("v+��qp�C��6V�+/]K]�zk^LF�;��Љ��|HW�O�p�J������8d�oN��,>�V�1����:��	��'ʑR}8_�
RIMM��<,��˿�������]��N)) ��C�'�eX�/ⶫ��~�_ɸ�&�C-�\l���R�0����f󹏹gUC3��+$X́j�m��$Q�XI�!��!�}ژ��챓̞3ҷ�"!�9�#����ߋ�?���ܓ׬津�O�"aЋ�:��/��hX�)�̉�h�s&�,�^�1S�E�I��ꈼ�=����ɦ�>#҈Ţk�|�x��O�{�����ǐ���p�a&�����%�x|V�ɸv�$D����a���y��g�j���@� ����c�y�U�g�������ؽIȥ,2 _}s���V%�ɛXJ�l%���U�/|�8ʞz���$��HϙP�G�;��<+Q�jXK��ˆS��sv� 6�%s�N��?s)�/�)5�frlD��xS��ͱ�Y@�6����hl2y�F�!��G�&�k��:��w��B�Ķ�U��.�	��.b{)q�C�׹w���B﷌V��o�y����t\������S�Ost���^/������I{���u��#Z�&�$��Ý�U��oƊ壖��?��� �wc�C恣�م��C���@F�J�⼜<_D7}e`�8E�C�����K���Z��.h؎)^���" �i����X���3J\�O&͏��M ��Z����Ř��H��@��f(!<QM��آ� �!m9�j$�D|[��󄹶��S=����jLN��b�{ӻh��R/�}w3��y�F$æ5C��붺�Z͝������#���=4!�6���ʪ;�a�,h�
ŒC �9c�Ps�O�ĥi���5�4YX��!�Zut���U���kDF��.T&�hf��W�4ES�LOs�B�fu7h���������JFi�]
�6�r�6�h���^ϫ�ߩl�I|����{����Ʀs�_8��:�b���k�NA�Q��������g�ݒ�,$�b�;;�w�331[qx����[�i`6_?)=�_��O<�S���a��0��w])F�1�+��u��}���/��?�B� �	$.-l��0��<$̟9'�=<���|���y��ؽq�t�\���X��w6�%�C�K^Y2$ �_c��m�:({����q�J��S=�x�%��/��>�����_�ɴU{�j�R߉:�ٸ}��+��-
�s�0�:�Ͻc��'Ob�.��6��Y��a����/"p��o�B�o�`aK#��'�
ޘ��~����*�
l����!�6��赱6���],��v�_U����T�\���chx?K����H��#��T�J��U��h˭��Ѻ#��DB/)�\/�ҩ��Apf,l�]�Y��[+.B�Hާ���������Zz�8)�z ,��tG0�|��s���c=�"g8��!J��(@�1�b�qB��CeHϭUT7��&���G�ͬ����k���3;H�@3,"/�&���[΀}��z�Ӣ9��(Gtǂ���'���g{T"����jTN��rxsW]6ɍN!����p
�3�?@z^���(}P8:7P�N3Y�:zLЮ)��*Uy��en�Ҥ�1�-�Gd�|MM%jI���O[��	��� ����`k8��i佑d5�b�Xk�mp7yJ0{|EH\I� �G�!��'��t_j��avj�=�J-�,S���� w�`^��g�@�w(���7u�5���0����N�'�6���|^��8�]����>�������]"�3����5�4o����!Vꩄ��H��,݁xH���c\�7�'�:��Eo�[�+_��糢���������Oo��a5�x�'�@�����+���v ѫ��?G�Nk�	����]����3�8�G�_���sFŐ=O|���w�+���Թ����}n�h\��({�i�2t��pqD��_x�����*�1�Ԥ9����7@gn�͸և9!{�X�fa�զ����L,����o�ƪN���ho��9@�ªJ��s�LT[�mpF[k��D_W_�x���R!�g߀;7�e�\�>���#i#$ ��B�8���-l�d��bLdMZXs��qP���fW�N����1�$�<c��(���H�:�2�Βgs�1���9\X	s4�A����.S�-OL6���*�_�V9+��e5
h<ĩ�,��<�U�̀���PDU���Wa<���0���i%�B��q�f�Yb�ؙ-C~�o�"o\R,��w������<�)�*���Ȩ��s��(Y�x���d�|Mߜz\Ju�/�xi��qa&I�]�fk�Ճ�#�'"����_�@mf𜙎M~@Mʈ�{tx�dz���zŻ9�} /�M{�v@���ab�ϐ�������krDx�Tx{}���+�e
3�Ƚ�Hj���3�F����+��F��������es�����)[���z�wP]m��$�`��4O�ו	k�P]��5[�5��� ��=/�Y)r��&,ؼ�5�A$�^9X�(r��r�w�R��֝�Y�!F���Οy�+AȢ	s=��:�ƅfyŠm�y ���$[��ٕ=���		z�����L��f�z�_���}�x���6Q�n5��?d�i1�^�N��).Hˁ��h�y?4r�tz�mƔa�{�뭨#�A���/ M���_�	��{�5�,����,
����,�ަ��{�⭬���(�Q+Șqm�/�hZ��0�}�����T�f��C
�|%�,��R���gލ>�aTm5q����pipr�!�^(���~��7W4�1n�}���Y�fX87)��)k����y���\�R��1q���,I(l�ni-��	�Z�"�dbs�y��l��>��4(�s��\�r�����_��W\� cV��`��$�DY�3`S(9^�K����ȉ��z���P@G)������Tm��0"�n�d]q�J4�S�-��ͥ}��
b`���	��.�8�f����u4=�:�EvƱ��%�#�pV��&(����6�[��M�+��W�Z��:��2~�G!��1�]t��R-RhoC�_�!��%�/:��.|&�����z;w�����k/qm�!�:Hj�P�%�F��`%#�熢�`�QS I�[��h2蒱��g��,&;'�$M� ��F��#�5FV	�i�B��g��߱���uc8�O�4|�z�886�86�@��;`�{X�	�9r]
W�.Jv��5j�P�ڛ+A]�+�r���E�WL�yn��}H�1��)=�Q���7��ۇ�LF�ן�6X�l �mήk9E}ￂM�	z ��)c���H�[r����R�^��X��k�������@+�	 &�è���ݺ���p^�bG�@�n�O��
*����H4�^e��:hs��a��+�<��L���L�?��C�bT��$\��UjQl{��
-�`b%H�<2(Խ�
~/�6�/@&�:�Y�k�M�!(�L-�x
hxCe�2�	�Z��97I,�ó޶_�~�IcC&�&W�(�XC}����%v�����oM�D�>B��T]#�n��XӪ&��~o��.�?Ҍ����;�B}2�Ee���K���g�q�O�l��X���疁sxw����tX^?v��A�M�G#���XPa� .�ȶ����}!���*���0����r:rCK�)��GY"��ﱾ=j���ԫ�"n�-��b|YS>/F5*̮�H�B.�>$C�٠��V+D��!V���Bi�p�R�pW��_�R��"�S~pk&�_��&~ 1�bx����?3����}Ǣk)I �qXuF$�6Ϸ[�j69n~_D�2�� ��폌Ϯ��׈�C�m��YB[�!~�O�������."�
a�Zу���T%b��I�D�f�? J˩�u�z�/v�����K�s�W}e�����	*��)y���.�y�}�5S4e��c��"oP����S����k�;�~\��!��]��Y�Amq2����-n���_�Ű��������-��9���G��hM�+���a�F�v#�\���'B�m�������+k���S�qT��8f�1���"l����77��l�Y�����dx��t���.R����c�A��r�Y��X����5[��+fJ
��52{�[Zug6���lu�V�,��z�wN?�����``�t�>m�wvL�������|������;B��zt�܈��M��r]�����������C��h�x	�O4��ų��D�:���A���4#����e����4�9�ɘ+�7G�U���<���i:�u��<R��dU��kPNk�("�F��g�z��}2%����,��(Y�S=r�*�I�cnR�p�?��'W��U��*��$�l燝k�w�ï8(7Ж[rv.Z�̵P���a1�*^}�I�D��d��aD[a�U{�� }T�.��*o��W���<����I�6�p��E���،l�o$�����]l64�t����"��ٝ�&�RG*��?Yܿ�ht��t���_��u����3��j�z���K1w�Μ��OBAv)�zF�zƻ��Ahu��EՎ�X8 ��ZF�|#H��S����#�L���	R���쏏��Y>)1�5��6�S0�3V(M6�������������ۈ�T�;�ی����ގ�*���`��Q3;)卓.T--�g�5�S���D�������2�����ǿ�]���*��?-b%pkQ>����h2o�hTܣ�����~��������^� @6��;�V�(�����h�>�d�
{J6��Ss��Ig�����锌�ʆ<$�� ����<r�=�E)�41��f��y��B!���G��cъkK�o)嶜φ]�1M�B'������Z�����5+�kH�<��-~b�W��������侧��h��q�#�	5[J���"����$ì�Q`.Z*��'v��;��s3���/a����!�{�����_T�FO����d?�59O�����UEc,�J)a���[/�y~_�(�������W~:�p�r�����"^q�3�9���dԻ��9����Պ�;�p��#pe?�cr+T�X��(��������0�غ��0�k7���#+ܠ��_�4��e�%%�Χ���ߌS\)���_�}�_���ʡ�3�XT����,�N6�݂5��{WFǺ��<�>�k��ԆS�t��J!��r�8�AD��4�g�n���_�^,$H�Nq�>˘����,1��V�Y��=֡7}�[ͅ��vcت:�".�n��*We��&`�'���+��՟�{�ly�Fn�'�m-T�|��`҈�1�<� ��_N�� �2%�Gn�K{�d0��hF�m����grʬ]m
1���$%�h��5Pߌ�.��0a+cB��M+��]�P��W���ZJ���@-�2�	h�=Tk?4Ú-1��O&iț�{���n��9�2oZ�WEJA�|�>����f�]��p)r"h6օv��U�7�K-7ȐO�q�~��+����!�%f�k5�Z��}@±�鶣�������O�DG���>>���'q����}:d�j3IQL3Z�t`V��.E)���F=��ť�s+3-���ٔ/&\s�{k`�֗�����t��EEE�T?-�6�T��AT���,�;t!+V�j�8v8���W�њ�ˁ��B߹f.x�:eV��r&z�S����ղHGh�z�m�^��/+�[}e<kZs���̘�N{.��?��,��]�A�����u�zi,qRd�N���K���z2,.�tm����b`�О�e�Mس`���]�_T�!����1D�{������r��S���;��L�:5R4cX~����O��V�Ω�[���6���8�àoAQ�����r|1���°����Yj�o�׸�L����r�z&z}��Ha�x�L2�8֒_;��p<�f.?=X��崚k�-�����\��N�O�~��F�]��H��cQ>���Y"�,Q:�Z��&I��4�����Y��s�ٶ6(��v�j��A}/�>`g����{���e�ũ�:������r�:�֙gVA_�z�U}�i�-{��9<�gF��(\�'�̓}��M���{�\�q�Z�3eR�7}Sd�;.�<~���`�PT�mJ�{���6�Yc'<�!����ߍ��/ zC���p�	N���Y��=L`&�4EPn^�D2��a?�H�<�h2iL�o�,{D@���c��+��|�Ky����Y��$(��`�l��3��(`�����7Ћ��"-K�� ,g���>�$��u�؞
�(��Y5iix]/�Ii���\��$�qЍc冽G]�!��·{�>D�P���9��h��;��4~����t�8C�����T(9�E��Ł��6���ppHƗ�"%����C?V���j�Y��!qB������C���g;˘�α':ƖH��&PH���1k��"B�U��10y��{�\C|\�G}��Y�EY�K����9��l��@�����:���(���g!���E8�@�?_�>�.U)�:q�7)>�u�Ż�s�N*�3h����nGn��d�qi֛8ʗoes�ԅ�-�Zg��;nAAе��t��
�
�n&��8AY�4�в�J�m���oz�(ƛ��e�Z�co�<�p����2AS���I��p���F�� �؏���98>8a+SŒ�r$�0�*�Q��Ǎ�J�ڦ�YL>>x:(�-f�}�m?��3��V��1��Xd�� �$�p��%���`�}��-˙���Y���d6]�dZ@M�V���iQ�����*n�~�)���� ��:�c�}����w
��F��Cz��u�#B�G��l���@&�fxsn�]^��.�������PF��0�μY?��C+�"�m���J��1C�u^l���IOp��� �OLDA��􆹓�Ip�'*k���K�Fp�T%�؃sj�������r��@AU�8O��7�s��6��g�;�.w��]�w|��a��G���H�ׂT�C�g�Yc�Nw
����9s�m3�'��@?r�;�,�K&�P���-{�x�?�5�28^.��`��ܷj�L%��Ry��<	X}z�z�k�����&��k��+���͛&�gv
�0 X�9L�wl�
���P÷��6<�cl|�W%���BE{-mqĺ���֠�Ck����@����J�Ɠ����׾���(x�u�(;�i��d�� ��H�ul��ӃK�Ljޕ�K¢��yDK����s-2�
�u�ij�ƾ�龪���Ϳ��>�I�/���;=PД1^�vgƶ��^�u�p���ť��l'*�rQ��	Rb�g�;��?0��M���a,E3��۽��AǮ�[~�,HS}�@�an���a���e����[\+�)�@"6�I����u e��UI���S�i
��%|��(�j��>t�5p��f�)�f,�K���d,9+��[Mޫ1�]�d�K,,.�Oշ���H��4Z���Z�x�₥ܡm�Ţ��� W�	�s4w�f��hoo�5�D���_�]-N��P`3�5��3���{��X��`�j��A�\�n��Ib?�nUn�d�O�;�$������y������u̴E�TSz�X���Y����4�6F"v�
C�����ަtG�
V,3��xw�v	��Zl9X�՚�Sǉ5�*��+����N��f��B�5�z�����=�n��5�҇�@�U�~a��9^���],q�Ce�G/���̤�~:�C|���� ���#�YOv�y�*7��&ϛ>��{k���m�CqƝ��s�y7������<$�m�k�iy;�g*��G���S�8����L\A�����{[�&;嗘����Ѩ�,RF�\�1ԑ�h���D_\�_p���=�z�\1j�T=�T�T����=
ܭ���W�}anc��"O0Q����͉�^oDl�4Ս�{sR���JXsr$�i�r�{���R�$;���ce.�`~��]u��KR	�p���5b��O���`����d�2��XDyH��͸hG� �����.xI�����`�#���҃��w߁�S�*Km9��l9S�������'����#�	�`�bCA���Д�����N�U��f�l ^�ʃ�Tu���4$]�p�Kc��yi���������>�����=A~�@y�5}��b}���h��b�o�ǒoČq&���<�K��7gb�D�6@�9`����������c�l�W[�a���\W��w��>��%�a�<Q�õ�g��&h�K��븺��Ҥ�����q]�]%��(4:N��Y?�[}O�-��ʄ��E�!���nq�₭"W�}��� ���e��� �vU�Ͷ� Rj�:�)�����Э�����k#9+�!���9�����N'?K�J��z�U?�f������=��	��QiU#�n���ħ�& ���Q91eg(���i���W���zRLl����I��.�f��n]�6[}ѝ��/��z?��F�q�Vw?��r�|���?E�O8�;���	$�E��G���?�1�('$�~ǩ��!*�'ڿ7�`]p�(_4�K�ax�{���_����2qI�:�*z,���v �oU�Ů~v{O�����t l�37��^�C؀�'�4�n[�  C� :H\�����J�c�8~pT��=���j��.�ԟ��	����]��-x��A7�X������o0�T�G��<��c�J��V����r�s���$"S�`X��;��c��\`��՗f�l���K��+�R�?S�p��f��� -N�C7*��ܛ��!�܄�ȏ���,g�ԥe>�`�g�J�.lm������BhV����5"���= ���}a���P湺�ب��o��V��q`�EM�r�]�x%��<��%��P=F���;N���k�g���D��z�����"�e��c"מ�A̐N�a�.l��N��r�^��]�Ωo�߭������J�KMrR�����
�J;����H駝a����.�Hp'����Cp���F����S���	�`�a���S�!cIzאԷ��k�^��~����'��f�M����T}�@�V
HGR���>�I{��և��6��F_xбl+"����Z�V���9e���z���w�c�_zd�5v���+!�����hB�K�����s̄2/ѓP��@$���F\c��p��{A�ޅ|�E/��k��Ο�O0�me`����0O�{FG;�밽U��V��ᝑm��2d�vC������;[G`� ɗ��H�[��/��<a��%��3����sk^��/��>�*н-���E�+]��-������|Y��N� �3ڧjG��>�6w��=��un�tcClg�&�_h�$|�*j�KC����u]̀L��G)�u����<�0�6���&�j�66�\t��z�-�\=��%����{���Z������f��iyV����������K+��)[��¥U�H�n������F�w���)]+�1����2T��8��"��d��ю���ï�'����%��H��|�t�F��(#��Q؟U������uH���� ���ێ~��#͓�S�Φ�Wh���}���,x�����H�z9gdM��`���]!,E�ߟZ`���+�$Y;k�d�Я=z��k����А������B��!�r5�c"q�ѓW�ԡ�&�m���X�K�_ݸ�=��68�	��A���P���o�wU܀=u��h�m^C��r9� ����Q��r?��f�����`*s[0ҧ�5�I�x�4l�p<��p�t�c��4]�=�S�탵<>(Gx{sJ��I�,��%���O��=�c�6)
�4��=�K�r1;�| Z̢����z�:Y�������޹/��J�:h�k�&
פZ˞������)3
c����y��.�V�R��j�Q��z§��CVeMJ���a1�@ �qQ�b8o6*����?�����@�ܿ���h5>��?G���`��OG�Z�v��e���$}��-��R�I�J�怬�
9�*ivE�ٝ�/,z_pPg_�
h�&�8��k'��d[�l���قC�}c�D��G�rE����])E+qi��+j/�2T(ߖ8�O���?*�Jt�������+����`�8F���\��_e����ݷ����u_�MɃuO����e3�!M�,��J�AL9�z�~'z��)v��N3���ĹB5�'讴\�^�㒚qEX�A�mc���^7��z��4����ec�u���7�kdB�aL#�@^��c@�z-��L�1��H@KHT<��yê�9�qO]>M�BwS�)'�ʧ�<k��!�4̂^�NV�d�dn���/ ����:�hTv]y����u������X�݆	��9�Py|��e����k)}��慅8.��Nku���g�$G�R��8�y�=�Lbk��_ݿF/�(d_�j�u�����R�]�[�*��c�d��m���LJ9v�zQ(��z�Tт�R(��r�S��m�Y���9&�_�����?:�ޥ�h@���ٷ�V
��wNq�-��9�������� ��,O�u	ڵ3N���H6�$Q�6�� �\՟G>��J:�)9辚Ϋ��2�QՉ���Z�03�,��3j'���jU�����^6�~�Q@I	�x�K�ƣ"��Kh�B���;e���� ��$�%��ŉ��'���%�c/"J��c\�Vv��U�	U���7�~�%�Un�~�ď?�ֹ'�l\�۾�@O����ih4���MS�cl�ie�2�>�����#�v�p=_?�V�G�["�����@P��;�z�۴�R_�MReC_���J�9{��/��"l��yX �M�<oA"Z�逛(X�U�i�\8���H� �oIy'���F�+r�����l��)<:��Z5M�胉с���Ag	��j�ՙ���N�
��ԩ�]_������`b)��Uh����9-�zm��`�<q�ܡ���rj%�iއ�d[u;���JGX��*NVX�;o�*���V.��K�����a��^���>c�M=�$����;^���y���_��.�wá4��yZTc.~�`-H��%C#��u�Q#�O�������[�cÈ�B��EA�֐n��~�٣�_0\��i?C������XG;�j�S['��a_\�Ve6�%��|K�N,�vqK�3�E1��J����`���jgT(��9��o�Ȏ	�ߘʨ4��ny�.b��$�Bx�ی��8���h�%|�Q��=�����>��Xn�,b�E�>"�c����xD@c��~�I2�f�XhJ[l�Qcn3�D�ٻ�!���������{#�ˑw��Cs��/�{yz���,q�&&��^MVjR,?B���3c��s_�}1��s�9�;Ɗ��)I0D_��d��O�a��u�i� ֜CJ�VP1#�@�Ok�"����E�L�]���i+�}�X{��H�Әn��-��I[	�襳�@]cGRPH]�F�վ�%Sq��s�>�'��ۉ�`I: �$<�L��v���D4��lRu�쏊\W˞g]�e��s*��r4ާ�����{f�����V�]��o{��ӳ��`�ܐ��%O���z'یU>�&�R��)+�� �&��=ޒ���D�F��-
����Ap��Е���5�ߘ������60$��̼�QC����I��6w�FTngҰT��k�k�Y����/��q�������^4&��;����P �pK_���*J�02��s˦6�!��
0P}TO���jߢ������>�b���
_����vH;.��8��m~�M��yO�(q*��m���r��\s�a#�x<Of
�A�%]*C��@��ʔ�P���P���]w��'�P���5���l�\�:��l�g��4��'I���W9@@�l>����7�c����y�`�'�"D,͌
��Ӗnc�c�Q{�r����*��\�O�B�L�}M��G$�8��)BU�>K��{��&	8e���w����� ΐLiP�Bau�{֍�Ov~���~�h��-�c��M��3�Jo��E�w�(֩�H��;���@�QN�a�A��B�C�af(IrX���'(�r���Τ�22S�����7��z�R�{������XP�f%.��ل�����mV!�E����^�`@�%�}�Gr4�+0�K�Lĭ��L�Iv ���m0P(��2�2��y�����S"����B�g��y̢�n:�j�������'ݨ�����fB%QPO,�K����N�����m�j�����t�CS�!���'�w�by���$�����g"�N�>9=��=ƨ �h=l��D>����t���X?�z8�8����
��cz�Uw��ɺ7��܂�\	��=����t��l�PV��h�Ҷ��8	E��X^49nJ{�HP?���:��b.�s8���;ka�*:�7$	W�u�3R��T�O5k5Z|��|�b13ԁpZ��+r���!���gxV ��o��k��Sc����mͣ�Y*m��˴p�V�����T:���fQ�o�C�7��z9�GM���|n݃��U"���4�֛F��:�$"�s��ج^�&)��"���H~���Ƿ��\�/�e����C���h�q���a|���<9�2���ܠ
�1h;��a M��9�6�s?���[vA���5 ���nxK!Ow������wf �7�ڔ���8��$�bw�j�&O�n�!=؈NS��e���m�fc9	�Z�}��@��Z)�{�2��/u'��fU�}M�w­Dț���,������UV���	��h��i�@߭�=
��e&s�u_#5a�FSb���~V�'0��7�z<i�|3q����F��(x����
���꽃�"Kn3��h��n7�|P�
�!��.����siǅ��)N�8�W���GР��<�ee��+w׍q4(�2u����`i�H�n��S�7B~� `	�m���PZ��b�_x�p5/p�{b��_�.�B[9�G���s����Sq�-�8ɼs�?X�7�q��w �s�*@��*��B�Y�LI9!�[ї̀mĎΕ�i����I����'��3Ʋ�Ԣ� ���|X����e�e�&�`]�>���s�t�[��2짚
%��UB����R�I��vE(�B�X�-P� ��f�1�Ө���C؎x9i)0�����eȢwI-L?���1���v��qO�k'C��H��4�	Mo���(F��8�ǆ�������M�y��]hiGF���V����N�:#Ј4�c� ��z�|�ehgsaeCl��烮��Wz+H�^ �6[��8qO`wiX����`�/��6y3<�h�9���=�ݗ���-�I~'�<��[IBi!QNu-v8/KXE������>��I�}���̮�:xj*K!5���Y%Vo���,D�_��$k_���%��F�?Z���5����j\줞ނ¶�zT��IY�]_�{*����9k�+�͈��Ju/V�1��j\�Z�������6�o��/� �ڋ�K�_dPLǎ�'X���bih��H�B�/���f�v/V����D~Q�Rd�w��0�|�ѩ�=m䋃�,ϵ��Ͽe�pB�If
zl�2jLhC9auʡ/�/��b>������%6�ʅ��A(���p�����16V$즰F��W�OI���NP�=2ȧ}���q�#s�9��6t�Gפum��b��R��n��^GX�	.��γ����{7v��3>�a%�� d��Fo�W�0|9�q��A��5A���f����(����RC�_M�^��X�FC��a4��ׄ..u<�{������&L���bT�I����ݩ��T����ل�o�'4��aM8V�fIF�3n��N)��0�O��i�>�a�d?�t��Z&M���_��s*Wǩ
Z��(5����V�y�T�8ۛ3������2��Nf�"L#��0�Lo�eF���k�6hԬJ!���om�?�?�q,�6ɥ�<u���̸�h�v�Z��_���b_ir�"���� �KHwD�
R�!�Y��	8����d|W��F�چ�>g�A�'g�bƷ�`�T��B~_�5�m��z�Z���F75�%�HK�����"��S2�S��1�o���H˽�j;F��""_�����8fJ�#��Џ;���=�~����/����8�������R��t��Ю��r`?6�s�Ǎ����D)˂S�9���~��g�*�B������� h&�/c]��Q����aQw�\��mf�S���>0��7\%Xقy@fܚg�e��&�C�'���5�/�ȩO)�`.y��O�N��Y��0�X��=�R� 6�i��S��nJ�5��d�&K=�D$�y��m�G�䧏1}��S�.ta�=A
�e�(b䄟dM��(�G/�0h%Ik ��jpBO�����{�ҋv����O�� ����+�i�>k��滝��7����M��b�$[��Av��S��D����^S`���L��;�y��cR���# ��ߖ�N3��q�pK�j$M8ݸǶ�J�I'xao�4a����g�a��$�b��E19�=pQ8�)I���s5�=v�-K*˖�h̻h� �I��H#�:S��/�;���&O2��A=�{k� WRF:O������3ƾZ�B����2��+��RZ���F��ݓإ?���4���U]��Y����-��T���#_W�
�Ή�����I���H�ُ4��;�:~�t5�$�n�%$�i���,G��
��o����+�I|�G��GO��tp��EO	s���5�W�7��C���,U��I[1���F�'-���W���z�+±��Gz�N����#���9D��	k���O�b�ӬQ���*6�F�M5Q����ph/{%�	����a�N<�"��C�`�)��ʯf�pr����&�Lk��q=�ᤦ~E<�)FP�{�}�����t���^O['
Ĉ���}���o��Fe��Kz)4\ n����.�	a!|�y�d��O�� ��H<�0/�|93�LH(÷ɏ�F�~
�[�L�e�BMq; �,�
A���O�ܵ�M��D����i�F���r������f�8j���^j8��|�b�'���*;�����pd�c�G�G.��,���\����1~�jzph�zPoZ�*��#jb���7�w���A�ॊ�����3<������� ��㉦ZaZU�#��"�&P�H���	�j{@(V�V��{~N�����s��Sc��>�m4H���k����%�ғ3FD��N�֕��`��W���{����ό5���8�!* ���7�Up��<<k|7RNl"�c/������"?;����p�Q�k�6���^,xk��t�H1ǯ-a[�~*[V0,�v�5CG*��7�[Mˬ2�ٔmnMq�w�\�DrN5�����EǠi&������#��1#��@2�?͠����Σh�}�h�w�t�k@��Omn;t��3�kú\|Pċ�X����dQ��|�
}��� i/S4.�+�5��l�`��w zוF�	˖�gnȂcj�3އ�Ӏ�����:9=V0w��D:i;$��$��3,x:���:��W����VJBnz#Ft�O�h��EK�5їC���;T�h�?�qȿ�Ӹ�j�R��D �q�����^�j�	��U�RFt�x�z����%�7��D��,�"�i���*K�݁�F��"��F�ż<���O���<�9�m���w�&��j��@�`Tی�f��.�-0Ys�ڮ4��f�%!T�����g��|B^S��!^�)^�
-��O���42L��$� �1� ���H�J�ŉ�S�u��~]W�4��:����w�NmA�I{IUg���ڸ�k�&��<W�9��������a5S[���\����ȳ�&�C.�E��;0�H�{jw�5t��x����I�@��-�w��*�W�^ȁDu��58�j����]ȸ�in��B���twuI�G���T�e�}:V��$��d�"u���`e~Dߡ)φ)�����x���w8�}w=,YG�m�l}�'j�]i	/�vO�OY��P�YMD��n�vEd��fe���)�Q���H#��%b]JƮN��%�Ks�h�i^~/LK������Ծ��h;�CD1_�@ p�q�z�J��{��wր�(Pz%�%J���.N�7�7�չ���/N�j���+]��
p��9�&��ӫO_�~*'�ȬN�3�I+��m�p�"K����_v[L2�T���#�,�l��0n.6[�=~~1�{��#��+,�N�J�Ӊa�ϩ�p�%Kx���C�6|Z�G��B�݇g�'�����ƪ���o���3��)��=�����7NZ�(D�p�œ��L��C����-���=>���]:ߺ5V�9��%"_ @�A1x����Rt<^E�>.�چZ:�s��s�ej�����{�X�!1�H��&E�g�a�+X�a+�����YA�[���pЛ_�²�yC4���A��e:E2�Wr'���('��&u����-�2HD��Vg3n�	H�\N��������Dq�"��jA�4�S��l�J��8aD׋3��K3?��� �|q��*������3,m�o0J<Sl��dK@�ѣ��25S�'�?B[ŝv1>�B�y�:����LݒQǕΝ�-�Q՞K�7v*�,5Yz�W¥\�?��SfԵ�K�*4�* �)��\���;>�`����ԫ�ܘ���c�s�<�b���}U�
({PrB��FY�~��C1S�e1:�I_�l�
�'��~7��`:���9�� flE��{{���oL�� �/�`qxT�u P|�
5sfpp�����s��H��O�"�$� $wBf�=N�b�u����d
L>��H�>Dtb��G�$��k�c��ɢ�Xhę�B���.�봙'���:�Z��Z�}�p>�1́�u����8��r��s�b�\Kmlc�k�u�3P1�@�?ܑ��Ai�����W��_��+��N>�Y�&x̋|������#�����T�< `m��¨�`�M\ֿ��q�e��O�����N�˪I�.n�y�[ ሑ���H_D������S~ǝKe�2�4?_@nC��R�:�q�$�*�6cK@���Q�m�#â����s�g]⭀}S�Kjߤ�y �S��L(���\d������֡e����l��<+��k�8�%�=��ԓ�8 ����1.�Z)*"��&EDF�i�R�cDA7��{���H�Y�$1, ��|�D��_(�րk��P!.j��O �i�Y
��fy��U��l3��U�@x�aK8�%k�|��&+q��Uk��.��4�i��s��%\�!��ݛ@�r#(��IJd^�$�e� ����a=?�M�Rb����"M�Ν[��}����G�dLlXD��74'�ҡ��k�'�����h�ԑ�۩H���﹭~&�U܏�vv��1���tM��d� F�Yh~"%͸,7(��	2�d'ζ9�jrKxj��8�Q�ˎ̙\C�j�&�@C�E���\Ó�f�q�A��/��_�^�����y���r��y^g��E��k�F��<BSp
�&�Gq쒅_	8�"M���缅h*2��>Յ� ��b��t������qDȹ惭�O>�T�q(_��v�ȄC�x*���=�US�lm��G��<=Y�4�M�+=��@ �F��U�L4���h�0�?���s��5�B��]R��YKL��7o>�򟮴(2F�E
&*��;���*���QJ-;y4V�+��M^�T6��j�>����e9w�t��?'�o������sPb�e�e�ܺ(�ь4[f�{�.p8�fy�&X*�X��j+I�,�=�����+�c����#�2.�WL�(��CI�d�%ҩ�����
�����8G�aL�͑�/�s7vBv'4w�2��D�ҕi�S��I���h��p0p�_�}��Tk���\����s2�������0n��~1�`��=�bū1�(Jy������Ÿ�Bb�U�l�i"�֯��QKNihXВ�6�� ̻S�*\ ���H$�I!GV���c^}0i�{كn��#�'ϋl̉6�,�q��٨Լf�v�}3�D��T ҅'-�"�CMS�dPں%I��)���P�v���@��{�^5�q��������/��X�#}ù*N�W��dx{+����2�n4�:�%��D�Hݩ�5�h
�I�_��L�I�kH��V�>!�{C%d��?a���˔���Sg�;;��ix[����!R����P3s<�/C���9B4�X���������T���%p�m��U���T�v�2��2Y����}t�&@��FY��H��:�\2.5M�������&+�+�e4s{$����&P���
1IfsP@f����烰
���M�C{:Z�mL��é��m$�LJ
���i�9׉hI�ݳ[1{� �8*L?Ŗ�O\�����>y���NV&�����r LU��rb�|w�1�$0S���sz��4Ȥ�f����%[��B�x;C �x���޺��쳬�w��pB#�h�G����M��L ͹L�꼉�����ǎ�D)<U`��#�v=�1A�o[
h_�^s���\�2hy)���ZL�s����E`hO~:�u��������;}�= L34o���zS��%"txs�/)���� �V���G�N �|����d����{6_/��֚��"��v��j�}]n��Sн�d[f8��j~[�4���x>���1��Q��'�l�7�?�G��ۗ�Լ��4��bk+e�)O��'#p�!�is����ppyYK���a�L{λb�S�fk�wVpm�8}��W O�Z�9�e4��N��̠0H���b�b"�<0��D$����OV:H�<�n�7�'�*�/�FOTB��Pb#�%\���L��XI  :�4g��ŧ�~�j�]C����z$-/7���I�j~����e�%�HwN|+�H߱.}mp���w�K�%��CUW��<JNH���-��T�1\���Y���0�Ϗ�ϲ�G����!���?ҧ������6�d(a4tt-t?֮;rw��a��Z�N�is��/W&�c�f�r�;�Fe�;p�m���e���
���2�+2dUw�|\�dH2��2�N�Q�w����)xs��$�~�x��N~؋�A!��V�cҥ��QH�,4k*[���"�Mt{D2�0��*~�˥$��D��H�t���@��Ỿë�<�E����������m��E.ȡ���@m*���aMI���Fħ4p]z`����8!�c`���i��[	"���҇�W[)0�p��?��^V�F���{UP� �6R߆��V{�Q_n�B8�.�z~�:�0��^j��Nuk�C��1κV^4�	sbq_�/0b�$�s��F7c��9(�Q��Z�	�=Ǫ]X�&kA�I$�O��i���6!n$���4��1g	�Aپn�t|��炪GS�q*�qQk4�^�[�n�_qZxu罼GM(uPVS$�Ip�8�DӪ��&Ob�Ǣ���Rn�@�hpJ*䇾\T�pY�1<��i3[�1���أ;����c������@A\!/W���92^��O�.;�mђNR➙"���uQ_O�@6xi�}Z]���:�����s���^uF���Q䙎W	�/6X�@wq�y����^�|+WE<j��;�(�
�7�{��Z%z���Kg3��0��aS�$�bq�q�M�H\#b!D�ͅ�q�60�(�t*JP,����Tk��Z���ŷ^��~��׆���D�h���w~P�w'��T_CS�ש���N��$�����Wp
F O��D��@[O?m���Z��ް(�W;�	t���_��k��2t$�B�Y�+PܷiXtI�n�]N����CF��ʮH������/���r��<S���E�p����g��9;��>:i�@��̣�Q�}�"8���ywjPl�\���uM?,����P��F��R��f�r�W�-�^�[n�f���
�)spR��mTg�Z_0*,��|�P+&fǐ]���p�.}�m�����p]�v�
=#o�|d���)1ѣl�`�0�K���X���o����!>��G����~�<�JV�)���Ӹ儭wF:!�� ���?շ�MD��G�`���.���B�"O�~8~m&�F�D����J�я.�G�C�ep�4�Q����٘�mcX�fov-[I�ؗ��au}����vV�LOH�6A�g^s�K�Զ3-U�֧�e������\��]�$uST��m?ye��~b�T�F�uz��/�6\��.���~YJ��r��$��R��@��f�k��/��6��U����	(��h�?+,:���v
2Ϭn6f�}k��a!�CtM��u��f���՘� �eE%a�}+
��0[�ۆсO����g��'b���i=e��״��T_��G�N�4:04�P���o]ק^�ٸ�/ofU������li�}V���$dN�&M%[o1oجx�`5S@o�,����ypPQ������Z��pS)���oG�� q�Pgw�3�D�uԧ]�1`�怹H�]��!�u�ޚ����	��w�4�I�����1x�(�0k� Z^e�s�hp%�������9�p�u��S���K�V��b�A��%q���C�W��sKk>���O��:/.b��)?k\��Xamq�`��~J{� 8}i�.�ފ��r_��2�NV*9��l��7�T'�̊Uް�a���Dp�x�m�=?�O�U%�Z݈�çMl���A�w����+>r��/��C��� �r$wrי�1CO���YH�6Ti�:D�a��#A1YJ5$����֋X���]����}ס�Ђ|=8]�Y	�u�V%ϐ6��,�;;�@�^��ؑ��19��fa o�FC�����]�#�Y���ė�M���8Uq[���R�e\�l�ft���t���@�}�t���޵�p�u�/�ѭyc,�(Ƞ��}�<&��	�q��+H��v�,\�pY�MWD]���'��ŏ!�����X�d��$�o���P� ��c��쥊��%�)��ٰa���uo��	S��8�q�U����u]i�]<�.�W�$����;�v�׭B�YW$�|�q�7"�9���h\rn�'����"�wMl�Q6�VNމ�Ir��u[�L�ɕ;A?�@l����,�8��.�@�@�v��w�X�yg4>ES�~�Ȩ٬���!$m�$�܎�̺~[!�{��Ol��hi����@�{����ڭ�\�;�O�,"��R��~��
%o��naR�߯���jHJmw�ץ�Y[d�%�D��H���Z	�%��8��֕�܋��XJ��H�n�8�N�b�8 2�~�g+hHww�g�^ F���S�I>�6'-��A�](SѬ:2`�%4��"5�ƅX��z�����Z�F D��jkv����M����F���"3��H�:o��d���h�!;�?�H�416�_W5�Ii�$�c'|n'�p&إ�1�Ԣ0��E��Ǒ�Qp�� ;�^��J�tX#�	v�y�܍7����J���T�a44����:�a�\�0}|���?���9E�C�";�)��&�f�>{�pm K`��t@a�M�틮�3{Ω�W�D�F�LgPjy^���sd�[�~&�	O��4��au�js��k�hT�m3� ��Y ��[(C&��r�
[FT 'KNu���ʒ#�p#��r�zA�B�K�šr+���sُ�"x��P47Ú�����'h�_�o=�?nV����Il�I�8�@��L~���hhQO#����?E�f��h$���� ^��9.������#B�J�ߥKN���d	p:���~uG��C���a6�RI�6����K�#&]0�}��z�f���Q�K�D�?����;�鑘9a�*I���].�)���n��AAJS��.�N"ؒ����J*6[Z�E�*f���05 �2瓯mvl�/���#q; OcI�o-SδȔ��A�[��0�?Q�<�dpV�W)���]9I�>��_�'7d�� �D�p�Z�;��=���o8��w�V���r:HJ�ӧ=o�HuA����E���H&Ox6c,ØHx'Ug���c#ّ*}!uH�^C|S��	'���6�|�����O��>��f��C��[�J�-��\�=�3*��~�v��lY�D��@܂���s�j�o_-<�i/���z���h�?�l�{�O�u��n�qA+p�<��K���dů}}�k쑍�In�o��(��j�(IgY��'��Q����ed~`�c ���]��P ���+��D
Ү5�km��� b�1�l�Ձ���2������v�O �/���6�?=H��ܬ%?���lӱ��y�C��=�'�m��c%맾�Z#'���Λ9e؟R�/�gB%Ƌ"��c?3������KЫ��q(?��ח�7�����m�ڗ���ᦨ��"��EMK��$]Ik&����bY��o��DѮr��h�
>���n�����
�;����E�[:��'Q������Ͼ��2����"6&��r�,���V���ܲf�%0�=:p��zD$��/$����2b�L�?���|����.S�����V� ���3O��ȍ���8�Xc�����u�0g8q���������У�qg��{t�zoS�N	��p�Ű��Y))�\۩`g�u�#Z�����3J��	dB`�?W|�e��?�f��Ҍ<P3if����옌=9_�gL�(x�tW@m'4��O�eQ0Q~�s).��	G@"�7W��^��{�O�[��`��o1y�tKy�F���b�]���g���y�����3w�|1�r0��t��%(8mm/6�L��9:Z#^X���<�|*�s+jf�3�&Y�:9�zޢ��MJUNl�������V�����!���M���l<"	.<_�9�ȫ�u�"tlv�{V�!�)p%fE�b�P���"�̈X�H����m����7��/sX��̌����E2�P3��gp�k�%��sJ�s�@�>�������E�:�MPF�g�m�~��^�Ј��AS���!��d٘� �=��s[h�J1�&o���װ��:��ݎJ���oww�1{������)��/�V���l��ԩ ���tn�>"D �@��[W>��'��3/m�;�_����dp^qW�7��(�b�´�ģ�\��~�l�3�&�m����&# �BN.ɳm��^�n@IaNXx��E^��cc(<��|1Z�!�-��2?�F��^s�,����1^�i��4�׶���h��b`޷����q%7a�XzA���ߛH|Z�e����U��x,��֌�qO�a�������=	�������	Kί#��Z�J�l؍�C�T��x�b$�wt�o��W����L΍�_7t�P��S'��Y)/= �B��i����bN��d�ƍ����R���T	�����N���I�c�m�D��h�։�l;�F�>nY3�	���ӗ���@"yʊ5�G46�4��m���nM���T"�.�-<ń�2��0�8$#v0�N@�q�H�G���K����7neK!H�*�����6��8I�"�� h5���`ٹ�|��F����s'd��)F�J{)�Fw��-a�B�Xvu�xpCu���'�Q�r�	���')����к;O2�ݝ_�E0��RТ^/�S�$��+�$����#�.�C�����edLM^�%�8;bV���0��So�o���A&^9NA�hb�!̝s>X�ܰ�6���;�:��}�ճ������R�b7�Pќ����]�?~"�kj�pG��OAh�Y��F|EZp�!����LM:!Hb�B�Q����'����X��$��L3���) �3q���n�OS0v����i�o�&B�8��eA��6�$�Vjx#��[9��h�$F�[�Fhk�b��8F+�KMa�����Ӽ�=�<ȴt�v*b6�$+^tx�N>wz���i,�՟�Qbʍ�~��>3���q�,���q�/"n�������}���g�E���]��F��Cm�5��2D��g$�&�)G_W��/�b�4�Kؒ�&wU*yY���r��+;�_��{~{
s��W���}��0�@B+�P(�:&�+Vh*�=���n��.#��"�������m�n��mvz�)_��_u7āѱ���$ҝ���^IG�o:Yu��}��~%�v��%�e�5`U]g�5�4�!���)�?�.d�C���nj#<��<c�r@ ������2�Q LQ��,`rC�N[�i@Q7ދ���O�j0\��s^?LT��H�L�8ã��ā|eTA��Xd�M�m����Xn	�XSȅ,���M��)DrE��\�X%m�v���I��Ymk,Im-Kv2��P{o�2�<cI�����k�#��x��B�0[�e�ϣ��<�p²:V��L
2!�{^��|�"^P�:�5w���Dm]�C�]�'��%fK�>P٣�M�ʽb�Stl"{���j��}�/���� _`+�lU�U��5	�,�1}��t9�0F'��@���Z}�Hi����r�-��<}�O�z���<_d��^��b9�������1d��5z��Or��%���Z��2���	��j�Iue;�������� �7�P��XR���BS�����oʽ*7�$Sm����U/��Q�^���b��:z�žk��4�̅��T��&gQ92�%Z�俕���4���|#�Ood;��'w��9I��;L���8
u.>'��1;�\XeQ.,���f�2t�7tfɾ������s�b/�[7G�E�Mx˜rM=�^��rl��ME����d�Нx�Q��:��%���g7K	�Q-�.,?��CO%:���*$o*r#b1�I�����(�/�)9k��S}��0l��1�m���.̨g^�d����p����C�q$w�T����Sʙ��쯪R�~�c�{�5sw˛_Z�?dx�Ph%S̺������F
O�u�݋Ê̘�n�3G���K���t�{�cU�B��^]�q�d��Wm �)� BV�R�����Y��x1��\%p���R�3�@��:r�i��Ԯ,��=��$�غ_P,��7�0�#bi}Mk�i	����/��=�DcP�p(�jؖ��`IW�B�	_��mk�>l��XG�Z��W�W'K���<B��ٽ��� ���%>�p���T��\�?a>���(����7�ѱJ/�GG�o� 1N ��"�u�X�Şk���2�>`�JԔ���?A��	��vE�	�༏�R_�b3Czq��%bG�4�;��sE?qyN/��2����=0v����|�6`)۫�g���lb��H���v�}K��̹��m�JӴ�HG��h��������\f�EoW^���$j$[�X���������v��S�,p�2so0���tN�#E<2�M>�J{-�"���=ZP�υJ�&��-'"�w�JT�Օ����6H55�j�Úsj˦,�
3'T��~�+@!�^L�ls��Hx%���`L�f;�M2�&�)�~ >w�ʖ4;�
i�N]��8+��Q9��w.�/T<讝s�`�E0����Ce�bq˭��p{�Ye���յ�i�q���8,��^j�F�%\��z�Nl�K�{Ƨ�� ��W�T��N���OL� �@D��]N
.���¡g�����58"������"\�JI��l�"P��(��8Ϗ�m��а�5]w��,Ḕ%�n�/	1+.�u�)����������^M�����_H����
5;�ˈ���7��`J�5�A����f�Cfl[�	�&
��:�$�G�~dZ��@Z��g\��K�\d��@��QV k�y�wbMކ���4�iM�?n5�nr��+4��%��0�Si|��������)��ȴ�
��W M�2�ƥ��;4k*��`Lԅ�P�캱�ɿ0��y�P|׮��U3I�JB�G�����%`�pmo��&h��g�u/���� ���8��mUG����XP&+0��-��^��ɛy�nC�B.��~?���4}%�����ۦ"��lƄy�������/$��ܕ	mGB�<�����7s~��������J��g\2!�
FN�f����$R��� 9�x�h�v���~���0
�V�9���x}X���|^{s�:���O�l��ʯ��P;[�8�(�d�*�+i�U���J0b�P��x��p�擷�/�vΚ<�F���)
��yi^,e�$�wWa�e/bJ0_]�9����ј�<4��E�G��H�>�J��Ť�b�o^�\čs��]_��j��/0��7�:,eo�R����@����$!^�ڤ�f��2t�Ue�e͙��A_��
��!.�_6��E»�QGv�D�����k	��/�;w:�x|:�v8dU�v�L]QRk{&`7�[��Z�6�b��-򽠡܌c,z�:)F:�H�ʏ��`�}*���|�?L$��!���v�t�~f3lv��@&6���ۭX�Թj��P������][BCd�P���j�����Tj�4p;�g*��zu�\�"@@ۓ�z�]��b�S_�(#�<;�ub�zB�A���n�$##�.� �.�V�A�ű)	L���y�\�D�^By�����]�jP"�?w��jQ�٧�|�����*��h'��t ���>�4��T�z�×�#S�>�����=�M�8�K
j���a��iR�Yڟ���M���'4���ʯ"���*GN�~(A#h2~~ف�����H	��k�-
^�@P� @�PQ2
����a���a�j��;:9���(׉�Ցx [i`�puN��i;}�d $��������w��$dB4.��R�x���B�� �8͊7�3��*�?�u��Į�� 13)nX�M�C�ϩn;�)��P��"마-4�-�b��Ќ�25|����o�{�F�?k6cDOf�_�)��4��.�I�%�������|���1MG[��Ȧ�SO�ItB������R�i�_ ��L�!�ǻn��Ve���h��ڜ����b^D�ENYw�p#C������E����o �0ʟ=1�e��\�4&�*"�Ӷ7V.���Z��_mق'ڥ8_�0w}�uM��^�	¤���z�6�5W���M�,o���<��h��{ߩJ���ˊ<X&��,�Ⰳ��Y4��r%����gYgU���VE�17��U�5���Ўn��m����%v�,�$C�a�E|��}������$���9�.D���~��L����~/~e��u�vF�/� �a!��]�P	.vM?��F�]�E�) �U�s�d8����P:��+�����\�|�{4l2I4�A��}���G��ς\�)�{1����$�=&JhK-8u����J�ؠ/ih�͛
�c�΁ä*� ��Aս���:�ux]��`��8�O0�K�a���*{@�u�nW^0Һ�N�x����gK�S�$W}0�	�aQ\Ui�5��jSׂ�l��bH�}�����c�N����5��<M��1�i���`�W�Q�w1��rb:�w	T�_���^��P=�/' ���B1m�t��p[*6���v����"�(jAM��12�e �ɬP{�D|�,
�� EE�X��1W~U�Ze ��� 4��۱~��M���e��l&YO��A�����0��B?44o꧚-��?��~��y�QSJ�R1̖^�����(�<������}t%��`�}�7mo��3�`�4�[����u�l�x�ͤ�����J��t����%�����)�� ��';�
w��[�P%�D��oI�f����
|(�>Zaʟ7"�H)�U�+��U�|[��n|33d�P�Y�5��U��Ib����W�!0��z�Y���G��:J�wx��|"�&��b �7
-�dǽ4 �1>~�ݝD�#���/N'ݧM2�qU�M����K9U��x,�@s�E�sA���j�i�me8J��t=��]��k��Q:�x	x��3鷷�I�9J׳�s�U@���g��A�#Mrs�R�t.�����A˱������I)4L�<5�k�XTe��x��d8��B\��[���'��N���Hx�:�	��q�l�z\E� ��:G��2�M#a�?d_�G>�E[�NY	-~�{� {�3�B����%��qo�<+��Sa���Fo����p�c���ڤ�&�8q���ӯ�:�,�vM�CukŹ�ZE��16�O.�0�����6Ǩ/�U�#t6��m�A���
���hK���udU��d���1�Z����N�z��(�Y��n��M�~�#�O���%�<�
��ū(�s!��ґJ�[�Ƶ>0���c)�����ШM�q��1M�,E��Oak��̋귴".�S�����S9�e���@O.�;u�m=Mm�5G�>�_�����������ͣ�k�L��J��N��)p����Kmc (:�=��qe������	E9�椶f��^�u)�ߙ��s`�	�Au:�N�+��y�J3^��ɠ��m��@�,��}�ٝO��\V�t��d��AxfcBF}�����E/��r8�6}�C�D��gE"�_�K��Ί�����z*���Җ!

p�<N��/����W�h�>r�ֳ�4�F�(T CSbק��86��ڧ�"�8S��2�?��`?s\�D�����a��6�q-G��p��&mL��]	C�m��T?���|t�gb����ϔ�� ��F�"�B����ǧ��P�QJl+*/�H��:	:�=�$�\0wÒt�'���uN�T�e���V<�D�q*�a
\ۗ fg��>��<�Pm5��u�����!���
�Nw<H̄�._�a��fj$��ui�{�ڜ�߸�@�	Yj� ���=�����[y�A�"C�{$Z�cd��s���BF��d;�qdB,)%1��x}��p��I� ��ڵ|��O�x"!L�(ӗ��)��<�#���#~������xڶ,���S�n��7�j���PN�x���ie[�;NN`v��J�	9E����� z󸢧>����~��,��{@H=`9�5���b�k�����E������FPƫ��2�aͅ�&��Bi� ���p:u-9bR��58M�_q�.�mf���Uk��?��4&G l�`�K�1�X���p�~�hi?A�����
�^Ju��[y=\N�5���Y@�cJ�fL�M�+�X`�x�� }����	s�τ�G&�uUQ����#�jz��G�W.���^��C���F|-�5��ݧ})Ϊ6�9����"�/po�$_��P� :'HL�<��2?1�P7{y�� �"����"�%�XOq��C@A���&&7�<��<�]����|@��&Kc�:�6���>w����������·ĭ�7�=��' �_�Ez�iG��~f
�#������NW�M�A��"�Yo���k�C�Ī\s%��ST�m���x�FZ��+7�#1φ����}�法΃�3����V0a�?� D�ځp���n�aݖ���ؖ�	�:O�:j:����<
@������Wň�?���$:4}�5����`6���v�1!!�����>��km�#}�`@(�PY_}e������v��`P���lAWf�X��44_1��TW�;Ƌ���;��0%��.j��qH�a$�~��]�5L<����]E3�Q����"u�?'h�x<wL�.(l��>AV�R'bd���ce��>�oX/K�-�h�L�]􋉣����Oٻ/��Ç���B�����s�}
�����;�wC�']"�@�T��|hJ�1ES�vʌ?+r��Lz�ŏ
m�&HXCq�h���b���Z+j�"��H����!?Y"t�ʒtU+�F�#1�\T���-�ŻX;�=�,�5J<���2ۄ��	9�z��&#{|��dA��}w�a^i�lwV��(p ֝�/X㶷���Kf��ƻ,D��e�G�G�I��Z����Ջ}��u�m�:���3�Ăn�d�2�4�c��h�y��kT��kVp@?4�����u�Ϫ^'܈�X&�5+�L?��l	W�jr���wWYUR:aER�u�D����ݳ�o���h1j\��X��!�񩚃S(�2�𖴂�r��C�኏���!P����3��o�Yh�w����h��2�+�n�5�7�
S>���@=!���܏!��;$��s���oz��:�[�HE��G�Ƀ<ءyQ9 �l�]J�M��2��e�v�`�m�* ��ε��2DT�x�ŝ>��9~V)���I�F�.5�`�=��L�]�L�]p�]��ԅ"ˑ�Fn8��N��E�'�Jn"���+�ü1I
xA�����2ѫaP��Lv�� �u@]��n��{AȨ�{�s]��㋑����+(��q*�0ѩPC���ca�{�\���f�.�,��ّin�h#N��Xr�q���;���¯Qe!X龞��5�&A�{e�st=7��I��\&�0\�0���<
\�oAsA����H�mtMs�U���
8�����
��o��t�?� ,��d��s���~��xz��0��ӂ��q6�25M�t�×+{��t��\AqUP�79��R�8�����_mB���6�V��{�ݔ��v�\��:�2�K/��E��W�������:I
/������ �\�W�/���T?J'�h֒K�V�LP���ҍ��:���">�W����]�/�9�@�Bk�h�	p�R�+-\3�Z���e�t�},��O�$4���}1_�r.B?������pZ�Β���Ru<����>V��D�uk���!�S��}0�6b�Пȑ� ^S�-��^t���tr���L+N�5�jy��i�D�N����h]/��˕�C���ؓY��PC�-эD�Ve�b����u%����qP�l9���>
�YTm9�=�vW��/&��"�3dk��=�ET�x�V�wv<	b�[��W�$�F�����r-��^_+\���ȱQ�(�1���G�[+�~l����~��K��ar	�|%�QQ,��e��_� Ӹ����j�eIo�̈́��B��q�%����t���wi�9�b�ou&j����I0A�2����q�����ٸ�Ύ��=ɮ'���S�%>���J	o!B���`�P���~+��-�$k"z�}i1��V�PC�������6k�ߍbC�����/���6���&��������_�}.9w3�Y�P�~�͍X�����P�0��#�a)�H���fw =Ț��~��Q�L�I�r�K5>�����|��P2b&�1�*��(��p'eE�(���l��2₌il�Z�}��*�]��sgы�a�)�S?젮A��|��>�����G�9V^fC�t�Π�埯Ҫ1\Y�q���!&�q��Z�o	D�4�0�6�$q���c�B:�.;C�##��0���'�mI��D=�Uc�5�<�Q}���5�\�e�ĎX�X��d����ք�o�x����qM��Ce�Fhk|Zi5���Ga����������dUI<���@>TmE	� f��M6-������{=�-j�C1k m�XD�5c�"��Uw8��l�S��}ߩŊ�0C�}��vd,r;de��A6�B�@x��S��<��w�*	W?�º/��d�pE�底6R;�|qKu���p,�Z�!W��$ ��C�ѓ!��@c�,Dx�GE�L���s�r�ʍ��d*fk2��5�A�N�%T�T��Ϟ ��5s��h���H���v$��n5�k�g��k�����u耖�!�r�1���0��!�ԲT��u������1(3�!�6q��i�T�pn����`c�z%�.Ӱ#��