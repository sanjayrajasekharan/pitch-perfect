��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����I�w��/���8!(K�/�HC���=�ΰ��F'\�ޭ�j%�Y���AsD?<S���R�Z���S�eI�B�\�pŋ���?��h��b�k�<|�/:m��h�yJD�(΢q��B�]w�{ <?��Zj=sv�7�Z8>/�l���T3eRiB%�����x�tW+���T.�ɴ�>lk���8������E0^�9�e���ek�{6�(�i��P��Y�>�֙�KHm��ŉ�%�X�ڟM���~��շ,l�T�Ӟ^�n�0c�.�������b.8��A�Ir�g��y`z�3�7��0� �[��أ��an������o�о�g?{t������o��Fz�ǋ=g�s�q�.wτ��=�r��rIO��Uj�S���z�*%2��є�D0�q&O���jk�8�]̈́L�E�S��/���4���#.�V��;�q4t: �@E�cn��z��E����ً��U�_�Qe��5
�RpK�Q|�M���^N8��ؓ�ݑ���Rs��T
d��'��Z6���hL���"{�4Fq�_z:��].i��Y���+)3� ��ne�+.�Ձ�������p����P��@�h�F\�ղ@%�sL�h	q��el%[F�}���Rʖ	��=�|��
�Q~�Æ�͠W2�b�3�WȖ)>�y���5�=����+s���b���\��4�X�`�NJ��*�x
�E�[�������exڗ��%����3�*��;T@}R|��x�ۿ���!a���?�����I0c��ή���&���u]OtXRsh�W��5V?Fi�&�^㲘�1�冉M�;zs=�f��UD���oLs�F�b�S��O���{GEE�Ä�ӯu���gLP7�NE�����^(�����(�R��	p|Z�S�k��ʚ<+%;��F�MQ�X6i���F��Ɲ7�H��6�iy�XG;C
ل^o�
����B��Fe�ߑDS%Y�~ٗ��&����8����Ȼ�6@�y���Z��¡O�M��(�e��Gd��'�+�y��s'mt�V8�n�<ǤK�J,}�d{�'b(9J쾷���|~�*�رv��� U������r��tR��JЇ��|�m�w���@:[��[uV9ޅKZ���h��X;�w0���[�:`�-��#��U�I��D~��)V���m��	��$�w�*+6��	�q�o�����bL�������g��\U��kH����C�x/��X4�]hQ����p�0�����x51�G}���E��a��JL�;�J2ip([i����XH��t�:�����gMμ(:�`@crlU�-5��pz�ͮ��o��ܸK��䈞ŁsUI�� ��s�"��*=�C��S�d�Um�	f6cB(�I��#�R�Y�)�h��h�a^� �Ʋ����}`���N�ԙ�SO4���]�"�#51#T�H��"Ũ�ᜏ��F�D�v�������n��bOB�W�|��k��*M�iO�`@e�"��VfR*�͞{Ј�D�<
��nߓ̀�QW��t�v����u7�K��BE���kV�X>D&�ʘ^Rp���$\�$W���&�����mק¤�5�u�p�1}�,Hl���ͱ�mi&w�..�@�kAA�o�7��D�kǣԎ���x�2�w����	�v�6���/��m\E��(����i>�@�u�}u�o'V=��bF�v"?<t1�nĖWy|�܄����2��e�d�:�(]]<&0d��Z�}Y�6�Y4s�+g��"�n���V%iR�U2��#���}�,�m�My��*N����v?ʕ�R�^�~�H/c;�^��/�g+�=^*,�eU&�njm���`B@��j$��Eow�P4�a6��!��2�@��)���f $K�A�9'�5rT���ۑB�P�DhP�|2����K��K_�:����u�O�4҈N�p�O�љt(�x���zI� ����uy�)�|p�	��>�X�0�A����I8�n�@��c���Q9O�6��Ih�!�r�M�2v��[���	�G@�\ާ�Lu�!I,�堑	��@�"4$t���w�y{!����e����� ��?�hgДR}�_-���z�S+��P�:�Yz��51�<QW�bć��عv��kZ7���`�'�;�%�ބ����-�V"^�-���d�P�^C������
����Cl
у�JI�����{��l�� z�ƍ��H��7�:�]��m��s���U�ѓ�PPL���i��������]��Ӿ�i����Z@r�aR մ�J	��)�4��<P�6{��]�~���St��X\���8���C�dGu�9O���	=���9o�=�± ��$Eĭo�;
S�j�!9�Yti�{Ԛk3J��C-��M�{t��H�MG�7�����\)��)���UZ�XK8����yhs%Eu��тO����bLْZ �זߺ���|�y�y������q�_��W6��huI�W��L�Uvq�.��Tҥ��^��W?���S����8��M1*.y\��:��I��]d�P&�@";����w�u$������"��M���W�G�����YDB	�F�50N��e�>[e��r믡���-y2=�{�֦�+����=S�����W`��/4��A�~.�r�����D��Ü�b���s��5&J��Hv��o6>�T�g�6��~[E�kk�j���2�)�]��͋��ǃ������;y�Z[�N��)f��J�Z�05�f��w��옱>ْltQ)��>-�t���o�l�"C�v��2��4�����T���C���;�{�78㚛R��V������^k71�x�|[�=R����=C�Aⳟ@�i��o}2�҇�f1��D�>]$/�����C4��?z;��ߴ�4�`"%9�2l� ��[��ֳ�_5��Rĵ�,�vܱ�2��q�5�l�
��`��3>,R���9�4�㼍x���[ь��>�X ��c�%}֔9���;YyT�6����ѓ���eT��M�YL]��t�iP�2��n�t�1�bi}*9GFE�2��ܮ�
���{�'�
T,���6�zd2UeosWl+I�$�0&�(��U�5M��0�h\zh����<i9�)�CC�̾�d%Mg��T�ȬJf�J'ARe���9��^�׾���*+굾���AEv�V�0���DK���=W�F��=(�� R�6吇�b\��he��vȅ�Jyv.,���"hA�A]�߽g������dӵ�spB�o	����u�5����CD�Js"W<�61.�<ڵ�~�u�7��
���{Ƥ�h�*�ﹴBյ9�`��s~���
���{�E���T��V~�1��_+�iSW6�`�X�̂�{�^��bw�?)EA@�\#�2(�O�	��)��P�Hx5�i�M()C�����{,��j�Q�p�8�ůlЇ�Bu���\S�,�|p(�a���s�ל�p�e���~���wJZI���;���fQY� ��/�띯�IB�F�0Ǜz9m����&qW�ܣ��e#��j7u&���&��NS�LY+z�oW�hP֊k���&������ԟgC.ܚ��N�Uō:�ۛ��R�6@ES��O��	�K|��$���w¿�(`*%䶼'9�q�4���g�P>�_��/�����1)�I�w��BL��!�56Q�Ǜ��d�2d"�w�QC�t�§8eF�?cWe��|l[�,ڢ�~G�闧aϫĲ�v��Ux"����^�uyimvS\�#������uǿ�ٓ���G��X�y��6��n�!T�߭���/t,��+��=����0��(����q*�A�&k���K
�2������;?>���i���\�Z����.�1�/�:�4Z�U�����'���0��ټ
Vb_��T���mP'^,��TX��x]!��bYW�����ꩥΥ�Fq�oI�-D,���9��$�_e?�<d@����I�}X&�Y������r�yh8��k�;N�Rz��}r�}���UU&�(k>S#������'�&> ,��������>������l#l�x���o���L�FF<���"r��"�8�t1_�P�zb��&�*��f��H�ϋ������Zy��zE�u�˽m���۔+��s�B~ ��F�tk�\����~m�T�z�����e�lNyo�(�X���J ��3,N��8Ƹ3��1�{����8� �Ô^ �?Z�RE�OL��Op�7#��;Y�Ճ����kk���	����q��S����a����&�=6ޟ�_JIt��޹�4���m8B�P%�88>dI�Íi�`n�}��n9��XG�����u6"Y�����yD�P��K���+���mb]�v*+�����w��tLxƠ�@��� �D�D���n����/�p+�2[;�ğ&J���wJ?4j��J�od9��L�LMq
��l��=��JP4�~���B�]j`BCγQ���y���%`ë�u�.��!���R Rvf9��`J�~țO�*�g�Xy�3�s�dJ�'A���钹謹D;*P����	@B$n�����E����b��?�c��B&���jdU)D�bɥa�r�"`��ratݱ0�N���I�J$�E�Y��RB���RZ;����ۨ�7`D[el ��,�WX
���>�E�`%|b���;��&����R�"C!��N1�^��`@H���ظf3ς~����L�w��乩��?oJ���g�5�����8L��@8�a��~�h�c��w����D��6�$��m�{��C~V(N<Y�������q�o[Q�-��7�	قR�CO��x�*IfJ�S�]e1/Mg��31�㯆;�Q� P2G���d�3�b&��X��T�����T��a�P.��b3b����f�k�h�<��I�b�|.֩�YF�v]~�����R�P��PS&%q��A
������{%��@z+#���U�$U>�?��}Ch��L�<�[��gq2�[C�2М���P��+��ܤ=�*����f���G�o�qe�M��R�E�&�3���"����_s�
����Z�d]~��CE<r�K7�D}����sz��u��&���%����:�3l�ڋ`�Øۣ�?2�|�w�����ۙ�vkPV�!BZ����H�����&�+[�eFn�ō�|��޽��˛ z�)
���	��α���\�\.X�����t�pO���]�Zg�J��D$�-%U|#���-�sst�CR0а��݌#�t2.R<��v�g�]��R�C��|�Y ���{:����/t�q���v�3�v4	I�г��ͻ.#�����η6��F�����wnG�:��/���m�4C��&WۍK	��%��J�|8A�n��W�'��H��d
*QÍ�^��NC��l����.I�7��ToE|m�gP��h�=}�N�6TF	���8f��6��<Z%�{6��� =^vki���!���C���p7�g�Xv��+:���95�6��`�:�1W��'���w��z+�x��{�(�3�梞a�����bo�p�Be��D^Us�l���3��J��L���O�;߈�\k��Y{\c�����
�Gt���s�hs�6~�_�K�����dn$q�d%$Ʃm����?�0�TD�}]9�������0*S��/���+G�\ԲL��$���(T�٧��d�q9��M�nSWۜT�Y�oe���ݑ^B͌���5`@/d!��$ޛ��%uQ��(q �O�MG����׆�(��ᓊ���5�ƽg�S���^�ų��֢~m��"݊|���KY�6Y����aEG�whŗ�m���h]1�xP����\��6���p�qr����%R!��-b�>_3sԃ��ܖ�p��4��^��B���Q�2e�SU}�kvtوJ��3����Y��G�.�孾�墵(��RVs'�	�i�@ ;��U8�E���꽃�E�7(�݁��xe�	� &��ሇ��{�@7� 4�2C*�b]��T����S1���C�m��u��(���C����;%��!�e�E	��m�G1˵�NGwO0��ID��/NP6����7�+!���')��2\�_�g� �_�9�� s���s�r�bH�);�]��\����}c�,���k��cL�i�.�iŪ���ʡ�@d�v+����w�$��� 	����>�s�u��r�6k��O��T8Ƞ lF��^�;�d��W�Bj>8H�
��*y�uB�{���7!E��oYU\kX>c���4T���@zPg#jK��}Oፘ��He׌���;`���3ܴ�Y蟢�G2̤�75�dMh��5�pP&�������������*��5�/��i\W���TE�����7ټ`��N�T4ɸ|��2 ���?��H��{(=g�k��L�����L;�L;��Ӂ��U��s5!L=�[(��蕀�B����4@r7H�T$͑�?a���x�I����4��P�����	��|�z����a��sQ�=y��^I�F���_�^H�Wz�?�
� �9_3�\)�oV>����ٰ%o���W-��z<��:΄S���ʖM0.=B�8�ެ�I�?ޝ�UI�$���������<�?�!�RK�̷�(�p6�����Ö��ft	І����1��=w�9���W�����������O��B Y"�:5,�T�x�1N�!�}�bh#�t�5I)��+�Iˌ��G�e�Pm��j]�̄ȫ$�1�/c���O@e��%F�h�)�O���6��9��gt�u��W(B��)z�"��<aZ�`!=`@��%M� W+�|��̿�4�
�K6e����I�9��_:��]�ʛ��8/}If�"�s���H�0"(d�\���%NL�S�{]2�f�� �P��g�/�"y��ى�7�U�/(�OT�,�UEQ��7��I�{�"���<.g���R��&��sC�G[&0�A#��7'QA���_|	���-���k��.��i���/Z�����^�V���d�_}�z���`5������_��8��DY��@�����H}�p��K�2�����Q@_��2b��2��`$��ű�