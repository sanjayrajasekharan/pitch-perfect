-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
jY1RmkZhI9noorLUIp0ECeoG/jwXSohavs9Z7UQ/4txqtKxKAnBHY6OMTNZULb9V
SdVqtPJTmhUPplWm6ib3Qz6K3O/r6qVW5X2xQlJykYujSPIuox98pGsnuk132d2b
wBHScE3+HcteV/OAoi/u3pTjaaUCBVV1riL5V4ydJ98=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9440)
`protect data_block
5O7s7gKf8+b2JvLkR4r9K3vX0xwvA/QjMMgCQjICkjUI4C/QFBHC9utN2rWwrIPo
mQz3f6qsE5giK+Ge4VZmv6n2sgJbzZvuChjPmzxiVzbrFXWtdyXphhOYDPF46G4x
Gi1tmxV4PFuvk3a9P1sdoHG/+dAyTtKtZK2te+kGNyag42Jjr/BLjH1KqueBc3/n
FbX6rZDziM0PnKvmNU27+EnB9hHdGnANpkPYvipUjZjQtT0MyuZeR4h5Urga0eE5
4GayeJd25SzZI8fB224C465Dd1hFHpaYjNVmizuHNZ2idr/3ijSAgu6/gcvh7bU8
1grzsZkNJE2/N5H9PT6IlfBvwvZH6uB9ZMpFeL1mvmmmelnR9DwQ9YtoNONs399d
iOnqYlMGMDcQ8fg5Jx2WXtHvixDhZ1wFbp6uhvB9A65Vh+OLIU6JFxmxhLkZn6lV
wwtwL8/n5A84wEXYcME6GNb9lAEiRF8k5tEvKwilYSyGe1M6+cGXbs5sYHllgn32
StY6akbRyqIVRTyIPQgGlcABz3QEyW/zZ7dum2vdBE2VV+By7gqLydFIU0U1D7oX
XkVfUjsNNycP1h5bVc7IOhFKrOH1h9mWD2H/jMWKaRLxauhD2gyRVat0r63UZmEm
t99AnJzuIC2AW1HVmuzay08EcvIcXDD7OAMFQUQrJkBTPYto9mKI5h+CG3qU9IyH
SApHtM8yYYURsD2LL8iRPS2ieeFmLpulHtBDaBqnZBSr0yBjsx8nlVEB1wwmNr5P
odIGh4IjYU5/uwjbxbnQgGJXZkqblDPuK3p3IcbcjaDJDDgVi59lKOu+4yhkjs9v
fBpVut8qzaF9tEP4IPAh0wkhLin+/niF3Ap5DRTpO+zWuyVE82HJTfeWEmBJvTIO
YlboYBzVrlcEo8+VRQa++TemvUhtJ23C0/cCtAGrFmLX4NAWKund9DPNNR1q/f99
rCZFTj6SGFVCmRZKiaRteIv7M5baClnROeJkL6kq1wL2sGNBn14qm+LJ5KBRl2Qj
X6ITntCiLZ2tHqI/y1bmsPFCJAzhmMw2Pr+HicTrRt4jYNo9d4F/C9ylRGLEJBHO
0dwq0Hox8NaCkmyiD7DOTCw/pMnCD1J6ubLits6tFob3G6Ja3ztUgFZ41S00QYwH
6u+d5YvNznYKDGvenHL50pj1MA/HhW6VHeXHklMcm/1DT+0zo36THK+u3CPwo69w
ocs04BJvBLUP2QO7yELVVZSrDhfryCbruViVu/pMIrcI4gpU5ewVEphdS+UnsDyc
SBcAMu/lwJAeGNha6gzq2O1TNhTxHN1OL2I8NY2dk5vUfMD3pDebVwIehX+KnLEZ
rou9ous5SruYXRhNU/DVFuNtxzYrbIEzRTPf2kWHqBTJGg/qAOjUmEpJLGo2ZnM3
IAG21wWHMSZEn+0EbuYla1y5P5hdT6YrWoKd08/XtbwcWbjHJrXNEj9c6OrTBgZB
x5l+3ur40Ba8gQcde+7sRuSFt7MJn8VSjWOP0RjQL5hZ75W89tmNmTrBeCEvou1O
7QpOURdUlAkDXeRHnBjct7TazVpoeWJqQy2ny4FsIjjmjdfP8RbmQcQ+Vzo/TYSQ
1jcU2QfihAhuZTeqpBi6dKw3Aj06cEdXeX2eSHNKLDhbd/wya8utDCKf8g3/wEZI
CpbsTcFzCNKIZp0h2k/cdKVQgT5H1qSXKKudfXPJgWYBY3/3SI5UCGy2E0404LEB
Z3xm8BTSZK372FfuVKaVNTeKbcJv8P/i6jlpW/t605bAcS4ap3IHMkd2ID96E/9E
KGjpBMhxv3qtRi5R6z6w/Hd8COjypdpds1v2V2j8naz7qs3HINp3e2o8XbM/hpLD
5Pm62MRb0cZBeZvETWpJnCc3RjOGw86nXYMPQDvJnmm4W0aUq0zfbkqYpSN6+7mX
GVBYU4klTf4YGKA3K8VVVaWVf98/+/ED87uybwRjAkqCj1MdAAbnsiFJifFJk2zY
acIZzqMw57Q1r+VkHSDHBLHdKB0bRdOHBtaLFif5yQ/bIAx2w9J24cSCNOibmvkO
8XbNUJBzz6N+otzPczisasWBwrqho4D2C/XCzOcnKJj9M2HS+TQpeIl7xGpaAGWc
ZugWWO5VfKYehaFPn+9FbyBPre/vlhkD1AOjFsGhJB8znf2zxviqW843iSNs70SC
BQSoP0zGvxD4N8gq79u6h0acuYJphWrpD26tJSPYAnwUOxhbSf/nz0kJQoKunLse
0TXM02L0AIjNPH52c+9FvfsEZ7vbpoA8xh5NTYOpTmT/tm849XMVth+Tiu/U4q9D
f6YpCrtZ0IpBIsZ6JQa/OclbAWJgbS0OSSJcCqde/nf/s5LhFHOYGyfmsKEpGkzf
2/ukz8dNIRMCbD9zv0RH8vZbxgcq85JhKDJLrL/zfRQFgO6A6BRUieXuP2Clu767
doEJfzGvROLDVZ7DIMtSUDBl4WH/swSGwF++ZOtCWdL4ZxtoYwRIgsFGvCXeCU7o
I1kuoev8VPAItbpq+x8UhUk+f8fRXCz9P29haz4WU2YHi/VWStUr1HxfwN2mG410
WYzsfBkxZ16iexpR6VE+9E+u30gV/HiGmM+KJAfuBT14Uy9SVEn2GEHnE0toNpKL
ypWGckO9oo4vdrF9hVzBcE3xTyMhlc0DURYB2T6qeWDxJqENBf8VnAl8amMjqfm2
jbwcWmepf83ucLnUUmZ/UtknwsJUCAI7Sq9anJcMvksGH4zM6EsKPqf0S0EN4ZVR
27IoKT86KsSqQyh6GF7KYobEzNl3sp76keoB0Td+Kxb3mX7kAeDG+oZfWSR/VmEG
6QNw4t2tGT+53UuMypov0YfSukL7I5i5Q95P2vr841g3fmFvSzhsmPz/uXmTAuHK
kWWPRnPvrOtkkjxs1WzJR5mgjkhFlh6WUOjIuX24qS2K1fBe6hSqunzQsJ6iYrkk
UIULW92CqH+mwDUvFfzWgdzMHSxNs6nDVNS3Tc2lVOH2rOaHvmTLFtTxVZ5/laWI
5NvbtGRxxWCwjgOdV67L2SM8S4c1VbYfWx3unANzgR7bXs8g0DoaEtIy2CPPkg26
hIgEkTX8Ym9bzm9QjnVJNKRWHxXDpZ/oPilbIQTPSuEhrxfvicLxzHoaXpFJ611k
AvcbRPHa67zAYw3LDuTBSY7TAkmzxNooxoHf9bmyXPara9suTerFyUdGDWuRtGr7
ooFiLLknO2/waHEqJmdf9txV4yY1vqGB13Bc0+E6MZi+gj2De/bZEoCBGioHcapO
dJVeGRP3uN2D+vP1OWxfy97kzVowzMwriP2Mje5RAPDI+W3thmF9gl+tsalAZd7O
KWqdrO+mIDydruBJj/j/y4eHCoZ6/F1GKm3fYUxBghCwLSaq273ugoGbALxLtxkS
gi4R9zHI0PBMB4NkCADdy2y8YYkz+/c+0AqHr/R7TQ9RJWmb6nZPHwZnrm+KKq35
/1GPWNGmwkyBqQcHfO6ly/NQWG3QMGlixCAgEtPZp+Enpx78c27cS4ni/EXHqQkT
lpnhQ4JHS9Ju9gyOHOQ6wsCpKJZl3JJtXkEG3hs3vRGLfVuIH2kq83na2h6TKPvf
5AbEAlh0G9OJYxq1ZbxwcAFWvGsXlidoiAK82kBZRG+dETQLF69GCn9i1Rut7vUa
z1b0XO0GuzxFGbXZbTe2JnGmnKoQAvgye5jJKPA2z46u5xdGZnphWAcQoLB6+r3z
rqwSxApXoZyjzpYUdT53+PjDfcDPBUWcINw/J380pLnfFH0yAwA3MfoNuOHS0WHv
uMoa5BbAhgmDY39rXYgXoOxX4VxcvpGQyvOejOZ+Q+yDEw1oM9HNhu40SiZgsi+E
weWr/q518hAOyzv/CDdHa5H6zDmtub70t/kwmE4r0zMmDmXQh0QE2OIj61rEIKYk
Ws6XF0T8059ya+WiD9kvxLLCnP54P1GxbuxDTjZmakIFgAU0yfmnVzJvS18P80WV
9lMMRXvRavIfje6YDtpdfCXAs18GhfE42R3z0JunUYKamCSM8ltXAPshYuvYStnd
k4RwZDQeaIqhEi8U4LIexFeUCd12YOXphN1T0MfesmFnVXy0ccD1xjBq2Py9iAnM
ujdLNssgkW/Um53SSJUO7RVGYvOpKQKOqfBivxQ84WT1NvEHHApFY9wOFOBAODPT
/ZuEWM+amtJ+Ff7EL7VFN4AegVPB/ulczePo+r50WEi0iNzxK2BvWxKgunsWqH8q
msRAwpAy9dGPpQaBgR4rlJC5uLGNvTTRzFVRjkfIGW7l3sSrtLE/3uFJ28js09gF
iTJZsth2oIw79Z1I13bbAyCXyrTM7JRrO9jgLamPASSdOSt9r8y44s2Wzee4Cp6q
8YHY0HXfnn7dm6P/Rd3nc93F258p7oFdVyRdZR9l0+BJkF/QPud4x+6ssGaj25Hw
AhL15SNNaCKTiLaGCudO1VJHgnCNBv7DK7Xt2XdpVg7sZXgDZiZIT0MRpuqRvgas
lglRCZgyLybeSCXG6TyOH/MIXQY28hRID5R/9FenYoBkFcSGdpoH0ZC2d3lh+oiL
yGVyGgQPeKxEDbOqky7ARFzmPvz46PDLc324Qw1o3P+EyypFxtI1L5YU9F6IZvNN
yDTpBmKDUh4oNUbAQTSZX6vKVQlfK0om2olj/lUh9uzXPZtOPInM01FEZnLjw+co
fCapxJxFDD5Q/LIFETsvYAtbnWl5gnBXXnmMWO8ruScQG8i9wNAzhtw6465GJIh/
kobK5rwvL4HMhLTx2KuK+2ewvjjEyJkmzI87EFs53xUuJ4hnjuwn3LNEjHiT1aFo
9Pr6vi2R6jjInDhSAHUh0WJ1fn9MAl4fkavxVnXxJgAaxvHjfRSt4hbMXN10Wvi+
NjJyeSzH/1n0vsMr7D6xtpu1nFSbGAsMZ5pkdym1C1wX0Zv8rG2ZIF4U6Vm1uHlg
RXwvDB8si51i6BLJ+35xVKubWFpskQhEYdBHzyrvXUGmQGLY13hLuLNMpSp8C+7e
XeHtYfxIynT1WOYMaZ1kJvtguJjhxkNQeAJqxjJI8iMkOqg6wJVUQXXJuk8rmINT
a/iRzHHDy1ZOZeH02EKQLZ89JPnmJagsF0elCM3oBZCQgHpwABdf8w0wkWeyJrwT
oat6X4CdqFxW1V4gGoyM7MWMyh8FQh8YSDtvAlXvqPpjlCUPPGf8QpOuM87ZHA+i
z/xQJg+EjnRdkRgxsg4Fn7J5M9OU8Fg1Yl0/UFAXdwH/pusE3rF9/i2Xhx779lzt
BNoQ4RpbgbYNDCnGYTjBppSJEQokHIe0bm4gNIoNtGB+reRoDq+qrmQe1Hjfy/JR
a1b6UAZ4LQ16vhcpWjHBCXsj3X716ix+K+fwv9UmpCHhANBAwgoSe8fcTRvY4dTc
yBEL+rrSzfOroDGJrn7yrOhGjowW68kDATJehBUoClFWnUbMrMjnzCVm9QJ87/6y
dfYUkczHLT0nkh1gFtfpXICTNMl/xrth+8/LFGvZRbOek2a5mqJ5OIRjYVBhKioP
H3ca/E6PkSckS4WoidpJU3JfF32hA1e48MouDGKfK2tEhKG7FmnK2w0adEFDzsq8
s/zWQVVof8ywRd8ecayDrUmRQVL5T+OU8KWHZiq9+cpyZTLqfwVf5/+bnhqYq4GR
arIdRFAaXKh3Dim9kXnX/OjdVSyZ7HNffy94dc8ZgEaCGfEfVkefNpFd78X1ibxA
myM1UpJPc+NNRU/AJtjQ71ismesw9TdLJHJtNF2q4+PqmZH/egoy+rYxFEvPm92i
7MULVlqtS6DyD/IkXldV54mCIMkbIvInWxMBJzsLtSZTb6O3QFrEDGw4BAuryrWC
txTRYHaeeGnCngTa/xkFQBbQk7pDyayZBeA9U6d7/RZWuE/rghIucDQ8ECMoCQuz
A6KodUupWxZWi8kez12T2pr8G4dgNsKsYDmDwTjhirAHQ59L+OofW263G8Zqxdq9
cSpv4Brj1xdfmMUcJHKGNhrpVpOZlspQB/dja0THhXN460Qeha+kiDnHm5ITKTnt
+LJ/8fztTu+ib/8uHHiR+yIlVRTp5VnSV/qCd85lhgnSRVolR8w5uUcIkUk48TsR
1VRHZX7p5KTFRsXxpuyMt+CQEjdbsZwA3zlVlH5oZ3UzTeMsZu9KNMmGK/p+WhK1
nNvrdLWagfGQB3Bl5hNKGBz1RSCnwzuFgAvS53xEvVgXGwMe4/KMVk62PQTTtwDX
5vH7QKudgOl51/O+RNsjeeu6hVSJMItPqK7aryLvSvSIJ19wtF53oPz76TJ5+URz
srK6SaA5wNpX/qoAI6aAdihI3K0dsa6r9siY0RWRUbUOgpVz9dveO0LwG1e9fhEf
FaY/xooa1uHybzKuUrmC9+HqtZAloKyeXJWT3HRM6Wf9hNJ+U111QjTrZFabKWt2
3P59+pdvjDXSfaVJarnui3DCr64zl8a8e9J2b/A3n43IgCJME29vxwFZoNDR9P9j
1Vh+NvDxeWbKyBtp5xmOcgJbfbQcV8vp+ITR+k+QESY+Mfw8XAAsQ3DJsaA7e7Bh
ORKGlwTAghtdXXjWyAUM4PKtpsSQEc4jsc9debzN6Qtjbic/mN2tRyPrMLQtjRtq
/39+mvrJaEelnRhj/UKN0KJaTzxySnNqya9Q+WNS/KSphsCP1VO32NTa4/V1AgXQ
zcGi+9jjAetGdIaNOfd3e5nVc4ON9oIkk+uQfERXhI5tB+v4Su6mbSHTGU88wSu6
RqhwQAX+VW0kQXMagCp+RABspDUlBWBgUHwizrHWt9EFGANmQoAIKrRs2ApXMgkA
Pz78QsTvZCA0n+kEN7y34jRAF+pUlmGvLd2D1l1QQrBs5zNsoa8NZQwtvdHdj70D
zNZS3xgfabUPwMALKoYKk+UM0xqYTOEIhlD8cNzrUlIoA/9rrpz+13ma01dn9tve
JVQpvfVhtNZCZdkX2Idb6ExTdw1id9mTmN6/QNoaDfy+fGdKZL2tMGFrD2ITKQOt
kZgMjj8jMTBvPjL6nIIgg/V+dek2nE40IRToAG7UeWoPsojRalUlaRdUP3jGgsF0
yrS3Mnapt7DAVDQgtEOKuRX2OOCzFxcljApYfMR6uhCry8mzhCqbOHTWXZsaQEUG
/WEq38OJnqVU/jwGSRzawjKh4a118qURg6VfZ+kCCu/TGE5SRlUu7wLJFbhTW/OD
eHso7EsFMrzbt57ANP1F2laa1KUNuBV+MOeZf5kl4hc6HiFTly805g0mocFSiOOS
xwJvsVCaOAdPxk0qqu2kfquT+x0EANE1u6ly9wnFR8J0MdIHfe6GfsziMNy8I2rH
Iaj5qIW/3g/RjKhAxGMvqTugR+B4ke5+nY3WvZDh8UuBXdOngV3ThSDVyv6KhZCE
FBRAXESx/0L3+Lxtx3FukGNJOX43z7F3uMxxcDaKI4LlDAHBtwVniGyjJL6hS+DU
L71JimDVq/EcBJ72Fetk3Gk10KLg1g9fCHki+QxXL3d//av9XkIkXEpvOdU1g0VF
6Y3aTHiayqE4Jqz4huMaoRuVN2Lxw4s5K68A8vL0kFLmZGZP/Y8AT485lKqilizA
UmIAuVGU0sh1o5wC9zyAV01dJ3cD+NZSPr8MOf015FUlvu5w+kfBUW8U8ZHdAXJU
lwJiL2bADePnIE7cFYrnki6yPvesrD1ao5MiwrbeOT8nBazjfu5lI+4l1Pw90JZq
n294xsP8fk1HXDFwLNb/bdHchSS49V20Vbi//LQQvMxl9RP/zx0Ak/2Dsf/0PrJN
MxPlPxsfxJIYSxJ2zynj0scqVdCTtKiuluoY9EpCwQw96qBh4+YKWSMLh+9nF8sy
fZqpiL/p8ugBEloaUIBu0+K6SUZ4ey/P0fRGcmmzBiTXQVzYky9VvjHhLAWgPy2w
F6N/K+spvu2eV4bl3a1L+Zz6H5G8oxBjNi7RYM7XTJGBzs1TYqHq3rrXGfkmdZee
Q4MQN/rHEIGecU33iMFtNofNmKtSkpbQb4AiW9iVqmfdsJ7ZqNDnnvuaFFgWXIsi
pXvdCQIwb6RbrA233mH9OzhFswog9505EL5wsVxKlrdWLhKzIL37s3aXRu4K8gaa
OMVaaI0LKQfB3xBVzG24H3KuoEFrI8IoF4QEN5Kh21BKlIX1WZxiprox5vQFP4er
mTwOJeE8thZUqb+Dwe1IITqtN9uGstKniy9oY9Mg6ZMyri3EHjfe+C/q0e0vZWra
4wkomePlkuiB0GpvlQzVdlVzEJRUFla3uzH9MtP3eOy4x11VtY8RtZH8Epu399zW
/jKdfu6kLPDo9N8g2NZgpT3Mcc6I9wVsNC8zMqzGg/jgKW/4tDAXzOlXyc9LPdbS
3cgupeRNlLy7K6sLYEDbCYHGOpWIUn2fM1FuPxt62QDf+8Yblv7BPb2bfEbMfeaX
qiIBkYEXZqKmuDacLO5FnLmtcD4SYqkrsPJduow5ONSuH0OJmzeFdmw36tmRjMNw
Xi1lrpRZmJYszcA5sEuLo7qekOvC0SpHoVyT5cGjmzwp7NwKtzGdvR5XBl4gECXH
9WDyCMao9gnUpYv9L0j8LkuiFig0OJUBQKAzMy7ji6w9Tl+2IAntxdvOWv13hWoG
BLfAdYuDb8ZzH1WoxyWw40oIhVNI4PNX3MkPrmUq9Po9Ux7peb0U7efacYc7eTS9
fYC3t4sd402E93W8wNyfqCMAOgQ6ftqoqNdboLQtd9xAuLh2sTWSwQ/xgcGMdzNE
LuPpPCccHg4dsIfJQA3THdr6N5zTwqyiGPsPp0GGutKtY9e+9WZka1fhGBzXzE9A
xR07k5GISm5uOiUu1IlXdLYqJQtDnLHuLiI1Co3sORFoydCGuSkX9FJBEmg/iwIs
Jsmp7HhiHatPGVmajvc4o8ij+QlHLBZn2TRRUU19yFTbcRtC2Vxr0z1gNc4EIPmJ
k5jaBsfwFDzShek7BbQN6yYyyzBl6cEtwF/ZbpaziMwmC7B/QX0V8UPk9UsEt/hU
gaxZO7a5agumQXBePtf5MogH1Siiv6TnFODZxEgc9mjIAh4TQ5N5e4LyOI8jlocs
P91YVmyty8L1lJs708CTgXrvwW+ZhxE99I+QJka6Ja1e8/ztzwQFFT/rLO9fO2R8
zWVMC5CSoGQac6SHfnp6FOKwzuy7pQXH5fCPnvz3d2CLz/0kUxfMfOjUa0FWD+c7
yh+89Y8HHYR4Y4BExzFjobWpFwsabau0iBKpAOy+WYQ2TMFteQ5JcmWngpuWrFKP
ZUr6zywmIvOfTczYQ78+sYywqkuh2NeOMZXnNnFIwdEYbhs2LHily5bWj44vgo03
YQ2jGn0y0fMwlCo8Vn29T92VyEQuvKy3WdLqjixpjmvAaEP9P3B/69qat6NqD2u/
6FRQCfdrfHsefduMiKlgGkKONgyl8QYUFLS+VKygVYPjXtUPVh/AAEpUAvqdbno8
cYPj5Amhdi12LbEyfVkTGr4MIVViadsQDTmBRISFNYQm85EzHDww/K2cRjFPsYta
CKIMlK0GZvuJ3dUFHEFdC6cmFFt37Hs0rs05RSlTdd1EZcr/fjnPgnBz5RIuEfQG
AA1M4BK2iVMaeMnCd9jEuZpPe2iXfJdC4ZC0mRMeLd03sacW2zCODR/T/78h0bSA
IsPEKsYQOUFJSbasx4nbGzVpfu/vITWfloj6gG+lhVSQ3j9GtXLwWAEQs+mFG3GK
yvMIAW2E125CGGDn/w0ETp5Jgpm5cPqcu+8LjMln8oj0QY6Jjc94pgXJ9i3XPwx+
m4bZV3TaCO2KW0gCYUYhSdvH6kXFSB3U9BnLq+mcddfdKdmohMZO7tbvzJm/Jcia
7GL+adDwYTUzmcAQXNr5nSldWT3csLGBTXbFywyZqX40eabXw3mdM8mFaAY0IuyN
CdKJyC/8VwGHuZ+3/HAQcZPvacfSjDTgMgTEzv6Rn9lKVMfXDThaA6qGuXn78In8
4Rg0pKr8Tv2J1wZEqQCh1eyHxxDBS6hLUa/o2/tYVFBlselJ0rQC2L30aocVE1Se
xzGtcn1nj9Q+93IEkDWE5SOXawtWx8+tMqoV2ScwaSJDk+mxNcq5lPISxFvwNPE9
FThZ0vRlbwc+DHslE6BRXCNAJyi9AI6YY0ZUx97KCuHUQcJSbEmiAb4ECT0KWSjO
hBHjiLlYbTqTdazRMywzJvHG/EeIF7DXo22ear9CNNhlDyoFLdWYVBj8NahacVqg
ciZsMINJoF+ibS7qNsmKxIWhfG6y+VAQgnNKYDGeqNvKqYltrTYjYnPUwT7avRoT
yrQMr4pj0aIjWo8ozhFnjjRLLwP5LivicwO1nwajlLWT96FYuNiUsKfKw+MqqBa7
AVLEohit7bcljVLgOKKIfrUlsHpEEREZu2jJT/s81A4Gq2okd//EYOpdSmdR9b4K
pntf/h3TsCh1hGG11VvMoY4uHpx0G1APllGjZFSHCfTlw9NeFkUe+yguUEwhIn4E
fSHzuVT/FzObdGV3pXOWEnbBz7DC7OPbenI2pIgtNI2GuZZHWZIrEA8h0VJMdJKc
ctZZC8LazLIRxEOz1ARQcjkmKIeeQk+f+JzvYIm645r0E8j4Owa0oBP8VS32Fmf9
5g0kzqyUSWHNazhKIYvsIRsXp1EwQiZS+c2u7UYRqfKODLYJu6pcQULKTPPwbvzm
IXSM5y7tYqe0N48hOGNSkc+KxtQDwgPZHzdSJWwcxFZpootG9ge+yYBaHXM3m5wL
BAaV0up+a2hLD15Q4uMaD1qQb+f6NL2qbpXwAg11ChfXCPpW38gRdZmhIHVXJ23k
G+l6ZXeXPWG7Fn4+9kO4OlLR5dg1FQPNmZ0Vw7D39tGxhR8IxioYJIN9Ut3zzPYE
a1A5xUfIFJJ/3jceS7ZvV9Wxyk2T4jjkBpZWeeBfO8K67iihkJfFdEitnlrRqxha
sJjgZGzxd9x41qn/xNScGE6mlIwt4mqK+7IMiCkbnxkCSDo+FnpwIIIXJFIvRyjn
VuZVpWtr38ACMqc4LeOzOJhXaFf/ZERnIFXKlEJMlU5+SeRmjBXgCnhKIi2SGsOa
B1kGg1tPem9DOD5gfNFWVYeKO/xEOLrTTL8qpUSzeJD+APU+QksqMD609NR7RKKg
UpRR9Nxkcgi/sih2Gpzyk1Ltp7Znb+koo553q/9qMWuiBaCvteraLInNf/5Dy3jV
xXcDypbWJVUjyp/OzUD6JwFoRXhk2WwK4rUjVhS94BIZYiwk2j+shWGKlg95baDJ
d/bEvNGakwF7JI+K2r7A+hPNS8yrRaFomXllbI3mrHRhKViCMdONGbMhrRQapw9+
aht3/nDSk6tiULTz6ORDDUvB/mZvGQ5HKIrBvf0BPy7HZeayoKMbNKFz9mqDn9au
p82CgsqBEzeWVwAfL/C+o5umFHelbjsz6eBjaQb/ojM4CnpEK6OexUIqC03ebLBZ
Up0mGgC8ujJLqqgf3h5L66YrOVqnMK1g5/52dX9QQMsVmalJNptLsRX9uyqe66AZ
JTxC/vQDWeEiUEZOAxvNthR9WVw82y2+tpEPnWgMvvW8clJrqoox7cpKSYkzgKDj
KYsT+4PVYZKb05+JBVdJFkM7P0xWRnP2Utvf3mdGjq0TZQ7rSF7zXvEZ9SzynjxP
mZbjMJ7c7+Srd513/65Rem5nTe1kzl078ZaqEJU95POOsMGt3UNkE/x88X7jhbTK
0olDZbzVENeF228gM7Mw//zP3IeAK/FG0l1NGYjr/GW0Fw4Yf7U1p+bs1gLljWst
GBH7UXFk7ptVUWi7doeAEJbN+i/2qrjAYwfiI9tn/nqk+SrWNvaX2pU4+mU6MKbc
O2mb5xe+LZkZbBEe4TVfDh2Vl7kikjzwTjFVd0YewDdxsUsA/T/s+hePzoRkYV3L
g0qadJ62NUl1zCfP79zCNvEaKch/YE6Zwh+ExfHorEOxeLNksleMGY1YkEJ3LEwf
wIRHq1bKR26wkaHVlbZ0XMEkmseTWfB9l9qMBpJgUb3/2cKtLXOcEHMx0pnP0jgO
DkrP4ZHvO4bV+/fFNjkvNKu+FEuOvyvT9rXGJqtau1NR9A/4G+oApsXhVewgxoHH
1OAxkqRHzmmlQp173CUd9oM6l8Wfl/Li7P4X/MPxoKcapad9pFtcBt9jZv6Dy9ft
7KCxdkRxn3jZ3f0z+pK60mulcoSr2izSQ4KxjHFan0o2iR4kdOrEvyTXQL10afNy
v92OSd1qC5wKuWHAKSj95Wd7fo2p/b1JNnn2EB8qiE4ESRIpdSSeqtHi/qY1gxk9
L1nS705zmjIZK6JbvXz9wbn5uhjJoTx73vqhyvjYM0JyKObYV6rJDspQRVdBou9F
XTIG6oUuuRCX2fkPVt0NNiphXIKD4+n4A1VuXHo7BwJZo3m0ab7X2k4tgZy44JqH
CzjNuSQU2BBNZBlIYFmo2RKtscGL+9TenUtuXn88MNDS/OZseP7vGyyQQiDcOMxN
rf7NBQyjcm3H0KujoeNOLsJPpQsylTsPrLap+4adiypNrXnJOw8M2E5H2c51bLBW
P39+guXTnwDfTAarVDwoKgL53HV1o6586A8LDW+dZ1x5qFf2s2ADN4OmzCtyTInu
burOciZ05ZGWC9PRLfkolR1prcfeBkNpzaAl6xEFDoo=
`protect end_protected
