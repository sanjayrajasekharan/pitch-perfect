��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki���2p$�/��tD]*d�4$O�n��������xู�Mf�!�H44�ɾ���#f&@it��Oa�&l�D�4P|�צ���n��D���M�2����4�n�8C	?��f���	?
W�Jb�.8Ӛ���c��F��!Η���R�J0L �R� 3zOSw�##�h
���B��!�����(kWo����(4/�(ҏ�\&¸._��U��7[���Ԝ��(�X"R�2=�id��a�5A�Nr4F$��TO�z���~H٥��=!�Ϋ���m0�]U�XRh �m��o:p�V~�%۪|��&�,�}�������XYdr�lGCu�x�k��'H�����>ce"[���E���2�1X��'L=�f���ƞ�GNɏ����[��ߍ�3nj��]�Dxg����_U��&��
aM�k�ik��$�H�Y^^�ڋ;Dg��ML������:-���ӱ�1./X��k�nR'�bbZ�Խ�۬&��3o �O������?�;��d�t7G�¡�
v�������?jp�;�k�.n\���BgF����/�m2�IA����@��"� ����L݌O�^���b����f�ѵ��Nj�ҿ�]ɵpmB��7���By��:�%��Ɠ`�StZ��ޫ���� �:7=kN����M���C=[F�q�(���>:>Q���ڃ��\i�͢B*�yP���MSs��Fۚe�X23Ah�v2U���W)�j\Nm7�,�n���#�����N��x+{6�Vp���ƿ��Հ�-���(�Ep�:t���51��M�)�7��&�/, ��=�������!�!��W"��
�VU�L伮�-�ݛd�j�:;���G��.DIywk�'d��@���,+r��sޘI1��M����0����ä�H����B��q�������jF�R���Y4����E9�=��ј�Z�C.o�~�� �ܧ9��z����u`��fL�p&��4:�2n�!�_|5>x�{x�dӧJ_(�e*$[�n��Q�7`�a3c�UV�� G� ��x.�p�$�������d�#O!��>*�S�.:����!S�O�ck;9�0��+�2�h�R�fYاhx��j `I��k;�+����X#\*��N{�W�e?��,��Y�����Hwk~�Y��);�k�8���#����Xj`�Qx�Ry�����أ3B�����k	9	��U����Փ��f[g O���o��u��d���8�$rZ3�K�}������z�3��-+�f5|jŜ� �M����` ~3��CY�]V������k�[oX�y���!I�$�M_:t�����3��ZX��j�����᧎�I�J���L0��*�t���\Z�(�;ѐ� 0��񃏅�;�s��aD�U�~ʭ����:%��d�%��'z+6�J���[A�z~R���7�Kd�����Ǜ�$OW��̮�Z�BS�թ[��/���ͱ��_)�$�YyJ��2-˼�@�&���c�C ��,X��U����#��\[�)�[�DP�7�d��yR�k�q]k���]%�����8=.�"���Qg1�u<*��6�+�&)��ו��=�	�� h�N��N��@�H�W\��b�ma��oQ�_�xA����C���� ��5w ^���n1��_)�th<c�<�k�7�=��N��q7L�n5fq��)ȃ
�<Ht�o��2����t�͟8C%�Qt��n	�qN5J���	��-� E�|.�~u@"CHO�m�͢�����>�* �t������cV[����L��9SD���#6EY�Ρ1l���&����bЁ�VdxL m�j�rC�,�n.�� V8,'u� GJ�����(l��e)J5_7(��ONLn�X!v}K��5{Ay%w�Aխh��Ո��f��3�cLYv�����������I�s���Ϊ�V��-�&�|7F�5	���q�ykE] ��Ԗ%�2��v���	���ϐ��5$��Klp�����^�*��0�C�n`jDj�g�6o�*�H�ˣ�r��c��`0B���'.��v^�*�ʄN�Jj9�3�������%� 9� ����	3v({l��$��Z?���v\X�"��*�f���AȺ�;�G��x�a�ԭ[x���,$���vˮ�S�dl�N�^��ܶ��ZH�X�#u�Y����5��\?��%�;�c�<k�9Ј��g���=Mp���N���=V��I�Xזn|Y����(<���=�?�K���H��L���Lk���f�x�7�|��ݦ�q�	���e�B���$
��=RUy��ٚv��M�{3,�<�r��tȟ�
�zuܸ�/��8�/�a&���~�jy�K��L����*$�0~уwQ�Rib�!8;W��#��R݈{���sz�YL����������îF,���.�tF����"�hO�UE7_ٷx��)ݤMؤ��1���m됄J�[���r�/���� /W?����z_�"���AO��gn��sl�7Yl��=�Н���v��-�3�k�Y�UTk��.�y�r��v3D���:�GWz�dg7��^+zo;t��)1f��@��XIZN_��+鏺[$^-J
���ڒ��J�rY�e=�X�c;�Sg9�6�w�w=���}�����X����l��Y�gLj���o�5��~4��bR��2���亍*XE�/�_�/�bH�S�F�t+��������JR��P�rHP�% ��'{�̹rhP������/; ���F�@2��bf%�yQ��o��3�\�s,h8�7�{4`A�ڣ�ת����m�Ǵ�9�4���hd���b>�f�QAS��C��n�T�wX*��6.�˻�ȼy�M=�y�_r,��3�Ml_�i�cY��L�6a��!��&<��6˫�?T	?ڎ��F9��6e#v��t|��sX� ,DA��l��t%`�m�)���a9VO+��5y��mK�=�3�.�H�(��#�u��!���������X�Y �}��9�� ���l0˚�75���A���1�'o|M�U޷�d}�5�Q��)q�G��.X߿�����Ɓh҇Z��c��B����N�絢��<4F%>��;�0�Lߖ�*D��[E���j�ݏ�����ށ)�Zϖ<�r~ �Y �Y����.e��E��E5l��sT,
i��V�ף���7�q"O�K�,��ۮU�CH�P]ط�I(��2F�3Fn��0�F"�F�ph̉|�zi���$]��@�p����@���jG'޴�00?lhx!õ���#�{�2$�~ONv��/�X.�5�Q�#�E���̃yz�޷��ߏ
�n)g2ǽ]�Vy�FTp��w\��"��9���`χ�a�J�>�Ht?A��O�,�,@��o>v��#����B�uN#h|q������	qU!~_�\/o ��?�Hg���U[����D��e���i�f���uAɿqt�'��g�Ļ@��kw���&���)��u�O������뻽�q������2�g�����U�9�Q�h���J��N7#|�]��6n��c&��j�wU�y-���^���"Y�����06�h�M���yzQ�(����a�bM�2l���bhū�l��w�~��Y��A*�&��	UϚc�c�b�&!3M��w�QZ��~�gǬ79ڸ���Hđ\W�������+Q�|�����?RFC��޼Hs�w��O����ա	�o��e���;��0�<@Y����G�
w���G|��}�Orpٱ_��Q��|���q�ke��XV��P{�+���,n2����*?��! D[��	�&�����n(���)���h� )��?_Ƴ��֝7?�g�ޒF�[F/�� 1��u)!Y�O�G�5�j�Z��w�2�û�(rԫ�'�	 "���ff��o�fy�HJ��Qb �)eA3s|���د�W]��?z�fw�9b^���
4��e�ڸS�Z�"����/�k��%����gɽ��aG�{%��]�Se�ȩ]� X*��-Mݓ]�TG�k�B�=�r����	���~p������ͫ�P+1�w��M>gʪR���Q�l!i�-	2\�/�7N�NZ �8���o��<_������pK��w��b�u. �ty-#D.�>c��z�^���ZAƷ�֛�db���EA�&�F��LL�YaϨ��v|��Cėح=��կ7+�@���������dh^j��-&�95���A@�t��Qf��Du�dA[���6xz��Ѿ�9u����b&�.nQ��OT��EA�k݄C;��u�!����y�w�Z�$l4�Bi�'���re�X�i���� �=��C�s�b#�Q���Ձ{��0E3G�n��Ź���S�i��;؂�/$�b[���P�~gX]�T$�P�D�^R�<��<��J��'Fp]�9�����{��*���^�2^��t�4�O�������T������B�_T��|�0���l������H�u�D� M#�f�
@�k��]�@�
��i�-����Iۻ��(剣�-�e��D�P�q�>
�F��9 1���:)ގ����, �Hvټr���;Q�k�E����D|�}�z5W�����!�a���Iٟ8+p��%�����Dc?�}'���~����Էl��i���Okך���[����?��a�LA��5/��vT��q;!���������*�ϓm��2��'`>D!*xd�M�go�qM�9�xA^��b`�qJ�1�Z���"�+&z�7y�o}q��A��{����V��l1�rZ@��Hz�:�6�]�S�����р���
T��L�{�S�����/��Ʋ����L��Y�b"�r@a��	��y»�!�1��?��`|�g7��Q8w�����Tv����9)q�R0g��ڴ|n��d��9�o��
�����ݨ l�PH��z ���pN݂9U6
�/��?�~�U!\{���fIb^�),Xa#�jY`0.��0�,m��ei��g�q�:�;�G�V�n��(jQ�]�l�//N��A�D��ڦn��ӭR�p� s���y�50œ���@N	��ۯH�S���Z�.��gt6�yQѪ+5u���Z��C18��$o�&V_�e!-V$� u���<"�\9��*��K�[	�����aA���]JH�)���w+���v��rL8ή�������m1Uny5_����%Z��
�(@@�q��3�L����BT[~�-0����kL	��̅M�~�<�z����������#ҋ���x��Teɯ�Ni��dfa�R0��$v:��Km��!�φՉ�CO
�&�T��k�z�[�Sg�`#�2/t���T���� ��@b������࣑�FY��!�����1���1�O�hj�v�e���@���6�Q��!Z��To�6)M���Ԛ�,88�ǻL�� �.-�Ȱ�ſ�_�1�g�m�7 �R2���OE�z&���4���5b)� �=G��*C>kF��`��������f�+���Tܢc(���D�]�dC��4�X qI͉�l��L��5mB!�RAC!:��\X�p�2j�o�k�`�gJj�jc8�b���ծ./r��D�o���z���}~/#���m
���=������Ǧ��z-x�*yy�XRQ���z8h՘����.������Ze$�bX,{{v�aT�b�Q�=zcf(�2؈�����)s��O�����jL~U&�i&����>��<�&���ߝ:����Ȃ�Z���kO��X��Z���sE�<��ziB��b�DI#�F}�eJs�>���̛�xK��.��������6쎯�nƕ���/��F��O��!j2�CR5���Qs��,22���N�PR%˨w6����ֹP�!��*��:���sҀ����$?Q "; ���ø���F��_�(�x����r�BE�c[�{��4�Q�v�<=��4*�0#��)
 �g���c�~��.��Y�i��Rp� ���@����>�Ӏ��ݍ�l�q�?o���}I�� ��M���R�� 4���+]��xx���On�_���+���mIaSK�=ލh�J�1Sv��*nC;�#K�4\,�91�KJ�a��7����)pm��B�1��d��e࣯�ǝ�֧T�ތU'�u�	�e����z;i�i*��k��T?2���X^G_���X�TL�)X������X%'�ݮ�R9'���TMΊ��@����	��\{ ���f�tŵ�NfgX�N�n��"��Ҽ7i�-��
�a�0>�_�E���\ �*�5��\73o�� �Aߨ�P<���j3F�0/���i��*�:���i7����
��3u��X�ơT����_�P����F�j��6��ϩ�<��k(F�5 lws����T�//�]�f������������0���V�CW�� 6�cquH�M!�-��!�W�J���]wJ] ߌ�y�4�c�W�/��n7��h���65��o<�Ҭ���'���
��" ?�t�Y�����OZ�gć�<$�/}��	��L	D�uY;"�/,l����&��P�C�(�TC�7�(�R���L`����_���J ^��p�s3N��sY�+Z֣lU�CfBHCz����b&���GJk�y�9�B��1{Ք�|]�C̷�͇n�JVh�3�S�ڳ�Q�*�_���:�]+�=���m�%����gB�թ<yeZK�o�����#�e<v#�]��|����uE�~:�F��F��8R�*����u2`��!�1?��K�Y����/սp�`�t[�B����b3iѡS��7 y�N�LqM?�+���݌������V/��� ��g盞�F-ݪ�9��1���ų�2�DS5�u��س�`p��3LiMN$9��M�X�Eʴ_�n+�(�j��m�P���EQ�nq�{~����H�[�8ouO?Z�3ח �`�����R���,�~��"�����h+�B� �p46]�{p<�������|�z�>i��[&kȁ�
}�%��EH�z)l���5��yM��OL��&��^�.%����$,��Ш�:������j��Z�~��\7~� ���\��"�@4�JI�0Q�x��<Q�#��d��b@�v�(Ӊ��<����k��3�ps-��rX82����;�)�g��3�o����㥗�Q	p���$)��Y�7���>3-���S��Y�p3A�ƩwpXD�½<�kjz�����������	?��x�Sդ��ڴY������X�=��mM�w�?�&���%Gɳ����s�Z�\1�ĽY���c�	���k:��}%lc�W���m��I�fr��zn��8ö
��O�:�˻�g2�Ԙ�"WĪ�H,M�E!�9rsuqg�^�+wA��@z���@���<.p��_���+c?��m��/a=@-E9����f�pkΪ��	�>��'=�2�Iר����Z�Vp��+��b�p�{E�~R�O�f�M��Ph,�|�)��y��͐�Zͪ��"��D�
�����2:�|�Xb������F������%�*��5�*�y��p���G��zd>)��q��f�n��W���}W�Q������;9a$����U�H��v��7�M�^���ЈH�W-Gl��AU�B5P�M�m��a���ת�ÓA�Y�#���8�-�؛D���-o=����C���j�'�ާߙ����]�TM�u���)�������Ʊ���C;;�kws%����25c� �#�'��G[y��O��WL��Dj%81Vd��k�4asΝ�|"�:�⑏ѹ�R��h��s�bhx���ͺc@�b][���ف�A�r�>Qm�*PP���϶tJ��Y�0A�
�4o���9&�n>��D�z&0=\y���xn�:h��d���I4N���p��@ �I��R�d�:���Q�7�$+�u�V�hl�ܢ ���WW���rv�9;|ԴDll����D�>>���^-���(ʮ�x%g� ��;�C7���a��!�I���s Tz!�%�z<4����	����E�F�bp���]xy���u�W��
6�>�y�N9���ӱ䩃pР��{��Z:�N }.NP�	m�/�����J�W����	h�Xitj�-B��X��!�m�.o->f�O������ǳ����q1O<�M޺��}@�עB��Q�!
�4