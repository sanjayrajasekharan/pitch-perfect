-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Jm75Sbtj2xAsIxzQWMYQ5DHrHFkjPV5rLwINEHwbKGxKHfPt7+idzreYG7vFPUWE
vzG8irUFF0fZP9K0t09efGCIXod+OJqIfnvP49gtx45KeUfARDIjpix+VM8dl6KH
thjVeLvGlNdGl1khMZIDu+Jvd5/5u9TlsThgZ+hOvAI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 12096)
`protect data_block
lt844jY1cedYs0/FHRcQjb7pIt8mkELoatBiFrqaaSUGceKgb/qjud1/UEYR3dvF
vJOe4MSiloEEq+Y93y9cuDnuOfTezTDCAWvO6y8onxkEEskHU5h0mVRYN3sJcpgs
kkXhzNAiUw6r99bpW6VVQ0Qqq8AKRwN7CUexVuXeydhjboFyQ4zizGZ4j9x0hfkT
IY46oR6SVuLb6UNdpcZGujOvOqg00J7rre352c11bDg0DhDIWDjOh0OtIwDxsO66
9Ux3quMRUAJA15y2FgX4B44uCwBGKL+IiqlxylHFq6VR5eHPJ5E4J3twkAtJhUql
Y7R/OwnO1ewKaSyI74LXwmpjm6ZK0CLvhlo7haYmnrYaW/BIKZhm3+fUVM9BMFkY
LdcvRCJ3zhVrTq9HzrJ1KEu8FvrnsRYB7yXdIj8kEQ6oc431e+FKWaz9URTcbT+K
pxPe/jO/EUG/oMHSW7wwGsGcx/hEJRCaPdAD2JzOaAE38XGbtTu4PWRixPFDBPcP
HdyCss/hPYk42oT8ylIbF0GKvQkHmQFoCAK6v+N9bw9Vbhe8GpO04gyKhEgy6K77
ceNLme+ZBv5ZLMTXpHhiiiYrMmUKAbR+rmiZw+2usMHMRBQff+V8E+AmYkYaRdSj
kB5bIq2uH+Zv1UzFReKytrHPNSMdL/Empi5tAqhIQLjRVGwFNwYUOm/rTgSYtJYO
rj+6uA9iOvMZT1Xpe4f7ZHjYwrBlqKYu/lJ0XXRqNNv3RFrwhp4stEucfoLEeGmP
7RyjskZ3IBhQYHg35QMXCZjil0/CqYPetKWamgm3H5Hht0pYictebUXttXw8Had5
KsJMDeXzOMuvjhoCvRjlxt2CFl+IxCxx/PdWZ+mwfY4HZHZGmmKjC3+RaQ8MkVHb
Zh78NWu7qE0iwlnZTfFYGUR62AF1aOk/lxZ2lBngOY+8PtVqEKsdvS1eChR64SGb
k+G8GoMuaF+rov5T8w1ChW357+1GIvG71t6GKyZQaVgOY5/piLd1XdXRAb1eKB32
WWSt+8lslZbdoS462BTaIiJkqc7pvkDmSDL0ILaAtIYKSAiXoLOfEhOxIUzidSTj
kQDXEkfXGvJb1EkEFgRtxC5YEHQwGRWoECxQ75FNpJNY3fMdVIqJ/3byzXbVIqG/
0i6ucd2KrcIigffGxgFm9wmc6Aew09Cda1AYnmGZRfBgVTcSWj1kd3fWa402sRCK
UMDtrYdu9xhm0i85S7sSXZvXdbbf2YBXZl4NiUDG19ybqZ6906MeTy1BcYImXhwE
2E8u4ItMZZEnifl9CkjfKrngtjWl7m8JXv0HgOWSk+kYxxdB1yzYQYkgEz4wX/Pr
sDKDLldR4LJVbjrMpjKSnx4EX3+d5Dix/NV9inG0Z+ybL6cU9hJD7AwoBIp2ypFS
X12rZhKC/xXJciFQR34uicpXETN8o9AknezLzJdVOF+0stWoLHC4rUTaqA/JINeB
EuSu8SoqKWWF6bZKZXUOB3w5NjVcE5qRTANl23I5T/MnA17rVyCiSXQURteOKNF4
AQit0ooJprbBmHbWcmsMitD6IdICG/4TDlXbbV8Bf0R5W3FkKc6X+Tt86KcMbwUU
rx3sKZdk5jz/Jb4g36KAfoDyQ16J4n0utRU1NFAMOPebrIw0ToF7mClrA+7z1I1m
hrO65vphWdUBMFxesHMHLpMW4xjhDA9o7hQEnQytmlAi3p9PcbxLQ81DyHD/rrcX
buKqR2+WPlbI15D+xMV/Gx6tchbcnNuILNizZNpxIz0PsdzlIg6kYF5LNqfgFQfr
yQxUE1TRAdYexBEtps4Ov7Z1qJtE3h63eo8X6MyvrVGedt1F0Z/ToUcOWRGqyMha
6r+J9SE383+ruXzdGlaajU1VM188bMKgewp3nmtaf45HXPcqwawVwkL/17L2H9V2
m+UTM8uLNmADgcqOKCKHoALL9yc7Cha2PPVX2JzWy7o6WHMnB/Yy/l9w7ntCC793
Kt2PbTzKw76lJ2qtasJ50qBNflZKl1i4fl7jvP2rLn2bNWB0BoupPKRd0S//2Zz5
Fu3fD327Zj7lRXfN58lIIa+8qbvj3nqYMY5eA4X60Rd4Ye7PyrwRyDdNsZiJ5Pz/
4Z4iJvx9xkxhAg1aeEsY1mdPnuC5fA3KGeBr5aOYPujjtwB+AnmBY4jFAEya4L04
2GLD5hOTe+7buuNvfF54a2oymTPlGOISYXsRYNdLXYy9NYJte3R/BASOH60HiaJa
4OabnGAPWFDslHr3BzL/BOuElRzsKbA4JbEvwKIkV6SXEuhIMfvnpJEjHnNxewND
pRr99PO8Cum7bWAj4zw58Ptu/o9u47FEZsP3YxrDSJm8xfPFLSmvyt0Caj2Rcf2F
andKs7Saavuu9RaGSFlzlAG7b2m4WOyUfz/+UB6IOLFanrNLuHftUOPXpPM1OrfO
K0poMcnIqNmdzVgrchrPcbvHY1zSuyffcegEVXSkcYV5v/mKJcds98dJI2bkDAy8
YdkorIx0E+i9Ylxz+gfmSX9QXFAA5WHJ/fwxAXtc8DmC7zXvjDw39y0Y+7ujm62z
MGUqWD3/erbsEZEPyIXuvcPI7iX/FsrsdwR27rUkOCsarKo4AoQlOm6dnBQ9iBtT
7zFbgQcP9M27L0TGiJm2pcNqRnxjchvmvMW81YnsPGMe7IbLu6pPs2dmVPiPEC2y
8bnmhsZRoopcp3LZgg1dUJnbBW+CevbkMf/b3okCXLcyrkcrFYJ6mIrSR7NG/PSa
xtxu0TXRj4aKGGziaJPCuEHqlz1Im6zvCJU1i+eLD1Qk9rQAshLPaxUyC0RhIQuJ
7Ut2v0R/y9FvEjzHNrAVRQI2Q3CW2NYkZ9BIHG7SilVxt4BG5MsuAH1ImnmDE8eP
pzF4seWg5URi4hjvqLpzhSXaSZWw73ZBeSMB1YVMHCtqAKjUPGPZAWsCIbXnneX2
0ow/An9gGg8EEHbzbuhTaLY0HudzhSZdRfb8ZSNkdfPcf+JcA1ISJemR/u2LIb/e
SH+m6lNpM62Na+9CxoiBILBEQzCGWkB39Y7/Bw1qWr4ddUA9aK6e3w+NvddaPVCQ
3lJkMRvb1H1oHWC2XmkIUIljWFCL+RABPvMqcubdXU3j7OeEjSg7NrkyoujQE3Kl
XKd2VXl98PWKohGXY86DAIGhtmY1oxXWUNBjfoz8O9IBi7bqKiReAhaWMYhmiZ78
5kJpPsqB4hRwb6pDgzh+trxO9dj0XUMIbHUT3aYpYUczh0wDER6a4VxCsPEoRaZB
6iBRwGI4tp/KtQDU1g2RQPjrP0EnEswZnUPJWuAPA1N9nQ+cQ30GUXG6CF3idl+z
V02i4mjgaOP0I1fMJuoyZ+mgkJI3C+Vb7lyH4VEKMyH+vCTKpvkXTJHhOipfRbOK
lGF2N/MJK1y/Fzk786rTGACE4RWppRsgsBBdGtGvmuU84nT3ujQXlmcMD/svaSVB
vimLP8vsPFVA02XMb5pQeCUoHfJVIRpNV8O1635MLc7adqTp8G7/3qUfdWEz9svk
5+Bbzhu3oTPiAtGGMC+7b88LjJQD9zVwVAHI9zXKHmGVu7BD+T0yugv+6/1WlYMS
sfKd5lNrFYiTY/x2w3LHB1AhGi4FEsSWBvXnSd3djm5LXDK8xXEFcW9DDFYCsCee
pCNabjRhe3rE/O2wqyJ9PMcPCWUlvvMKQdkIbI9hxcFAENgXazRWm6gbMxnLYQCB
k6eWjLUc2NAmSLpYpTu7Vox5wmH57R8MKE7g5uPHXNm9Wp0xsOq3KoReWOSTLQkQ
KEggTYEaI3taLL23fLYYxjuMIxbzGwUeFTGEgngPYdHMLINWknFBMHUBRIpFJJ7T
03CRzLpmPlEZdCOkLcmYdjTMd4vOqkfW7S6aW34652Zt/+WdvKvDIZfATpPFwC6M
POZTywmjxrb5c7tXHAJo1ariBH7LleaHI0n6Ne8JnoPWYX6tIgM6OgqjcHmV7MFL
St5CT3xZRzefphpC0rcHDqiliEMiENpAqRIU06xFh34lU3Lh/v6WpskgsFzXjrvP
yCsLy9sa5rOK0PXFAh8C9vHPyihCCRkL39aHisKXA2Zl+kVfO9fKvtpIPSi3TouF
Kb0GSRDDQDHCc5BpzPj/1sHYuTRoifkVgPVHxBhmxR9r4ohnCb5Y3U6i9uWeSfJq
o/iT+4UptRRv0Jwnw2GxgCVde7kpvIMiUcnE8iQDNXZc0J/bzSoWPleOLpVhAd6f
Hkacm4DBZlhTvkKuglb+e7RGg45T0RcD8ydvmelsUvXFW7bhhNVOosPpqwZjubuq
fFByrWaFtaZ1uqA264klkwgqDx9Pr5q0Y5/Ej7IEE6lEtR+35XLJ5xiwaUMu4ZEr
ioT9MDHqEh8kSgifjtVOjQRty7QE2EkNRc6hJeOzwS4OnW1xiBR3FLIDvfFtXnZ/
I/qL/jC7ztjm8pNxgAT7g4bpnQDLU2efCgfw0TSo8JnZBsQJ8yW0VZqspusV9+Yh
S/xDKSMVqW/FI/8mmFVjG0P4CYD1b18QuBcWhSGJwuD7O3vYqzT3dm7EwY891zhh
YD4tmam9fRur4ItPJQxHvh7Tb0c2amP+VNXF9dc+bMomhu/Ffe8tn0T+XA+8Djsv
f3pLyt6pqwvj1HsEXGzhjxgsQQIwoEx7Xbrtgf686z37AvYKL3KsaQfNkMAADsXV
mLZbAEAXbGlw//Bc03g3/Y4pQoV9ioFKSmYadrnW8hLxP6aoHkDrL35ukTFWnUjE
kbJkJpK6gKUPsC91M2dUIKrFmIN/EMggMSSjoNN5WkIKNPmF7wEtbT6lGVyWSrmm
ZkedwMCSFpMasBKaz4w8+hN4r+qPav/saoa+b9MVHKn9FrS/MUcm6MtelQ0RFPhR
/LikTeiod7VTn6ga9W2EedkHHe6FqtZ5Nzh1TvDtBR+BM65KY2gu7LUJUZl7+0HY
J4+2QxpH2aOlCWfORWdYY49hFqbbOzM5E3dZiXiWu3Gyk98YR8jCEihRjAfZWmBU
VNMLYHeCvaoLMz+iWaTWD+0O52zIZtfxxGU6Dha0zXHCS7ZdwKpwY40fERq8hSem
6bAl2jeV8O2HuxFcSH02AuUN3iIbLq6Qh+GQV1ub3eDBnaGwCdLC7ICp52Kc0Dlc
nAzVi7u8q0LQKpJG6WZeWcMTcK1DBbAV7Q90YrIB2jspQ4wDxobs0srRmHM5owD6
CtCuo3LOIWyFPSe/oSXXGKl5btiiviZlfCP45LLb+guxATVwa9s0xcNpuC/yMtEU
cN+wLcC/CizQvPBMrnxpXl9QNzUyMNOepnAaXMn2EbU0KScnq/dJztVoF3hn6bMI
KCPBA5DvatC1y/fLcxdTdbG/LJAc952cikhdKn+U1yv5UtY8mEU92Jrfbowwq9/n
MzJdClg4SDuyDC7VGCFkiQuCaF26MCGx+HzHYSQ27CDbuVqyXa1tuYnYipmMlEbm
BR7IxctBlmnsrKPVEh1vgZqbZxMHvOVhrRlc0C/GbQh8CLpVzHa+WO8ptCIF8UTS
4WgWxteGlEgWKZ77D05JDEalhdzfaYa/bvc+xWhqydv6dlCU/NKFA8HZknqmfIKL
wbjiBIS6Mkq5vKZQqrtXOsLnQlUDlBACrI9VDe5PHObZdryZVF4xkDUGDiaKnSeX
b2OcBcSbZTxVgl3On19fPy/QRLG+rv5yKNPcPuw6dVHV9UZy+y5kPV4++7zHbnlA
GBtuJZ1UBVIgUtCIJA6WPhpesGXjNXso5XeJJFOJ4A+srAmwMcEtRxCJhYP9UCPR
ncFTz8VoHdbn0np/1rdaVAMzz5FVQCjdkPmx5wAnM3cQQ+LWc2JDWv5f7mJQawws
ciABOGhDilKxrxCj8HEd8tbNS2C0vgQ798PwNhMOqGE9x6xgEsXgK4awJQ3iPmUn
EnKlpP4RbhIfgKWbifETIJuJgoWdyIPAcHUHZvm7xaTHVPK4B5D0oBUX3EU7SJQm
nOwbYWwLQ2aOBZeI+Ut60VzRXvjuxq3kevh7DPiR1qpOSysHtsDX9+pPhc875f18
NnXfcfQ0BkcpoByhXdOV5/peJutrFRUyXbyptZkHK8PB+PNruy9R0dFS7Z2UJdm8
xRbfZDf+50bUzHp1pXMRLQjzxBMc//lBI5WoaIu1p3pq8vjfNH3BnWMowUAfA0DB
6wv9etxWrgmlg3/OzB0NPeaIjY2ODrSjh+kqZ80c5Cwoz+QhejTeT4AXZWyOsqH/
OWe2QaoyTkcaqaYQ0iOUu0ZH602I0k0IvPHD8wZgpp1XeeJx+Z5PA+0jJduQQ9tM
IMEUE7S5dCAytJiawDaH8tssvZ4ArajPnEcjgmO+725XqhI3JSEL5bhRwZKzqlhx
KtrE4gOSvoCDnzX7ZkfWrm0T77B9agfKjchWf3BcePgMB2ZU0CMWLuJRyKwHyvdD
H7Wk9wrvA6p9dI5NKbZ8E9xDRGQxNx7zi3oWC1NTYbLnIMsAqj4hBBFNeiedFCpQ
oPugZFvNSGvKI5hzbaOusrwfbLU1LHOwPM8MBeL0Xmc6F4ykOAlZpJp0VGmfBcoS
RfUlsvfw1hFbwKjcUZmusdlrM4S99SfV3kdZfnGWMhITtcdCGzWXgm6CYliZxSG/
aMU6/HGu8GVFn9tvtT74PG9YofqbQGqJqk/6jZR1DLmsEcdiDfkDJGl5bAxwgE7j
LnUmb25s5GvdJK82hrDV7oClFIW+rOrXn1I8WeMCvc34YXfQ5Ye4C1UTxSXNb7Pt
sb3uV4zRH1DjP04J+FLlL9KV0UBOp32ZH9WreKxeTamMfhMWgASNULWn2P295nza
Cm6jPBgyDXHlaw0SBGa6HEaTrUw+BdYDCyY+OuUzwkgouh6S6LAm/54lqRuo6A1u
hzADM1lX9ngyJx2oqKR+0XgRljk0MUUfZkcZotKcrUI9pvS3E7HFtVSdo09447Ak
D7ydxmRgH5gEMxjk8nF7EQ/U68xjiEMRfG9ZHPK1aW/ASLibW9FW6ZH4MSYgCsGW
L3N2c+xynOEv6LWnL0iMy+4+xnk/OunFdFX7PZfcweUvRKMGQNhDcof2sw3Cv98m
HWvu75sgo3NLvf8/7Sn2uqSNEzoHcm08N1d/Jfr2BJjCR2hVlspeda5w/BnwscCF
Yl6gk8ipNYr01lXue0UsZA9RW5BYwQZjzemqhBzXWn9bOwdfXhDnBjJMbUm1TigD
XkZrgLkgCrWJ9go7Q+EnB3i0NJAhBPNJEJSZj34Mncz4GCq4vEOj6k5f6JOxoOuw
3Y3kFTv/WqZhra9BMr6471cS72yoCm6OXePm6wn8uXu81yIMFkdwLUxSdAtokk/p
dYknx9AMA3j77EpuZ64kgf0nPKByXHSjmnLZUGpid3+wJm85P9sdr1ycEFD2JTro
HjI++5GOqIF4au1SmIQ4PHPoUd756noK2Se0RC2qWOOPM/rE1DrsQ92oAVztKRFC
xmLWgocae4pSRaZ8sjEC5ofuG0f5HLp3eQHJaUeEC0n4/8UNOg1HonM2c6QKqETE
P2PQucSGHxVsI9z95RtZ1bebpp9Am3AqxoLD6I8vNFD62DHHRiofXEXgFgJWF/ur
wRz+lmwwRKWOO1ElccGse4OIIo++lqhvYATdfkM44BlXJrwIsUPYa96MGU6UEsa6
oj4KGu2TH2rz/jUapO5fdc2Fhi2yGl0glzdNJ7SbluyjGFgO6ce8uwsKoewl8OiM
mXY0y4H0YFzAjQKkW+NxMlsP719hrfhfRL+Fjse71ixwj+4c4noAGQPOitfWmNm6
AurBkAdVGs6zPqc4uRBNHYy/pxnF1OqCpR0ZBA/WJAz6OVZkvyldc4qDp/WW3UJl
Qr7r5KMFe5/nddW5Ocgc7q/ElmPW5818tSTP0e1+B8wuoLWg8cekOdES7Ff0IAl1
zhgAXGX6/3omr/Uehb5B97xdRj4NtrwLOc+/9pBMOVLso9ZSqCMq2TRcyRZVsw5V
Ns7+Gf0yoTfcbHKWG/sV8HAV+fUaOgX1l2vkf/WD4uJNRw9n7HUo3EgfbN3+RPL5
B3zKAa/0cDTsmE5ek5K8krHcpRZLRRfZ5SDpb//FA7nEHbE8cv8ZE+Ur/DqN3g9q
Mg/QK2yuVLSdNbC8fUZ30BD3S4l3a9iKgntQFVGs7vMsfoZRgJ8PFSNEiWT3Lqes
0/5NeoahoaBBQHChfnwWXs7zUoH4MitQ46aypH5LCiHkXoYe2glS7StrpM5dQ1+a
H70Lo9bKf77wHKEei11NfOlGhKy66fekQeaH99O1Vvbam4TzttpSUiq5N45Vz4Er
ew/ZhlPmidskhW5HjYDzZqWw3ePMlRKyUK/JGBWEbPUgkSlgXAYvSun3gbJP9Wnk
IaM9qV0sJDZCqN8SBLqsfWM4YbZrGL1yQ9nDej38ZAAsX8QD9L4sq6U+qf2bmqOE
a3HKTVwjHd4G6lXoZcXBwQUPBi7BeIAsuS5zfNcUSpq6hPaacPQcA+W6+QG9og40
D14xY/nVypstMm74YR62Jkvo/XOqhXxWlVWx7L74oZ13PPhgP3q1796SA894GeY/
HsUQqwEwRGXobH1poV+am5R+yZJle+8NZe9bE8gIxFfNjykGq/5vmftsRtGXhsMJ
p/V5mHcBTPR6mR1LzgBAsBEfRPImJfDEvbH//yMgY3aZyMnXzWDTgEdGPNJfOD+N
OJPgj0LgzekJKzQhTRzao0vYBDUUqjcUqMZT6pNbcsfS/EQHWRPZ7jfESbgtfaJW
mjYu8RlkGKjvUVWy+eRVqTVn+Gj2OjemJ75exnSQKizD0OVd2fwOKFiDBrlyvhD+
Mhcz9LHVT8Gcn8oMxmU2UKthnl9vIT9aX61VcwoNQkFm8IFSBLLlrUOoCBBYbBDX
zyF1LwrsMw+AqcdeXjIaK/8a6SqgRa+fKpmEN9VMeRGnk6/N4NFvGW3MTUdzIBbC
Pg/pByCNxmXklE90qlFmE/5cvhA90vuFCYCeQDeFC2eV8oZZNkUcAH714IvgF4r7
kUf//XyEcUKCGkhecvDfVDhuFL/CWOoEsMvNtQ4H2yOzFvjKw97pvftDMq2ZaW/X
Y9Jm3wqxdkH21qUZbEUa4tlgTRZUFUp9TZjV8W2vaZNT+jwyxYoig+vU8u+GUXx6
sNZEznUSNFLyFVQk90rYH00Wxb8kRYh3HEM75o5o1Fqoko1CtdullJJkWEvNOe2f
sejMnA2BOS3yPdkDZ+7B1logcT4LVoh/a1CFWu8ujDZIwagPUwsXyEKOZMVCW59Q
/P3LM+2Io6q+lrS7S1j91dq5iPOcyqH00EWkSBuAkoDUqxwrEbjrlDYVobB6+au0
l0aI8G/btdEt2EeAhaTIrnjXKgYzXSeAuEfd5Jp9+XVcSqZ3bL/4PW+E2N1whdKE
hScmYgp2xgR9EE4wcKoEj1vNQsU76xAabelyE/dZy1bocYSONB8rqKHRF0SpjIyi
D1+UBi1XohhJ2hqMo0kCG8sfxGlXKUMxThANAp3qLKcEEQWBXOXn/AKivWZYoREW
IjEVQa9KLy5Rk+XoPYLB4u574EDxcJnmYvAQI1Dg4HBCeeO/ts3Rr1rHCoGDyt4n
4ePTevmP9hXYr3YX6xNFP/2pwwrHKu2b/neoSAhG9kzlMd6k9/kk+jkIadtUX21V
DaQzm45o5Z7hBtvfSFSbErfn2Yyr9KtetDfGh9lnDCF9kCteddj3Tbg89rO3Ufn5
zIntNDvRG8NyBJsNgOphqEJZ0fXdxBkdXyL9UCU31S0eGy4aQ8F4yaS7PQVQc3SB
Wxslc/+tRYsvQ6KRknM3yxsjxhD9VGIJuyk4SA5VdmsrrTTvRzHFkfu0SSWhh67h
Sv6PSM2ah6oEtTPX9MIZ12k0a+62T80yxgVx90RckDDnNvkEVtgeGwqTuUa51RSl
qvbfXir2LHw8kVXu9AR+suZc5nGP5fUmTo4/fpDWbeN84iiPlQE1IF/bEp4w1qIQ
7rTgMeicoXGSsCYZczxaCfVLaOlNUnMcCRrfil2sVmT/+aWbzgpgmr8CdLI/QOw1
wTUP6x875Jsg4vHkiG8ISRz318lDum5kwV0GF0Z85M6YCViWmYjKEzJxJmUwNu8y
Ykx/6WSfMIrHd7QtSK9FPNix/XM0SNhMN1x7J2OabQQXDf/VwJSsR8xIW73qTDtv
i6ERApEYUegAhjxu06a8qx8nRjxwIR0xpUQeXKibQkQd0E7xKT7nb/H2mI4t+zfk
ECux0Pt5tdmS0WQpheNPurozVGlsz9C5B1wrmnyjWXa1W5wHLmXQCEMbatGnVbnG
1BvXzQCOvfPpMJywVR/bJELddmWSnfeVbZ8kFTTg3ns5SZZ4S+f6ASjnYTry6J1i
IzV4Q8Ppb90oWAcZdYTHLN96veyk8xVz2sck9PhP8yXvJzu4byn37YXPu9RT36RJ
wkrtG28ADam+XT57fjgH6ghI2dwl04zCU61W/ajx5G1Dg6HqB91fZIOfXhea7fQj
TSoYjEthzbPpAJxKrk5Cc4002MMJD+xHoP3Q7VjHIAI0U4hwF86TSrDIG269Q7lZ
GoaZC/IUNgVG31fCy4khLqhJ5ZlCFywk+uGDfes924Mae/NhvtVjOWL3AUCa5RWp
KOdB1cqAy0zXDSD/ehF75YxL2cON3rvr//6yRF4NyOT/qdWxhZLQGlyfoP/hE21h
72ehr8UzDme8HhqzEw98lCwJ1ot+FCD525/cbfPtTFBMwcYCUlimKOqPAYYNoi3Z
ZexveFtkUYYeGszavdr+rHnqXbClP/8wr9iXB8uZS1vOcdVm54fCpuXX8+XQgxjh
5I6lk+yAzaeEZn11eqFDawLIumjmIQGoNbcS23p9fmoVYflXdZIZfbRy5VFj+PRE
ZAHegjdum28tfrg7mlYv55qbl76jSsZtgQhxlvCbCRJigcp/AnUtWbkbbgxc74pD
CGtcK/I9uoOMW8TiUrtH3GEWazReYgVXkIKWUiUSGKeKrZuNZPWhwiYktCLJrAfy
YYkjU3FUhhghnHiSildOAGfgqNFh6k2gS645J1r2O2NwTgCEh9dMmqxQHHCJm2Tc
D0Uz+fVwdIWW5KZ9D3vs4d/UMYFC331xJeO9RdXGMJTp6h8AzYL8/ZrBuhZiaVHH
hG8+yispEzo0I8kR6/x1mraaMeli/9S6aC/+SDH0uE5XtfyPnuzTe1nVKKeWtnOF
monZUI99EmC7p3aLPVJNoTtNrJsA9K4jYY0+exY+gFZc7s11yAOMcbc2wtFqo2Lj
Eomki1DwqF0z8l1KtH2rX7OjhdCbYxnvCFJSp0jxPOb+Fpb3Nf4S61IA65U7JS/u
4dma516Ly2QvsryDnFUNkyA7OxCJc8LEtYRViW73xJOra+6Rh1xHPa5Ilvne4MiE
ipGGc84i8VQCyPxiMp2ieqMjChgh+brn2qwllh5v+CYlogg2N1Z+oZWq+AUO1krJ
69sOsNbMZFX+IvYVETFpkMWhiDv7fuA34JTa6WqxQgTlI82pvJoo9pJaz+nTzLnv
H0iy7tDHkr3C4e/PylYaI/llG4ZnDsu/i3liUuSNNybJhDiVkV7/57kCaOW2Ek7R
9OwqUN9rBKopHu7Xy8UI84zC8lcZB4xAl7Zwlv0h5s6O0IWmD0hPPjzux4UHVWaj
B8uOPpWrwWDB9S6cX3BFipYHg4iI1JSIk2yZEitebix2mt0cpTh4njKjsBcAvEwu
ZwUCiWBVRDEhQgQw93L2pe3UsAn5AgH/de6javSCmUwdNKnr4le+wSqLXB49zo4m
x8QkQ0fSZW4e38BQFKkFKt8jqbidv3KJcV6/so5KOffxGaD/EJVBeOkq9qzDbih7
LLtDTXdukJ7QseeCoLhbC8T5am07OqFmvVwpO/y1/plpxICSy6dXFNFz4N+6cyuK
4qC3ImATRNcS4y3TWYvcZUjfy6XGJNEepgh9rrn945Ic8VE3y7AG9gFTniqwibUk
tzOKKU7K2I+bYwT4zardkmdpcAzecf8UgjCkf49G0F9K4FwdEBWKf+auoFsD+jyy
RvVhMiUSaNpA9Hgxqp9ScVwUdfDh4GoXw6SJoHhtE8nQktkbtB6tVL99biTSKYzQ
lCFDOMnm54svdOtlTx7NB5v5ak5VtGYckhHIqnIO2QoY2AYZBTCminBEOeegeQZq
bqZM5UdiNCZVnK2CgBn+2hL68quiFWpSYWyCtccMio9qV+5yHoN7eEDqgw6rMvBZ
PzfZRa7i7ImsH266sUnyMDsw5mFYf6i4hUzLHbtV2dJ3pRTYuJKoN/kwzEcC8vqz
kWVL5Q7cpGDr0Xv/iD/BJtX++E1U8rRXynEbta3nr3QyOYVE9DiCtnY2F6Kg5tBG
Ql8qL9Bcyco11+nUdAu3bJmRa4/MWQzt3F9tOejF3a4CkRsLrzGazBuPXhXSknVs
c7MmHUhwP5QLh12E5cyzmvLwGbujwxHxBJ/EbdeAzX5LlPYa2BudiZStx1xx9MbC
P0wQJhlsD422rSCWZo5W5lCRMGnHrpWrT2GbhXWbKNpgRvHiEMBh/KC5Dc2xgwGA
7yX+FeLHFcXCExyGFJMWka8NRJV9bkqFs7HrbtS/jwlwWCOap/LU3AT23Qrul3Hh
ksVmSa+rrwiPkAfAg1DbZkj8dYTMA1+lY6sO/jSHqqzsrOa9IdOt6e7mwV+Rgz0/
ARNoE5czZl3gHHHr+HvNr9Wvl7JTXCOhIOZaTrg93330KzQS153X+kuaH/kDHi6j
JleG8nSy3ZJSaWcpcUwOF2SSrwhkcCIQ3WjlZLLKLe+7X9Ct6QuRrojE5yNvfgSr
ICycXm4EVBzYq25FD0QsuHfDBfoz+pOkdlT87y2lZwYxF6p+L3XDfA4Ui1zy3P8g
ngulVo0IsKmJaVDC+UPTsYCerXlcAxMZG5yge4cKCAcwb0yq0ek4QSMFVmstmRIp
6O1kB86MDRNU0/8CTd2lGzHWuuH37dQFc8IuU177UPetOyE+UZ0QzXL1E7XCNHYb
mtu5nEuTLFRkn6E+W+OBZJ/udnNcwmdUYjgSAOsG0QHchFeABFw3Ge0JjMx6EvSM
r26fr7oFCqkYL4Grgnli0Od8+HpVXgtiAWUApugS5N27o3i+MjIf5+jSy6pxCmQI
MbXg7tlsMvWJ97Lb2kLoTUZ2fLh24HWP13wTf37OGlD5CoFYbNiQ2loQbJWSxUAk
k5Gp9Oo8p3UhnqDDuberWTiNRSt5+KqWtCNYNJDUUquxZsxMUAbH9NUHa19sPkLA
Vp1tJyWgNQhzgTuQ6qk4+4J4LIry2NRBfK4xiTBOQICxVQX32y/roxjIOvvpM6Ie
jjzzVhaX8nBpTaP5z/3Oi/a0Hr/lpI2twX4OGLkwa+MfcQHQG2P19s4HLFdvrNHT
ib5suyCe0mK7yxdQPJWcfx+HLmohVlXwzPa+h1AjfLG+TLDwsBh7twS4ibnv9GQb
ndvqxfkfORJsIbRyXpOEBTWXq2K7PamXFv33nECv5DNbmiMjciD8ml5yShpeYQ2p
/ZTmE8XJHj0m/RcTFuNd1c+d6wYq2GNZ/ob4dVOj8HRd1dVaKrs+nrHMIFwPiw3o
JggDEQqFl4U3YY37jIIDgT79ngaARBsxflKQQn46Om/igfgYQP+PQN9GmGn/REG6
2t5YAbTjiBKQZizUH//Mw2nre32UT7qUpIui9a7XbNcDIMDtgN/YxYmGpAqgle6d
QhKmwQxrn5ykxHVbhqQOAFC4517vhvR0/wLBQddmILmJlQ8tE3S2BCo5snloPVa9
pS89HfS7El/EBTVJCPUpvUuTVL82OOZcmcfIR86X3iXwiLc/0sQlwDdd70FpxHxT
dNm8efhQnY4Qd3c1p94uyOosU5MzYOjakjtRmJ9KluzT7IMcMK7VZ0wfFnkCwcnS
4SWaiSN/mFhms+HzytfAA+Mwovr31pwtp5NxdDUsfsfIMv9Ead0qAWDf6+20YJxa
l98duJwcPfkZPpcaKis4GyD8XxhqD2ROazDRFAC59tQpA318ENUFRfXHO0NOo/vy
iar9K8BALtRlh36dWKPNkfiH4rV38xiAe7E+Ste2FHQInIJFdRax0bCc1zpEXW6O
QpCwFYzJ9IN4WmiBqUfSE9nX7ktmt1afQnwLAWejnIQmelrkxaqdPQpSdyePHs4B
EVg5hpmTShUq/SisERoh2CdXRuvPW4v51wkb6+S4ZvtmyRfdqy128TFiEZ9Ecsh+
4B5oWSDc1iQ4EwMZea2V6ZlF4cuSyhkUsR5JoWZzkyhhGGbLrzEZaIilIh+fVe/B
cs9M8dUDN32cvXKQjW/d4RcRPJJSYpuNZyghNFsYR3w/+wz6VWHnjN2uBw7Tg+AJ
p4d98x+nuZMmCosxnNnuldraE7PXSzDUbiuoi01YTx+IIjqf/Zg9apHs8FZNg9Cs
S0wRB+WR/YetdnMKi1V+mHcROM81YfBCeUZC4b+5zbR/fO39AqnoYUDajgBUkCe8
LjzgThBvB9QlVkB7beg740Rsv0tLrFd9JFyQNbbV5ctGhrEApa4RYvx2uZzCOdvY
aPjoq8D2n+ZpDc4CyUubwPk/1F34MDd5L9PAcWzupFPBjRP3awqx+KCZOQPvp7d9
Q5NuryLaFqUpu4FPZph5Wpa7dbUeCj9lu4SbLhywOeu941IU/UuwOLqBnKshB9dI
UOrNhhtWPy56Q371FzDQ9wuz7wZuk5HvUoQ/R6oN/AtbN+ZIaMsKrCMOOaMj0CbA
9yBD6o8Xa4zDM6jPRnRy3iUyQdPnf/pVgIRo/FqUw2So/c3m4HUXoI9eMVGheM4i
uxuCaABqY1HXYwZQsTH5PcANlwS6K2s/pqn/diDnFTOHoLuIiaDgFk8j6ZjkiKJP
EYff+SUmM+7qMjSJZfxHofhMrUezXQpKOX+5hcTkYkTfFV3DTOTC/hpYlsLKiDMk
TmhjeIdotOtd3hJzdUTxC+9dD4aq6zR/X7eFHr/oqbBBqFcPV124MQBNtKihXbG1
HRvGu7ntx5TFWVbI7XbbdI9ZTOPD3DSuQoJ5gVRYJgTMbUgBwOT8b8v5uxxgCkp5
1RNoMowLWNAx4Xh+oJ9VB6op9KPzPEJPbyKcWYNiEoahamAzQs/XyjsfCSchLCty
2wd81d5qAyKV7Z1hmh+weGr9I+qbYu1JoRfDQE37yd2//AYeqJ2ZMfC5CuzEMpEs
nNxi6tMPnDdYsx2RlX0LjqDYHF2YfYskhHqLAr4AWqlmdn9lDm0LclGspzmGhAbc
RXgIYPafzhg/sjsa0bjyZUAxSQGKD7zH9GA0UK0JTGJ+IUEB7fAgBHyrHXONKWnO
5gVksJ5vLFV99IG93awfVbqDQ8Yc7L+/TV3KqbYLJI/Wb9YBUkxdmvRaUduSqnzf
eT5GcnIsgYzNHTfNOzRXvQbZgLNxtvtNEWp8aFdt2dglwA6FRf9RZT1Vm61lodPw
h0UaTBzBIjOZKIwXGE+/lpeWnagk+H1LJt7GdNFvCnWN4SAMyW/GuEpt3/QasH8p
c8BQTJLg9R2Mc7+u5tmPBZ+wU2Y3sKUanIIk3Ep4w9sOpdloVyKI/pYO+juVwkns
iXhCqIAnI0N7BXVYsUCdcKzomvdVfWvTaZuXqI5euO1aowoLTUv5z7W8qtJFawwu
kh4bHawbRXxF4IpGmbgYv7Kab8szeNuEZPoJN/k0z8CFJreYOZcP65MKN6aCcslj
KBXsKF+IsEPm6/If4iMLjtOQncR7TcRVgTwtTF7IYucAflFXNAz8dYr9uv/ctW8L
EyCnMBd7bO7jXsWQJnxVX/+YD5fzf657KGiWOgkbcgB8/DPuGdPPtzCSYsvubAwQ
NvNkR45r9d2bJKPl5a5hGazMwTzo7mwnQzUDmgLVMyrPqbH0xKi4GW5kasX81vlk
Hf+WkgeHboZQ+JKC5XRnKsxJF+FvMI2j9OTPzZD44ix23MF2DudReliuP7+LcBBG
ZJbJcjdT/za6qdKjS3PoQYfhpzdsPVVMC10I2/SCtOtFNn3Cr6rL+JqX27JtkxRl
qm7OId3IEAyMz02MMO7CrIu7ofau04bwH6zrwKRh23lsWsPTnuQWYEHCDMYOG0E5
sQYIt1DtxPvIBkd+hM/cnJmn5lNRjPULAFCaD4HDamSkHy8qspDT/lSWZE2DDxwX
wkWgO8RlDprDgwJ9qs00yYSpB4c7EVF3Okp4IfA0RS9+7mD0EPMiunV8U2kBN7qv
`protect end_protected
