// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Zh2LSGVFuLY8RRWMyW1mDG9D5kSuA3O3XADrTn1b1lWpxUlnZYSIu1AplAb1HcEG
L47NNivTUiH8FDYQrJN0gZzcY2UpSH21nzWKqNiVQnZ3FnJWiRhKovwXA7ViRlS1
wRARnBlBvzMy2LDhXmAtKrug/2DLvgCI63GfkrDZfTWaz/Bu6DqNhQ==
//pragma protect end_key_block
//pragma protect digest_block
XrrCv4D0wPbt1O/IuUW1GKll7qE=
//pragma protect end_digest_block
//pragma protect data_block
JoQvlxt6BDLsQfGrmDablahmBNXanWebI4KN2498VbFRytt6bs7Z6BsCuICjCn1u
9JuL9yvYfGiV2MKjY1Iz4I+JgtZ+6ImLTG+Q2FA8fX7GWyWJVJgNDCOXAQ2CvdnQ
PietYNLRVLNz4uf4cbRUKlxkaExG8QdodLRP1qAaToJsws/wRd0U5jLmD7mQPnvc
dI0Lm2YA3RCxbWRkV3lw8qwutx3uDZ/ZlE860C2OZNwn9dHPjDGIQOrmxuefvHOp
iA7YwTAEB2CyZGhZoT8pLduv1WqOIV+HLn5qUQMPhzjuRRdoLeXWkI6zoK4KO70B
cjEBk4KZ4vOwv+sLEKPPrCD8AhnJwcbQqbr33oi6UxXap/m7s7FRFHtVZI8c1I6I
ZLfG3j7LFwt7lp2dtJ6R8qYm5Gop5cbg2Ypg8tTvHVanhR4pZXfAbbswNUYYXYKw
qP0EgWENEy7f6YuhvfVIMFh4p41WIyk0k2k+NkFvZXXcTrwJeKIfokNqOKB1e3/n
9a6nG4qVk8tC1ZLf5z/6Bbw1SXnVjkqwzMmPGz4dqRLhQWlrJd/CJza3FHeyM+yG
4xCXpBG9op5OiHB9Viidla57jfFestx/5jgQqr8cH4HRz+yZ2lwvwe0nF+aiw/Gj
TOOLpOy8OPJ18wdh0ZvLU4ayfu0t1jYghJf6cSPQkUMb+7ChulXplKz5dobfXIJB
s5QxBqykZbPJW3Vk6gmTYSUbMs1xxWO/5cQbgXJoq8OpTBpkqV4JqniW8pTKGQq1
dEy99Tk7b5h8rhlTuKTWaISDSElWcFmWD4IHm2uDt1PBv21vAobnhiPnu8OPgG29
jwlb6vwk05unHQOi61LRDDqh4wx5bCeAxDIljLEZlRbaIYjp0wv/6/HsVm8QThX7
MiJeagiQmm1iV65776dg/bp1FlQ3ykkM3IZ3crshbWT270lQWE3RdWlOjogjxC4i
UW75sJEMi8pM1/yuv4YKsB0Vmc4nQ++OGnz6m57Dn5orTj4iFl9IUboKxtQhnFei
owFIOshF/As8gL5njrNAK+pI8rOJZ2ZPNjLfrQl25Ij7ZMWFQI4UssFw7uzrsvzl
elMkHu/VAigI2WvqIgZKR2CzDgOkNwy+Bn6sAd5ITiwED9vfjYGW5mCLubsfTpgi
sASIG43oJdSJUHbGNYOj9FN21ZccgnGdbJNiHx4qopNTPqGbMR4jn2wKgXAx24+y
TrGYWxAtlzGJWOTSLGk11z3E91CYT//nz9+XDBG7yTsF5yypKqNmgHPw/Mpovo2I
+yXMCZuztUYqHV4ylIWlPqEVssqgNTWf5tD3Ipv9VQTYQoIUsKlKdX318MWr8vo9
MEZ90vVv52HZV9OVLQBPbxJwK9RcEGaYh2XbkteS/TGZEcPi97yVgHDfSJNGYmhF
rdW5BzaKaAO7+2TFgy80Ns9bXZezZ+Rr18JZIXgu6HBLX21YNKIzhOSdl0+MwDU0
Lhq6yVisC+qR4P8xQJR916pUZZJK8hnkEAHYq7BQHQmFC0x3rA82hUf9iDLqtnG8
La6OH/QbLrl5HnZIJazH2mmSc5X/ZR1s1z/52vpqZX4c36NMmkTSSOQZE6slQjN3
+4mzJXKy1z4etDKQB+3tqzHFJuaUhBaYcFUqGuoDpKXTEI7D7DS2Q+uzMAau8rlY
nu7+iyNd9/4RM89wS6OWKAxVtSW1vSyK29syjwLa5aQRo5GAejfq7LKUtd21b2xw
KfX/e22Nj05Co55y8YFlnMJE2/EPouvqO5RaB8o196SRoUVRaG5fKsMr1XXO/XYg
sKBI9620LWbe5zcbnGXNabgVHXswKiwWU1YyrpEyaTJSd+2SxxrYDSQtOyoH8aS1
cgKAQ38qFpzA8nJtC8JUdFLjyOY+7NhggDcYeXEb78Zc0sPjVg06BeR2af6xDNAq
GYt0pLOw3wF0D2GRogL0bHRdh6FsH70M7hi8hMS39JNP6GmDKCKBdEuR1lb/m9Kv
Q6DglLbuZVneT1+n07b9OtyYiRCq91w5AjROReKbzbb3u3wvovvTIXc2PMPp1k+O
5FcyxHUpmtRUNAstebIpia3GwgyykY6FJksWsdlucENAT6jkYShCjWF1mxuF0WOh
RlmF4/pjpful2oRB5ASI5VNLsFqkB8dMPT1znlck2G0NGxEyaB6OkhGyYxLKzZz7
CFaRxguVlKvAvFzJOhHJzwMMM77niBcbsTLCyHMqykSoWPda2s86G7fMufbDUKjR
/q/qGXcRdtQ3jzqBIWtB0WTMHMSg3MLDxe3I7eHn0iEettn7Mfv5OEF4yARexnLT
rHJY/EWAvkcDAHghnf0Kt9fYkYf5KVfeO1AFgFLkSebtEdZugVfVt9UGFAjxmhZa
jiIk58EAa6XlYbCT5RttSikvfa4MSrY73GtBr7IorOFM2X0fdhdzdj0bXPRsMc6X
zrOzZyf/dNmtVdwvi4xMEGXH5z2DjqjUqYrYe7V0rWZNjjcVV9S1vwpdd8+eIaxF
95+7GEPGKpjF4aGuyG98V8ssGrTqBwWjRVJBcXaEl5w85ej2WhiMxuhBMXhJiumX
SK6PaZnPr/AzuBZY/9SAB4b2kDMwU5zrZ0yCFVz7Ji7Z1L/ndyhW6Eh1a/a9Vn3P
ZMuWD13SSgN1r0TqVv9GG0h/t/nfnEN0T05GJNmNc6OAzc9o3oKXagJTmB5WlUFK
LZkMlbu8QaB9b01zXnGVNwXqfimLIFnJUY6f4CsxVCMbommTS/SZGtauEN3eilbB
Hf9ee+FJE99mWP+3jDoWIhR+hhg7xTJaXaEx18cexu3AEfbev7hsw/jmhhWwKxU/
YIVxo+RD6k+1kA7YlEk4cbpP0F5r+tmBRyNjNKGivNmNAX13TiVPYIrUfscJSOxZ
8p/u57DU9JWRnidkLdFLdYTrrzzyMd7xRtt/RJ331A+vaybkiV0P9jdzVfdMiCba
hcQKbuWeBF7kARqseBkYt6OeyQeaTK/VyMvj4aNKXLzFBed0EVtrXHSy24XJR4Nz
NN3Vu3wSzNi5mU/NQti38uzOHSKFQNMvyxaAVRMCYdFbi0+K1QFUGfNSgSUwGJFV
TVR8/a9us5IALwCt4bZLzpuKSSVbkY3E89vt3aW4pUliH8uachlPMUdS61A5s3SP
+qPa29zWeAZaa9aEZTcX6PXztiDQPfm4ZpVZ4plUaWyFrsODl2srMzV/NYIvhGkt
mx7dHJ4CFwEEphJs8PkkLjVeSWZXNAREI7S2idBF0J/kAOINKvh4U4PzreHV7IX6
M7MOBuh92IvV1u/eTMRPPEHV1WTWEWjgl9dldsUbhzFBg8dVToEvux7wHrO5OEST
X0zTlqHWbaKYx40gp3Npo9jHfLq9Sjs9XRTnb9F05MuYx0YXy6HgM9gG6e4wxbf4
Ckw3oLiOb+Ke/KSu2N0SphmzGvP4+3diz+oc8gE+wflrnd29qsZdATQGNGHb+gfa
L6NCBEJzyXHO7JJ6S5uuuAfn+C4GKI8dY378xLLN72Oy//JWEN1KUd7a9CGwuGMR
+Pc8MzzBvpZNN3hRKNFNhwbsL9+2VxJKAkuGk1KH9sAYMKqHTFumJr2nJEFQLY1r
TwlD4NupkQcr/pVHBNAwWV4lGtVABSB3g/U+QOxAAzJtS9xbhH++lLhM6z+3fXbU
7r+ibaX/sxcpd+MikbM8sRKlZrluelukMq6knu0RSw8RcU+A30Cy9tY/MaKFkHRr
wRrcxTcYPpih7NNjuDcbjZNDz+YSr7AfrNNDlTKGI8qLENsC5oxLPMwuQbjfXOUV
CAsv+c/ckhWhRvF8QvwwYgHxKMr+3nUGcjdr+6qX8S8A5SIS/s15w+KFE1iwWjT1
EPq87vuX7vf390w0g9ArcoR54e+RgMNVKqwJSydaz1Fx1FxgHcqtn53Qur3h/x02
aGZJCTZRycWj9Y6DC78h7JwVrhYBQqG2VUuGz4HWZEa51bP/kXCmSXZkal+23nHf
V2sBIWmO9KxRMDAGJkfdBLG/FuKcD7cLnIpFJ5E0iL+kbfeCgD4Vv0vOmGjXHEtN
EBv14pRbr38dccgw5Mu4FV9jUQdzomlynG9/vE4B85MFB2a9PbXpfNKNFTtHMsmu
9guTkOxIaCwLXqia9nJoTE8/n2OZFCMj1JrG0n3J22hZ+d4P0nXjtTvqY5XChA7o
Nhh1X3S5pRwoJ5V3UQzurzwIBbniWrqCDGqi9Z+pPZlj3eG1VGj6++LyImOLhEcQ
lkLD5ffK6Z0o5jf7PFpB/SmXsFGHUVZDWUXtnnIE4VrpwwXgaopxz156Bc4ooCys
4xfyfFtG8tPPt8hdoL+UkIJR4NeAKlydOsBluZ1LLRHdBCvyyMhRuO6o8tpw4Lyy
3VbETdvoXYgSzsCwt5tqJMsUIND0v7dGXulEkQIbP0m6aXpsw5Nmgp8+RquJtp1O
2ZTD6BSQ+6TMHBuJXXaWEVGvdNCCiPclIe8skVsYlAsPkPEkZ02MVDkkIsActOBz
m9scOZEXgjMeeD+61r6i643xDA28gaYgelYyhskDlYS3Nz8siOo6BGYNPSNHXXZe
QiiNfN8n7o1rUPU/p2CD79FQOwmy/fa3QHIK9JlS79UFtx0Ph3bHVFAUc2dTq3wm
mbXMb1fXkp6B3sjF2KKnUMyVbbAHUIlMYEIhNGJFbmtG+dA1cV1lSNzhyEpVVgh9
X9tl9UGOtr+AZ2QdB1pF2NgElaZ0R9CpkQj3RUVzEBjBVmWvn4/X6xvjKW9RM+Vk
yRcpDMtjGJ5aOlwGtyQTZULRFgh735cIYMPr2z2dkZQyhwKSk5iBB11TKuwc57lZ
oXAQbdnJUddBNxGkXOTp+JQBWwcfBVFH7qTO1mMn0RkH4yvyaDRtGeBhlu8N+kYs
UDyub72fKaxBF6h/mh4Yx8BlLx3dIBJNDGm7YZmKm4QCiRYc/5ZaiswKWUQ8QJgk
vRCVLxsA9wcIv5bghfA+XsNfI+zfvtYHzleZQ4VsktYc/O8rmU3n0WL/x/G3r54Q
K+WUz0Pr7O5wbQ7P8tmeZbsv+g+DpfK2d5IkNsVscjwbqk4j3wAve0VQxrvMT5m+
WIICTtts/uBcT6C8kC50zbgIvXQw1D+KocH7x6aP+b7r9YuBeKu7/I9wGd2FBgd3
hNrZO48R3zvkOy7sqnHOMWZj03m6J9hrSL8+/1LeicNF4bvlvq9OHR1IhP7HiglR
PY7E/RIqIe2O7eLu6lkJeyvcCB2EG7bErKzZWi2GNxVHyw8sYsG351YxP20N7p5c
5+YLRNKtrzy5OK20GAxpdbi0J2B2NTJwN99QQfm2L/f9Ydh+obcWDiqNvIU3nB8L
+/46cmdau26UxgezMM/KX5a9Hy208rOUqsRIiXuXBGSuIDJqr9YtsKq7wlB0Vzlj
B9nXC3pMvg1W6qrz0uFnuXc12dv/xKXdGmlU6v3LzD65Ndfb7k14KVBSzH8qQ1TO
EAsGQ0eS1/skvqwp7zDw30ERhCdpZ9Hjl6MipvfpCRnVszSydYGT7RXv7qTEwCm9
RqfCZXUHtl+ypC/eRrWS1UGj6o6Tw4XQrpMneVlVRs+egGbS/NuwUuf6xhFUNom8
pJRlfODToqfw+2oY2xqwu3midzwq4qDykhk2Oycqr85mzZF3zSRmnTD49hVgBPBG
fpU3+AqChtrCOPZfBna5T8c5dBxgEEm5CqibKvexgXDhVXKsAOsnPcJOAuXwDQLl
IuPG+n+cCDTohJ2TxUSQt4zu5vYfd6xfvxYJw/pzSeRFTsOVD7za1dB79SjK+c+/
fm0U6M67csCoRnr2bJO0mOM7i88gC8ylideZP7S7yMTbdddbJJfEFDWSdUrmO+o4
ndGczQLFg8N7zbDWwIBkXm9ivx6j/3B/Lok/TRW9tMWlJx2Jb2prOhvbajgQM0JQ
3iBlsp3ni+XXQuTRVsSXkOoS6rFxN/1VRukalR4EoPb9l5o6+tcwocDkJtCMV9mL
csKPSe7oMmyQ54v8d1vsYxa78t6c4IXZ3+4HFmS2TAankrbtQHgThPsJaEISgeCl
ZAD2XZ21qgeBPh0JAIJDPKegV7FGoc2JYscFkCc3BQ2Ym6pQEMlvoj00BqHoqV6g
fv7QnsM9jetlBGqJfnX5NUSW4uMHBkh2EvS+zvWClI9U9emxzMsZVZBb31BDQTFs
N9Qn1pOF4+nFQ7SAQR9oUsvJ4w0INEmFE1xT7q4X1eBc539U1Xu0XdWOQfDh+FeD
BEMauYlY+1M/GwJecs33kVCoX8dw7Pj+JyH792l+41bs6P4+eSAtaULq4B6ufmbi
bbbZtmxZKc0s4zw+ZQ10JAmiQ19KL1ytlHmnnzs8NRZfYe5StQBWB0qgSV0o+6ra
M0A8Gx8bsio0T1J/wCCMGlflYz6ihr4OgsRy3sSjq580/3eTbHeHSV0P5+UGzdtB
A210VWNMTygbx+/AomvM+Hzj1xfFBKpFjZuDt9HMeqjBTtJ+WnF2hinisIaay4X0
kV6JqCxYbUOhrJqAh2+rSfXxxY/F1SCJ+rE91fipcWpJ1v4mriqs0PVWtva6IBN5
QklGC76qJERuccx+MA+U8dYKmXo7gHlIrdQRbZckRkwkIcaAN2ArPBFWExYsVdLq
+qlnrNkf9GUJ1CeqbHUTTASFgHGiTArrcEISw3DByuyo+6JM+kXcxbDH2mBGAS+p
H72wMS5+PKJu23yymlMf52LoKjKCex2/dN2L0nTuUQExn6D0+zVeWSLZk8Tv/0YV
Tg3Tdd9+kcPpLbdMOu7v5Aq66dZ8uRKBM/5Q4pALwKpu/7Xby0fxe5X2Uzr3keCx
jUN87hV7WQmulIytZQvhmN8dKzWTLegHNYd6SUIcCmHw6kQ09F9LlBUaL56a9yl/
DLDvjXSfx41IPFo4JziQ5GSXDlxZsgbA54RJ1znddnMBSH8vVLjMtyJDxMnnNEMT
OWYoFSVJnG0u/ECFAKqDDtpQEoyu9EYb07rJbIIsPDdQp+H2c0wHhn+9jsSvdM2F
hrkpAB82+uuou+QU/SBaIPZSEzjrCBBYP/S/BByFJfDjTdPmoGyd/plZhPipsW4B
76/fRVoscV95o/VS6ApMdZEoNuGi7dAXr5vVl6ofigp5b2Z3vBxLnaiZxeLnmzZp
5FKfAnhjG6lRIYNZdSJ4Vtt1AduxdymutE+3itRVad8z08D1qDzx1B0hYjTfoWFP
anYSy3kRjJGnVkAfLt9pes4t1Gm8uKQcVsTCblvpOIitjYH+jEr6qXZxRmCr5sB8
+C5nOY9rtvLDsRBMGG2x3uQJR0mVJp4OFTGHubn08JHa+mmW0clfGUjVQdNKQWNs
ZYxnrC2MYEZ+uxnXFh03tkFG8yyJZRKUd3bY3ovoLEBp6r+zd8gByvFNUDdBLblv
eC2oKkt9pOL76Z5NdwDMl4sRjnaFOQCeuW3JeuerjLSb20FPONAaX9DIQ7frnljb
AIhTmnDhQNVTfJa00eSFATtO3ZfwHO3ei5/s9O035wxCTik5DW1ed3H/Q9f6YlXg
Rck84O/1Ujkiy1NzbOhA3SKij2B4wBqd2X9sM1X7GdmqDEOUmbHbf/JefzetQ6Lc
fXzz1qAZFsoEYj6PnsZj9ET9nmhdGeTZha3/5lobPq+Z9WAhrCoBzbeiDYVUnSZf
y+7Q0KWEz0AQBGv4DzfGNBiXLtS7d4lf/RP/W3Eca8GIHC06goNg2nu6CQ+oEuMN
7ZxYTK+2L7JQKBXQTsMA2HFS5Du5+FGQqM42lPgU1GOSTuQRNHDVu+qSmKULzozf
tBFVNn9UhYWSOScQxj7N/HciTMljrgZwBX16Wz/+f4gs41no3vJW1ZGGO4eVpcLy
VjomkEkLD3alPX5BJ7P2dxiqFyTg+1wQYqNE6M0BczPqQHZdbSmRkGEMYp8gOMRa
nok4mzhrvk+Neg1wvXnda5Rv7yv9KZkbbEmAqdt19ESq3ynA9mgNBOu4C4sLMEqP
gj2Kauaj5E2S+AQrtZEnNciqtxzD9psXVM00eBGEahBQR0IYJfezKTSIE/p7AREd
SNbXlWrp80NNGwdNM/n02bvOHBWJuV8Vo42h4F+mVrv10SQBrNECh/t43RCDlzUy
O5m1dbFUb1tdOndh2Vn1Q79bXOgUJ/fbkBZilNWn6qubpBxQM4atv27CL39jqjKr
H5tZXuiSc92E35wPOk5x35xcmyNBThc8LmSJt60kZ2+lzrMB1zioh7oPpzsLvpzW
JnRO5B8Vu0UqRvQsiXUaXqjDBw5OG+l6OTSjx1r10nIh+dZolIbSfLHPJCHjxxAG
ptPNJi0VQRWPChE2ehSkC+1n9vXyniuBTXWy8/DJpiw1WXIry2LQ9dS9XPXuMLK6
knwUAKdJJgU9l5TP6owU2LT+Z1DNXvKMFWcbF2Yi5tVlnE/EfuWN1iixotGXIN30
E6XtM2fPvfZxyGp59C0NzgzUM7+XQX/elMAqPGPk5+Uk3fr+dJIMDwdSf9uCP9S7
vmDTeLQ7M13GE8dGctrCDeQVLlS21ST829k3IVHyEMEUXBfcwp6irIQoO+Kbb2KD
nPAQ4znnKFWiFulCXYsNsgJZ29KCxh2sPUHSY9GchfzJe0dBFubhlsGItjajjPd7
tcr4Y+ln7+3BUtckoAE4VRBsEYqNtE5GHNxOwhR1LtlSk0PNffLujtgjWvNoGUxN
qdWx3sBqHJ15j73us7Mo+z+ekAnnLCQxam0xr1+XIN0yyxm9JfLcxLeJkwv6BvXS
B3YOkaaoiuJeviQZtB571avOveixpifSpSAOr9gY1hKK9cPx5f5IcAc6Jh6+QuDv
7SY4XsSERimopXDu+Qv8/LUlXC2g6QXvpmAlnWH6f2UCGRz+1TmyuBeB7p8lf9MY
0OHbYkLuFfa5Xi2jtd7lByVgJZp+u7NDC+ZPDzyK7CawtQwaVSJv/v+rz8w1FAYB
i2Qg9Lsmt99KCPxJAKpt9n4Y/UYSRPL2wA+rYzIm77X7ovAfnk5rWnFuFgMw/c7e
gUj3Q58P0rOrIZ66Ckp9Kcv9RcKcMQPRo4tii7RzEA4QJbjk4c2qdYrj0H5hcGrB
we/Jky7eJgNa6sf3ZFcafKusTxRfUG7wulG1I3Z+gZOWEm0bznD0/n9f/RqWUQxR
y4nEfV1Ksvb61pxa0U8U3nkFUdt5EaPlFdzkfceKozBLR8BgKEn6ute+Rj5Gtgo+
GstHXrs0Pq3epkoMVwMPvyTE76y3BWl26hei5BbPYD2MCat0A3BzziJ5rOwyeRTN
ug4MDqc3NpkrA/D9j6HJ1SQzs/GOZXJZObaMTmtAntRfDyNi7WIhtUpr82IyGTyj
I7eW/QPrv/f25pCH/SM54/YgD0AHyJkBj0w1LPAbFERcD4kqjAavfu/itRvRVkJZ
p0+v2TrRjLjQFlzQkohsormNNM+6X0FlKhNbkwBvUAm9A/QrL8Z9zG8jzp5xkaVs
iRB07bJtzA4KUGuvv8h4U7wFCAl7mqiXdFHYpu4PmLbPWgg5pBZyUbt1HwAUHxZJ
nyaBwVsoX7VVaIsf4FVKz4nfHSwMQMJlPbal/ZAP3OrB0poUh7LT8DrOqSakBt0x
99TS9W/3CT36Z8NNVNT/yMdUxxOHE3nM2Yf5ImFOpGOHqjpKOA+PXxUIXoSdKVQk
5j+xxYqfB2clV5+WKjP9JUMFpk1fN7ah+W71FNqaubqmYNuzZwINm1cIlZST/lbv
gMaqW1bMHA11Ts2jfomf4medeVZK0JOd0TagexYhf4FQIqnrId8u0CsZlPW3qLl0
zuGeXILJa7u4xzeTYx6jmdnQQvBb4uouhjKFBAGe3zwpvFoVu4s/e3U3oVG/G+fD
omFqLZXaITucb430yOGoCgs9Qto2sFwfGEff98su8Qj/Y0h4vgN2tx0Fczsho5zi
9LhFjp6uCFuuLWCrtN4Uc6x2znlSBFwhelZ63/DXzaYTYQtwxUrRM7fUTRv0QBr7
Iq0v7/a700kuv+kc2GqqUv//tgvZ9Hc062e0GadQDKyRE2PVYcjLxu4mtuujOHCJ
4ILi+h3St7L4LQjjTPW+TAAEpsSSTjPpmqQGbiFXVCGWQ3Q2vlPsniXj6cxOJMt2
3zGgc3/10PbJ2vp/Gm8xEZUD/Qsy7FcnaOjXQbIV8Tz0RqkWQZmljksPxWH5fxUP
H/filoZHRl3o4A5pH5PV9aqIwTWVhl+58lauc5U24AKikM/p6+/5Tmab3UcY6wpL
pcBxEbDnmmlSQ2YJPN2ApPeMr5bup72umocsHxbU6YkEi/ZK3xRGLHMq/0hdpTQW
nE1dq4ezJXS2TjtYnrUsrsFIe+YLpu9J54ePCjulE9s801D3yNmzoCZEd5RK6oes
aJ5WyYIfGyFwDiYxZgUlS+DXR9Nq1zRt5sbXnVhNtWCK0WP3QsLMIEAqhnn+jexj
BI+m6wySOjE/ffgsKrRBRL9Y2JbctCtWbeTZMszIbcR+365IprrBY0U4Iu77dZ7w
J5dceO9zS0pl3NJpIiZu3rU6h8T9af3fkh3Kq+b2+7PcaFWK8rQwiH9iaLj1RM5L
nggOcZ1wqBl4RVHBtDNF/0VcicD7dHREHujT3qNx6NZuPkd27BqdjHst0EiTbKc3
3oJMHpq+L7G1xO67D8p3gSQR8wri4K27rCdvXGNbbKu9BMqR1hcnNsGmNh879Q2m
6KDxibgbJm88QiHEWZGHzSnLAMNZHrzfN+zlr+eY8tebuttWTmWTE0pfN8rm2IWH
jjA8by0QMOhyHiaYOd1iS4EalmZaXJm/YQFwEDR1Dgxw6OHYf+4feYY+vmfRQWfm
ZkDg4wP6h5eUlJv7wmnRT3XXIV6Wja/A2z0yfsP9w/Igu5gSJmTFwo9KWtOQAdsX
BU+AD7cWgIS1lE9jE5174u3G3ATvw8iJ/IsWY73JM5HzVZ42O4IedSfoKWmPI148
xkSVYpgKvoLncQmuzmHI8fmxNguCJoPElljoYq+Sny9DM8EfW6PS+5MBoVBC9Djb
GjOQohAH7SiPEYbc/jNv5IxqjLY7/Js/qYNDrQglZHmCDzlWKtmLDa/jxR0usGGx
fEYnaUa6ZYVmEoBrNKZ1mLQpA//BKNhPTQYV8QtIF7ALmpv6Tg5Ogbl7kSeVqX0f
xuheRmp8Xnr5sEVKK5xnnoxVTMPWJuNA/IWKw4YpB/xv4xvnVerW3jZTQwAUdQ12
0ZkkqF4Dxvf4Hzwuq2c82DnTGyZIQdDAR8ewcsXec/h89Q476Oz/1XSNbl7pxXKz
p3OHIGFWBN+GfTvU4UHqglrtR+Sonv3aWIAKh83BRjAmXvUl0HlUnCB2UrQDil4A
cK4yrujvz5kiq5mFznqJt/a6sKdsz3rRUqQCao45+24FChKbkx4spYZPVn+pehuQ
F0JJii/3kqE1LCIjz6U9ruMJoqoFTnqSBWlOdr35v3fnTzoqJ5DArOGDEBTFTyov
6l4PJI+ujFNbRulbcSi0fdsllEnK1SxS/X9yWcYOssSxKs5uhNDdMMtpsikhH4aD
m3EVztmtVArlQnP8SvUtE1FMBwrojHlZymOYboMWdvXsDySywUzHcVIub9WEV91w
jYOdLh6Wp5uOg+OsL5IQ7TbJc3afps2O39kIv9ZT9/o7tU7irVh1vK9XCrRzpRlM
lwebZp1i1ZMdv5momshE+HSsdf7Y6UQOH0Ljnl1Z417NseKqQNpsJjXYSDPcvB0W
rr++Nk7IzUjjCEug7q+/yuQab52osVOLg/sLFmXHzD0S0vUz+saPyAD3mjGVNPLA
J+TkphIKDzz6WrJHJxSQielnItdkEvpBSTu7ChT61VrlHlc5jzSru+yTt4zIsQA7
znlZZt2XLkVlCJ98SE9FHZ1wJMC5euEcIgZuK2B3OB7LsO1gcgDHLukTzLv0qYFK
dESDkOAnus7O/9iEcpTUerWdVxlihindq4I3GYfMk2maXRt6SkNPoYPJTwiag5vp
oKDAeHAOBXEPh4EVcLzyaD6oyNEooRrdMAc1WPseKdC8V30udQWs98LrGvW/y/n6
dSUnJLXr9xg+woAv7doMbODj4qE6m3/PH1mVaNdEzKDn9opErTrSLbesYPqSfzJK
4VbIe4S/fQb7aVm/EWAWfbMiTfT5xILZ/tfnyZVrG/3EJJj9vjv89nPw+xpcBArY
nXxKRAi/Jas2ofgG3mg60bLnWcDmceqhQaIEXo06QAJhf3CSHKeYEqnv33pKfPwC
1jqbUVAo4moeBq3kTpZy6fPZecA7Q1zFhA0T6ugb8QdUDYZ3dhPDunynHu9PsXjH
Si5txr993qGkjznXE5yka1LGHXhSQtZgLS8p+OYpoQbMo9j9wfkzIPH3Ra3P4Ct1
xumEG6tEZCavgkl/Ewss92dD+R8s8iR/tAXlFCjECfLYFpms5MsGaJVQMyCUfbrE
EzoeeeTMHP1yqPYy+BEZjxngXSUpuZ32+CzvDb11tkEy6OkDHsAm/xXC3Qp3zblf
Quvt6rB+Hft0LDIfDHG0gR+BFrTUC4DPYjq1lhIbIMr33crQVjBUx/Cp9AL0oc7j
r8dn7swORb8xEHYQSfdlajbyOVe2MvdCzTaKMOA3IO0gNyy2udwQJqihetPzwgMJ
zG4fK7B6yoWoIB+Fyp8AMDmr9+tfK806ndpD4E0bIE1+NkY0r355AMFHf7rU3IXj
tb+ZMoJYxd4Jm8/Vid7gJfC/Ei/hT/gkEHczE3MAXNgm2ImUxM/bmTSZUmWoxKFM
z5v1dWKlC5CCrN/y9CrfsgZiGYKGQ36wxfYVO1wMeCPo0xbYsVN48juC27gSJOYb
SmTz/ePbb43/5hZYimsZNF0guiJN05C8XU/odbc2OeUabzKuXbmHPl2CWgxkMNqM
Y+uQOse1d+PVX1iSO4Q9W9xKVYwr7kQ7RHWX092rUGei12yvEnx075U7tt+VpqT1
b8E+wJczy6TUBZ+8okWEbhOPFCz7S5hJLxaTL1h4BVWSO4XPizhOrjieAbhqU89+
5dk8cTrEx+eQyxa6ROpyacVBCSWY6Z5UuomcEr47uTm3a2YUjrpzHPhJOygFB2Fn
UJUZx1l0GlTKGurvsazgzNeRp3RGP3/6ZluwfJdE8yI+jmzd2kEalXz7q+XO2XQ8
5crWfmRjzrDlvbiUX2EcfZt9g58B1wFU1/dQ5MgH2znz/Vq/q5QCK2LMHusezHjI
eg27KywSoBhKO/8Nw9ChBUQREj+hTnBiR3IbypeJqqWI3DN5r15nMMEU0XBtqW4Y
TgF7tFTBcBQFJtFHxkyJVtn8Cs0JnWxoTIUbj+zshvKMRLRmUsPnMlvBn8w08fM/
Hm4crX2rIpde1LdqOGZ16V7hpEEchjphYTXAExcMex/nW6BP0ewQe5I4AeQGwirP
h6JucfFyE8+DuBHcVYaaR5YR8OBCa+Yrd/NssBMXuQzTBT3m9UBHIoacZgg44spp
FHlHDA9n+qhG6hZXbehLAmgm0C5Ym+yZ4wiTh/6rd9NJ78ZShbg3FCAxMu6I6wiY
UqtteeUOTETLFEl0HjXUOV5XNbDzEcRl1IhdONJKw9Y7i8LS4Ez/7ls9qvGsirb7
b7xcdOptuvh9l2EXortbAunJBm1woyChKDtjYPR0p9Fyp0svoTs2uwplS6+FWw0z
UfRqqzIAyl90F6kj46SWG5J/oFaKbhAWp+uzJ7vGAXKrb80VAH1fMHM+IaRKgfbQ
CavFBt9GVcAsmG9IvmxcFsdesC/LGBs7MJ6dgdpoJNM0tDoHreptITuTAdm/COWA
rQEi/iGKy/Id96qJ7bdoH1yumYetiaT/FGQ9M8UMKoxiin1icVfIP1bM27BuLNfU
+k4YcEo9E59lcnEKRdNFh7sdDz4ml34ecmFWRBeB+w/zlH3o8fkCo66O//7oRdhw
KN1xWKyS1poson+2f5mvlfy0Hlxj7+Dwk+8qmMFhwleuOZ3KxMwV+Vi7pdq/a/Hu
H2MFT4Yv+jrjtRdhy065hP+jpzd5DuZW577QCk2GC26kxyFEZTX6I5p/mub4Ci2L
+95B1VC3QpyTLNVGLV0VSDqlf4/WcQ0+cdF3JFXIBbvRoojRej+oEu+5nWK78IVL
FwtRiqcvd2xcaXSUlT6U/2zvM24hOjDGyZW2X9BT19wgWYJppStxE+hvM69IvbeW
N+HDi7Ai0Kxnir7Arf/3T3wlrXxQiuWqrJlWYV+kxrBHxGv0gfL3xi/OnzGBbSqi
Ien829uURavgtDYZ++u4cmj+GBt9B3wz59HFJ8LmshucD1Yjq2PiRW0abtQNKLT5
oaAGe6JyJ8IxpytNT8GMXueCwpRXqZbqVEtAQrIlQaqhVfciDTha7rlyro0KAX8H
RpFjVmr0ywr/p+vkyL1ukI2Nzo9/Hq5HQdxEjbM3GK5Ra+EzLf7Gja/gz1b3v2YD
6N6om9cKfhhFDpla1nw20AV7+9o8PbEArNwdFcC0sZM7mracFnPp2LAR8q/JLuQN
5NRcc2ZQ7Pq4ej3JFuqjyT0Q+C/xsgZBDINiYaqTiKvhAc3C9iFE5QBPgbLwNJH3
f4A26055r8nSZ3cK5RaVmHAYaljv3sRXAjXQv+2HMN64wKpK+onHYAtcP0nT2eHK
JltEoh4x9nS6RFMG64qgbALiJ4v0tDdCAroHDSkNHbYjLVWhxGxNS9SByF/gbhtW
2+tnmYErp8mpAGpZdVa3D6NhsnkqKp+m0D1biEebxpmWPpHV7QWghZH3u81Srnge
2OkUp/EPBToyiZLrgIgkNeffZmvPuAhCZOvP/Gk8jD6dgWZzosnPxk+v9rxT9brn
qDSOQ1hMfrcBNsf1oa5BSi9ALveZFb1mhr1ljkP83N40TcPkP1EzqB343zDma+0x

//pragma protect end_data_block
//pragma protect digest_block
266fhzxNI51Vbs7jZjay+OIHtLk=
//pragma protect end_digest_block
//pragma protect end_protected
