-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
tsmfd2NdcBiQPzNM74axdT8FvUGgF4qGPAF28MN0mf+huGzQ8MrPKEmGKWIrJxLG
U4ruKx2D/eThrm6fP6MhUEUF4JrF93xhRsj/R1TFVATFY3hZzmZOC5fRB77J/aaW
VYUUlfXYasK8GxCpFPjgCK5s/v6WQqgMGKnea2HP4Ww=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24112)
`protect data_block
rfQ/dGI521s947gjWR/RubuAdy2O4//0RScq3qBBTQygZifRUzKYdj3K8C7kxLIC
p++jePN1ZumGhkXAnEpMeXnYkFfsZ04xyKv3nVUHpsq8nTYVCsVJdB4Z091+bEYz
4FBLCS8qyB54ul33X+WRzbYhuRvjJIc+Q5QZ4OWKkC/fVhhesjo7xQccxtW/yAA0
S+lkgJw4rYePg5UIv0+7456U4wAzViy4dS1RsgraGPQH2mK1QB+v69neJGgAfVIh
yK/y6WBPR9ZjPi62Rw5BZ79QFDEf7kBxuF8N/Xk6TKkVtGPKeIDRteIknBmPJ6xV
kHFOiTy+O61Nz03+qMTauVgkvdgQsRRhs6koJXMH693ef61kg+haFtlI7Y0/24Y4
booY1Z9bOe9dfDmmNzFlqr5g5s2a6nmMow9STHFzwtI+5rSjVNZ+nbjBhoRVIPPa
EBsMSoeZ8XQC3D6mrxyZfAaE70ykJ8dmd00yqERcEHjKHKSlf9+FaznLMueMN5wu
HFHUVkc5y9Ov1icAG1jP+BWmocl9wGZC/pZtRnzI4VzzUGTYNLMLz2XRJOhx3cdR
9Dui1P2H7TYa9M7AQten+3SfsgRAqFBUx6shBHM6NOo1GQTZbrbUiWck0aKiKMWR
s4w93pD/tMsxwnR0hz5jVPtuxbC8WRfhG7Vz+hS3JWFSAdC/EYwPO/6rhFIy2o6q
QVK6LJERhgmmGfEStfNlvXeYzsaOXSEdAarlevgVHgLEP92BBC0RhfOZMRb4Ojbn
nIRKiYCV75CD6J5dauEcYrahilpGYYKKzghI7buOVLwrW4Oy2Z9T0ete4dXfkTZt
d6227Sd2dFcgdA6FVBL9XeJZMa/FuOEthgLFdklkkd4mkUkXGTfJOdvRQCkcERsp
iZll5VcLPGGwVp15Nh/kewzMOtGKdpgkPlyeMpSJxcW7UAup6CY3p5UjbMf8oNgx
aSmI7vyKEhF5jt5nn2Mc8mwB8/XZESKMM/5FadfW13PGEcINxFSnOsk3K9Wp4O6U
ZOuRLVSf1v4hiF+cHlLASzhGw3AQylMKeg3//sqPtISH5/zI7Wl7q1j2jsmLdjv0
21O7WivuTCzFKFeW/P4lBIC3QMWPehnnwtFZVzPzV0lklerj2BkeZhQ+Juhql4z2
qDCCV4O4B4d048hnAj1KGnUnf+j2WxkqnyoBy7tcHF1PHdSmH4IVq8hQwn8xq6k7
CUW3pk9uAUA+TMBBXRI9kaRJXx9640mHPIdarM1k66SUMjPH/M17ynJZkHevDdn5
nWTWCHuGgdprx0GR7Oqu1og0j7ZEhH8fzqFkxoySHtRsXfyGQZyS6+oefbBP3qU3
gAoo3CSUm++plH2u/0jO4E7Fj/efhAVtH+Ks1ddFpzpxmxh74KAnbfdSArXjyBoP
6dCP349D7IpLsRjJZ5Lj+KPATajoQia9egq0+UX8nxRJu0XOyLbuEVvj8G4zkn9J
cEPVZgWOdQp6JmPldH0bmlHYX6/CNPT+ub2sbQznCCchqUvjBuhGJ2Triis/mDsa
W7XAl4JpBjsfYnMyQoTaomtFmVTluPj3UX4/3FNORhfAADQbxZ/Pu3nGuXvQJqs8
FsqYC1HQrGhIFAbNp8qcBHKtgOirsELZYkhyHw+s0F/PnOUHcX+WyZYUyDbhZk1b
MBiONQGG4QC2SSYLdGyZMHMq9FBiqWvD1daKEIrHTxi6u0t2PJmQDGcWE92NHrsD
TjWcfaF6uTcw3WcWksxINxVHZTSw4y0H8Lrle+76VKPq2pcNtgTwqIJ/RWOsm12B
hDKmwr9Zqpj/X4CI4S2vIPx17P4ZA9D6MS9/CBpr3ITpRRt7NLqweXyIpG6g47je
f86EtR3Er6EAtqDcTg0CufXJf8yQXOH+u4cdWEx4ZGEUbmRvNDJVOdtOmbJrohPR
AAGRfiHybjfGyLnlf/Ywx+y+JiWRpUu9LH1FgAk/ETmfnwraRc2c2y6goKOJL0rH
zccbVuaKKL5Pma4VeFkIh9F2Vyz9QHFnq8q2eVZLfSPvWCF7LaE2DxZ5ul19cBgC
PndvwaX9f1gYjNYpnI24jFUidQL0nKqxzNI3tlafOcYmyGpiqL+NGEjA/LZsHhWM
retLFALWB4CN23fi/N0XqllAUq2iY2CirOZgb1TyX/zwFbyzLIT0q8NHb9z/+4db
y53B0VAZ+Lc1nghB5n+LPR0x8SSsjls6j/dbvXgfA0YanXbuw9v1goW6nhf+W5Ua
Jor9XyOo5jOhUeTDmpATiH86wkiXs4Udpqn0LH1CCblWbqz/gFH+oNFiiNPqu4qy
PAWc87SgFxBQV4G/m/06gJGEb+vnGm8QAFBScqjzgNQgZC9u+TEOqBH2pm9mHEUa
RJdx0WTGGkvKEqgKOPuR2oK/rQWXYGCl7EYuD3zSLFbG35EaYP328rF/3rsoi7Xs
2tComkBCoDKHp+nMbtt47Hv47neblAwqTSKie5gdm29j+yARKLZUFjit8LDD/tm6
+l0HHQzMsaAIHhZ5y+qbZmVTU0zLWNDTURO6Fm4YQhn9FQ7I4GlqRgoKGWelr7Gf
Opiax3bocXoO6mJ6U41BMNjdmVKlux382rlOppUIHMgvsHT6FYdZCaRxkMZOY4I0
td5B0GIiBWjMGnmrFfdvddl3jiKOTfxUNpeEwzyNwfNZb/jjQX77tnEZlhP641u/
zFPIxX77Y86EOI07j7LILx/Vr0fYfzhBGdk4P+ZtgAjdu1rq/ePSXIEbP/+Pbzko
pFD/SMdO9PbytCsX/0RhRw7x21W5nQZPCCezQa/6mmQ1mzKUHaqrCajgWOOsXwvp
ivdu0JuNA/L36dfroA3F1MZBxl9m5tmLsBBI6nqdG1GNEDYg6l3gH5T1O6YF/9xX
Ag8vgQuxbpcqNXJpQbrcYmYsVdXAlJuJSS4ohUxnHj2L4JI6ZtY3vtKH+fmdUuSM
r3l/KjtJneFR/SC84mPfE1qNM6mKSe5Y7PWFjnC75PyntxfSFunvTuyW2KYnus5f
BXqoW8I8On/EpZ7xadhRwCUpoZenGCzeEnhudX78b6TlwTor45Pe8P8Oq241i5Dr
fHimDzR2+Xp1jEvODOAkoJ0Uz4O5nbJjCgpQofhxf7IgQPpyshatMffDfbMNPpA8
edegMxKYSnuewLWjM8FNpbBiV04lbWlBt+73AtwFOSMYgf/FwY02ZYHrjwF5c/38
3lrjJdG0LZgLwUY+gv/dwGk2bDbkIrptL3RmMvufE7jvHBlaGjXwmCWIM/YhQhcH
uC9zXnjc1LbHFses+buz8yjljNyglOKcJkEaPYXuyjiEsuAtV59lOrqlQNXhSjVy
0sfdXrGCcvGawypBSU5LK/h7TTAEvb/p7M1xXRcZi4DKTCqOXRoAxR+zeOjg9p5H
MmIwfAF+gMezrwoaqtJ6xVfh0Iftx6MA6hO2jVLnD+JfPk6SLzGaKvLFKIWHtC0P
QKrjIC+a8QKW9E7tz1Mu8Qx5bmpDaz0QDVnjBfu1Y273Songzu/Y6OQ7uSLzPRpH
ukzeHa3QY6CCBpShY+ZzYTTRG3ncAi/fA4k9zr9xv3fxIZmGs06oNycikNlm3A/O
RxpHphYHP3RbA7xMarXiOMFUGR+Xp84SqdfwR+UpkAa0jzfXANwCJW3g5CZxcBRf
VdhvnwMj4cPZGUo+wVtwJ/81XycEX0KXUFh8lXjMsW3FBx6ANnUMr3di+U9mdZuw
MlltN4CZk6c9UuOUOyaACDZPLyjll/h69/Mj7eCYUuLTR9qROUSMwoSH/L9iShPF
dU6Q0qPUEnVgJAJsB9XCTjbr0ymOtz5V6l4IvMiZvoFZDgYQlMqjRF9ciZBNOkXo
Pil0oQMMcQUlTY3bZ2H0pIJp671HLn2Oa+TpwfNCr3JEcgDozjuuHOqcRHVnv1JM
hgEHhWL1TAv8W7Pf6QmjcDFD8C3ESJLl9RspF15HkuInLeb35NZO+Lit4/AiMGSD
F9E1I+7MIxiLLgNteiSu9J1TIZGHA/APVlqTfETuDOuiArshYlZls2V6vJhtc0Wm
365E+gk0ULKC9VLzheWUft1YEKhL5ZzOSP+Y78MWMvmn90eHDTNvolNaNaAWf0tm
nE1BKGLYxZ7yfe09Lq0+zbPy6rthGxyK/0xzL1Mx8DTU/C0biM3ojihy4EmxCm0f
Hc7IH2H/BfbpDV57/m8zFDETTFZVsemPDAd3bouGmQrOFQFGJU9lvfEDI5wZ84kz
geM5JwHdihKfuuLs+gHy+at4fLLpv4iJH/SJH4HN9s3y2yY4H17ONDR01vlQ1xXX
zmoz+EGqn771ptNV0losRNRpSKz1B+FvTBBDVMpMVMATKDx4l+TOFHv2nPwPR3z5
4xYM9/EgiNSlHB0C9zFlKBCUM627HBgTi9Lttdjxswrx0qTyCH2czqkLrhDms6+s
0Rv9OguRDU7bnj0yIdpMSqxx/1cxA/mlditdTieagWdNhVgGhJaStqCIYqsQlMBq
JgaZ0dEKmcnHR0ocKxUoqWpItZCQkbyo/JcJTmqMQCbNpFcADd6/uKC6fwhn1B0y
ZmrDwB0YoorF508RuV6oqTIo+4uC0QEE9+ig0sdyRMg/sW3nK6+eU25mEjtZz+7N
M+Jk7YlLSKXM8CHJdyuA0a4o6R72lNoRwZZlFpP+D2/lfimqZkXORnsEtR25UIlC
JhbpXwa42hkj2EWxKgQcbzlDv3pwauej4125KqWtJw69nIFzPoRrB7lhl3LuJ3A0
57+cIUAaRYITlVa8Cer+3miyf0HwLJA0HYyftXyBmBiNr1hRWJZPdlXPcnl/lWf4
zTYuVVLuKpTcUL/E/u4B8MXtHlSOUvoPf0Y5Qi9n/3p9vfjSSroO99YZveFY0s5J
+aKEnbow8BDhDQBIJ0ze3FrG36W+fZmlksdN5pFek9U12qBeUTmc/FeX7Ml6peLf
kGgPLRQ2q2MXMLAAwLeXd/xylk0MOlBQkFWXu19YxhrPr1rrvRy6ob3asUBsEnBP
SzKBmyhQnVz9CL3rpVRPzJWQq9g8b6enhYOx55ByWeN5FDq6lRodwznTFWYxfK4O
/0UA22Ng1YOLqGsVkJu0xQvA8dFHAQTuAn6NMIbtS8Ahi4aM/3PF2RTBH5w+yQrX
P9FBCElZujFKaxKywOCCe2u21GHVNt4igi9sZJUEZKOVGLQhO9txP5jkEEj2qOep
J2HGpH05finQkT/C+Wh1wlAricI4QeQODKYekeHpivvi0aT5kCU/ZTUb3mIJsbi5
wijH/aQBABSYVOi6axlNazFU/dL0rx7uf0xtpS4iPfwO5RV9yL5PKtnPDCaf6kPw
sqPtFFvLfyIPDmFqtGspAK4X0jji6CVWqlbl/9Lv0gOeWzVUs71K7v7YAxbn9/hP
DOGQbI6KBZnTa+yDeOYHgPbE9YISH3/dcUrWQBM6zztwYNy60eo22AXFcCLtw/qb
Dd03PMN4sGvJgDaKXXxru+juFDlfWEvWDXO7CIhpD/C1BeZQC9UBaiaY/6arnAP5
G2EGVwLPpoa5aagI0ma+zlJG5ybYeFudPgFTwrXT7mYnm3R8YdlPcULq92f1uJIk
whbmw7ixlQkUoh6wg4B1VR5rTr5dAdCjjj8wR2L1CVoAE55PrdDGSdoZ1QXwpcT+
dEb9OeZpVlN9nxZBirhmKbZ5imqMdVilnS3V7RxX1x9Dk0ejOkUd+XhddzhuEbxP
3mqkP0rXRZyiNjx7lXgBZwO3WuVTdKwCM3/weduWa083WmpO15HFhMSS/JKlNIQG
q0yiGS1PyU53kZfXEpDnU8irC7XVCkh+zrWGh4doJ3zjcVI2ea7HR9CXoNETWsYG
65DThm0kj+hR7+aXp3YrxjeXvaddKR8ft9HdVhFJqVXZbimmmJzyqU9gQCKqZJ7a
VMeazprqPm7lW8Y61IdPeeGYszMKfDSh4O/DDPgPA7GJXea4i+bF2Y5s16MONVJi
SeAaQmKvj1aVKtruwAtX0TriRcWENY376npJaCxZeNW1UatN/BTJBgcvXEWugD1+
F1XJYE64+m7R+9xvzx6U7U5ade5rdxhV7rXkTKXjTArYxIeR7SsPj/oEcyAd9iMY
merPNlpUxkne7ZnX6A2nZ2P+lCufSI8joo65aZcuMmdfZcICDkjKK2jSgWJRVCdU
J6s5UDmnff5HnTkOChVoTswudACnmvyXj95Kvi3KAutDyjnWbeDuwaIuc1WG4FON
ZEHSK1QqHeM2NGJDI5wa1p4joNtWDpWzoDydHevKnIoc4IprRoBDIXKhtiyKA/K8
gX/VjE3zAmK/UujJ/mwENZatNspqCE0ULLzrfjoyDr40/vYmUvIhbNq/U/2p0Eqx
N0fmcj4ej0w3bqrY123Czn1q/p3oRSonXCHwkXtRrWa8Iflc/gPMnqaNea1/fNsR
7GqVE23lIA3yjNkMVQA8aA0Ft+uc+JmEaFJ7jHNKopmba9prE5kk+UfWW0IComdW
FioBrAqrj8N9txUwMtegh2oxJu4yUBnpIjfBm2QcdUmMHJGZfl0OjereHQRMV3M/
N8zC/ui17xdukjJtdYoJgxM1vahDl9IxayUyyGw2bSVtb/vqUICqeQmQEN+d/+DU
tA39WObEkygG8j6a1Fr/snoNSEPb4KDeHRPOvbtePlo6MSUehe2g6sURNwhJ68KU
OKFF2pZ6lfQQ3E6DvhY/b+3Q/KtDrNn9AdQ+0o/oyXoUgpv1tXi5sl08c9YmgHdK
X6Ix3ii09wqEs/Bowho6R02z1iVMWGEiekl1mNDCq7r+8hpETHDnc8s6EoHWKuPA
8+oMUCpj8epq6qGcIuYdGiEvzCMBzxLLnJe6FPCTAA+13A6d0LrnfrhpxaUYuBwB
WRfILavJhOhdfWCl7LlaRb9IE6jIfPqYSJ0z/nq8L1FdIqtU9cuirnaKVQ7wAnWL
fUtXfX1+6n0VOd0n8lQHiEO5jJA8A1sLCgQQV28pO3OHLgoF8x9oTjAsv3l7Pwcv
2XpwQYTZX9snGWTudTAUHbNssMwL/VHc+q4Zzm04iaNNZ9VlR2om3leHe+FZJiBi
TFvLKZTyoVHYSit9mgZRDXTwvBfAFdmZTMz57Liaotu0SIQo5Fd/uAPveh6ymvKE
BTyz6qoM5pJXZh0K/c/FHAcoq0el9hX95Zx8gkfI7AzxgvdRzvLz9e+r7/GmIDUh
ZoDxXpXxOmKj8ioAOZOG/jtypVw51enJCgVRuZsO5PhLgT12HcrF0XKHwNrcExux
UkLlvqtAxI9x/TEhy/1g2ufdm1trPOl04bqjJ34IWNg/p+7hs7pnrv7UyYxxVFQV
4w0bfBVv/g0pFSIG3o/9Lrir77Ubp0lXRDnvC1wF36E0HrnzulmV+AAThoL1QSRn
zqLBJJe4p3xqb/JvvNGCXhYR+oFaDZz4xhwVeSgsWx/fSI2LeOubLEEWf2cLzFQT
jijReVRTMrT4SIdO+eIqeGgTYGuWaNtZ2R4eprCFrCRL72QPAX54FfKNPFLZuoxO
bK6lk73a54VpSHfKurhU+yYrR2CAsL5dBRHjFb4N0gAUVyL5KEX0t127tpEU28r8
KfblEVLI2UgNpdiGkHZL9DYqhEKFE1tHeT5KQUNX0BhecAA4QRBpZN1gQcobzN7b
qku+fT3/RBzO2Eu5HHmQ5T4eHkzlGlwWrwWpnVWGO2UYCPVr5svfWUIgqOxoxCba
G2oZF+ZWkenhJHIioLIGhiqzxd31gaEidFxgEVaZh+aIZYQ4JQAq+Ud/qRgdsUVN
UP3GKDz2+f7U32dHXXAsfpDJMFQoGIu2O9+QQ01IiD59sUOOT9jmPsZL27XA5hY/
7Vi3/MMxAZPNemNJcZ21GTehFLCMD6BjOjqRiZhqdK63WJkunRmipnAljpuSrc9h
7V/KUwJSszTEuS8XPjWK/QXpjrvI6o78h7kzD4bpq3VUUgdT7+Xo/NEefs23NwvJ
GR28FkLkIw3fz3zNMTLmZjXe2Pda/+Gy/VTA6jLMy+vFiWAl6LVC2S3fm17zPhLz
0Zb/PID0gXAiAZmu583tmBCvhfGp2hZdafpKeBot/1wLKA3ttNEV+MFFHsmdL3II
+7T1zDs6lkUv2Fett2MLzZZHxvOEJuW8o2us55NQwZaaEG3QCwhwy128ILkB0uaN
zdt9t3JOKCNjkbjHZ35MToT5Ptove3p1Uhu8UpwGL0ZiR6hffVZCZa1PprxToLYw
lkRRKuDhl8uFJe9WAKOq84Az1LpElx45z0d7APRK1/QbWZ0cqlLYh/3GXnIGcDJx
xcvK7ooWJuFGd0vfBakiNI8mPSmbTaYt4b5V5sSHJsenhDAoP4ehsxBkJ3y0bV4d
+pP7m/a2cdmBhRkFxVSL/QpBriCbUh19QlN0H132BWKqN8oSNhrROySSCWKFCIEP
KnWANli4hXj9DuCFBlydOZIpZ9++L6Bc31ZFP3NttlhJtJT37HheLUgK4fXaFNLS
tTATpru2sl/MVCZvVsdUMj5nEgaQzslFryAooH2Ux5nIdnUYcfZ0YCIbeH1SnVFk
Fjz7CNVtqPhw5mtMerjmGA1mksjkOVhVjkUDbnsRKTd/XYbS8pUQ7sPcvy8DHCz9
bICkrJaM1lxZfNuGZmjIvxfkFCyIaVj7MKRIu45897J6hBKPuckMLNfFnoTQ4LLz
iwFtJLxNz6fT7szRSNA6/bvmZY79TmrVybL6WS5BscimAgtwWxg18VxkwZ6qmTCv
udnGyQG+VnjM/VcCsKcd9fJQtXj02Q/ZeipAruw2EbnMl8yTPDJHZJfqLqr/LHmE
tF/m01xfgpj7fVDOSD55YeM4oqQ1o4gKy7npnp8iAOgFD7cihAsZCAFJT7o4HCKz
V7LeQ3wtjl8TbVQw2K0SPu6l/Tpasbmv3bHMCHK5Dap5uvhHkVdBKRBLphH9kuvL
XuguzVFRIMZB19P4nSMb53GfS20IXT6n/gAc1esdSY0LvTQsqXMoLDDf2tPNEEES
JkLBunqbwh73bX/9kYUjH+CNK3wfXMX0NePXswKdjVgWPP1PRqoQIi+pUBvv5Zl6
G++4QEWm4odHkXRcCrGBfiysNKQnl+3oY7NRw5ABTdhV6e53W0dFB8QrPvVbrX33
v5ZanIA0k63b2fKS6eViOH5AfQLlCyrZsH2+eynhge95bMJMS6jk5R5tgFQS7ZHn
H77M4Jq5XD73fHRPJE7wuhU389MVi3nMvvfQMYSxZ1Wo+lsNsZ7FCysk0ttkMQG5
NF7L90frAAr7K+QfOrFFdUY5IxzWxf6ormiX/6LG6xfNzp15YJGA0oh+17uzdV69
1PK75IkJ5JuYtxAf4pUTfGbX4SrOFTA6uu0OkoKLuI2DrhlvXletbsDVUTMQOwvV
KG/ag0YjCrQ8ZTP1mh8lPFzNNleLh5c40ev6rCTi3kVFpqsgVMadNHdB/ztfLapI
p8cgGP8HG8xYVSlGBFbHfWGKs2Y52ckTgCIBay1QlW6rpioQM3CFG0FeklnllIli
y6h5afbVdnzDaV+xqfCF+36H8X8QNMd1MubcjQ+m5LvhROal3WX3fU0C3DKADwcE
VvYzWbCf+L0zY1uLJ7DFlHnhB7jDKlH49CJ8ba5fGDLSHTu1NCGDennloB3RZ6yA
f+NlXdBItXQLgLgpg9WH1hFnM4LfZAN60mq9x5zvWG8oM2GYZw4VUcn0nGcYSRqt
hcc7Tjk0Sb003YUbAuncjIYcTD/B3GPFeqcnROhQvCOVA6FSiDeMUE4RaDBX8B4T
IHHEO+Kb+W31V4cFipMy7amCzE/q2iX1jS9AOmm+7JjH8585n+WaBjvraS91vFXY
7OKDsHL4ZPxUa9YYAE4AizJpwicS796P0X1/dDYFzXKa9f5UNCkZZRoVL5EH6rP6
thdU0Vz6eMzOC3GBCD4ANdZ4iVd5AVe+nv0vF9zJVbqjAZlE5bWOsi86Hz0Badey
e/KbLRTmCPINPq52tqrfhYQ2eAY3EMKqeunfqtYcjOoPFN47K1MNVsLFktZFEMby
pOFDhC5c8mpSTZeBnqgRdRejWtfdwsCjBPuhgTf9kh8v3gpRp2JauMsGH0IxpOR0
7pFsKzAlcTc+lkrw+ueK5KMwuxpGlk3jAH4ITR8AoLS6oOqLot4YmvIjixCR0wDI
8pIGMw1IYtMObqx1VWD7YI2E7DVOjZ4KBMim1gNwve6S2OQuqtESOYhV8RP+Q7b+
9XJI2QGkuk0QGYdRwkO8YC5BBwGYXlF0BScbif7aY72xZrtYEy/+ot91/3CFKQYb
pfb03j9eDAfyIY5EXx6qDNYR0klLWs0qjGIpW8UmKk/7BzSjyhzSCQQwrvNqyIKb
8z5nCcewmFAKIflLUHIkiQ6FvZXzOi52DuOaxFaI4PFB4XIlD4qWzJlFmV0En895
NQw5TXVlq8ipL4SS08JAq7dfve7sS18ZBIctbP7/x1rXTpvUWQBFahdYkH+B3O6w
/zJ6z6HbwCTVxKFNYn5EYOg4Bfi/u6qJb2GUknLf+Ols3L3We9di5MKo2fix546w
3HVhN6dSrEfvOhskt1tjqoACn6tdxXNwitTMk/TYA/umsM+Is9pOWUGdZLci1Q4m
pFUytL8frrKFmXzfO/r0FXHXJS/Cn7oelb9cMCREvJQOg0HHkrSS/rftKKlMXIWQ
D+EmiH21nGeYMRPHgutX74DkoYC7UYwhmUYgRU9n0GAiYLIcUaU4WS92O8w7UX44
6aj3f+PaHn8ilrrJpJ+gKnwz4XpFOb54d+apVdTM+nRx3aZbASq4yIYqWUKn2TS+
XKVHPB/AwTW0zHCDXf2oA89ykR9Dpst6MfNw8dMjKh/e79v/lRLOa9EPY89RCq9W
5NFQKQoc7opqx38trZniawlBa/2Q7eyUqp4QDmbxiN8/zjLQroAJSowMh/kpImJ0
58fyrnx0czEilx10tieZbnsSg1uqDKK3uMy4d8li0NwVMMVKF6Lc9gPSTI3fNAgO
r/50i9ddaiVvZiwfqws8ApWDXgsuN78zWFe16lnSEcTQirr4PDvlCwBt6CPfGnV1
npS+GEBJEnx/5eHTPhKVLmaaGIbW9V7fM22+lZ6jcgamLge+H024uHXrJPSHW5YM
WrOqhIJDVg+xIYGYsUaybB4wewEb9HgozLkS6iXUefb0BhXvpFiBYBgP8NPVBW72
u6tst6tvrEH+T5GOxT9UQVxNTSDp3/1CcZqN3cXquvQ16E2lLu/xEQEkTFOKgmpo
uofwrFtaNqJYPH58MgH95qlsy8q6d2UhrFzNplRZk6PS2TAnlVLVod+ud9Ck2I+A
VdN5w9Go+fO6As2qb6YiXLMWYkpAu6Ys4WoNjTVaJnQBilH7CL4wSwyg2bKvsO7+
nrOkTdoZ0TDdf2QxrJCU9MpV5CQOu8yjnqqPtMj9zWnGILZoVbYOQFEa+0j0R/ML
GmnIZBlHMTeBVHwoE8m2n9v9QYdYL/KPQkaduHmfGf1+pk6AXrYc6b2uAunCHCcl
X60AIzbyihleKllBe5mMf3KLrKaCPmzeegDq1atUencaPxWLL4gj17mk27re/FM6
Zwmrt4gFFvfXJgNZofjB6CTTshrYdhx/CDK5hBclMFyr+vTHftmNKqfadtBJE6xc
ZYre4jnQAEC2OfUZQ8h+Y+lmQRJZcbeeT1mU0zc7r7ic/CzYosgvJBn5lrmkqdrQ
+ZM4qvSXTKJ2ejxQg+uk6Ea/Ti+mM6wOqGVJJSD+BXNN6t5nXZ2IST01cJriw2fH
XQvF2hKbKyAJDhLFdPq2vY4ABzsZZpWBJWlBnktTBQJp4EbLFT+uVlyPOSvLZQAk
0IXy7NbULHxHTCKFoCc+MbB45g6AhQdyQn2f2w/svPisp79m1urYbL+HOJXUwfcc
OE1q71o3kRcXFIq/Vtl9Sp2PNO4FMu2MmjFLSU4Kn+AffTSS3f2h0CfHUjPlr7+r
DkUEBEnz5rBUdd1mCxGiq8CcQHB1OphAXF+gJcpX4k4Zvi2rKjbOExSyCAL2qghD
ThlOG8aX9IaFrnAsUv/UGG+tOXBPWZ7KbfW6175N1gV/2yItocZ9RW2EaFen2dd+
JJcYfEaEQL5tTf/qIkbHtsjU+FYXcJ+SNAgIBt9Z7Q0J6YKnox8iC702T1MYTQoO
5wAZBksKM5fTLMVQ8TI6aDvqTTqcoSy5ZGcg3OaZK9kzgsJ7NFApy13djnNXhThF
8ptWWOcl2Cy5YcZ1FH/xj+jSyXYxDRiFEgfUMzvMGQzvRubGDyzBEryFMawU678e
vnKKOD+rnwOocwa3pg01315ZoQNgKzTKyLjARaZ7eVFm0YJgSjnxtcU7XyDTPkE5
g+cLbdHSg8Ppl3lJVYg57K8bCJWf+Wc3jzUEmLcXjGeg3HmLJEB3ZN5j2rHR7Hd5
sH7NHH3nEgJuu1cgPNEOWbjj86JdcUhUWgtR1NV06y97kpjYnlEpywFPqSZb/Aft
IkPtGkN80rJvQtbKKJ0e7yMo22Zvr1KYwM1XnGHo26UzSGPo5xrRPVk8jDe+fiG0
QzEqDsAfl5qmoMbYz1mTb3nnR60FlBNIjFLmQgDbsLyOASb65OKpNTw4/Y6eUtZ5
9CnewBoOAHF/qWlGiew85WC2DRg/WmrsazTahP2s5F9Jbjl/a566AFDHhUBQfWFw
ATHL0+bLeJP5KJds/dl7e0wiN9T0QumYdTQQaBS1WaVMjxWIeUDr+y4SSTMhBBTn
yqSkM+061hLPkL5r3hkRhuOAqwiVM5/lNIPKHB2u9uIn4jDZG4aQ/x6mzIWsp26B
+unS37UyhEZfs3E2SuuBTg0aoc5F0vD34JaWyiZEuCewEl6sp55k4XjkKCcBMpEh
z499i6B9QjIG7Rmp8ctsCEpufXQZKeG4oFTR7Rvud7KlkXgJjKD9A5wBGSeVMetG
wcnkbw/AB8c/EUk4A6vZP8ot3+QAdsrlzrnC5XrxKyaA1chG53v1UPBk+aJtStYQ
FQDf2N6t7y8H7hXHEo2054jdS3nAHX5nANF8hpDsJJnitU+Lm3BGoUPgG4zp+8Ux
akiGnqA6tUWObz1GFH59JqwLKMDYP3VYWBoUugohscQhhq9cvZF6vlRa4IhpJlEF
EgDcd4WBF+PI93e/B82SNlfjteinzg4lsv07lwtb4xZCLEKJMMXep0H2Nenm9SRN
KGS1xI5k0pBNEHKJt2AG8EC5vD40H2UC85by2MaoI2aNH69h5Tht+iTPNvmWU7ah
kEGWXa49SarmLabsEv5mhaUPDJS1QNHS26pG7DdJ+S3E+8ut0eQgmBErYrtfWtlq
UiOoTcWFywX6u38pnxodgsuEgQUmzVeva5iFlkvv36QY1SrGx33loZYu/s9WCg7s
briZtn5cXld50sqzUIlEyn4KNGcFBcEuZ4cl97WvDupRwOdJohuntmsmUI/qjtoD
1/0luaswuja505oQr8jeY1gnqlWr4+2F2EpFUjhyVpsGrcEGum+Z+MsKT/LPE2aG
RGFtbABFvo4BIG4n7iLAT3aUktbV5HuEjkp35+ZR6wXDuo8/lZS4ZyHjePMk1UwJ
xctvats9Dr3Ik1RktdrPvAFs0tbTHQrLjl0w/t/yYjmUYLtBtnYbyVAOcLV3BZdR
Db0ff5YcrANAwUNwhkDbGrffPXR2YHBni5DC89DX25at8gdwNaKOYC+63lRYez6D
Sb/cIIRDM9DwL7bsG82BY4Jwl/oyFjWlvGKrLgTS5N+4xB633feLwQ+HY4Km2hbz
Uu6L0L/qBhYMwQa85AjETbCMRaMTsY6VUe1Qj+SBfeZCshW19+2cR/kZB5ZVB6bV
9/kUS1N2kJ7S8modACzlQ29F5djvRV/C0IoGBiNyWvma8UarAWRW+AxB/idWvbCO
NbLDCsVkZ230UaR4BL28P0VpSaXMr/C54awhSIdzF+lHeSrzO2Dx/aNPt9UnJis2
G1lFXDQSYPj1LPZ56jqfz7WUwItgrwfKv7TVOVIO2rqR94bZGJRjiQRVPNQIp5fj
jNcpHSgwUjfOTYSDigkwI0wuHDmqmZbcVxYr0irUyNIuGZ4XaLw4bkjJgoPSAMGy
+pvsZsHL0JhpQ5xhE5so69GyXd2foffotj5dOGqhjOeCTLkyIK2OMVXg5ASQci35
qMbopZOxXLXOFvWpUnGKgbSZ63mOhEdV/jnRz2aIOW0iQiwpdpbA6J92ykGrVVZ5
+0TS4fLC0x35ZMiBkHmcI/jiKsrceUj4a0GmVebMMm6lqv0HJf/lsFx3IWeQbTyu
4INmvFzZUCQpiM0YG8rYBUcJofP9cvIR3WGCjnnXRu/60F4gNDAisqiokAJCkC4F
jFkw8uSxCUytQdHDcpj3Q7LuR2qA8kR2qaEWBXt2jRhi4lYK2AvrS4lNF4GVRkEn
fES4WH1BvE6UyOjmrhR5yUpNaVY2iL1HAMIaiYXmzH1KFeYxyQHETKRwh6CqgdbR
3w6ZCpvCbI6Ii/mCS5Wt4yYZDUzYGv0W6Q/LR7TCP6xRGCljuWlw7LNaayPVV4RV
xH/Dm5bxlaEgtzumnDA21FH682u27OpYz6Iw7KEGUIovuVJz/cs7+0CPvhjVOn7c
TEWBEG61932ouI/JB6kdf7p0pjS4MyX6MAxgNQNsvTLYMBRmasZDA0Z87abhrtAf
EIKM73wSl12GjfwrE2Twlyghr80+toFmOzEXsY2b1btaP4iWjg2lvZsoN9E5NG1w
J6cKwWv1qhrlJjaADWR5l+XM5bl4NhI/yrzTsL66zcGD9EdWq3Kat3fMDumHrx7V
8lC61m7S582be3keTb/h7gcAmtL168XECJgHBXuVMII/yoODEfG+ziOBNPoZc4pd
37/u6ZqQ/+KpmZ1fiJx7IqBktzcemLkThmrx9bPEZCpREo+84EnSiAJ/an0Avq61
eLv9kIE4kfaRWmee3/od2FPn5wrKFYXtRj2x3y5yCsaXw0jyac6Sk3xjdzidZ1jL
NuT0/k+C1n8vrR9mJODEX5VB/2fgj/2e6rl8K0sx+KnPhZy5/vGtoGJLLc3O4QbU
KFjqa3Nt4lasEwN3HgOnNQjZ2mcJpGNe+oAMbRQ0UEeUbymSo++OOLJhHioS6wR+
Q5BZDpOhLsTYKvkdInz/Nansu0wCV05Hh/yizkpm+QNasq7EHJnZJVLSOMV3QmE5
a9KvRWWw2kcYEXlUVjnHhDFGr4Da6lq8Emi/I3w1iZBoTrnVoxf8YqBvpu7bdsFN
VNTXYmvd+9eixeluKe5O34bQyRO+hAApv5IzD167Fuaizd3MHkotrzb6dyQYBWYJ
cwqlmEW+3LFMsFAnIytTb0cy2zyiJPtRnut15WSrvJdaNLjTetETC6hr9V4+9rFK
B6HUFaRRfFMiu439KcOdwvrhMcLIHZkd8nHEIAaw9baspwmJfXR+2YF4S6zM0i5H
Xg5A99ZnfUkMkKUSjNYVJcADu+6YTJH1PwyuQSYFRN/oAdhoOoxtcloFu4EA5Qa1
7Jf2dd153abNnlDZ7Lk5Vm4yOs3iAePY8A2H8gKrU42qhMfVEjVMmI4jxD5C5xSt
pysm6y6A4cIiz7fEu9lteinywtHZCl6+XCYfyfaX98bJm6oIsFNFRPKqWghoayfj
Hh8JsxorVlMff5I0o8ztACZEKW9mZaqJVUku3QV1ziaR1OGRoMw9+l89atFZDWmR
mZ/6RB524Md2kHyQISGV5JnqFFGm5uEusf4l22yfw2je0XGi+2TfSz8/SBM1lRo0
7EMcCN+6XgnwBQO8do7RZwlfxo5A0e9aSqgRrMR6lxribPKZPi0cR7qVcztTO9Af
cKJ2dFeqsZ5nzo706fdH98eqUek4+q1PcAJPv7BMzAgDsHb721ACr8kNQSzcC+LH
k7LYc/9IM2o/uPAy1j6OFBcD9PrPsU6xCLHwenKLeT888VebHOya0yQJJWSGmIbn
dTwGeTsl5o0nvTlD5IADgQclncn7vNb4HxhLQe/f1pS7GI8+koqQtvAkIpPq6rWp
EsQIJSxHjetKQGBelESbGS/3M2/SYce80cGimhHjhMmg6esN/hkUJ3/BvmCj5w3N
zGW+ZA++Wr5WGsGIxVtC/UkYi8WMV+9deUgdmR19W2V6Gn7foSZ8H847ehR/uNk+
cE+o639+hyVo3vTaYigfwdKIMvqC0kXtXqzkLz4PzJVxC13R3ip4LSa+aGduceR5
tixou2V6lYE2vxr1PXwQxnVIRDw9IjHhx2JTjIfCJJtskCFxGKof2Z/yhpK9WbNH
Q+GhbDTNzz9AnulZ0U5ch1mtiFRovQ2PEhFr0V3bi0YVPrqDnEocJ9Hro/carIeb
2MctAMoIE9MAUHbLBlAaPurCmQJVHwjFCBEebxwJzOowacud9Cyo6G2rKM0I6WAB
7bwSPfrkRQceqeaiS0sxiULQzh99tRoxTGx4wc9WXyrfP+bDFXLc1sLt5SZ9gUqK
Dwe/TCvjU3jPfrjPBQQms3670MxxplDbBKmh/Hz/Z+FwPCYQud9+sUi8cYnEiO4y
bRpc3ehjjsSGyff0ZA0vq7I3O/rZTBmZCB/f2dZVgTyWvmyp0DOjJDiAS8LWVDNP
hTZBuhSKkbOHpf30yiRg04bscd4oGDLyXImkKR/LI+IgRe2S1uWd/kjpEG7p+Aq2
qWRq3kQrkZr8Ad1677CxCccH9yMqLBoij0+s3o1MMEXOa+CFYOCP06HMxnERBuEv
4zTDTyXD+p+iZOrDsr1ygfvWaKMYOQfubkbajiMPMo3F9ddyRD1O8FVXGJuFd2Y7
GDfWn6+zVsjtJbtR+/DnDiEbjJ9uU2SF4cyXF+amoxkJvv9KWzrLg45Gu3vWeaeF
WR139mzw2/JEmfkA2nbzAHKRQ8iyLUO4/EiBp1qJZk9jXsdYBe/nH42FAfrdUEtA
G/V1IazdKzrqXF7muw5aooMeFrkb56InSZ+g+ECCCcxfC+ivb8Dl0anZDgmv47vt
HyPADDY/4dny8JDhmMvv8MLYvPGU2+dCIZg4fwkSfLcp/N7hRg0enLXneNZ7xk+x
EfyMTmIlv/O2LjVfnhHtS3I+thsbpzu60M/oY/tfFLeJXzh4kmgNvfx7xSy5CrYg
G0iHz7XYh0sNCZd6lgjvpYj8oLGAGYK6sGhMi9vyBxwD1kNZBFYbR/o/MUr2EPPd
pSPc3+tNPWEWiNBXRer1KJXPyCO8uN26mEfH2ET/UVhwdwuNcpss0e/Y2A98nE55
3kWLZvcQ1CCtAVs6sY4tuVu4R4tKKX9Pu9aPYHrgei/4RWhwC1MtzIyY0XdU1xhi
Q4Bmuz39CmYFP3ULqCkW6OU51/p30SLRG83dOcAZkgTK9yLcN08HGOrt5x7PSTI5
orCjc09r34CAUqBCfHBu0G15aaKUAz1NZ2XxT1sJcNEv6dfZoH3cf5m7nsbsZJjc
/+8GgAdr/rFvjnW0BJhNtMRXbSn+Muqqqu9ubqfzdO7VJ1CfdrmzCmbcgvk51lIX
vUWm/w6V/AIAWMfkmBq7aYrjzKzV/ZsJQ57ACDZGocjhcBwCqQ8esXNEKepuoLc+
zyg8cg7Sm1NFg65HVKQs9tqpiREDGw7r1TLnPr8JhiuF9zYI3iv6yXQzfFpiMF4w
8Em1oXKzcny+4AEaP9/7OOQCIJReA9iaKZwx+s7P/P+VzzgOcZNf8ApIADUfRaPm
GB1vk/JSQDUGz0sUF6t8IB8RUGJX8aK/4mv2wLL1/MwgvdvuUDGIe6yHgHEu7Wt9
xmEarm0NtZtjNbHIGmWAfafhHZM2ejaxaEl/qKnk0g1pLJgvj0VEL24Q2bRRvyAL
J1fWNHvPewowdrvQIePMVG02gKnTLI+sTStpluqmKe0BzrWhg+f3TNlrUq7xZvyu
pJ2h30bbDUIhKRij5yjLMEd5DQgoirOQ48Bn6H8qJj7EAeLtLNWXyh82b+oa/swp
jzpEedKH2KXSeXstgyRP8bbxEnogBXDzYBGalKS5LJiMc13gDxwBeIelNbwor1dn
lbwEj7GIsUVbrCSmQJtToGvKO017AwzCvoGs9m55h+xpgBmoSAMpoezYjhH/L9p2
V++KCADl7rhHnuAdyAMHM140qKQmvYihzWj4jypTEd9poFYQlGKBG/UvYOp90XmP
L4/pS5Uq+XPFhOg/9oXv1RqUqB2oIOIKSlUT6SJCRPzULSJRGf5LzMYt9r5EZpJR
2gzJh/R2lRBbUjjH5pBmpuCwAmNyXX598ASOxBcsW5F54IqP7fmh5I8ce34ppVwf
AYE137RwpgbpknLqVWSHURtyRlCYXCIakZiuMyKdaRLm+SXOj4Q36IU0Bx2VClHg
EdfHrFuJoGOok/ty6w0re2vwyhDWhEwJDXfNjpNMb3CeUGGyIHzH5ELaXMWO74g1
F3M6XYkyw8KP8a230m+W26+LcCK5RBrDMuQvl1mmIhACGQCS/qcE0jEXsZ9fgAUM
lUquCQbNXzHomjIwDJJ3W+el8XLL1BEXRJClm8OAu4BLlSR2k1AD9YC4S1v/8+HB
S9a+spnJf1i7Dk/A1Ii4IBgCp8DZTMWh8ge92HMG5rrmn0kp41LsOgusVvzemyiU
PoqMudehicSV2SwdEs9ebOb3z85KqnUavDCZfc6sELQlpIaI//H/4RjcySp6OIjX
pSflU77SwSWrqZH+yMXMgbxoGtQ38a9vbY0xPk6xWzgg6HLwX/osFKU9PFNiFKcD
ZJ0w3jEyNOcMHd7fFd8jO05csF4DowLM4sBIVZ1jjVxUpXLBU6f68kf4E4sJzrt6
oBNwu2RhBt9tBzHol9vl8txSzWuUWQxk5q53xPn9pWiAyfP1cxNnpRXVlVaIHVV2
YdsSsArv1XiLVtmH2Z7Ktq1+3q+cmHtN4DiuKll+1zXgdo9hv603QtYLkl0VO7pp
/KBPzYCNkDrG9YpTRBVP3n6e+jX3/XTLLT1oxiUDRihaIrmydIYyTvHvKBCP0L7s
fT7JC436C2Y8g++j78V0tNUTiHMjYxbMaFGPDl05ruogMZ+cAfZ+t40M3+7IANfQ
UBlq4eQsrG9VlQ90GmLT++yGLwbmd41647IrV48MHpLFbE+augWzxFEE/YwmIcHS
tlJMeL87Chvr/47tE2Dpg8qUWnWeHLBOSBCHe7B5daoohrwFss0kmcqqI+gNrcMa
9otybwDmdatHY6JdCpgYcqVDFSBHgyUJsZPZ1kqJkPX+P+JPNoCTqXpKqfdlZuI9
SIjfsx/tbT61gY/susrb5A2RhAfxgv/xzro3W2f0d9bldIjU9dmXxydzk0wVTqOt
gjUW+zv/bfmPqEc5S10I7ojZe8u2if+0PwLEN/DHY40NpBAN7xo3AD/FRCvglab7
LtQt7o2Brs8x5Cg8O5rAZ4Vpzjezr9po0bsxwrAcWpUsQWtXTH7OXbMFPo9S1Xw8
WEvHx1V8eYpC6LMa8Ce+exkCTNWfnn4TkjKXB8l8syyowwsDeJL8Y7v0QR2Ipdm4
zrkoQH2PKn0GRkcWOrftgGIo3I2TBtzSI7C1JojeEwbb5Ud7AjgURJ+Y/DaWDW7K
cFp6DsWvqhIz6LL1H6VNJTR+FHCtGdgkdym0wujll0EvkjfhZ8EcK0sky7SiP3na
4M+RRjC6f5h8b3pOJK3CyTHsZd+Bo159qqDjmcpgVb6Ks6FuVcDDRM8U8I/8DIxV
ePOLP7YGgV9YxtZsQIzK4z4QHvHEdWxCwprF5Xb7InIgKZClf5Zuzw7IKEIeHJmb
MRPbJ/4K/C7Ppj3ZEukRv3CT4OojpyfI7dFhzEL1YKm3vTn6fjLXYjIvn3elLpRN
6KgK7Pe4KF1UjqPSXA7vimcwh7yM7VUqmvHlVmJ96I+EC84ODEBJ15+QjfvcKPmd
3ltql5EMWxO66ln6E+d5VQuj19b6iSP+tbhsbl+Zye/9eBW++5Tn4H9v+El3Ctkp
+2aI4q2U4/XZVu8BF4dbBENvTAxW3dvTpwGeCbgm7G6946XnBNqmOqw6Exx0YB4X
xO16S2iskHvlsMz20FujnlWEKQP0zmN1psMpA6/qKGBIoJ1o136Y0pvDKp/UjSCE
0HDNUmLb/oIOJoGSDKh6fUA226nNy0oNTawAGR671/sJkUwePb/OOakF6ELshiB7
PcqHA/rM4orRUHjBg9qRp9D6VjQ9nXndHWUhby+smBfu58ZI/A3OclHWH5UnSRM/
vko6DvgeKJfWzZxhaif2VilSBLgzRqaXrK+HkiI6Smt9LcJdy25koEfe2zvY9DeT
1wvgrjhB/gAA9IcXtyOnISrolaWOH1QxIeTMaFDJmotf+J/SiSw6Qi+kOKkElI7U
FB2bl/otbOmvglIx/AMa0FQlz1wBXpsuABQopqtRiCxIV2M8/ZIPdDZS5NupJWf9
6nMjCijiWUwPf4FqegLp+8kSw+HL+ikQN9Gk0jjh/c8UsHy2bZ+zIeoC5yD95Oky
VlZmmZxD5UJDGtohimzZBaliGr+FclNA4F1Z/kCm+1i1d3kadEBtSU+fALvdXkuy
v6HMrHEE/L2y2O0MElyTBl0sVHuqbYF0yujGahl3JLxG+TxnsYuyeqgcLIjCAwp7
rZWu7zQfXcGjpQknlwbCUyR5NQDhFd0w6tN/2P95vhYHSwpI4i+PZFyC7g4/EE0n
W60QASdMgNFnm8RCa3k1NQi5zEin/iZ0h4UzS4x33hwTim2btIg337/jGFnEjMuQ
eE2eo8ax5HHC/QhTd2F+QZB+QadYTdeTcw3rnA3vcgvaJbRmky1eBBFuEEg9EFq0
3hZ3PThBoCWSVXFFekpZOeY87QHXBe/nSWsSsXJkfNFmH8K76rwXAmTygpFEJEAc
zMd2dNtnJfXvvWspn7tYA/tcvMsjItmGclKFGhhF8DxRWQIhXArK82Jz0sPYl5fe
5kMZiCq69a1ThwMPhKhT2Q6UQLq2HzqG2B7a25Tk8MpXJn1iDCVAOdWb+Y+3oOwm
Kmho3giiNq6fgNqHk5YsScDBw4p4ikBac5d7legJVgtP+KpOrnELTOHCiNVSuU4J
EHUJmieKYv++yf9qT1KT/cE79cwURxINoXdM+SWAuayGPY0KZG9cEoGfLxIfh7hY
NZWxL5LSur/YCFSiHdEIXvxOX7qqrwmSyTNHD2pssoSq4Ypk8SEJryAUW96WP84E
1SDpeNpkbG7nPfvbdl8nrAnH5gqTWjSvcunhXBS0S7EYzATN1BhVkXE/sfJzzrWq
o6CurtCNnSm4UF2GY25bltAApkKnDbS5uoyaDGeTFmIBsuZLNPJ3F7gNl/S9xO8A
6ae8Tkfr8JAJRf7ULo4tfPUheqCQ94sNF5FhuvyNctgWdx6/GsEgRZ5W5KvXPoZO
wkUSYePFDLMl5Zioi+dfWN3wZFeHrvQBZsBdlybSGQH+y8GLQUoXF4QT0pkY5rTS
e1KKyVyiRU5EO+hi11SQ/xEX/Fbsqtxa5dDVYy+Wn0nzvA03RE158ZNN/N9FwKE3
O0plj/2eU8F3oOJZOTSK3e8LRLmeNQbyx8KthM0I3NwrWTEkxs9C5LmrPpjJeXKS
oyiheBXJZAwyvChEQpPWm342mI5x9kHiVH9Eg+rtI5kwB7BPx3mqvzD1CrvZpNr0
gQZwhCDO5iuxr+SC0wtS6SgbK8FRXqGsvXIfw21yWIIr1KMefB3Ewh//hNDc1CNr
Gx2TOq2tTujr536hPIrWQGMwpvOncVcU1dftmLSywdhgHGEShWepQP2SD/uJ3c6p
OHOcKJLonqo4AgTur2YR8aUcyKzKf7x6RhmBb0TsFvZAUG2rnXoAApiORiKefjqG
/lwNUVCBSQM0ZOBi0/ubMNwEv2cAttuRDpJ9Rkg8nPJJSj5zXcI3hhy1OlMSjD6R
a8OJu8b7DBOq4tZ1UAEVz5ba66+thH/f5PI6j5+ByylVfWA3cecm1AzfDUYmfRvM
zplS5vPG7Df53HZTLOMMpPLl3jePkOsHst6xpB1crabOHOW0sWaLuow127mtRBx4
56KCTUMKC08DhgKyZnp0Iv1A7G0XBNFz+zQtcKtGuto9gRgCaLMuhdp8bJx3WND4
D7xOLmzIOBhRPYKAEbuaZgoSUTSl3dqZDMFuOklcdGKA848rrsIGFPfy6nnibqAx
Czbnlrw7RZ4tC0dvuoswtqCfZl2tL8+RGivqTeI9cGFq+1aLPPEFgHnro9xnkP5t
+NMWceGchqyRM3GpFIeu773pEovfE28bmqcnb7Kf441igLPzDni4grx0dq+AudBQ
nlxvOEutAWI9kcriG9CUTEMxpEGkAwmzFGlZ65BH+8hTgimFK6iHC+Uh9XNmxcDw
1hqS+4T9voWsmrGYJSLFlYIKYg/sKaAHYivJbcfVF2QlkhEQFxn854Dhm3wxEHmP
f1YbLCDs+ceYBDgwcNhrnV+UVijZmkrI8KkTX4G6dtXuAt+sFQouV3aLdKT6GXyz
W9OIcuIqGgXn27/2nQEFr60k3yuu9mOzzi19jvEXVuNdpEjNuCtcvuQ3hJdYoBMH
dQpEf+xYkQzRUcHDOQSqD7gJju/0Wob7fqtsQfwxbquSRXNUw5X2FdFFMRfzmV2X
nxV3TSktb83pjgWw40+8lh0abrcvZ32OS2CVbtKKq48BJ7bSh2XtHzttR0unLfdf
QalwLktBnQkCCve//e3Fpy90jG/SGzSMqUvaA5fFlBkvkxI2rgOOqzjg7Ett1cpO
DPttEqKW0tu6EQVS9PWxMPnDrGSYUu0xHcktl8jVm7EqwsvPA56t1BfRWcss513K
xfILYdD98Ua/tzLYH50STkecabYHKLNeYvKIAkHfTu94CxUQW4YIG5f415DnWEMN
s5YQmORHKZJUOFBilmHJ7oaZbY+QxD5ahbkFFjeED9W4sEKVwOyRxCy8ITlpa1MT
R86MYXkV0gGo6mdd5021yEl4f55dbaS485kfVbVerV7Fjso0MlWgobsfcieNSKl8
BDNP6OnPbuYyxyzllJWlGgTqYTmYuTZQicHeZgERTBaysdX1OfIvjvGSZ4AOA2hW
bZZqfl603nBkbQFPGlRKhvTTe8exUO+2ANgU9xiYNDksgTzRWgQLDzyahUIUc2Ji
5ouTzs95tNPscMG5EKPJRs3usv6MvgXt+oUiCyvaYE+ECjtTtfwSzxyRsuUSdazM
Yc6gzw3ZwsXzARSCSGi+OZ/YFsMde70VPU8lIs9Kpwh/bowTzO1loswKBm8YcwY3
qIsTGO4wKS1YmHD3y6t+V0o3DDNhTGhGTqvqCTT91TLA8zZcwizltSz5l9/undld
r4tHUx8RNEwn2t078Mh0uw95zmeEWIHPhOBfXwP2sOQ2o/x8XrD0PnBGsjoskUdl
9AKMFB/SehjJCbcvzPtBJwKanBpl2ir17ttvG9yHo+yt72Mi8uuIfqql4mI22J9Z
CHdqqW8jKY09Be7RDMKQkjw4ql8BcdisubQ+fG0DfTJiY/v8PNVaK7VnTcotoLbk
h5gUb0YU4KArlw1b+DWhFrfNDlK8QbqFnwc3EZaa00Ph//q5nkad8a3mX1coA4cL
nMz3qrJUwH2Dbc4ROopRIOxnvRpTut1ecRt6AdnIlDaPCucpYuQZL5uIwjQ5SnWu
Rn1exQRzYD9ykx2dtMKJj50k/4+esXVuSyFYznOoM8+v3Gt2jTi7/JLkKpzIGhUK
XyoNCW19qUBNtzNOtMZANlWpVSFiJLU0wLQpVd7z+KflF92Nv0krcAcZRbTNvTQ7
gNqgahGtm4v84CICeuf8suRQOqMFwYJxXwIdaZjQhEqnS/IT2GvHC3PV3wOEhm1S
C1v/R5fo9IsdseKSiZFT9AYdBfVHDlpXmmZBoagNFfkxGUJ87NDXBB2sNPP8gpb9
UrjFhg6s3mZfZRTszdlDPpYsKGb8K7LTo19NltxJSeGj4uXPE5cfcnVMBDPi/YtA
GRcuYucRGBqggAhhRiEc5b0/lgL0hAHxY9VWX4AoJLNYiD2mCMKPeX24+Izm8jeA
k/WxRj3Cje2do6saXQuLS3f2YbdpZhDBalInYD+BihcjVvHk4RU0b/WgLh2uRiIT
RTJXvTfwETcdlsabdF25/MQlMimw32HFjCasJC3ePeouyGt0VR3JGYun7EsQizcA
a/HZs5yNH8VHo7AawilQAqCucWRD3KdOgHLQEqEfS/GANoG3F1IpF+xwsGGi/wD3
Elss3FqKZ/KM0hAYKeAasN/aCeEHln+rRLsN5Hl5UUtbfoN+McQIVSEp7PzbS9uB
sG4cBgvchf48/Sm6pR2L++RnBrh4YkkVs8gPvYgKr4jZMpzhSW1UnxanY/yDlDoI
zo0Uhzjvj5hS24O+oh38rsyga59jOtFugnCf/I3A4B2GqHVohuD4xSfposVdI+wW
j3R5yrddV/mmfXLvJgMUsY7UbdyMp2TnLU4w0wMblDtojRGBR11wHC+xKKBa49zT
SpdI3tdAsOEBITefY1iVnD2MI6LQHD2NVo9N42nLmX1/3W6fxnrN3YCxebJxwvRs
CPhAwrJY4eSYAsVU5t7polYE3AgFgj3tsQgDsdIwsC1/gGXBjJu7Xv0a+/5KinY4
CCwMla8EiOvc8cv67EWPbim2zbQbivgBdntIvGhAQ1N3S6Ti93YtiMywTvg+Jd3p
aBYM6g1P0BiPCg656F7eonZRO6sxD1fAliFfbUehWR0NDrao/sGyHjyGAvTDi66M
Vihh8wTn4qXrzzOTK343tAiIlnAvQ6bFBLThUHmWwxlqj7ZPpkwxyELWr/7ii/3U
SyxZz8GEcr6hlgMfFGdxUjvqeT6pSh+LX31+Go5fYdr4lkjXlivd0CeOMy8DtgCA
S7/qaU3tvH7xO0cNL068i1XxRIuSBJHBG6NkL7r3vaP4KjkH1QjiJgEdwidgDysM
kWOhG5okUrRoc9mcuepjnBXFwoz6anFgCeJtJk8+0Gyv15BK982TRryuwyUNtzLd
QyoR92Kne2dYrwRRhvEdyFhewJzbY4O6ojoBgxlaAn3gQHEQhfxdDwBZ7mYvG+4I
FzRoWqW2Gu7V2O8YRZFqunui1sndNcaglSvZSQlR6+68LR6zKJW22mzUJteKfMHY
XUdynxsHZarpCKM/Xatu/cR2PEChfLPSF+7opgWXTvKh1kiXx20IA+z6Yg0vEdwR
bfDseXSF2h9ZFOxqISP3zIvCG5gh59U1ufEwCSDJGvTpUjxnRjm/YsxXKDEqnEmi
g0AMwaba7P9NE8QuCSDYzX0ldP3AGbp5EjE23BzTFFDGpp+BgUJPoWnPae2t7rp9
snIF64t1jvAfyX779JyNIkryAV9GdrXKpPaQDDWscjKu4GDynO3F9YWrhKeJkBdO
sl51AZWdq/7Yi7gMcItGzgZoDS5QK5zT6gmje6N1L70q1TbPU/U3h4cviPVIUcwI
vjPGsJvN4yzhkE0SjtCHSCjueVsoRevnYPHprRRFtlDmNWN0dkYnnyFg2Ohth+7p
n+VvykqV3JXR30s3mX7GJiuUOFM2t5FiIyOos/ycs00Mz9zWLy4Moz2/uNgKJKm1
zd308bQ1BLOGOJVOedweIpKFYQjSddJqpjMc6TZ9v0A88IK9LlTlXgziHHYA+vFP
ajOQlLt0nmpq/4bZj0G4dQeluJifQZcVF5bBXjBOV/JBGOCwWNzPl94P6fubS+rs
1Ue2tdmOJVsC5KMVwmkopxxaLrHAEtsAn41t5fWyMrm1yHtL9nShjCEegbejsMOt
r8MIl0uysWfev9JIL0aIoPCtgO90rEjFZSAC+B1+KCTPy2T7ohdm/ZqnOLmWsSw+
3ZGc0MTPAVrITOtxsjtuoOtzwCBUEhH7oT5OJ2ytNZSMoUK4iJGBT+Siz85KAO0t
GnJYqBI7VX2tqVXjfKCyyYOqeb+r7LtWiJ20JjNU2IAoyTfkvhLmZjHwprj5Nk9V
Zd5UXIFqVbGsAQNkjKhXkIKl2F3x1rzX+wHwiSp5BHp9Am7i3RXUBOqvAnuUg0hX
P1AOI0v8XZvhg+PqOuzRURDeqphH22DYgiPzXJhAYjGPestpg2uuEV4jGiWrfbso
1SAqot95OgGGz75tbwlAhzom8bOOD2rkewTVjagV02trKj4xEyOUSf19sXHYJYoL
zqrADkkj7q2Zr6ElHPB3Wom0nCwy9QhNH46PnsVsriyxbT8LxPopDCwPQooP685z
B4Qi7QAqy+Cig0FEMKwRsABPMmgLuXMXz/C8YBF9tNLvQsjRS/8q+L7RpDLyIMt4
rzHCrl3chVlTRvNsQ3hqAmaw6hmTFLN3UOPGCD8pD7FmBJpBbIbY1SmI80JvkinJ
/IQKZuPe7VEVrwXDZbPNYEwQv07CsntETW8N4G25ehaTvmeyze1131i8+oqWrqit
PgqGIiC/6N5Mm89qf6UmgAF7s3kQLpslNn1JVTELVLdfNggoLze1MK4qzG01ve4A
URi2OZxiAZ1TiYWyIu/022h1A/PbXjzn4jjMDO3R5ypCXbI8VIDK+P8qbug6un5Y
RaT3+mxeic6hoWPmeGWeEFfu4sQ6SyRqIZFxu517KSeRjeNL4MOjhNM6bim5q8Vs
/XEDpEroyeT39lHpVsHS9vBCPx4DQhiZ6noD05bByIEh0GeXdIdmX8Ytuyv3LVWk
MRCaPA8X4jZIzzbVrfPVNyDZ8B4HSh7NgSoK+gyXkB1Iqa0USc5bLH/50+bFDn8q
Y7RlNjFc73GBVmjhiX5wOoq44qjTMqzke8/yKKl3oqTT7PMa8iCJgLotNqARdKST
Izcu3IZlXlHLJ/Yt275C7O/naRkfW5S/M1bMrKz1Ry22uq79DibodExZzJcU84yj
gztJ2mEysJWF9Ka+IkCqnPTxnTwWGmGHo8mNgZBqp9j6mhiPfe5UO143mQR14X8L
XXWMQBcCWKYU1J/Y37zOcqt77IMZIisEfe/5tC/VNXPoH280yEHAaap669HzVHzy
CqgXJHC4/O3L4bxK9wafjj9GHojMqCtbi/l49N7j7t9AOiVGSwuDpyfnHNvNsTBj
ApXrbU/f4HJaBqAec3EWZ7zes4I7uzGyT9NO6VgKicddHDZrKkmWj8plV3bt2hMD
IET0WjpETTprS+ZxtL4p0RI+NjRxs1FArYetDuP0Yb6ziXv/iiRI3jzgHA2bhNj+
yq/a2rK0sGzKL7JPS/zGB+ifK6Anh6U9GKw0EB+gFSAZqOa89sckJheDld0wBv2M
SMvA+7sfPyRvIu1mKhjut+fmlsY4rLBifAxxV3VK+MqavcR7Ytp6fecVJHeXiY9r
4h8dCTOpXB+7al+T1Mq8tF/nfSV7mgcCguiwf+1xIS70poELywYqcr3Uw58tc74c
osJ/2si+MlRRdE6U3AsMNdPjEstHwpE3qHTaCLkeVetktmPEpAFDbMsTUWe5oSRA
YuQanPXofb+5zcQQLwWl3BxK2XkDf0IdHl5/gzAPZi7um/RQucqSRKyxexMjGXcm
kelYgphhSoTKY2znamz0qDADiFgJ9Xu6KtZgquE741bGnMbRsOHWMkN9IR+fbXqF
hsq8abf6TA0yNBn8DnCJ/IH4ypgbh+30wsedQEBSAJ+LOVSsfp5bKJXubwiFfW7J
ZFLTo+P92IcwY0DL243KlvAk1mjwMAKcfXKzflu5pgrdqZFHu0U1sxeuAt1Gj+nE
l8DUGse1SThusAdxvVh79aTyaDbAwLrurffGQx6cYaFLFpE/DXXfbP7xKkKvf+KZ
irODeW/pTPVP1yfjRTuLORs5X9XL/6y5f4rgsQX2fUx2Ye4WDIYzGou/HFw3472Y
8Mp0DRvheU5X7FNTcmN59XJVpMNrWzCo932g2TQTcB9bLNIWdBYYA/bzT4tttpU3
1Rs1NkEdzhiO4TOIg4KOHoBSUb6+YeT6pM1T3IEhfiVNgTgk7O+7OB8pG8quXYwu
PSqPU//yci+37YWKUWNK7jS4YeGc79j0Q4Tle5Vl7tiHY5pEmUm3jWLem9y6Unn5
TiGt9KiGDR9GtrNu2mjJlr1VYXKR1qDYJ0JqkHTkafc0BeNyeYTsrHY+6afdJ5dH
xtICXqpLEAXHYVuAyBbLkwAQXBr+l6GumOKzufVVtTW9FD3zvklRev7w8wQvYvm4
BjX+4glwREq1Cle4oYOhgVRD3aSDy1ge4lJ0mWRgiqmNNQJNQfCb/t7jN0QVw738
HPKW8yG4SGnlrdAgz65gEeCarmuJZRTVUupshoiAF1nkT5UkAPg4+1HSCwQ65nQc
YGb731zIWsCpGfwUB6JMogHVmRXrSRMwTWYzGMmlHG2x5ei5rS0wO0uxUwOBDOTv
9JDiOFR+LMIxD2wbr/zOm846RbxLWzFNoJ842A874/d3tlTTTyAIsT3N5uZPYoqq
/qnsFstHjZnpERA1s9LEmN58DsobhP2Jufq2escQc5dgdPL4iZQsKEyVYYKJwH/a
dgwrD9/VI1hqsTgrgw4ZH/+/zaRoLmvmPva4tWVZ8u5VQp4S9dhY3BFuvj0/VhGs
N/P59PzhZLJtbELQV6izSRd4lc51+q/WqQNcu6i0mu9lg5VE7msnGEikGue5VnjS
SUYl8EYFEbGCGA3vmbqOriOs3BH/TRXnVumLNC6cfrgBVCXrAOiBmNlpD9/1Ag2z
UQhfjeIpSa0UG+EONpK9c+CxJ1MdFbbhQbjq01+QFCnl94HXFbEoEaesB3kF29vb
pnElPl1SAoVSUuVH0cdfSwpzrQEuDHupNMl8DszTht137RXEWGx6DHpjOclagCJx
multWNJmm4dlgaHkn8c7jPGB9WMKXrbnCnjudeabsruoD1b1V0/T5NSCx+Fwk9rf
/ZpAMIlWAKbGF4ZHaI/i5pUyFWVdeLKPNDvGfNco18kLdpyzFX44GITCNNwH5+pZ
NBnzd7neJqxuCdfJzuzIgXFULn86m9xjNYeOS5RGjkoiHeUl1AKTX0GKKY+978Kl
YWKctzHBvSI5LvJIfzkJRVBMvE6tpSYspL3IWwRNKCdCEB+x+D4W7h2Rt45YOJBy
HMP9nliiOLDxuFfZzlL/SL3tksHpm+EwCqB/WTusg0kXjXMfSMfG5q+Pmt5NJUE3
6ayyUD0+LKdTSPQNSkBq5rSZgHVRhi7+X2wdoXiu9R0SpOyAZT3fYa/P/tkDvJbh
hFhArf+DM5zCVCB7NPKN7fh2EOCrrXDSwnxT/ISo4y9yDpg+lDZrNu40rMctwq00
0SdjbIhxoaVvtSNBochT/VGoojBDVOtaxEkG3dv7Izf1z1+3tWSk6xwlaU4Y3o0A
MBULhWH6kDZNACMfbpQFB1vCKmxlBSAXPJL/ES64070+mOrXtg9NrGg5tJ+NRpFY
6zLlxvyXYmFK+/1FaUd2YgedJztxnjytKY2zUQehh61yKvx4aQY4B108hAAD//ER
4hiatfxFKZJ0Ah8VAHXiFO8OFK3cIJ5qzJKDGrwtijl0b8fPQ/RxL51IMzrajpVN
/KPd25Y/yjqxlU1hSexB3EeKGTEjmrHTSbhvDg/9DY7GicSXsjpVlr5iQT6fXIjA
F+VFbRvKDza0mymoKvjYo/1BCQw9vXHw/AKExUMUF1m9wezjKVFHr6xOaWiDlDCa
Uay7yYhhEKZ85i/LrGl8VwyxCiGu2/JCoPlJr4VGG+fe9CqId/nRPQ5HYSw2clY0
LrMKPgbbhrAw/30+hoW3/CWDK+7k9uTWE/z0EOwY1gm7X+RJHt7fExuHhNuxFsF0
aqXx7YtFqlirVDOkmziqn+pMw5+bRb0uTElnFa/1wHGW9gtmU6bQRrfRE+0VNmcg
SWgVs7MZinoZmKKPGC4lG088ceyJkAr5g+ICTiUTtoS5p1k0DjoVaujjw2J8IRnf
HwdqyA7UuwL0K9eKrqxScejBKhf12QGzvJrnSzc61doSnWgmj2V2S0ANBcn2Mz5L
9NS3nCUyqd8KPGRubdQFikReWTmF899efB8Lri3NcSbsdK7q38IjZAsv7iomrICZ
6KO3t0XnuE9G3BBlOxkmA7JgzXv9iRx+6V0VdpzS7aEFTRrVaWcMC0lUcxSXHXdg
aglf18Z/NIFRifI7Tljjtme2BcROcS63iprzSAa7nLrlpzHj3aKGekDabTr8FByb
coT2qBQZPY5WmdFW7x1txV0W8ddW8fruNjgh1KJbAq+8pS0shPSiiH5Sb6l4Ucjl
skjvqxd8z/lrO6l1NjkZ7Ax5ubaSCeP/fTThR3meXysRbdzlue+DSkNHUJK04xMW
29yQl/M9yFumn07DtILRr+AUY4kuzeTm9bj8xYHa1x3H+Mo/PeJ7zaOThLBuiqWM
hZZaHh4kWV4H8YR80DkDfb1ANaYxZ7cQNuC0EW2kATJVpFvWDv7L3jdVGQFIiPE0
+EHGM3Ea/PPkhvo/CBXazk9BGYIhdeoZcbZAYHT+X/EtB9m+lY2jwU8YF5TK6yq1
xj87T/MjiMNMnufy9zIZIuP2JZz72hOpJ64kmuDLdy9dXH0xF7Ie+Not6hqxYrH6
JN5mcEYI6rM3NK6vN3o0Pfv0FOYmHNf1AaFzvnyQ/ucIV/J6H2sVNcNKOZMU5a3a
NHQzjBJSFbJRhLX20Ey7NUEkebnos/XNlZw3yo3zzKxJRgor9DWhn/f62BF0L4t2
XUeEJhHgKcKgbdyCy0j782yYnDhrz+kGyZGS9cRO0o5H40jO7nqWc0c0/J671PhA
zuYywziQz8Ui3+t9lCQiOwixweQlbFPFwElkyCqpuhzIKxvmpdd03U9LJlwFFmKq
ZNNpyPbE0KJTnx2sfpxEDPybi8JvX02tNrmvhno8BO6KO8qmYmXlXDG33uZdh+v7
kWBAzcPquQI9ydXPdNzCZ6E1Pg3N66E70qooglrK/XTGCboUgeA6hNFabuXUa26J
lTSg2tvbhuYw/wJihS/tDQfGL5oil6Gft42Kb4lOCrNRRBUEP7pCsYXuvUS1hqy4
jKKznxubiknpfGE7fcn/MYyuIewLw3QeukhmEkGk0t0rpTyFf/InN9V7cCvD5f4n
jchpGUXk4zzNO5RJ76AtqThk4em28AAuksYVL84AfyCeUkd0jhltp17XxC8oZmiZ
wcrYPgG5uKWrhIirBGG5yizTc4byPQSQ65e9rVR3QFzXjjqOpxg3270gDne7nvrV
dEnHx9AzwqmOqNegOoNtqrRSx/tTCN3VTlIeu8TjdMj/oplwJfZuppXeMH8TQ+Ze
WLBM+YXsAUl3g+TMLSMER14ruDUtSJuGvIA1FTPac3xswBf72dXPOk5fZA+6gXzK
7sxBKmkKpkP4LCzSBiGEnEnSyzjiiRcu1PNOIDJtU92NrtOXwMXKoMJdCwOwT802
w3ElV8rKtm0BL8Mg+8uvrQCpOFSsNLZKZ+2YwIsEs7/22ns53V1qpgyBXxj0WDmz
kEiUqrWUyyzbmsjdeCsvHbQXHnGl3k5bKdGTKuaepm5InqXxOaWpM3MTy3wy0eHD
Y+fbFnz6peLjrxLf9UQU3D79vlQLUemPzzR5Coget5agiveh0/cQ8WyiTX54L3i3
i1FkWZbg7Pz8DmrOSJezNwM8WQXTDvQzN4v0ATMKdEJPgOV43AuwTV8/Uq6qOZ1Q
aqtdMVvtwDkJYfiuZMGC7LxPEX15qmQv2gOu5SA6cRclCvTzcSC7jLUevGYIoB2Z
QeAPCjOSTNdf4lj6+g4VVPgC/cVMR9yqjdkGjVmZXh7qjwslCGOiLBJBKID5qrxn
iu7WHpEHXbZr4xgMLAS+9W4/wvCzbTLhTjUY70hOyAurxZ3lyduJ5XKT2pZYVaJO
9KuxoxX4jMUKGAGirwwPKEeAhyPuHhb2ZJQ0ufZtxlSIWpUTIudO+yxDw225Dy6j
ntikOf4REChzTl/koVoEouboWNfyPY57WeNULifl3J8yF9CkcfsPIgTVwm+TFKSv
5V4swK55MNjxZM5Esnbk1ayeDvPVZ1JVPEKUcIx8xfWN0BGJIjEJqV1qo6yHVjal
nOhAx07f+E6fVAhG0ecenl8gu6Xt9p6/ActDA1Y2/apUS16Q7NbHSmGN6ajAgwj4
oPV0VIxWz9EwIwx+CxqCiT5u/1eCD3drZjPtQ+e/fRk84ZpICwgvW9m2rslavNoO
k1WV1tjHYkx/2/2P0lmeEPUDgTzoiQK6h3gMzLfU2gBg9Dg9x9YW7wgSBpYTqAOl
FCx/VVijBRHKz9u4fvyKVYVzQISKLcOY4ZiYup8p/XlmtSvEAv1fyYRAVB+vOE7f
3p4hDwz+3RoQBI/8kWI+khMDV4JwXMhFZs1ODy+NeimH1yQ2J7EqjdLa9w/+c0FI
8pLKVCG51mxWdnos6IieOg==
`protect end_protected
