-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
aHqO+nTZMr5/qaZw0Uu16OunoZWtUAso2KGzYZTbSTH5LEorUc4F5BjUmGfbgbO7
ANFsxKIEFOWNSFsrUQ5AmHKTxDi4kJ7LLU/kDxy6vkbDK6VTyuT5aEjTFSs03/1k
CEVdtvn9hIHv3Y/IfM5MzupfHRLec/ea4wSMgbE32FQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24051)

`protect DATA_BLOCK
I1DRe1n5G7IYt38c5sdDGB4PBn0zRFO4Ov9IC4ln1BNwmIBqczKdPASJRPriBrj9
y5p/sllUoBKXAhzog7A8OG2AMTxnGPtPwGgSYVjRyXbmN3zJUrE15yIFu4JFePQG
BefDuUB0eMQoLG+ZCqFRPIo4RubOgSUNRLIpSiZWjZ2gdLJJrPSXFB77oy5fZFGD
hiTgqBtotUihKd0Ry9SfgrF/0SKm0vNgoCzaoJNGNHrnbiM9R/qpRCIlW1eWbK3G
WR9CoIUSRAPHhFy5/Nwf9HH2WGrQRsyqU2PHorj9HPQdCjonMMCTRgztvd1RIO/I
kE8DfEaHVHRt3PUrIF/xEUowesVef1v403tc3pnETqfA+3ZCmwkfqSbfSAKhVlkL
tXRkjQ/DbfBg1er6t1YK9xlY4+WIoObB87mfnLqKjToqWPvmMaWhx/pu4OH5BYOQ
H3uFLd7Fu+qbGmMLV79wMERqiNrm+kvRsXcNY1MB5KLTfPn7KtAMs99ejoi0UEu0
cFy3JmfmlKomWLDOJnt0CF17DaFcKcbs/IDvY3y4q7AMeVRNj+8vsug7VRapH0vq
F5FzTl3zG92dvt+io8jP/kvyzO+HeTLjKUi7FK1iW8nD32aw5g4U7YPexm6QncNG
fKSiHbr6YSnnnXvrk5iQJ/o8S/c7pC+WhlWvNMgmRnxR8BRXDEtetNT6tVDJBE5J
jcQ0/hHeYPYBh1yxTvS4DLQMkfQF7vjY9WXASQ68F7AMUoyxv93qX38FmQqNY7vG
WEiFGLo2oObeoFYrZ/pTH1souncnDjtq2t3BxKT2GChx9Sx9en85/ljAPo3KlXDG
I9UEe8g+or7QCNg0ptoa2lcPPyqPg3zKM6CJkade2TKrjyhxc0zG4S0T2DVeOfIl
7Z4sEYZjjYfMdClIbpKxQ8TuI3uGx3OJVN5YQdeGOaHSvhghrkUVzUFhbGd9T+Xk
dO/MvLxWRXGTKawaR3WhaW6Le+NtsotoI5E6aBfwPmmtozqJ5OdM9T+Jni3x6uqP
51VAuxRlRVeyarn9hud66tSMFv4IbbksbArD18WDvlGWVa8pKAxjtzDlF2ZPaB75
Z4Avbh1X1ClA+WQHS2c+BAa3a1DFr/wG/lDmhu3KVB5Uy7zYwZ9cEwlgXorZ3qqJ
tTuEXmmhMynrohf8r3eA/PwnxMaMja7pSKT6pruZO8N+5BRft8CQq0U0u1Vmk/9X
9jOmHliosuTU5AjJd7WemJswZ8905ZMJidEl2tsPb9AZyGIGhS+wNK0WKrmmdb1G
X0+8zjMp3xYzL7jePcENne4+EXYX5SUNvroOaqJHnQRL/ud7Tt8YXdH+TQTfOxQu
Bnr89UIHOK6zEOUaGPoI8VKZCB+eRs0hm9fFlc1K4ZQTnon2XC/Y7U/PCIDTSpCt
HSdKFb6KLWau0axRHOh0YYYAmm0akkWuQExMram3/npHcx2mBIfCpdi7gLHamuZD
rBYycg/LdbVXIOON1cKcjlMC5vzzhtEf1YKdFewP24W7N8vhl8y5H3vK2omuTfjm
242DaqqNmJ1f7lAO054Z8VjchZaLJ0lXbptSOMA2lbNimlXkSmJo+1ZFdXA1BIji
vwS8T3rar4+c6Inf6zxR9Rbp/b+Uj1rmVXKK6+zDyJ6bFgWRO3CUW7gTO6tWPERz
b/1CLqRloJ4VD6GeQIOQh40eng+XoQWEeLUITZhJaOHohF8l8eVcj4O17PR6XIes
QMK1CtG8Mju6GXUL/NWY8+2c5msGAmqT9PE2w3oM7/xxWZQJEeHv7O1hAjf1TBWT
HA+1J6AE5fYy3/oZcB0jV/87gxw6CqmLFoqJ6dYuJL3c7kjl3kQPaduSKqzqIaax
erJNq6uHcmJ68zhZTjNJQ42h9R5LUMcDa/jJscqJ8SRdWszCHAFqYmRUpmiESi4J
ok9HVI7vXOKrlBBuLX9lUOkTUOBleHSt12Lyr8KgiVTu/MKnA7RBlASCWwCtkIBA
aHOCAQdT5+9PAi7n75P7SLi8btCsBuxIgvF97jyD4om9mEJDrDk3L9fnXvoNtbxb
v4ED33uloIBtlbxHWDVJa4XRxNcG4R/nqzN4mls/hlIPzGccNw0E9qltoW5CloxQ
Y0j51+62oAzvKGVFd1bRVvGgSBF+tT4cLMQnU0cjipUGlJJ0h9g5NsRLDFd4pyJY
TVfIuPfFlNgi1Z9XR5yUC/hCm+wwmpc2R05ZhhWbp/jZhxXX5OQbMxRTQkprgb4Z
UbcXTjmlfZWrRC/C/JyAn1dkOV8o2AkpW6hZGOLCLtLhh5ff8/JjKHE1ksOpgpK5
TPZwKNfPziBWfqGYVoBmpoQ+4u+kqWHBG8DwIL1D2nXrrUeHZ77+WJ5g/0NGBjA3
5wt/YIh7nTYtklldPHGkuFW4d00g+7d72NAN8435hofLLKb3PXdOHwaw1RF4C9Kk
TNJCg+qj8K8brsQacz0FSsojZgsDV7Gr7FS97XST+EcGPz9C1l/k5n4LWSNHaHKb
YoO2ytkJF3nBYI3Ojq+YFPIKtJZsDXhPnhpJOhXmSNH4kUk7CowIu4Zdv2xN3RX/
3meOCy3+dISVgCbIKqTZuUz+46MRGNWqztrszpUprBgoYmk3+hRTfPg04PJ8Wm9u
TrlQBoYlaG9zTQ00N9nzHatv0Fey/TiKstKDVJTJL59e4FcarTffZfIw9FM6I6JW
wtbENXyR0b1IxyCRYkRQPrTAOl2bH7/AnZZLiSXRGWzStRLwuBJZTBfZaDs2f8tA
i1DekJYMaVKcl8fUVQQc8TenKk4YOtGaLChfbM+WvV/VJ5xV14AR8NVMbyUV8wRR
NpYhw6KIYWVAslY/rnJ+LH9CzpZBJXjf5L5MeQHjNIDF0up89FpQgX/e6NOaObA4
69vc6Rt4+iXpDxxvKjoG7Af7OT9evrdomaDgLKnRvrCXtAzVVtOX0xkj2Hg/xOBd
9O0kMX2UKetNv83C3XEkvc4GsjrKF/lz7FvN1OvcqRKS+n29vjCR4k+GtPbAPFIc
tjSY51VgSM5MU4lIx/9xcENVp/LgzNyKVmGK0CS2Rq0C+74SQ30vGD985R7yVvyi
HIgoCYKMWS1opbshqJ73/pICmNg7GJtZORAxk6noBIiCx1ILQMAdshViepL28qzI
Hj6XnYyjCtMMQfdRF10ehABp/bmuI4HdBOaZXD9eCwhWD812hMRq0OrvvQ1ogRuq
iGRFivftYJ3Uf6qSfrRLflD4w9oEZ35Fi+OATOsYYN64ZglaA2AGK4lbxdeF2pvz
lZeE0FSMQPkljhTWGLeOpqWUbHYiDUeW0qiun1nrf4OgTfD/LzYWZ8Vw3ZGphCZe
Pc4oWz/cYgWtg9lM274JvXgqXwvRWhZ5bfOi6mHSfnho5rS4soXPsLMbgEzqEnqO
bI8myucMSZMAumlgMcZ4RYxcCC7c4MDikmXpcMWYJLlanmzSCECTkuMXQdSTVcJA
EKD649l6I16lkOSnmA1MKIAa4Blws04MFZw8Qmss37mFki5vYTHVMGdXvgIuLDqt
xh3Zf1zWtMWSQDFw/UJI+Hxr1Ld1A5I/IC2Q4q51HD2dUmA2Vslc28jzaCqHK1hG
z5QuFSQ0gTKEWy62oSu4HUFaxzYzkB+qY6yU3+sxN5DNi52lMMvCAIU1cvdAd3+c
g7fgUVH80prDb03P5EmqVcyYjyqPImDS7hjM5sddmn7iANQDmT47CE8sc0lXmOTN
eLvJhHvw5Sm1K06Cv8pr3p2Ho9FGAkLKpU9GWAQczQK4wUvjL2zI5vWr4Q1ZLilR
V8RyB0b0eYX4ILLLax3jrt6j32fimO0PoiJ9s0EF3wJ+I74ufcD2PHVUGBWEtaej
lNIdImS/02aoxMm0b/ssbmBkqhxDPYbI63ulFT0RgZ70ZkxETF2jRkN7IpzuVpoC
n1My/8ItGElw9Soan5hyE+wX0GOvaXzchTKAfz0NBlMOFER7BEEBar3iscQSgVz/
E8QdPIE9qAbAyq1X2CcAQnuytdkDfNFlOhTXJObrfMwmh0K9dpxBqiP3Z1uVMZyU
Z9lktjVzOjuF0Uet5axiRzoJC/d891hUeNVWfC7Se9+T58oEKxu0Jd92rvPxgxGJ
wTGXkcGvOp2/YRwHF4lyOUpdhCEB5lB5mI8zGnbXwh0Q5bBlABl3HLDG16kjjoA9
b77mS3JJrw7KaGqm1ZHtWAuu01lTedazD5DkKjHGk/vc7eNlU9yukAtrEvfonH7U
XdxuzN24gDfwKkPdnGCSkgD2+gZjacJXnAwgg71PQRwzV3fXpat4FEQ81BenGaCn
O0IX9rhdGuwCghkommwpvHrc/pHa+4tca2k0SBYsQ22QiiHQrVS4rzrOc4leFfRY
MhjqrGRN7usxgki32Ubk1F2v55uQqb4BtKiR5g8cvU6EUqYko2ROF+W1ib2WlMhI
wLoU4zPf75w6MT9j2ACUYb/anUtlgtuMl59agGdlz+TuzyLR7t9ZqVq+tg17wod4
DcRzoMBzlNp3b/VRhIdDSB+wPa6yYi+gwLvdO6wb9sWESg8DanrgZOxjXQX9rk3k
DldB7+FCqBhw6lF6kzLsVS4dPGDB4dJVeHp3C/zIB44p/C/Q+IoubPhatwrWJsNx
Uq7nlEvz0JNs98WjS56GhJVU6zxmIVVFWydd2ZPtX3HmyaOk8DrSbHntKurzEoJ8
3hn3rfmEJqXBLA4V8VPDXWQNYthm7JyfKC+ADnxDCwfuuHXUn3hSgib7MD7ec7By
ghKekcfjSZr1cRod7XkrJHm7wPnvzaIbdEqFTN6dPUfwkZ5KFZ/FmZBuJjSVN8g6
xb0suEnV8iGqn3pBgk1lTdBgW9U9eAP0Z5qk5oLDSVdgghoxphBQdjCR7Q1DSsd2
odrtxSyNeqE5TeBr1i6G4R+OJMnm6ulAGQAxUFOoSVibmcdTbhQyDE+LfS3+MOY9
L3vSP500IWH62DwEDE8mRiHkOPpakiNyHO0e0IBswopLvFmk6GQltxwlhdwRZZab
QITnEUGAG0j1vq9UyJJmWT5yN7CgBhCl/ZJ8hVCHcalhqGxdIw8vXWfoYCOE+CXI
rCvKLY6IOsyM3ZRvOJOZmgEGYyE/h4PLt8Blqc9FqwJD+jhh56BGx9kblCbtq12F
vPvanKG4YAk0gM57rlDCC/2+vpIwHrj2DNpm60tGBOAoRx8PMRciCPkwdj5eIpXa
U8tZGbzkzKPjxMPg3UPggVQJaVoiOnLRh/FvfKTWtmQdLtn2LFlobIBCw9cQ1wEI
jfsAtY4SaKgFkShsFykc9bZ2HKKPjKrlQuLoftBhgpOTlNMpyBatnIuFJ7+zo3cY
QzxFnK5lKplLLe6GBN2h0ZRoOLcWhXj6Ut5i1CyF5sU6SKjP5WZIyQyO/SP4B3B4
u1Mp6Nd6P1gbaVuWMSDq1IpjV/noYhduSqW9KxG8HOOjAwoXSBgEx/6HQ71dMMLT
goHvMfnatT5Fj5ZwJ0wr4meWrzOahDdzQxrAUD29Bn2TNVqL287j0ATQvOJOWMSe
p83bBqFHOa0NPr+Z/4o/VwJMnoTF2GH29yguQZPibEvzdPOyCKHIqjcdQOSRQjlW
1Bxa9qpHihmpMrAKqG3673qLalbzKJi0pZbft3/wj2pDWg8CpNmIL03NTWYRSv3e
/hq47V7gTc6Ew6HdD+36orGlsbHo49fdlb4y4Pjgiq+TtR/vcexvjRsUXhktQK2r
SlR25UiDi/uZ6x48+xPGCb6UmT3L494lS9dspUsL4lUyBpU5toJKrrEv9pbVXB31
DlVnSt/fxFDRALdwZdItyFymQNdtbK0YzKd9PmUt1+fCi168m/VbfTqpEc1PTbxg
Tc3VdCJsHSBlASlSR3j8Xtxz4BHZ0H9xz67WqD5+M7vRUugIARcyXVz2cj5itxxJ
Mlcb9XJCmX61VtfH+PWB27LHG0rLqmlw2M53Uoe/jFq9M1NE6ndhAWo2XT2hHmvT
szgpDTgL1F8TuzVR86vA45qyU0OkDF0MYIm3MrYGvLWWi/WUSAq255p9tk1O29Yk
QwwdAsByePn2WdHukM1HxuD2W2F6P8/HhY6Hp5g/Q5b21o6KJ379dtP4sK4lzqJw
q2oUcBYSoVL1Cr6EE7vi7Xj1Ka6UXO/3GWjwxn2gbglJ+PhtdOWgc/tAKg5F7YJz
XcGIMCP4kVkQaR3YhLKZnq4GITcf4Q+FNJc071G7WL0hfnuEh7T0TvNg3CMipJZd
0PyGpm2x5svlMkEHqNO43eIx1yctKNSanhiBSLbzGhZtycSI2CpieYNtJzNRmfXW
AJuv6tYxL4Z6zpI/LK5E592F+ToeC62MsMWqk8no7vtVsZ8wwQ2Q+v4Cj0eiOldy
ao8i/aCCIzwuY2BSVLi4zXWJgH4l525DUSDXm9MztsKSQl6cDcm9MaJsYdzcOOam
6IEaTg/R7D/vafIP3m8mBFp7geRyyTvKFsSeOV7+yOZ4cn+dxSjnZal0WGTen5Ja
sKwkGFQByEazy1bVrCiJWV3YLivFIPp6lZ/YjmMddNWr14gIOZzyhOXQHl6MULCr
luCR85cNgj9LDLiquN2dXQh5Se3FLG106HNXavgP2F3gCKVF8y4c4xKs+eB3655v
ilWFul6ri7bQtxmgxmt+qEZTvxxQgpw2011S4Do6qf34qZ3E5k5Hvxkj6R3qo45/
hlCps0eSi/0I+X5LZIis1FIrQ11aZVys1WCo0O0INmvjX36jWGylRGH1n46FeXDa
+2ULOVOy8XP5vjh8SGCtwKXfqVF/sjoUNV4+vGmfbD2n0vDeofz1s/ig2mLVTg9I
eXc1t8lEelFMEkIsDI1XFIoQx5HF3ntzTG45LeX4BdjnV1kqN0yHP8eoZZe3iAoa
67uc6nI9KTBxwZ+J9tkw2nZ88qxQXI1MSOg8X5Xp186cRGa0FeSSkV78UDLzfENK
AeVMPb2oII9loaNaXGpdAxyr2c/qJu73aoZf9FpVJiRnIyX+NhgcPm0Mu1Ec5Q2L
CDmoqP4KwIP28P7X/6IJAz8l/pk4sqaqemLqc1oY1BRAnYfY5//r2Rj2QlVxXVA9
PqNnqWErU+SgbcYC3NVGIH9eWMoBI0zt6lpEdvOyz+0qWEA3yitGyZ3/T0ErzFUU
nYc2mXnZ3pa/4b5Y5qtwb/idZx7T+2QzlQMa4Xum1lDiZsz8sWOcTG+9tSeZWcxf
EjEWILouC10v5lPG05aUvrjknMdhCaJtIYN/ysKeqEA+NF7RKM6BFujCC2Tyd+OB
1wJwWg1X3+mvUWYOKJdyTI7PoONpjIAJRMyuKM2poHelSwsJ25IjLKvXHVOxh1iC
uqSTwNUm/ae/TZytuKTSlPxtXyLkbyU7p6oAUQt3xnsirV6BqpmL8BoRyzXr45rP
vNg0VoJggAqk5z8jCIZS1ZM9GrWf/irQkPNIN6i8qp3HPsWhFlfyfownRLDhZxNQ
g9Equbm7iS88wK/wKkgsXnWqXGOgvGqhFMiRHGcvZJyJQLpoH14mNR5UTXXIh8Cd
583RQJ7pR9Hc8lJQn3Fq3acL5siri5FsYHOk6GjL64qhRX1/TU/fgzK8+1UsfTNc
iH2pJEKd+oA9UQ2MogvgaRUL79mc1fKMNd0wCucV7vxdqqOl48HXW94a7qVsb3UX
NXyvvnqHF2K+3RzOyD8AjbjwrFVMijM4GbUPCgizi2TK6qnQnOoumDadR6QfKBhI
CJcG7iGXe1ZiNGRYLntinHmQo5i0pTxtfU6oRwGc8aMsHYgSrgmuHpVm6wASUmYp
bfqSrDNJUk6d5UukVh2O6B5Z5X/JzaMTxUZ0s4CZjDTDng8vVHf/A+7IbUD30O8f
tne2GrSHv6FcCyXOD0+FB1BTmr2/zfiATTPIwSeCPrUhMEV+3k5yVyJQPoB2ilYz
w4vW4hYoyzzdgHI33Ltvc7u9FJSv5j8AXP++bZGYVx56so9rchtJMSsGUALzBxfF
/DUAvV2msW+wEY2EYNjYdQJNXLXw+I746JYk4rrBEtU9N5XGwzA/lA9QOvHYLChf
qq2mQLaJoD2McT8ZaKt3IXNXLm1gWmWyY1jb3vY9d1NTs4usvKVyciv5XJS5t4Ym
g9Pu/PScc7Ay1t39IdbeUeWvyYyFFPDcQFdE8c9x7Pi8AbjQCM8lszBEZ+PHdOAn
+PqEirp7hoN/Kd4wrNm8bwM+7P1ZIKoDcu6nmwT5F1NTD1QG1cy5i2SBQf7uYNOt
XFYbF5jxkOWfiMciYbINXbir66IpKmIxPtgcQ9kGpTNnK8Qc8DJsuwb5M2mQk9et
zSn22rJx2BHzBO9E4oNDkqazbFOqhF/0B2gRw2nRh9mztb6b3gnGVI4ur0hj0rTR
2Xb1J1PKmmsB4h+oWcT7dMwLVTTFcVQwXwzuSi5IfTvdYZdQv82GTTHPH40hDAcl
GCKuEEbNGVrB+gW+VPbfAKuvSAJM+pYJywa/zf4QaPsPPu126ZPeX15SHekhcCaW
jcEPXKfjLt4h5+/kD6Pu6+HOuSewcfTTyRBMq2pkKhiBOYOJlHbVvncDIoz6gsSw
E0VQHEFqvn92xR3S2e3j/P+EpCcBX+MjLZ0UcNvW4iWEpCDYflVhUL5tNA52slkI
JRpanO6r9b0ERndGi1/tVTFIFKxsQi5MXtBuQu+miTVJSVZg5g5QscPFY85Yomp6
l6AVMDgFno1iIdXAA4ud4M/nA6ZEQc4iF/C00ZWFnpPa3x//3gTIrSBAqBKqorPp
/Nvz4uMvu0wF/x5qecTST607HQU+90+z5AlA225+I0p8Pdaq1TobGKCbiBpfhWxb
EnQ2duCDRPPk6WvQf1bYO19cQGSiFz0NurpGiR8a80C/VxLM0GUIl/o2N/Sb00DD
HVOTJlVJFukz/+NFU5yGfk7Nbfaex+HqBY7OHVakpKEmn+SOL9PuRYJXT0vlDRtb
DyYqKq4/GYkJvu9G9+wSGbDPneZZCuNw1qrR7WRigGQTc4fGjWab1DglJ4NDtwsY
laB1l1GlWW2PW8hhYGo+A0mmFX+jhYD3y3+SoOWVLXWNnYTCBVBKXjBo2r6Y9+vt
vuPIwoBpxrIuW4//YpEB2DqdZDoce6q7MGK+i3OueokEqztJjG0HsMZCR1eRgEhD
LdmLShkS6KFQE7qHVJopRm7DAw+K2a50x9B7BWsNeGiMryicJ3KRYAFXsK8sxHRD
m42cUIyGGbZ8TdqMUjfCyBNyxaDGzq/5Excs6uelCoilcqL1tSC1aZU5Tz20Nq1v
aD69Jgs6/y3IhLJOtl6+91GTvL1zPBf1weRSNXsh6xp2+YTmH2veEPh8sw2Djwe7
DkILwDlSy7Ssb/gaAdnshYY1WUiStYRiRZkRULj8KrszN8cCOzsRnyDR1zWZpYyN
h2SzIXN6yoZkezvJxnTv+VLVHRdgQ/W9ZXElbxzrgnO0uQPYJa8mzZHMYgORSQbn
XswshQIVjtJ8GPfb437nqR49C1LrLpSWG4g7zXhvK6JGVCQYrC1+jxYSpcqdc5jq
l/lcuuwxMezuYqUOqK7bi7TqNL7gfxRWI6atbQZG2k1TccsQNB8dAhEEOVZ3EKXL
0pa172BG4jyhXU+piawdfifcmOWwcX8Qkip4Heh6ExO8y3WNRAem2UAHW9sgCDGy
3wyv2iei88AwQz5d3bwt03hnkORsCaqLhN/VC/fhggUPjvDoaDJMOgTfkEArwDHO
Wc741iOspc1qNPMNWhE3h55RBCzD72MUy3GiT5+yoHMsGH682Cgm8z46Kwf9io11
bIc0Afl4zxusAN6cYAxOpwe294HVeF0y2StTCCmQV0FQwpY/XYOGShG2hM+AXePl
aQuP0t5Cw4dScUrbrH5i8DIu1BWVLHKteRqXIgFlqpFUr/Dfx9hxn/saM2uqodr0
cbIG2I8Sapblajqd0eW6aaIg9g7SifjkulWc8FWhWLklIooFZGsA4Mxl+NzqshGs
bIRJ+M9DaW1VAk6md47e4UXVpwuB+YO1cCdE3UniWCfzq1vuoXuUG2yP85ZZ3vK7
4Ab2wW32WNpNo70T94KlP7wTYli6328Ktt7sXLFRIjan5VhOzCHCs+MEndyBe2my
gMSd0Bd8cjM7TGEp/h8uGq8ns6T8OG6QPnYDd4oHz3rzbdijMm8SZIlEp6Ich4kj
LLh/o5o+oCpNJOfvBOVdDDtfH+B1I7Ye1pQ2TlmlUcGWeCckgo+o5vEmo+1vMx/l
TlpJomsUlVM21RyfLpkWwYw6MOKjfsFRwl/wcj4vMLZaJblleOfXO4jEkSfhOZwZ
QOSjhHPqZFzwyTJftPEWI8RaEfa5PhASTfD8BUtonZA7gEcp80wex3WbETwf3Q4b
rXnn62uAeah7Lcaqbfl18dZ4WL61+AN43cVR4N7dm4jIszbutoJ5imb86gRjRRm/
RvvWZbDB5hTHO8pvjLmWmZN3n8QbjUZaZMkzPGNtm5epwkRjgLIju8/Hk4i7LS1Q
/TMa1aHSHdpR1qgPg+BX7vyd6ZyEbH3lZ5URjRW+bNB1a5fj4Wz3vJ6Zxnk40pE2
NM4tVleNIC8hoPz3ehtx31LbvT9v1QXOlQiLmsPO/kWmaNbIqRpP4DsjmQ1Zppus
02JiW5oFuvD+oGCRmFqKhJu8TLmL+3rKUm0SJ/vuJ8ST5zF1kollNQVvuQvsZACo
JvL+VBgfJTqXg5KZonmhkjbVGFMaoPJMN4PMS+VY7bUtYh9LbegJDxt0lNe+5HJi
mcGi3+gYdVu/p9uAhPWEIkmDHFH/Byp6QhXH+/kcd0wSRdHVPMm7Gw0HsbVx8H9r
q+KlfBKonSaP8yj9RGmCyrQzx/xXUvkUSQknJ95mY5wMVZ3L/6WwaJPy3oNMWoKJ
qg/xApvMyWISws1vTn7fT6x5+75LGPPWg3nKysxdINSgv5UFiehAw48OGMn4zGO8
jzygXHcnjJqBiPbUoXbnjr2UxVLTbc5VmSH+ke6GchnQlgUecWGBZ3R5fzDH06uW
i8Cq+sG4k9Yc5Fn0sJRu5QdQmyqxf1o0jEhCZvPwvyOvy/JzgyvkUd3aT1ydCotk
pB4kb0y0PYJzphDN7O4rYI0D+9XV+PgXsbyi9l6SnVf0cgmmjSPoybgKeJIwXR8F
/W0UXS9ugoaJmGpYQ18zCG10mZInSeYh9Twyl/pE+sX0YuhTCCB/6cQoXxj8HpXk
F5UwTlmKrXeeFvOxSuif2GBZubQFTx+yHOTDTCvjHQG4LN8Kmp9PHozM73gtinO2
lf02CGkM2dI+Youw6gBY0ur8C3ubjhvzbgTeZxLm+Mpbi9m8wGLP1Gvwh3T3RwhL
m3rv7cwqhCuaNn0w9b6IJ87THTWCz0yCg4s0iPGa/7DMyxp2O4fYf7YGu37sIfuR
aD+LTSNQhXj9NKk2yJPgatD+LmNXk1N7o8mwP2cmC4N03CFv5mi+i0C+DZ9ahlo5
4UzARxV3KJ/AFnsjxGFt2IcznBiaVsoRZvMR0Do61psvZLekDrPVdQijzShRf+sl
HNSmhva9PmeJInmg6X0g2BqLOMM34md6UQ1oLly/+eW/SAUd3s3QJrtJ2/sBjzje
Os0VZOzaSnB8T7cZH+B7RODxhmvCRvhLQIyPLNWma8hC7UhSxN39nfwskicmDLhe
2gHmchydiZZ46zeqx6qI55sKU3sVwmDHLg0eX/jN1Zv9WxQgOHSn1E4yCYntRyJO
XAiwXNzfkh7iDd4hn65DfhnA8tULqSWLUNb+ItrrYjzDoot/PFFx1KTdOHh5ACx/
x5jtRfpeY+CgW6YtTxa1g1zatzrRysBBWb8DxmICXQAhvHafOINEcwEsJE5X0pCd
ZrwPWOI+lRW9pZn8wcAEx4LkBJIPkB+0F6GJpv2XIu3I+0XpBo6ulMbCIwm0P4jN
aaz3+JfYEVmkHdKq2GJ3ShuBm11sYkCPWiyLJVz6lIHbiKu9yL9yWOxnLAnZiPi8
FGn0JytfRyTggOeNwuyZr+B1PCsOUqRt+M3OgDYQg24piAkuFkJlMZ7KycDv/QH5
wgO80gy2CMgH3/JZlFe8LEYFgDbMFeyGqSQ2YtU46Udxu/6HFS7t8IBl5BH/VdUe
QYc/LWonVgvj7lQw4Sqv16EnIs/sA9sqq3gP0EoPDlSJfv90DAq0NujPXvfv5MVc
QnBUbXfBbi/cWy1bpFhD9yY34GSHkbkbgXwNcWnm4XFyVp+k25oKdKdyBU46pXcj
fXNiVEN3BEVoc9bO/OOR0pdWaHSZdAxEY4NtHcVQDVWVbWq40Vba0VinN8xA7pOG
iUA6hbDNSbDCHEnlXlKVHe+ns+fOCin/9FMLRQmFyNYXR/gLFZa+fv/LlHi7jjoQ
PHAQ0PPuq5teoKIsPqpf1oRm6Q+aLOyOxCXhPJtNG02uYdSDkcrOYt74+d/btFgL
+jO3C/+7bre29Mc8MGz9liXNCpN1TLQUpz2la/3SQROg8jfbfNfhtwI7QEYcJJZu
e8/BFqNchy4YOmORd89qas25Q+j5TVVeqojuuh6orFoF30S/t4cuvcnz9Fu2x3Pv
qHUh0xHwDVhugxpQwhKRSoXukWcJzrCv0B1X5yGIK+guDc6jC8puJ2VacXH0b7GR
7h38Vzd2uucxhkzhZzXICuYaxwU/+EQdbY4wOyoIs90eLv1CzQe4WCKOPDGuyoR1
mMqMm/p19ecJqaTKVdMFMgDSoZRt6WxPixpvlNRvY1MGezjBHyzGG3u9CsSko6Va
k/kweTrvPweQf9qCc94fpZ9w4GHdJI1yzS1cCWqvC4C9r5I8t3NZdCldMX8kBFY4
FjRCbmfPWCrOExnb3Eoa+N7g5SyfmZfCQcFm5cvZfddyjM2FqbJVQyFFHO2mSJyd
NkSm2RddAjau3xCOUkTMhbzlbhCXDOY07WUNN8JhrMSrDUO6m9GAhQx89vHdxHfL
Bto/GmHIlQ0c0wLY3gNW/HYnxkOEVKg33v+clO3CstpqJ5mYwRhLeIEQwuJaR4De
7/+OIy9PIlEzuHVVt99Fym29fjjPVybDclMugChmDlB+SOSvyOMx6ahD8/pD3ivh
UcuFwutI6gBZ+vTa3QnxDODw66KJ/d0mIchRiNCRM6NsoA2mbzl7hiSwMfaU3EVS
FFBR8wABgGTafx31olRLJPFVc0exxOBfg3cQUVaq18CcViyQt0i1ORYpsVNLX5bn
b2JDfnHroNMayY1NuW1LlIpY1kSIrsho7xE7eRdJt4x3kj6m5xukrkgAr9B8Lz1a
40TovpejMmhNT3e4TgUAsjLaVjSkDiwZpwzur8337Aml0xXVFeItC/8ZzpJn5i05
5XMhBGok/VB0euWa6kZcZqytXFdGfgA1YFrZM6re5XIdK5L3h8Xr6MQS3tRMerGZ
oIeiHcNTFAVUilY2OpHSm+MzE/Wi87+aAFt2u8/437tve9zD7Q24JqeRCdgsVORb
JReVpbf/hD5rCaM+A5PpYwqmjPDmz7RDiX141N6bIOnYJtPINqML1ahWa87DO+St
eAXk4Il2Rd+WOTqdP/TklD7u7L0oWfv2DePv/5ERaMY1D8TMRHep33RzPvX/ZFHt
8fVgU7CV/Ba4q4/gCJuOdt9YGL+fBqMl7TkMhJx5QhB7SeIP2BDdWIqxVb4MRHPP
XGSdVT5xovG6CdeuxIXgT63B//S6UeJY72a1bgm7dWdI4SWVu63kqdfVbqXhmRMJ
SSdS8UA7naUa5KSFv6zcAOGsbaOXN5/oJiqSL2Xm/tYJ1bDI4H25fNfEktrswTTF
eTvw1y+HNVYUTczq1VGhR0wQ1n7fBVmM6vtO85nG0H7J12NYBMev9Gwr8ak36Mza
t0AdFJduKquIgfaXKGReqmc1bmexNdSJejN77Lq0+CCvjCg8ddRBakZO9WBfu+gN
Wwzfd2Ufg9P42I9pRYIbPHKd171ilVH8kNmGQnD13qPIfOiGyeXQu6BTG3ysaFZD
gXVaQ4xMgs2WYVgpa4CQ66sfmU4KQMRoEGDgnflNd0YMVTRcYn/TekvOgkfvyIeu
hoHfUKyy8zmOgjPBZ27zRF8vRksexl/wfINSg7ajI64G9bg6yGJO42b/YUOCFkNt
tIcih6K9zMuY7d78z19E2BEdF3wEL8VuZfbu9mWJWIKZwFwyabAYwkZYYXQwb9e0
WVayXKMTSy6cqBthmS4+LZ17TX8hsdw/bOlBK1BXuu1xEViSHOaBnDRTAcUu0iCe
qYUMBcletMWuJh/Wh4Zm7JjDnrKKn7Kn0RCIcJQoPk5k5HPEGtUXqCAUezuZE/iA
Z9g+kX7c4TZB7Pv7GWQ9+HM0+1XBKdbqagpaub5GuiXhX30C7I3lQhQjwCIf0dZW
m8IPTLyE/yPhcHNsTQBlrdtgSoO4n0ljUrzHeWWgmfBcJSaYO4nAnH1iNIjEqr4K
T4tlWXKtssIR5oCS96a6a1D3uth3KniufXslMlcWINPLuJuL57r/tSzwKgVzIyj9
YdS07/wy/SDftleatdUZL/67x3u+vz1YwJhbcRJZtAjYHw2OotTdZwsRpgVKqxY8
TeI8DQ3MlxoYoX+gx5BXyorbU22J6kgGzxjZh1UJoXcoL7jURVuaKz1HyGi7kA/+
VyDhV3hRuVIFcqvqFzX9uZu9dOs4BYNZMeouVNverau//N+W1Vtz4TR3ROBtxmqt
XWBcZvpa90oCOLZN4kOX+AFrnt69dXIHsqxTL/Qxw6D5s7OzWGaGWStWPL6KLxjS
zlLIUv7a6fp27ARjfL3+bjcknNMX8Du+6Inph1BUr0qz+XRvefJXkrbCZ6KLTuye
tjgDAujTk3WDnTYOe4F4oT0B9gvBvjx+iJQjNq5+7h4jSOe68J3rUZkfVqtboFON
eJBJj4wrurUl5aKUxtKxGnCE3TfLgvDs5pSGV+67EEnUdov/HdqdXw+UMT6u8A6s
QylNbWrzmI3Xv/pegix9M/eyq5BU4h70D+qghEDOW+aHrxHgC+mqxTevtr/Ejmii
3DXHfANJWnK1INMIS9jhrwZmP3FPm6g7738ghgyaxwv7dBWdFkfcYE/GWMFkLIFG
JWFWHCxBKLLHLTbkpOyEBNPJTtawKFHLJUvAktDOm6CVlPmGAxDRvByQrA35Cu/c
8+rwXDfo2quv3cUZdlhdPA6eU1UhbZ/1CmXxkYZZ9OQuY9HuyUUvkZMo2rJo2J8k
m7UjkXXkMyCt0zxQaUCYQgJ8gz/D0qbSHVX+5PcWpFqJoMn3PjuTyVLASXZLYg5A
AZ8Jq/In6NOtKbPVH657gHVcnYERmrZZDnjvNB0/GkHo+uX4Qixt+8jUCxSAqlK+
gn3Lix8pT0fERltORPkSxXCTnVk6DDhB7X5ZRfqefVtvDab9hUsJP7AFmZdlsVnI
Kxh7ctEwe7ndSFcNzS2vflC+svUEdOLTl1YTjqm9LRVzNlS3PDgQibwABdl4WQw0
18kffTSwW9UuYuX6eiBFBeCM4109p3ycFV/wb98Nhb8grQ07RG1vsfCxCwDjVZrv
N/LnOAoT7TmBY24TQaLRhHzEesQK05Kqo0P1bB6Fmq/9IPIwG9GtafGHJD8u8H+r
Jn6+C1K+oiACryqnlEsDuzqZHjnFYI8dJ7zwrfNInu/LXnvug03AZb46Fqo8jXS1
TxwV6TRb/CgylzoRJluoQ5TAzlY/OPW0OeEJpzmwIotJ0hBb9ukqnWst+1Mlt+TH
zowp+MCExFoEHOw3NWprmeiqtc0pj82v/RQFuMoc/MJUULbcW+pPVXhkx/V/NMZH
tBkrgKPhmBycxvJOA5D8T+iOeFCz3gXNqZCcaQXFnLeIppehSvhkWTu2LKnG6wqd
unSSOneNMZXrPsdKYz3WqhxIIp/HNhagyayxFIzfipnA2xYZIxEgEYq9N3aG+w/F
SaGeZUfk8qwe0RvNXDjPTl8u8TjVXqJJr/AcjH/dTpNkHQwikesVTp58ENI4Sa7z
QyVqZur90KVlCAH3r7HIglKs09QOK6SEJticlfGfDnsDi/rOjUvQhPbtErRvne82
RD63NsdNlzyi+HF6KIsSztBA/BVmt+SCBrOShuRNA91a5edCJvyKVDTXxEQM3jZj
5FYVbnX/OqbXgmz7DXIUHmbEQtw9EgLAKBP9vyGEGmeOe5qh1UwyrqlmtgGQDgzf
6GzwKbLIS5zoCTfP5MCqRsHhy7dL4X5QYbF8knt0FuqiDH8XEAevUqMFT8foGE8C
0jns+9cnIhIlmZ9znWLF0xDy9EOJWd1vrR7d3BVXIYA2UB3jI/qR1BwimmqMMTsM
Y2oWrIs8WSrU1Bo7dc1Hr6HbL3C1q8XPlVOtAGL4IHvXj52330F2iolFtvBZJCns
JOmGoIL/KyvI7lCQnJhtauMIfbdwBhUdHDze98Ob81cpNx6oopVHC+/37ooeIFzx
ASnyWLbea5XTfCpcZEj3NaCBw5SjTjeKkhoKw7cEzZcvQ2jgJmhqnzykXX9FEqVe
XlMbI1HhZzodkrTgyoab0r6OPoBZbcRPF9qzlW3LS1AC2PY5ca8SP+m6ru4p5949
Mai8JRcJ36ABV9lW7cgom5QdE1JJGRc4vMfBYY9zxuPgA13FjDCpZFT+SLL8z00Q
F02YrlIdJLdipzxT5dBZqt0l1o+/WxYALhs+7VtI8USe7ihKF81okIQoFnnQMzCV
1zOYDFmJDI0McEI6M1WIDmJ2QjI0+IjXr+ZT+qAN6xJzgZ+i5cCqwcccODbynqvr
NDeRq5EuXVwIzgykZnXwNN+VjqCIsLcy7vVb4li+4ouZNLRiHFxz+W6co3KVq11Y
R1Xdxs9XSCV4XFHIpZHFEZ4yNKjvFgkZrkI4Gl/jDhDhtjrQXguErnu7bPHmaY2j
MYEBlnMyCB0klFXK7vaB/2GSewmgyIu4mfAvCqeqnLg4CoBG/cgtKqRqE8NqDMu1
/ogr5cX4QYR0G6kJJAff1k+ciPZPqpJH5EoDBKotdQHjX8SMbBbkhWZsLCBak6QK
DKeoe/9ahWWvzU7lmk+wRNqcjFi8HzUGzjXgtddNEndZSiXQGQS7lg0jwfqzewbB
uBO/sC9EHtJG/22G5wnvePCqu5PXiLFuyLhRjvU1WwyokV8Skg7ORgS83y6KhcnT
qVGVQlbW1e/qieM+PxvGrAMv1leMTVOILafJDUnLRqf6uDmw0wQhWPbIlWz4UJYF
mC8ngxbp9C4z3CLo3hRWIThLKWuEczmaGsrau+QRSfaa/4k5SOzkLkFn/tIYG+n0
9YGIRSMMO/39UITcq0JLE7Kc+PC3jaUyc2ZrgV206Pw5FREdpY0HLa43RYsPGEKU
903HQCtH9uCgTGNPTwByW4ak7KViYvmWjTeTWMhushu+lspdHd21CXNWJR29dcXG
HU7ElYczWP8Cq0TmBvvH9JZXt0G/lKjChJq27SW0BZb5XV+rMLDaETuT3v7Dad38
ZijcPBaH52h312v1TcHJcGryhlwaZ6sHBWobc43qDngHXTuHHWPk404KgtnghkN4
II1ZhCFNJV/ysofLoovNXh7q28xqbVLcsQ97Jv5CSQSFHnNeWNhqcSVEr8qQXgU6
+p7warxLqNDn3l+BZgIMaO7I3a70hZHBay8nalmyMrhVFmFmZ5I+6+zw7CXLi4Fc
a0aTKtoOuIzSv+0ufl1ahTqpam/LDKQ5bAwz5ft1ybUT5hXz/9ZWq4BHF8sFz1GW
V127jpy7hDJEcyxXaUVr1bdZVVVbsS3xeuzkLMIA4WW8fXGDPfeSwjp7X+8nAqw/
XKMFpp7703lLRrSBaMk/KMjSWgp68cH6mMg4dbJp9wR/SwMSlm0Z9RdTPfJN+76V
HBgrOsq12QNg1vngktLyI6WRZJdhmR4w8oWjAZqzyIwlYNAMb8jcfaCv6Mqr8o1d
/8XebpKh+ptpwOuRC5XrhmQlBfRRQqnjz8YIrZw4qH9mNS6tMrmxoxY1rR4MndQk
vECUR/On2Y0b/5y6r689Xle2+eYBE/YeB1/h1KLf9E1JphtQPZuUCLzchuh3P+f8
JHidHgFWShnCLMZIDaODpfGnbee+jScOCMF3Oo2ehF8zIGyud0NATRFqSZ2CpT2D
JUIydXmXeJhkgp5Mf4ocvgeef/9F6R8Ge0xQkWa4J2nKfGbdKTpMvDvbm4ETVkEc
00s0+0G6eZqlXqqKDkchw3tAm64JF5isxPJmQeyvc764uzwD5Gvq7DgDk9OpTG57
T2A6bfSkwIBAYrnZfRGKmF7n/KNbCD8f6BjiDQ2Ecg4/hKCnQprfHH2IzlVwhmNl
rEYoIZI0EWZCwmXuwq/COgieCe+6IuCK/8j/Zlb9lUjVay1KMjU/SiUZtVjbSy99
AOtIQEtCxP1EP1fjWoyFrXRcBVxDKO//OFwi1WuryNPZkj4Pkw46skrGKZsTaYdi
btin0oFGPZT25MWpomEN2NdeX4zReQ+tjkpmufvFxALx0zUTjfmxVeGjqTLbSEcE
gTUhQ7cDquPhgLRtFGbk3gekt9zOVJ6jlcWA1cFY7CjaDV7W4/1Mq3UYKRCY6GnH
dAkyaiRipDzwZ2toof0Po4Wknf3xAsEJvRntdvix75dy2mUe1gv52XWDydD9iE11
3Sw31Csi1Ntb4LgmnaFFpfH1evc5PVw+Ny6KItIhsKILDFspsv0Oo/BvA7CaTTPE
KKcC/6rRwSj95cM++oEAce1u8g9rqMiO/6AHRfpr94U4nKnZOOTdLIipawX/76w+
zjxMptFDnilo/IvvIVl2qxowP0uCu0A0SiLEfjgQAf/EDF3K6fKeZ0FYySf9nuDd
J8HiP8umdnvSt/njC5QmLJCczRNbEKazY6cHgBLmRqUMty2NOLqKvIwGXfyhPvDR
3IToDxRZXBJQFM+cn785n/RRPgIQTv5huUw50rYVW8pHKzQwq8JNhz/gMGVrLy1z
dHkCJGHGphnjcDP33261iDqdbIXaNwMOIOnxDzHPXPcaxh/Yw4zaZtRwE891xTcU
XI19SpCu1RlpSx/vY22s9OZEMThPm0qLGnuF9UJzSm8kmnBakJCpB2F90LhEDc/i
YTHPFZmm+RDjrEeaR29AgW+Uk2cV8cRRIVA+T7QQ9ex/G3FzXqxjcfLfvH3XZ3Y1
QXVqbSWqz04gn/UAVLlOMPMio3upEcovGJNxWYdcStPOlQhm1gKjSGZv9xMNY4ag
cYup+lvsssmtbCx/LGJ5+3Lpebx0oDwMdbkWFdSHto7VFPoohyr6IIhupXDYRsY6
7/nO2luG10R83vnniqw7rJ2jiJa0JknTVwzVSlTPku0LoR2oRyIJXvaxRJcvjBd3
yW6ebQDfBc3M6CyWkpL/QKck0DXEi6RxipQjm33tqW/UEAZLVkOo97bus8dNrwOC
RCkYck/aiDHoWAmUubs+1tA7e3+3uuFNzDqruH3biLUVzgjVi8Buh+8/RL/iCcbi
A4Sitgd3XaluFFwT83RhyyZY4WBjQ1AZpkTaDVJ+0GwuR+Hrx7HUnVOYkXfKYmWa
jP2AbpPhZ899nXYJ1kIjMhZlRJSSu5xjhcJQWGbdqW2z4I25GRinm7mTPTvsEF4Z
DFdOQrTSFt+2S6WudRKMWliHZhXCTkTiSTbef2nNM0bU5A0JpDO4b343SS22pvaX
KSVftd7wBRgb9saCy7E6aKYYuHRP54PRQ1h2YpFyuznMTQbe4BaBPmFLDW0Lg6r3
wct6VxayRzTRgSqXBKhKp2etStIN7lFD1A+nsDGtdsywovsxzEX1qh9Hpe6XV5K9
L1ANyYUUJgC1NgsmIlOUG9k3kg3A9lghYIpE4F40j8x1JlhUeHp5K/cWAQKnJKuE
BERVDia56sniajTCAHukezGRQc8VIOXJVMuOMUzEuBdLLLqKRrCGLNbemtMxOFYB
1iSK+xWMKFZZpDyQQ7mjH2IIDY6ghvGPfUpnRqDYLoKYF7CZcV1emEyK083mOqtR
gAywCh5dfkFzp6Imy94JslOpQO1tSEXu/n+xoxfkmzGc9BWUympllACkmhxSPs1t
1jFuvij/ZFo9Y3TwFFGEM1XEEYvJfCnq2qsHdu/6zUEtclhWv5sh8W8mDWkvmxl4
GUpEaRp11CSGfPU3ih41dGtNPlBaB2d9oq+XnYfsscgxeS3RIihf32FnmUJV8sEL
7EJFwY41L+grMvpIheAqsWl8L7eJkR+1avr5NvlUrRRsQKaSbdAq4fwF/9Dy90uQ
EmK9POqR1MIEcDvzPn/fXV3rbGwyMM/RE3V+LiOU349xNY96fTyGuwbIo8pXCutd
0yQfHy5iigEUWNT95MclyxNsrrDVGsfdbcuB3iWieIkb/y0Qt82NoUbCGU2QGDmM
JpBG2EQGyx15U4++VBy7Z1BzEXg3ctADk2YfXAg6Htp59AOKIfLqusystNke//l6
xIyqPbAfFLi3tysSFoe9QBmtwXTfi1lVK8v9+IcM7X9oYVJxueJYE8kw8Z3yQV4x
SIQHU/rbyPShU0nfpz7BLubb1HNxs8Bxe7e65Ed/mX5F4sVdV27rpc8ODem8920R
SUYOcpbmHfTxp/OOfpfWcxTfoEQMA1L2bgIdcIw7bGp289vKLmwvUNTBmym3jyAv
Kv5fUGKQdaJ5DhY2Fb+hjnc2WPPlIym+wnyZ5qWiphDfMSQtMIwcfag6KS9FI7+Z
xBfs2b257YX6YKER4+It1WsvJInUXYZqP2nwa4uw6riaUs7ZeqvMxPDuTCz10EIq
45YWtg7vX1/NITejKY8p5F9foIHfpW+eLEV7wTnxBhfUfkTxiN3I7FmBfHD0Kklx
+SyIhl5E8TFJsnNy5q3Bh1Ao5aiRuQCATuquKLnCxqMXIQ7UvjkgjeoWi2F812UN
Y5Lfp90pDbvdCFNmbeSrniKsidOdyVxGvr7evJkBvS0vc4lyekMwHU7zUTWtu39J
vZvs9bmMQxNb9l3b/4rJ6Jq8ulbmAoJXTo1IPi1iZbWBOUO8q5R+kooaa0A9vyK1
biv0vJyZloHn2SwIHPFEXMHjNP38SHb/tRM49m5gzPFnj2gWA2pVaCSH1djfbrd4
8+vusHyXr1ZtHmgkCtWAPkU2/m5cPeKbNwFWYI3IeaTC5VvulI38HH6sl74xDzSe
dZ2sgEXWj++YDb1+2B0OywWzYgfp5Bz855ZLckwtrkaNbslWKeWddjqSI/+0VZnt
+4y3cLpnmQGwIr/7m47BrIbWUeOI5m+41z6sOzqpJe8l0+cF23o+uIEMKYV7mIrf
lWx+tLAIc+WJLzzVIG3/6tj/g4PSomayXzoD29bX72Ft7UEzm8FNyJd5RaluzYqn
eV01o20GOWlxeyRF2XuqOECFGjDuFMYsu2wzlj+0CBidSNmdHiIgXcIZXWAC8Imi
ZR2LNoS4uZphaztoJfKl+Ma6DX4JeNHedcvPYZv7HOSy+jg4gfIy/4DPm3cNCdOC
skUwwDvjRVjRLDgRnjoNHpkuV5onEqSbLSNrGwk55Ke8BBVaGiZM6fk1W92XxCVa
QtaLu4TgEF6y+9R51SqkZwKoDNTi5cgK/aTN8tecio+AOCzem0e15WTnfeQmq8qc
XaBtQfa1y9qVitmETaaaK/LOVtIgmBIp2drhcZ31Mmj1q1lK1w8eRF9R4nDI4rEc
iyDQngUo1XFpSf6LJ8Db/Q6VfbG2emloZqtl83Z2lmTGjD0/6nTm4zsNE3fDLvP4
cItZy6fwrX6ElYIW4HV8atoDM1DZTscuylLLt4g5/I0PN9QZiivNI5rUEh99HKob
uEHr+zkR9qp7HftAAhmVlmFOFsyOR9cIVEfyA/wzLQEaZpw53YcnZ2U7rjdP5RGF
KUGsz0y8bXwXsxK1DdqGDsFuoiSw19z0Ib+G6cskaMJZdfS9asv/tAgtyBI6OYDx
NCX/neIL+VMaX9rfGv3muDdVgfEGbSD9UAgNXeUtSsdPfASCEilAgYCT31bMzy3g
30XrioAf5ZvmO1I84SJoHSCeZ0P4FOjZIUOTgNw17QlVJmRyLynBhlLtBLAvMNAS
H/y2H1YFpRjcVgCiE57TTi19s+vfZMnzMLXPBJIDawzNruXNL8Jq9mpSVQSxOpJC
40UIU5HZmqyoyHOgIoMWNzEaqwDmA/CzfAzkgeGlXTVhm4cxsNXaorZJkXZj3aNS
swVcw9EpHM7nTAb/spLHibZnfInQxQJUZrxOby/cFrvvZbgob5wEDm+qyq+rmroP
RDGpnwJu0XORNfduGdjebXrN83ti9UMqN0At12cHHFX4lxgjEZxvaqWhgU1N+Ys2
EKADmHfAF/a0tIXZpJ0OvLMJUARP4BP++ycdpb8n1p7rDTiP3q4MAmCH9JlVR2yr
+R7tANXV+EK+ST6g4KsISJdsF2yNqvuIHVdeTLzmVj8H8m2DQmIhKRS0kv8I9ppj
/5J08L8QH35xmEY/1iiaRMRhjBvtfCkrnEkSvXSLPp90/RmCsN6WRVIojUX3olEd
fC2/XRn5j5NQWUBhilAK21XhymZVwW5bYftH6rAf8J6m0lYF16mIM9pILRQbvpXt
rbacp7sFedOuvM9tiQMxSHbs8+7NULrjKV06knH+9JX/mR2twrvS3fzZ3gLR+JY8
aMSRmwLKfqPlVEA8tDAXpdgLTpSg1f/jCYBmnEywcwoT82eHzqtMIRE2H448EVtV
j8PnDHZp3JFsEzfM5cQOhTR4sS1OcwjZSljCQ78rGxjF2gGtj5ASQCgNzkRmil6y
oVXXjXtcpE1EqYd623j5+Uc380JP7+diV2pNpYXeeWRcNBn1cf2ygKG9ow/CC3FS
LotD9n0MZNWWj931Rp7hBNbuMHChswcFjTtC63StNkWg0HewdAzo+4sOR0mVPJg4
sFf2ZHpdrY2c+ptT/Td2VUbMuAb9b7p59p5ZaEiig5/7XqUWuSubf435w49dBmK0
AajNi4PKiml1GzRI14k7uwyS3sFXMe1Q5W4N5+JczGM8WAiN1xqeAdqjycfo7I0g
nl4GzA0zVWYkl/xqZN6r0cReyNc7yUB5/ikvaEhLsX8AlfEZL8KViqnzcBA61yg+
1kMtSvVy4Zf4XSJaVwG51UllwNlbakrhlAKa9+K8+zdPsqcSDDRP8L7S2/2OOctC
KTysvwExzd0EoTx3iVAsNlOGY6mWdAvwplLaunmy4VufTZRP4wTqZLsCsQk2xaKT
CK///KmH1lOe2flKlecG5eslgriyLUxdRI4zMmLyU9/iP6ofE4pZbaqH/2TF0qUb
9RPUdWEzDLxdvSKngSdbLtZzmRY2oeT3eNIj59V+5hF6EemMs/du1XKAwX/yOgQw
fw2lfVKlx6Ly3DiQxiGM8WMpnKf7OFNmuqY1Z+9rnl/ZczgowMyYIxEi3bVmSN80
Kga8l5w3mDJqUl2EI6tPUSr0Y/dCD7HgaUognC9fGTylPeLiS+FpjDdCllx2AMAD
sXobzH5t8kVSymhyUizdnS0KR15FzDvtJEqbP8Tp53Sf0p0XKmfNVMaKbqjAQhJF
R0L4o1wFEzJXXisejG1/IgcWxQj1vA4fnYqC6DQDOsUqWhYfsbaXvl8zUfGwKJd4
gxsfzBZTuS6ZA7WMNoL9751/z54Yi7PaUSt36oIiqjaKxnqeVXvguB4bx23A17X/
4T3GK7bUvVoFBrHTLZmEmbkvnMdCjUYNb7wgHJw/xR0JNugOIbb62iSzozPEt+AL
zJEifT0PmGSMkdn3RpiECT0KjPDCY6uBV+9lZuQNi/8ZSlPJAVR6fxiy4db3s7an
lZJXAAoQyMBdKFQMgmA+zZuvy6YscyARTsRXpTeudyfSx5QxynFWcE2Zatd1gp3Y
GXuBR5+tuPnRV77iUtVKusd5ugJl/UkqWS5eP6THtvE+9OX1eSBFC6e2KKZ+7Iei
W40xu7VDe8+OVIy8cG6NlorCa/QT2gJwJK8oVy8LvHmsN+kBObniObRLvw8WkhRm
HCwJ7KiU5wOADcMN0Du3LagRVFX8U9RsfKF0z8FAwqQQ6G5cmO9/JWHVpXGhD9sc
OiCqlH24iDlbZSwAbgvKhZ6Lhvw3zO1yKI21rwJsGcqXdofy1SZy7VpVBEsI6KFs
QBjst9+1Elx8go4DVpy/y9fRTpa9DR/mcmRcbj2hzrlGPGsjEKWJs+yrURGLcgop
cF4rSKoDkA711NScPg7tlTbY8+4j/0GztaoGcqyP7CHiKZphYJ+o4Hcms5J1YP3z
be6bemrLu58yEJ3tKHVTou4rQEi3Q8dkG+SlM1XK75poTO7zFsKc+8xgIE+cPex5
1SiVd6yTwfl/o3o7m/6UevC+tjb1HSn//qvMQ7SL84YWfdPiWXdSL6w4DVt27bxp
URgddJwECqkydHluPpoy+xtpAMQTsjLFLPTGk12xH11bOZqsS+cyQc7zb4ayF+TG
zTDdmMzOeVsiMXLc5PX940y1iLrWV94FWl/KSfj42xHBu+msXTD7D46IDoV6HR2S
q76vgqBnnCKi41A4NgdW2b+OmrrbT3+FC3E37QG1+IlvJU58ZVe7O42+jrTykT7z
bodYNpXSkTLRgAbjNhyLMKTic/kqJAA9630vPSc4LN8R3ayuWXIW27j1lBqshXxP
svEUdGq5MR6lZvKXiAlqBuQWzD5umVWvb3dla9L/hX+3ETKkrzj36SHrIrN/YJyF
Gb3sty/AsSNMrspUAhmG3gkQqddEC2awkY9uNzr2/iJZpwjPVy1+m1MzkchSrNJY
FdkQq+G6Z9cuZEXFIPBVTcSpsEzV4y/Q92KSB5tS3BHEeaIWe/0E7vb7NcrOYRET
pKtpMEewGJKjuWieFnBUQh3aQHB2NPGQuAY9owmif5VuP2SOtjbEsB3y1WYeFDkx
+VquUYJNX+K3os7wJxVCI+7wEWJbTimT+IcpcRjZNF3XPPtXKeKMLf9hKwnG9s1B
a1nLEGquBlKtyQH/MmM+ETpjnyY+hSXrX8TTuYHwxzJm1zCgQ/OSLxSDWfDVerwb
J0whcDvErhK1LaW0WfIuObXa++oTDkD8cWMVIRYWyxaS63oKgXb1pzL4x3yGVe1e
ECEh2wLojN5TeaV93MDlrWCqVb1QkvWPEi5e8ZBfA7BpTTXeeTPY5QGCeAvvOGcA
8K2e0F0uFClZG/84JFnaELeq3VuyY67+YRioZbYWcGFAlEIORgy7uB+nBa3GOVFA
ul9VS6l5QMm39jyj0UUxdlX2IYrrpaSLLAa2e/QQ7jr1bpEuZmWaD2+ykr9Frjcy
AdRxkkyOiywj1D3TCAV3DhmQ4gFeBnl1M7EWsrjl8ba+FjP8lS5zvC9gJFupGhIE
7ddUQpgMuz68svGL4qEYV2xulXPUS0v9C3xoaIZ0GZO0OoH7KhgM3h5LrnMQrUl0
1GZYunL4a9q8wTkAA0mvUAv4IU35G55Lmj/4g6W89e2/94xeWryh6s/SqBI1MgEx
E4z8bU5fBwN8J42g5NIOuqiym4ZmdKf33sOkeK4IIfIF7vXjoU/Q+cECUE34Qp/X
4XsOsF+uP+9GrvQg75fFFUlWBLiM3AfbWKIrxzF6GXPjQl1mc2sX48pB4xC2bTtV
97ZIsEhLYy2a8kbqO65VkvdCj1YzJ3bFACp7RM3FzM1BPyiftZPL0AnwF3bpTqck
GY6G0aP20XCKYHEM7Tirsk5qzhuIAI6ucPKaum+FNI9WJS1ZXjEi82Q3nQtorfAb
er0HeG4mAndXjRV8wjqkZqSBilaE7wB1brs5f8486aL/UQwjJ0T3lBHUTprZ4lXO
kQLZfExoy/4+GDYgfI/TmdoHoGX/lvc7+sFPw2ZbzMTb9MQk+U86W1Y1jeI5oPPW
Tjm+Yop3mFS0mZGGJqAlxqf6C+u4UIOdRq4TJZm41ZC2QeeS55/gVnMdKlW+fB8Q
rXV6g39RY7rCCDhNc3s9BmNC91IqfiZ9MqvFdsIAGvlKDNN9Myyg4szgzg9v3M6Z
/c7O/qzfPEAgNoP5+dlnprTY/7liNu6/ECYU63HOgoq/dvL9kBU3Qxl2Qm911fLY
lMbPwcVUbBMhHzxw6tH4n/f3Buv2kVvyDtoLGl8SbZ8fOHDNEnIhTtplzENzlesK
twDc90aYancj6d4iNicZDhTMoz+GRfTiQdKWj4JJR4IdNgFS6DHptTyICwKVR8Ws
cGnDxSOvOUts1KuscUHzDIoeU/UrJT5jquU9njhADR6DcaWLJI0Pwc8NNdG22Szd
H5jwLVYHpQWy7nLzoeQTNbOxIi2BBay1OOgAm5KvLxDAuH05IYiRJ7bizEOYgGyF
DuXubLJTbRjm2tv+YpMewe2p4+I/KibtYcaa2kbkGnRivN357Rc8nRe1YNxrqR5r
EtmYH7H9f/tpz1cqT9GorZ8YzEHvfSmdxLZ4zmMRI+EhOV73KPuMerRKc63+g4EE
WKhvR8nzTWD0K8bLfPojDnrsuCxshOY/Bi++I/JUs0Ll3iJvDKuqq81GN9H5yapc
YOTG1udiCafIMUQpN9C4Oqz9tp3VHZAKUJissFOqvNwNWTBrkeyOW8uxQKB94A3K
5NrH1KkQSAJybFKOT99sLIZRTIb4IhKYArDLFx/zrJfynKxwrPUTe4Wd/tYl+cVM
tQlkE6B3h8K0e2RyQNwIXmqbUE1nQ041j9aPP9/NLFiPPUCdbAqbMlYn4Yx7ZGYh
wNqdzY9PrZ20tOJfAjkkxfS7R6s0fPMa1tR3AcF6N+MJII1ugwUv6Hh009TsH/SZ
rcZ9w5fsq1ty3gqJvHudYvADWiOMyHwZZ2f8f2xiaQDS3byI/YPQLcmvnfMt7lfZ
Pgnx6gvFLPG8kgRGJ7hzoiTRlbQ+Iwi5xxtzLMMj3KhzvbWUJ1sqPDzVeSY2uhei
YvS4FLWePud5rEHtJHHdU50ayZzLXBoAFaMyVAG6sPicSrAN043Oc0uwnpZfKYpW
pkrZ1Z+TGmPLxcA1/6CPUCEhmH3BhVSEx0Y+WthAUa4z3XcpMsbuK/39eJAJw0ns
YiFSiam4LmFTQjZxPGzQJRTEPWeWzRo7F5w8uYU82xKw2AFugZIWVlA6ix4cKU0E
mEK4DD9wDCvxfnM4ZzHBBrR8OsQIK/8cctu9s6qHWr0PKwLZRPiRmOkPMaLz6ueD
DfuQ9ZHXytH8eOZjRdnMwi6aJfum6X1j2VvDSQPsmZ5PtBYJ1rzrv6KTJSldKM0D
PQ9ZO3/xlH0+UNYmUdDTLSYYjfvukhGcuDECWhJnSpyiSVoZZVhl90GTM5fjKxvA
oGpexsnn+OB4wCDJKjprBdXUgIOxlIgS/7rH5CdX73YRtQdmmYFXtqS2NglmmLwx
WIRWB+nhEy3abG3eERMruvyLR/WuIWo6v5j0lBwhAO2AomtPxrFwr1MSwcwu0hsJ
85InaA7zSyWgyd2AdNmtuVfrlGfcKOh/QK3mtqylOLojTynp6Iw1cBk9hDtWlHdB
QprDlHVkGl95DzAefsxaq/ZpubJQnC52XALHozp44exMuSGZBHlofF7kqbfN+niX
OJq9+XsRYV0seNrgTBCLpeMGFBnoLhnAbnwhuV99Fu2Bcb56J+TsaRx4U42hMShy
/iO2mEejwCFZ0NwdmroqCGUTeQL6cx1mdh2IxcgDz6eRD+LnqwSQaEcBIZSnrpMz
/ADoaqrUH2Qtpt+dRkZ3JBv8tIgr89grRbPm9NxOG49XyCt6keCjH2PddVvK87dm
pVFSZXBrnSlOBr1WGWuIXd22bWFtUFLOXnVVjyYwy/LpRmoxSmvhqYRkvAhReTUu
PnvD28klZVxjrV3JgGagMuXhUlVxdz8GNMV49v34bSzYyF9KvQVeOONtmxKhUsYZ
R4uij1HKLcOGRcrg/KhzhecIBLuTMtCDaWC0/4BMn75QejhVrawDN05un8B6nKuD
BzNoyGyuQ/+kaWgRRZEy/hFD7JDj2GyKRUc00pxOTwHddati28gjjPUXot+S9NLU
NtGKceZV2WfwJdq9kZOeets2sfE3g4ULkWYgF5EyIPCHrx2lQPM8Ja1Mr2UC5TCw
PAfWd4AvwU8CuHpDNRfwzIqKhz+FK4MBEkpikn99qwbNZ3rAtAKOuuCmOHCqvqEa
fq0YBh5qDSZSzrc2SAlwRJggcqnxIY4bE/65eJyKj9Xkv+nvFCF1evawmIcEkt0U
K3iNDQYNYBXe2pKQ0oXEq1HSGaKYpJ0nlZRqOqJLONAoDdhJenlvc1BlRaW5uK8E
+rZufACEojOEwl6Zl1NWlLihng2PI9POj/RvvFtAoNURf+dqqTjonPfKNG9d+bV+
3MSj5VKqBsyjvn07O70Nfhxml2/behujvbU5WbP6Ug5pOl0mCyCy0pysd1IKzmKo
WmWT3PEVp6mOGV4SqIZjQps+hr0XGyLu8dGb/9re+6PVULPY6iattDe/5L0abK36
w4Vgs/T8wVGl460FqWxje9grU+qjBIObyNAuK9l50M13PLcjCvQ5eOSyJ0U63ZW5
vH9O+6LzGx5qRzmeFDa9ONfFN9Cw0VzxaK5GwjYW0/Yq9EPeAxxJayUOiC+inuQa
4gZkew6EhCHyBnvcpVvTNu5ihveF1cNdrYsO8OWzuhIwQDvSf+y3Q20+lmM74ACR
mZ5mpsn2FL41r+MhmlTSoq7sk9QTurOlbuVQCuEBwCQkWy110k6WhPFaixP4LIp3
ULAFsHB5xzOnoA3I8a6uhHe6HFq0UEEu7xHccwOn6ZqAiQFq49iJC8Qr/a3NLy18
rnJrUm2aQ4tMyWRS8hBsx/Jx/oX5WEwRy29hzchC+2mb4/ORNWiXuKgVBpfgYRkG
3SGwsXOmAl0vPq75N9wK2TPjFvplPTgwHwYZc03Ybb2fx7G8e+m7fHW6o06qkAtp
ETPsTqBZJmESwFeJtF+XBCEXMuHQatrChYi+LBvHoVbC9wYwZfm4qXdBbs6kWMrq
fsBr9Q7j6VXHEaacGEfCiwz97kKNodc8mH1afCP3PPf4Yj5FKAGZuSuVWSbduB3C
j77zXttJ078ABSrQmn/J3svvAxQHBngRa52aQ/ltCD1wTjlQnoEqV3wJ2C/KZkVV
RIm7fXinqxGCs6Gtz+75eGWnMBL6yLMNwqbOGHQM5U+nFppVr3Q5hZH2tg7ft1p1
teDOfYtkcSMEFMEo3l8JmaT2iMX7DpigWWaPYOzMfU2NdE+qIOt1atb8TzpoAye6
w+p3kxAwB3eC4KJT5qna1Fl0KZTRMbmVJkbzwqkiRVA6414VRq0d4xMQ4moq0lJA
F1jKPiseZQIC/uAIkjwvMwZpC6A9cUyqtnm3B8Z1O6EzTsTTsfDLNSc7h0qXNslA
m3GLY03b6z7uxsQ31Be5NQVB2mrSs+tbyYnFcA2DlsQZ6dxvOS1gENYHbvGE4I3v
KumEObQYd43QQJUgN6xm7dPkDGWQYkm5+1BBfbKbLPW5hcngJjRDygVXb+4KIO8o
6uABcp05oNr2v/XnFKSGUmiHzi90eWlOcdPLfYwwOkHMJ0m/yj2riNEs8knl+bF4
9zR2iL69H3MK/5RO9bxfvNaf2ryrwSa+iW/aqs2k1mxSbpfwdqWHGuTYeHrMchLH
iQQTzhc7BJS06exyXDzBMdogdBc0mhvXR0OUdinbNTfJxUcfY/zAsf9XykYP5tdL
wtT4HLGdxb4IwGWsLaI2OUfL6lz0wxzWAPXOM5Zw4OTwhiZmGcVyqahaZqDn+9my
NJNOGxzOIkyPuLM8qcChi2yW+eLFZ9svhZa88Tgvr6FfO0kaJo82LZ79GORX1JS4
VbOxJ6swmPgw/PiMPVHf/gpuVNaApjzdPfti4llEsnEbpyh5moAHFpxR9ipTB4NK
JSFasD7BOw1H0DAN596VeQfu8EEmABrBkCPALxU7Y6RPf22yfLIdvg86gmn53eAD
2bSBb/IRCXDG0qVfLUn9UCZRFBGyZPd3dVtzLYGLFssmnxjLfoM48LKjvPPS8NWW
0Sxd70RlbUPfPV7uJA7+WRnlCMnPEMr8luL2IDIQWICmCpZKij5BM9dX0pNlqjPD
6xo+LxD4P6xn4j7yVReUbAAtDOurSi/k3YzXpIxWldz5slN5vZy1IqWGLeltAomk
CQRAJ4RIb8/ZsNDowZUL6fcglsJ/M2fsLNtP3eEjRE18j6v09rclyG00rQRgv5aU
z7+LLu8FuwFuvO0L7T/eW7gV+LT9jDt86LRySE+q/emh5+0heWxgYACkf+rjTB45
yQ0ruxC3DP9CEFnI8fCR+Z5XQL3U5PpNHC54+g0P8ajQ+OAfE5XCRPW2ORFJ44Ur
1RHCr/rJMN2GQaxd9wjxzgnRYLZ1fiok/OgJKK3xvFWoqdF01eQ6bSN5fSvOHBAY
LuUNd6d8+ErURltkiDV+Q0gyog5zE6L9PZdGjfgu5OV6ZLHucnGJ+Hr9VudsjuIK
As4ozwzmg2erAppn8ZKTZq9Sf3vN5RbnAdK0OLstirlEwqROjuaVr+yO46VIFvU1
kabLkb56zzhiD1Ml61ZK2tpGSQvPiLzEiWcCzVKXTQ03rEqg1BBYe1Dqaz8DaYNF
6LtRfESH8XjqTG2zylw6NReBC9H4PQNPIlmkUc642q8f+HFl44Pw3pOTyiYO6xLW
0fKcEcCt+sqAjwR6A0ROpBn6hcty3a2iDT0g71vzNYK25xcmR4ONeuNj6DTcv6Ym
eMbCflzlqXUbbwgRtD/Ru59WEPDTPv0zb7c6yIORZr9zgoaA8CzjDMANxZfkNz3j
iIqxru242RSTlIG9NI+WOKuvT0QHTj4vCFfU9YLU+q6aTRuqFPP3iFl/nLdqlejQ
wuqewZEDdSwBYV780XvT2su067JlR4XrSx4evq8Flq3ewq+DBnOBmsDq1OU/zw8a
7CZ9ykAq6A62fGfBoxAOXQA7+12pBhbC4mchqVICO2vz+cCMUKYjwHLmTIEAubfn
NZUTXOxt3VQ6YdegvxpfjNADwJYxhaQ4fr/5Rm/KQxpmIRi166guvMnPjxEjq869
5EAKCF6e14q7JaSsxhtoBLzwRsX2VR3GQwqDKf4K8Zv5v56v/AR+gkNKSV89ewZQ
U3um4535a647+xO7t+0TVw9j/reQYIlbzVGcuL5LZXcslB0/yQDJmu14od9ZfAF9
LBjWZygSExC1lPGcHT2VsL7bqxy6tNeWya6g+50NJmNIN/3BumCquR8GiPxAY0qc
DGLMViMtWGZ05cY7jG0Re5XLAcGfK4XFrvSNOjQxkms55/s7mVMKiQ8BlDVYojid
t/S659eB5Q58czPfHD0r2sefanrPndG6TdPwd96BuDEpjqzUQfXwTaflwIugqMq2
B4x6y9z+Qz49Puy5bWQZWWFppeY4w5rLhnOdhzDzZIUmb/yUZupVOJcHWD7L+rUK
N2nFRChsfKHZk2kOp93roQoZcnkFiLSrqr+cmQNuO0BIQ6Z7dDlnmZrZfbW95PCg
LuRVPT8+AAtUESHkIo5s598OBCKYQBgETTzeu4p2sMGcUcvSe8YLviuWjsKxIzMP
wRs54CdrJaOlUOhS5ST39nAsD8QsxsPuJJKLItvOvKQer2S2G5NsDbZLnESBjypi
koMfaW/WY1cgiFeKBksyVCSMkTnNx5038dfZxoY/GdzmGZkoQNQ3dnGJ5cBqaseI
0QgIMRz/aN0IUEZ7euCIz5g/iGFs+/NQ8/nHiVJwUpkQ/pnBrCY4jtR83xogm57o
1aHc8n6p7z2SmmPapLbPQpFo5P3uCuCHEGaiiUtnYYmDTZuzJZl0WutBBqX7AjRQ
OIz0w/Dl7KSAUqEU+Fd/5GevxsDIQuR5Nr0/0S9PmfeBs8hIi/zasBtqUL/u3X3i
VHdxvnzmpY2bpABeiW87FZ1/q6NSRGYkHQ/LocGmuaxIwGLkMNefCfmE1wTlwsGr
B3TWvwex/CV1ouJCLCERRKlMwBE1iIvpp//lzwgjJcdFsiY37rHI7jIm7a+bx7IM
5qUNcgWPFmmR7t5twmenKqf31Fag7qJwRBR9bDRZOYfemFo1/0dzgqbsUt2Y4rtI
U1jFWG6CG4S/w6ArX+xY4F6DzkGIk3zk6sW1j5dmgW7cnGAk3LiHBnkeoxyw75Ro
n0QxifruqJUytAfujNIribgU9VxTw2cfHIdvK8/GRpEMPFGwyxHNW6pvgNa0huez
mvNwMzsJfENBDg9agBOdnEq4VD92LCV2iR99NC4OQycM5+k2QkDUscOaayVp8ip6
b/FMStBrVh6rCT5dkiqnZUDe6T7xpTDphgr+tTUJSECxtUWJKDivoFeJH/RnJOdm
hq1PQhn0h9wp3e6Ut31fkCwkNMgmcYx+QUxtG8IpfM4=
`protect END_PROTECTED