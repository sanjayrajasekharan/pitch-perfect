-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
li92qjkS6nbPuVWK3Dk13wwHHEhrjq26VKrMhU7ftRJR0r/Y31wDL40R+r9OoZZA
41Ta0IJFqclBR5kYm9882tImnwqTS79QQq1f+zvREPGs4QCnCINlmqma9ccwMeBx
AN4t/nAhuMdfexIbLTcF9RFCgfJER508N0nFoivMOt0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 44000)
`protect data_block
cMl9QEGDbEFSSlC0wUb1BeRpZZez1r/e23P58V5g3ccPYI1di+DSC4yQ2LTZ7dVW
m17KbgA08kyt2/yt5rmih79hkAS9R1bcspxOC0kn5Mcg4jyr0HKyslkVYMSS+lcr
dFiPdTfch6PjEVO29Zq0SuxfanDgVzo50mAjXcf0cIX/SUB9cSFTd7VyTEb3+/EL
h+Qp/g7M9ZA6RzZfF3sUB2FduaEe41wqv3Oj/GSiTtibW1BkUnfvHuI0NBs0S8BP
HQetbKBGh5psJFk7P8NezzUceeZBP06V/JGxfXrNtYX8IqOt6ctu8x5FD6d37vN0
JEuI1llwRP4ubsgXs4tKsl+G6yYsfdk5Y8CPgzQGxerrO9zdllcH3sIzU1esHapC
MCygAU26M613mw/5TnsY8UDyPDDQJi8RULnGlyhWZfYa+CzAgVwf2tuxlJDpaCPz
hrstRHXiAdTg3nqTfYU/TOydPGZ7ZDfGDqIktqqZ/hMWglco/4zuD+ckA3SYXM2v
q5T7VyyvM8WcV2m1U40O3oNCXtgbDo2Wyx7wjdduYrqYg1S24qxjbUI9uZzbcDNT
8uhwnT/jOfhmU9MYuy8Ayd+MFIdsHpYPBDeLfxSqxLIJpuzpt92RNmLmZaWdnS4v
ahdLr9ZdEGtkhliW9REF5YQJjbrCTf+j+HIT3n2ruPmSJ7UmZS0B5TTdIIi0IMzI
rYPgpWEFFNdXvg+uC3gFVWXVFGl0VYJflKP/g+j8UJltbRXAodeTE19TiMcHII2S
zgTzyVYBp+0nxL8Ln0eaguxiC9YbDWrdRU9yWwGCEMOXTO0Wmqprj3qv9BisTD5G
Qy6FzhVjsQN7LaixgDELlKtVuYXWkumER3s2zqZOOmcniy6BNIK3w7aWN+ZyE6fD
34S3RVHKWeSoLQbPJl44SexCJX5gjN/NpO+cbMXgb8mpZ/VclXtd8yZqNlAoZZPp
W/NNh7MnP6xRbylw/OE+SpB9t7+nsG3XKG/QyDuoBCAfr9lYKsNRs5H8a/QWSnFf
Y1bbqaNkqY3Rv8eERsYmmgQDFW9Qw6kotjPLiFdtQ3F+JJKbMIIOKcBMiGlsCfI0
3gtgyPzaNNFabq11sMk0vL/XbNCtf25gdCALWctjAWi97QXPAyKYWzd9wQFgqFUJ
YlRlG65mon8aYZ9hQGRwWsvVWaLF06ouWIq4ITQ42tWANJ/m5S2PgZMavl5nsQjj
tNNGwgrrfUd2mtiFMgtO8kLSNmtgm2ZkQdquIKa8ws7w9ONsewDCRs3KD99QTZGe
RGptMJE7o0kPNegiBXVdztSbPmPw02wXg9uqRy7r9oCWFN9VvkkLB46bFj4oYKJg
FmlhF0v/jjmPaDndfoDzuORmPXGeCJyEANMqTlp1nRVES9HdJOEqYGrInNCKmte6
X8ZRLw6CNBcHJgkfn0VlfNrlhMtovFxSqNMPe66cleaIvHaZTTWvBN2kw63aKuRb
CoCMr77KU+YSeneVd5whIExT5wCNfpnWmoEZDRY1HFTY7Z6WEgb5PqP16JUC1kxK
n9qWRnGPpNR8w4DSChnTZoxpqPrQquEfBXpNSa7DIAqhYS08O+a/JZh1tH48TZFq
9YMslHEaz8/hHb4yGotDTGC/NP3ovrF6d87x7h5k2qxXo0zZewxawCFwFzla/RqS
lcBZT2wQr5a5Lbrfj+Vfv+pmf1oZLKarpqF93kil363h+qf90Ydk0oJvZ9FTzapa
YPT1pZPwxY+6YncqaTi7ChGORmeeYbGs3LF6aad3mcPzMhEwhZCmLUcZE8la4hAf
cdd0CenuFTOAzvkn9IrHca2Ha2Kt1+dviwLkcEgr1lfCHYxJYy8afOJobR2captv
4L/CvJDDtTGI8zax51mN3Z/kUhcYo2vdqpCUl8bDOtMPW3NmDTxGfD4jicorzrea
WP64bnHXi+5lf0QwhjsJ3ksa9esoItgY8Wkmy3HDch/gH9B2flRIsoiaTrSdgcu7
ocwydY3MjM8ms1t1q7YnXiUwr/7ZJjLsxVZOxNO7U1f8yaTv3Y23eU7sWOxCXcpJ
l9Lht72simM2EMhR1A76dHK5FoG9HkEwhdim9i73H7xOx+2329lrAOlAVnQyIz5y
UIqrAl5XaI0XVUTb91qTqno0mKm2zbzJq0kWIpwBQeIb4FTuz+0Z//MY4Rs1OMCL
eemMdnsMecrKKOFpRcGKLy0n+BBLS8Ds2Tyr4QrOgvGfpxuLbI317jeZazdqgnnd
7Skv5plJrAIosQ9lJkyUDtm5g1b/BOpsB6UZ3/3G9YMcuK70f4dz3hnXj1vtyDDm
yQljmdw1WC05pPSU+NqCGfviM376gOa+TwgvQGJ75CfOuF3Zok7/viEYm3qx+g/L
SD8FtxzsEKWEnkOE3Og7HTljsxPUMAlLLQe5X4D55hj3JjFEnIYIluRLZSMe0h7p
Y37Fz2gyQj/Uc1+v4x3MZ9MD87XaVsPofIev3HkHgPpQMlqLBl5ZBU8XTs1QY2Qc
noExBJ1Ax8Ro7azW+yoVLN43LocMbaFkDWBLIeQn9yvPOBDKozVxhkHzLcuyrSYT
4Hhr3n/pazJYYNoXxm23Ru6Vh6A8WSaYJiXV8er4djQkDX/29Nrj2CkfJLs0cP+/
KOrNOhou3KHxyTNtz2UfXpxymWpemXkoZ8e4PPM1DtZ75GQVhFSfOlVqtxJCVsMq
NhtEJqiX7Sev5aWj/hrg0B5/51JMWkegM3U+gYc/9e0MCGynFj9ro4hCreUQUKUU
GPWg3x5TWp9OstgJRCQBIpTK3t6wcC6IX5tdN7zfDFQ8b4Byt7pOKxvywPY+RULw
YazGIy72gIsc8td5OCs4IuMotTmfMMpso4WuwpcCU8LPzBC+iRxSanD/sKVfN1aL
bVtYTeK07cHLpTsyS0HVeVsLVZa3r+qubgVcqJMXwjIMnzsAM8VFFY1eLNCYe/Uj
AqjCF2BnFYMGn5hHnCYe7hmIA6PS5/MzgAImENshpVnyWAWQeekd5cVz3Qm0dhuE
+FIrvoBEXtem2tDwo4Ay5WpWQDzOd3TTyzAjG+mqhT6ktRnJgSu2KdZWAjgvQ1I3
YAQYcX/5R7niuWvUcs3RfaiSIc7oPecHTM0ICAMDDZVLj1eTPimGlsV8fEY/Q+7s
qKjBdMD/L5BTsdLTUk8lf2TfBAuW+wm/U0L2OzsE10hoi370wdpOG5jtrtnvM3vx
jlUaT6643gQok4138P6HUZdooAXcoaTrkYn6hgFGTDJ+0umQsMgdwhpNos4lLBkM
3kcRO47ZoGYXFOZ0M5yHJaCRfAYNejjvhwtbmqCC/yGBQEToL3vVTjYeFqRyBd2R
o1FxcN1HxlPeIKNHfEVC5O7VvFRiN/tsWJe99aIuGt0qLCK2xh3/Yz5RCzKIVqW8
xbmpezJt+FcnFZG8w1HeP7Rh5lnblHprwNfMpDgg4TtPmlZkVNRpKQy9zmrA7FNR
pE8hA166ezMBTr/Xp401OAqSQfx8hNNPJbic3mIM4L3fnmkC5ZBYAUL4FacuYa96
xuwKkfYEh2fhWJLtZtXjVOwGURhDA7Uj1DEwXxPPt5PV2Rq3j2UyZDU7vRQN1xg2
AO83vWAVNOCfVhMuK6MQkgZhDQQ/9NuLL0Ps91ZAy58swd0R7XNf+MMfEzIos4+c
clBwm62PsKplZw4vI5ywK1HvSgvuAxEstl0pZorU4j2pnLh4tHQaQjpblVIvzYUS
TnSL7tzJ83aqV5kBRRkVQGJbp/yOedPAePGkBYFS2xH43ffyXqZ695wD2jjQsuZU
OZeIiwLSwGxhucmXm/rDJLJO9MZkPr6aS+TFvFbb9ULK/pSiqyUHEwVY3zQbgmGd
lC6OdQn6Frjl78yhA7n85FGhmZvILPPqSuJE/W/RARRVtYKr7BUuiZv5+P4YxtiZ
8Hd+NF+HUzNYvYnp/Kxpun4kP+C25h3suZpErP7A6JMiOePKo0+Qu+3tlsoqY7Ig
HLzNecjwYgfLvYBBkRVvxRa1Aln3yLlvpwhj4+GFgRW3eL3VxTlzA9Yo6erzu5Uz
7hnd7glZS4059j+U1DPnDQu+OlT8spEoROymJAoUUcmpPoL/cJUDu6WldlCy4YmA
TuR0EpyJmieQHhwPr4vR8TOTKqiqUXP5mXMHdvjrYXg9OlhdXZUbt/a7uHiZDuIQ
D+0QwU55dGjmmNSuXPDZJnduiGJ2VnLZV0enUc3Fl3edxbUvZLXeRbXUePfeEKOx
U8yo+sodyjHEhYeU10ObagoimrxC7YSxpny4UhTBdzGWDeIKqXWWnww96soIArz5
DbNDZK3E3Z2ckli1Nv7I40UsDEPZxmFguvefkPYmKhzRp7HvlTgVARHBroTccW7N
a4esoYxRdJpPeSjDwqCaQSF6NaHDsv//AkRLNKAIBU1t0cnJoY65omFixiXdWBnY
GmiSGY++q9pt9ZE13Z+WejeUnDSUHeniRAaQjj9UIuRDt7Si4eTS8+Ra/I5b+0Qx
goWZCOcWUCivh6bD5i2ZvCluoKn6/b8QoxDA7LwQTUulTIk8VLgRUCA4ztTz1X5p
9s1qBCKpAefF17ZSIYGt791XDJHdOndgi1phxDIkwp/ORx5TXPii9imslC+8KXSR
AX4C7isVkjOhEEtp0kqLApGj0vXNDeHzNRxByxSBW65UAXXgUFmpCGzDUiXi746G
5zFsLlfhznPY4KUlxFSvw+2Gu75pv/Wpq9fuPN6wwfDOhhuZ4BZMW3c4tGmXjzji
fB0EG7riIY3BJxafmMvmr22eYiQmhGT69zkK6SNMlGOgM4rqRiwKRlCRchHHXql3
G3kF8oWhZthlDM8zZM/XgGx2WWYCa1qaF3vC5wuqDyYdTaOsBh2N2aoYrGgr3UUY
0TACN2IPUdgO7AWhZ7oxKieRElSOkY03uTrxhVL3lZXojIr9Gl1PG5SOICPvyV6T
8GXG6zl0isXZ3amOhdcq92FoeI+MfjIRLKU+kOrCsIbD5zuVs9NrU7Jgt5RgEgJY
HR16FwBBv2IYwBQMtrrFNkX8aEdZtcMKg2fVJiFRezYjP929k8SfirqKswcKkKaS
hEb1+RQHSqoxNIOKKS5jTNfK8jmtpj3j128B4rwXo0+N6s759M9mU+CWI8h9Y2B7
CcM/2ddN9iJryvhc/BDuWRlJa1EhFcskLWNCMJSeN8nJ//TEWDaMWHhVK+aspHaJ
zgDrG+xE7gRoNYTx5TjHsxUUz5TohSA8jPFh+Jd4G8/Ie0jmG9jId0B/vQaQRUMt
nkZ9bQbP0tFeH5DVqVUDFZfutmQ5pU4EaxVGPq8rUVItv2qo/WTe1qqIMTaqb7ta
qjsc9lnyGO+Is6Gm8cBv24F/Ng9X8dO30XhSqDTuq+zKPaAovTY4wOltfY2QNBHs
60qSuOkrvEkr2OfYHSrfDB61FVvF3mgsSqYxVkVjlEOJcwt3OBvtdE2H7o6Y9RAK
68zMQ/gKBbO+kXmHWoKFXrDEMyFzdHHjE/6G57WwxC+GYG1JdBsIs5R4onsXKm3s
SVRrSuwQlRIcg1F/yMqPNJEYp27wdW4g6NLwpVUVr+aoje0QdqcOEBd8zOh3RhsF
LVOJtkMEXKHiZnmCDMMGtWY2he85xIyGcrPKuYmFZIX5hUF7MlriUb5rZpIYaSsu
uRuLCDcoxpcMcuxZjaBX7GUNkMQlhL8mzsMqkMGR6p7wH5LLYZP8rTJUyoPbth9d
QTFPrryhCifzJSoQ8dUic26uyBKetTD+LyXLrQ0A0PGzkZwXNEB7mgJBrcbFf92k
jbTA1GpkUF2lnNGQlocztMQ/KI7A9mv86JtbkY4cHfDoT47ebHEXKy24UbO9JmVm
5eNBDXElaqKgJpmn7BeEaZxaqdbILz3iutmPpWzgdJQD2MpAJovZpNSrJgeehskJ
MBBYODXpucqMq9VlAh/9ymXJw2gHHTa/g7V8oP8RelF+NRNP3h+Pg+rIkxyRkrZB
XIF3/bbBhIGin+zv6g5X8V/A+5Yy9i71fnGF24V5OpduA6mT+kIgTv96zm6k0x7Y
TkxnD2cTaW2w43bVpCMZU5E42YsSXqbg9k954YhyLDzEdoPECFJcl4CAXBi2x/W2
UKui5Hws/vLUoJyHmsO5usYEGIz5sQsmKi2YcmLIwjdSTnQMAQypRgtb/mBaa1tc
yZJeZqzWabm88ISdbf3zIkinRi6P4uTRzUDWOWJhPmTuAL1nwtNnmU5e2+sOqrPu
qq5WTwE7Z3ucdg0fqRXJFuIdA6k5y9JLmloBLU5ajQkPKn2ViZtQmuyLOsexL1XK
FXF2ykiwnOy3q73v00uwESH7v7iZz1LeMoL6DDIR+FqhdkId5BDSL1GkOjYWxzkU
5H+39gVbz+VEa3yodUElUjcyBs2zdy4tlUYPKKRBcdR6cl/2Tcu8F8P5I/997HEX
ypw4xMsKpNsQdvS4ITxX+qQ07t4k9xPr5QSR0kQn5kddTVqS6bUCUHxJuWGp/mq0
oRyuegrHbD/AOhuSuyCARMU+pLZ/KDcZ2Tp04XefSL5qko1TKoR7rdEWC+AXkjWB
gMNvKOFKHMTQhaUa/+JBWpVYfM2flgEWdoXQ3SsONkj/odNHBZG7jVd8SRoY7ppa
9wX5XS+FcVlLHt3oDmdtD0hi2W3yJCGDWwHhxmBSk6eDbgQeY4ZcNJJJr/iVcINR
4RoJuGFt80ZVCMzrZULGYmuDIXUfLrFSJk+oCrZCdCSQVbV+zxGTMZMPb6bNRxxN
ux1Vu3rwfYifYFi7JHKCtG4YDrCbQN8cSV+2blipwBGVfXNXqNRTZMZkHGm+aO2X
KrM0D2zNAHWvfSQEqRhNXzmiV/uBgflZFKDAf/Xo5zOI2jCeodN33odN80M8Gono
1f9hN16nPuSVmlUyevz1+twb5tzbZQ/NYBGFS7pIA9yOPx8z+gUuBYkF64srhPI0
HlBQCuLJyykYEgEiRKDQvMwLONjUSeA9bf9QGQ9N3eJzM6zWUdG3pMz4p3d403JB
eF8evcpQS1StP+8vxWcxyg5pl6+bqZPMPqUDsq8zfjK3MeHKl3k3WfdpcLZ0HI6c
z5bOeWMfR7frk17RSdM3XqTObDWM5R1GCDHPQ16aiPVHsoF7BIZD/ZaHckx82KTf
yftXVJ/OQRepXTFGR2cD0kkv57mpFj0/7WH2TTNeE/I2ZtrX2AyeNn6IvTtpK479
o+QIbXMhb0WUSQ0u6m4fAoFoPtprgxrmokrXouKCEIFSBmE7koqmaxuBwSrRhiZ7
PMZehVAZ4Xy82+UFfGzQdS5iW3Sdq868UFSXjENCwfarfCdmGs/H1js49Cr4Wjog
15cBpf0t4hTSpbjV5CTl9PZdkbeJEFD8+RzxmVtTmcogVTACmHiw88HL/rsYOmW6
F3CnPzTF4exkl9f3+WvL1CEFv2o/oLbgPM4Mdth4uE9pj9dunDKopmiWJHryh9E/
y2Eg2+QdRtsiDCuhKs0nCIObRaMFcnQiGoPi5QqjQB8X1CXJO1ShK/U9W5XNYv8v
iSB+/SlPklEwRjEn1xCzwgj2mdYTCjTv4wzIVu+MRT1cdd/gGsYZwvPkrVogSyFn
pszKjHUwWha7U8y8S23r0CiZDwY8V7Pl0l0XUVENV0RaOYiFsCWOAkI2gpjspq2w
eRP8ZuOUjUrPgda+NV8xI3y2g7f67DCO35UhpXSaCGo5Sxe2wvJX98a21NA7vqyE
KzkYFlvpAETr5fGhiCqphCdDuHq0faeXmOKfmf5g6C9NJHbv0ikQBg8BhwsMgvXe
rwZXdKJQeaDvq+FcCtRfm8F5gqkIQauDEZG+2GFn4ervg74qLoC5CCF4BOjt+kQp
dCn8eijtB91zTZ4Qs6WvFfN6GRe4KLPkNWUa7Clfxl7iu5GjwFu1F+HULFYlitXP
apjEUjQgim3/zC6xd1NvgB5FU4PyyOE9WPirv0nP3lKmo9Z2KvLANo4AqTc07LWP
QMv4TRT+xprbgohd7payuSKHFRyWVMIksIsrbH/FcloaAQMoQlwSXc+T7xrL1Vgx
Aq34sQIdLKfiPbCdDvJgQa0R2GWtSG+4qSdH7mDiL3v82C7J/y9nluO6ZhLSElT6
zEEiWNfT+B0KY8jtXQcwBzBL+Rya1UAM9BSxYFWx8ZDTXGkuKqt5NnTVBChyr+RM
VW6xm5jIxiEPmcPmeo7hl7mJsRq7PIIgTiOTwR/Jxt7DtsK0YtYuEwtZ2+kvn2ZQ
tlCx4yam+esNU5P+hixV4T1subwjJkd61DR7SiyO1jKHB0xQHFrJGsSzpGbB6GUC
0NWbO8n12u7hINCaZ1YhMnbkJujzyLRnqHbl9FjTdW3aN7vYyNVPTDzoT5UuUbwr
Kx4euIdg3FuGI39ds09GtTzTKVKGSTgFSQpMZ7u2Tyk7Mvjqi2OBiIbKG7GF7E4x
50p4f64ojqJK6hVqn3rSQ3aaHGMWXGP/X/SOiEaDAWyhYNRWI7VC3peTj1WKla5n
incCiNWcMHXDB7a2e0HdJIK1FitHNeI+vn3BhluBgyjA3Uy1+VYPAbZ8PqrPR/Na
QhmQ1sJr1ARliPpp3n2B+6rREGZzrURdwzu1k/zvfbtRrmKxpUswHAFqAEJL5Zu/
LPWyvwNMNYNADvl9BCf7dqhpkD7rd+8JgAhkWT9YMDtOEInD5fP173vYKryc0SF7
sIM1pvhXoMqmNyn8lor8UtM5A3WSoSoVOInfInnkuLd0fo81unmTFEtf1SWnxx0A
3b/Dga8G/PGpVScNK9meFm/vxftAiMlg/LyC0juXv+hgyJER1gNI/V1iTN3qmKkc
89+3QkY+fjh11R401aeDajuLmX5/5Fhf8F8gCs1eelNXc2hF9UmSOY3MQzrRFB4y
MmqjbvEb054dHOupubwp7z4qS1joZuhBsxZ3oKO+vY4avX9p3G5Ods5Qn0ibjwj+
ilpJA5ogvy011fK3P1akwnVN7kHttkQiVm8sCJCZ7DHdcgpD1FB17JoZYTomEdHA
J+/baBOsWB+aCtjQA4tJaUDKtbrM+B2UJdSo/Lt6SXFqsYUuqp5WTJxIOWx+C2kF
w2xXWLBV3SXsrb62OmsyErEBz3VQJmmolK9f6xI+W16dtyqR3UjAaPC4OiiB+I3m
Nn4AAJbOLf1EV442QZi1oqsdDacAV1uk0Yjh4jjNNS/Fa7dKBIIbqFLcevNxkfNY
H7LmINDA9WSUzCqSXtCfA0BfijDojM/l4JA4S6zjOeJ4ihcQW6Im212+bX93V9Jb
eApXcCsnTbCBAHxvW5FYSLDkgoF3++FY9Fjc0S2uww5aUQzefDE2AceC7SeSAqxi
BoX/lMro9wUS5fQrwCtn9b6NF//B0qdNg98iOIDviobn5I3NFBJGDRHQ1svDi0is
RwzL8GAHT/Wdo2QmbofEDXJX18ehdMMJm6+YBawvk3eBIucKihpCpvZMx5Rfn4oo
9u51Q08HRgZ3YrY29/pybJO+PBz/Hru8PQsffkLmL7K/WYbPWzNhk5g1OSS+BEie
tcuc5+yjlRIHy45K60AWGESxO9H60ZcpdBmltMgJqIWz0ZdAKSN441NiwzOVxc9A
BFCokJN+pYAXp6XZiNKKK0MWlqnpU6nXgR5Yf+bW3yYSvGIdR7FxLgNrnFsK1IE+
76mWqDRS2VsNkOSN58UwMB5hcjBC590GYX8G33RlqvmsHMZsHslFj8h7Ir1On3me
sT01yFztnJ8D/HtSeFyTEXMT4IlcnYnhKWA2UQsBLsMPGdHogsJTtlHCc6UdCA0D
vbGas6VpwHp0NZcdksSlCcZWP7NMPhxq5lMCJGb6BPxSOrAwSSdOyhmCLnrmtLZf
ktafIoENDpTz98REnCuFWFmfRSwlOVyVM0XOSvkBm8cCl6ncd3sVxCxQtiTbZgRn
AvgUGLX7nZrDR4/Fygy+o76G8vMJO4g72bW6JHz3B+rVUqgUHyYPfhOUs0+ciqfv
YQbk+tgj0X6vLIyt+Bp8Bn/RlRZwu4Lj1uK33rPu0NCBGiHXc8ZdmFiLc1+z0FTs
h2NQ/+N2+3ZC4K6bskgzJLSKtCFC+hXeG5hycNYi6X6KI3Miv4kzSQanOYv3VDyQ
3e7A+at++WzbAvbNyqJzgEJMCCjURZ3S3X3MX0GqqUxcv9C3jAdszmCD86lRYTcO
ZE0ZSwB9nlQeIay9S7CBmym0tCUYqcCyDwICTJRALkRQdx9P43cNROFqW/LymSaQ
OaJXHpfWivrLtNclCZK4NRiVbG3awH3vl/5cjaJNTwRhwuXBEIGMtvVHNwo4V+MG
VbjxkaqIsyh7tmFHFuhPrffs6ZJmUD5Z/cxipLNECOl7/pJHdA0tHkdgnmbK5tgs
oMakrHCBjFWzbYvQ+/lcCqCDaTdktnheUs+tblFxTjMXimpN2Zi6QTsSyf/w5uJl
AcnNLpV/D2byfFwd8I9qH0QBUNpfaQxZlZaVKpuu92keMxx8biPaM3Oq7fT04GyH
y1BVjWxXrYxzvoBRcc69zVHJV1MS2w/grP4i48wzpagTtFz91PxXVqvbAd8mtNae
sJRczjbH+RiOU65zxd7x9+BIx54S/phGeSBTCwwV1VOOW5+FnQShIselnocrWvMT
dGArp44FSOJhMoBqqbc8XnS17bC/Eqask6AHgDNE9j9zr6pBJhPghOJnLnfoLfTq
RP9AS20I+Zs+ROhpxpIw7YnGq6El0GrrHZnmvb7Gc7SW3IMm5o52G7qek8MP3qXd
1ZKZsUxwAyWu51L9mDue3VpFfVbj4HnngGo75s14SdTTZevV9HilAM2+mVa5gqpC
tq9Bbhp8LwQ7zfHXjz/9hLafKsIi83UdsZ+EOdALbpyXm7raA0mN5loMwg3a+Mxd
mvpYxGQ5+xnX98G7BGOjtA2AxxX41Eqp7m0oJjZEMBIzif36QSPl3MM/Ul0WKtYE
EftAvLb5qoiylWFs1HexmWQNwq0Ey+nsNxgjLpXlGTO+yefnNRMS7zsQCGEaGOam
55sMoFSH6LR5stRSbiTl3oWkmlk9Zla67yTlswEnBv2bpmjSOFDycnfRTCmLP4Iz
mbpK6h4CAjb1wE6CPiqZunLjmiYjDkP930EqJwGuTgRKr4qV7Jj06d4ia7ZPvldi
KiOYAagI+1OUsexeTqpQ6R8K0VarKxQtmk3q6iSH1RFAIhppJpSBaIgR4tIgEdmi
m7kEJZtit/ZLqvxHpoQ5ca5uLjFWZdDnyBEVtJVDA6H7n336nyjE3SRT9mMKSM9t
48fCOu/1uk4nKdkkVXiauwblwXQe9gg3em4TzA3B1Y4IA2eknV31Cc2eqZFmo/D6
QlQJbHH/qODlov8J7Cn7gBgJty7y93kNZSOXsOi1CfNAe/hlMIWQE15iiXVRqtXU
ueVpwZHDk8K97A6WUkzXXgT8EVXJvUxrlrf7VhV/gv4FwS/cTyZKmLMHcCeiPiUc
qMU0sO+X6gGV4T9ii2GGapVMcd+mbndHHGrF/4pn59NyAX/1sSuDjUqHp0pVUOG4
QnqSVXDwB6QywAg5psikImcSlXvHzXSL7N+rata/vtQqcwjbyYmoQOSItceT+RT+
nUFSOD1t6NPsz2HmBG/TCPpQtPunmpyANy4rUontNpYD662fDvX/G0nH5HbdAyPx
tArXzKjmFFnLX91pADkTmnnAe97ezGcdSiVe+ajreg03WwJ5Ejr8IzDfChTVy0ip
zM26SLTlmblUS2knCCfvAY6muK8CFm44iYGPreHgGhyZ2GVZeLGbi980Pvj0b1mh
rHmPOxHa9kS/IwCABO7qWc4nQpi3lvnLSDIfWOYDAQPkQN9fyF5cTzzaf3NDoi1k
Z/mkKKWs2ib1ux4qKUZYgguQjaqYKyWqE17w1YhPNSGU5ne39tKA7/EVES4nl6D4
c+6RGsZGQpIxRIcuRemC7WsPf+3V5CuDeKJAzCr6LT/Y9RoKJVrfLEx3dJFNFDez
bHPOqMBhvjRSVErQ4GrxDkW8EYfKuuOKrYKsukefXAEr3K/ONjjHLoLYybnL9n0L
hxPKthB/7VwjLMZPP7vDfIDnmBgKzFdnVBKf+aVEVmhZlffOtOc7hIq632b5+fBH
YmHf62mW63DrpaFnw1dBYWhZg6A8ifZ+6F5OO3MfMdBJpALZj1dqhVUWKMsC007t
84uKg4KWd2YzAi2MJnFSdfdr0ETbEePUloWiDYZAXQWIblJQksqfWb7BjkiVJz+1
N+sw/tl5fcJAOO4p5oloAzk38wfkBP68fA7VOWaibK+uF2Uj8m4M8B/So6nLmCRp
NdCmgs/hwCKrD1+GHVXTTzO7row3uy8fKy/4IPYqBA1sQhs6AAdHxSXpcbLrrM/8
ZXoGWQw5gWkaoEPYIeL+/ihFSCKKbCidHWXGAugqVMiiNHc3UXJ1n515sbB5h5jD
1VxUMFrMJVyw5RigVr/q3KyJoSTxB/UVHp7rqCStcDB1M/4pEgIy+WBRmfcasq7H
94Kirj0M3DzDFe9f3n0RSv7t3aInW3RtqrgP/WDAN5rDRrI0L0WobT6I3dfewKOs
SpZcfC5qLwzTfyBhld0rlbtU28tqEPIjLRDRwJWbD1KYuPnMTJ6ruyKNKV3Lrs9v
9yLfqRIgqI6Pqn2DcPL9HLHNybtU81GbNFjvy3z2IqLjgyfajJBc2L/oG2bg8LGN
cNrANxjPq+r9SCOCU6SHHZlm/ykDajdhGDAwhN9c0v4/x6VV8VMwZjZt7ATLdCQI
gGcv/i02a4ZomkEhQSdhl7Crku5A5F2YRmiwg0k7/rySluK2qnpTwczl1Mo4SOuI
eLJThvpGkbzw01QUnyUjwVqhFjWR0ed9taPMIogzQJPxZFjLs286V8SytStiq3hA
bz12gSo8vCu6q26DNmvoz5c6p65oHpYbzxzeFlZ/dEV8ribADH/6R//ndBQ1qwtA
/2rdC+v3fOE/yNHdxAmj9bepKqlzpGbWYeveQ62h9auk3aWPqMrRCzfHX5XsJqgX
u0UYgu0+iHds4OGJ7URYff9t2O0h110GvSaIhniEZRurvwpDEaFqFfLxlm/Hu8Vk
D/iiymWtXkfKlkzvZmCcmdFNndsmXT05mMo7RJtNb9vdBMks7QQZOTjaqHh2WZBr
zlld8IB9bCmiLiKmWoa33lUJks4dSY3N4hn6B3faKMFlDPwnrzP3QNcxoXX/nPhw
Vk+01vhG/BZ21oDtfbnwA83nWKWszhh6dBIkRAYR882y84vGgJUpwESRobuJ/reZ
izXqZSXzQoMUXymLaA5W/w5Vt6SwRxAZkHmbYxUyJgsS14fqMGk7QoCQUO8+5+HA
li0vBQqRyBAwRlwb9HHmfei+wbPRl8BiDz4DgUlSSMqaEykH3sUkEDjbV+TeqlKr
JgD9DymroQzYs0+sI17JJlP87aGugxeuJMK5fd61aLs+A/QJkOXuv73ZPLzIswIZ
KZRqvZqT5p/RUrnHdk3jgf3qXmn7cng58wgfUMSJ4KRvj4xbFP/1nfUB6BSEv8oz
EqD3fRWOHAi/3EhthOPifLsUfHyLYFNPwOeVgPyv1WqS7EDzrT9fSkm4GDui8mjA
iyiAZBXSyILFGrlM0vbxe3PK92JhHSwlYDL7B4m4Z3LOXFfbenn//LGzDIasyj6s
NkW/+iJq4mYm0/4Wm0zrKihftWthGPgkI2FcOn8uzs09Po2dwPQ5k1OP7tipT4n4
9/OqwCCRbt/Qx0f0GWvZaGO7el4gf8+VLRQMGr/UDP+Qs3VAvroNjbpdGmODX03+
b6w5avMPiRdNUdtV+6VRH/k/YRCwiWGWeqaAQEaqMLu1x7aZQc0Ag6LtR2zKnmce
7gqCMa6Ng/apws3spiZO/YBeyO27QKq8nsJjzW1cRIJs+uJkVz9Z0v2QwvMDrFh9
fPgjUQks3vHtg4+PsIRkEo3yIWDE5IpIAwpkCrNFizjIPtD1DodiRgsVRcPqSOis
UkPm9OPjODTx/3G/mnjrMYp9Wu3Nkwme+NQwlITRuCH2aDYYyrLa18lkUpCm7C8A
E/LXzjAY653qaqvRrfZT5CHLLOi/1oPQAzUJps8oDuWrsIVZsJfl90/5eAbx9w6i
SltXDMRdy7+aaaWJTVToRklNWJ/LGQl+Ycvag6OlFbjP6IGeocITI8rNtYEHgDYI
CZyhK7LJfYuHm76dkuEWKimDUozHPBw8cX/4jde81/GpaUDnP8Vi3DOWS9j+wiqw
tZaVA7WH8j3ZG/ZicJHKhBUnKWn2TBGEXEeEj5d8UVWtfddsmDp6FNdY+XcumAEm
6EALV3LYuthb7zrNiql6qB5XX08RqkcTAJJRoCNgi1sp0CEKYz8x2RxNqdq7xUEx
J6wjexxycds/iZuP7w9RVMjbDV+g57tTLMaqK/KuW9rJu8dOYMGOoIK1OsFDhtK5
gqSRqtcqWq+tm+Bt53+o794Z+sMz4gHRcNWRqqwqUKHqdzXIwhR6Y/KLWZjhVwst
86zEgCBUvSv/3cD2+akMDGy+J4E0mgxf/UsogUE85ve3kpJHgdKZz+na5ry9LUGG
avBxnSXE/H8XzE6Gi+S6iRqE0kfhnJoI0BKtZJC7WLm2qtYYaldE19vF0O984SAB
/vrHBAiAHez3DYwX7EaMYnZylqVH4qYsYY83UL4Y9wqkDuZ//vdahd6TBomymfuC
XDo9iot+mv7E2wVOg+t8LxYQIDd236XxT8YHKGCsMYe2ykRB2n/kK14r+8WBc4ZM
3PgED0GnkJQq61c6WQf6Q1RSSukvyxoTsZK4pad5ocsHOOEP1U3waElsqqQSFT24
T9N3WT4MAjQ+rnzfsaTvbJ7/yBkp8FWqI5sbBcF8QWmJrVDRRgSmJm8o5ojBsm0/
thPSJIAwU1RMfj0RHU33IB8nhd6MxQh75UXELwo6vAeVK9OMX7FPWpJW+9XWBZ0z
QIbCCA9WP7+bQUby2Yt4utJE5+LXp3XhdX0AaHipVc2Z0GnGzMmGikriN7HbBAgg
Kt4JTEyd7ejj9Xm4FLxUhnRm1xkJHYhmT8c/zgtn7V6gV/LO6sv+m2ABeBxtxqC9
9TepwKjVJFXJVBCo9nmAZtU3uXg8k5uI3oBtSSFBRL5GKWkWi9sykhdbAUebqU4Y
NhtJGpcR7zoZ1hjW3GavTOuPMFUH/MeevGc6R2IQf9XA6LPhkdsi4RTqoGRPhUOH
7mdvkDUUsN9+1TQJN1msnLphD7Djca0YRrrGSF3oLBPVTTcZPjm1MYXQA8uTkA3V
gLQuGp0mmYX2WCWAPhGzOdEojJG1/2khzmvTzLHhBu8nQcHE2awmJmJzf9LdbpNi
ZEUslfaAGtEaKN/FY2TLvT2F+kVSQIMs8JmhwN74dqE6W3h3iqcMsOcmPVlDhDac
C/dAd0MnZOhWyxIXAddYuojL6d/LP2W4If/adCyo8QdgqupH+hM/xkK/c8MJ6cz1
hJH4KH6oom7LuFuN1ZcJMm8q4wHskuupObnOJJLFKQ5Q+cIUxjaj9fBPPajwjtWf
3BzcD3LAVhtJkVwjPKT/2I5xzXSvKe0g+hcPszih+GPmuut28DsEbAvtldyDmC1k
4HD8Mn7xeBT38Y2QhxuTSSUkTOBD67Bos0OXbg7+Of8vUSSqdzb9SdAhPxIkbbTa
QaUzTs8ixYWruJKB70Dv1E8gEmbY34DzQdL5nIy6fTTC0r8SDm8lxMGR/r9m0Ykn
tAtUIBFUfZ/fEtAnYy9cDqBDm6Vj3sjTg9d3QJA3UUrqRPnV6tTUFQV08zsqdXF4
x4K9ckKaIuXmuTeiFQgpk0DlDEVVI6tHkTXuPg52vyRKkkcBkvI53rejcsGYXaX3
BIs4s0DXX7L3p80TyBEQsRza1q8idaz7GdOJzJcOF4yLsec4AMGE38Ai95PrLT2V
Zcr7dNBNRYCvFj1olh8RoLfuh1LVlwokocby2GFHjHkhQeY6N2HPh5Rn2qH8AxQq
5Xa/GIk2iUhmd3Vp+aDlwjiW1DeR6xwevZh7ZFdhREJ1jK7TSo+yGRtyKNXKGfZY
gzLAHnX587DSdhyZEGo9nOqtSOZrYPvJwZgnBfefMlKcJjCiVzpu9Boja1Q54KZH
AkCqzFdD5kQLdV8UTv9EolR8tU/3O8/iDrj61qq9rlZVKWNvrp6V0A7qjN9yUBRu
Ti7yy9NQRgG54b/l9hvxo2bN5PodRG6fehSQJ+kh3rC5sSlE9bGne8nunDETKAA5
Mb9ufoJjsmm8SzH/MXHV42SGnxgUhvGpPDb6cBoUfV2QYXkFa/E5FCJ7FjRbe8Dn
EKwgqjLH+jVl8mIhEKQHxcD2uA2DCDltMeCAojFvIxGVV4GZ2ZLJ/F6m1VJ9y9cB
0fvjMnkNuEyW8Q11O27azW5ZWX8qz4ivUosoULRTi1WW4FS1Il8yibtCVTi/Gy3/
3NC2fn1YwM4NlCwKn6g3r55doEg9+/vxPcHyXYK7N2Ll3fziWEgf8Mc7IH6WPfYH
L47zFN+WOfAJ4VtMnuMudLfR650G7h/yz27wCCaofOm9MpEZbrIBiE9IP4qfwkF3
QiUtWelSarDL4LBd9areW3QGG3w+hZ/A2FTSa/XQKYPGTx+AQ95o48oCVua1ipFT
K90tXvbOtPVt9d/HPMgpV2qPLr26pHS35MDG3lxRqxSsNF06CSNAeoSggTFvOz8w
6TFQlJ3r/gcedY//vaJhfd/VTpoYRo/XGQy98EhVwO9EhofkASAQZB9Kx4TP/WHJ
sJkTLEf0yEvTZiyswy+VioIKe/qsYd41VmYbaTGCvEE6hqZWhgw3iuQVxh+h/69+
0GIrvB+YxJHCGjkjI7VQ1oyVS7W27TucjH2LwCwBmtqFmy/41HNKoqxH+fzdIjFY
Gkl8pL6mVF5+i482ZnW7ZbhkKTwEoU+EWOE7X1ghUbxOnEvqPMPdxy1UZkXuE7cd
KjACQg9bB5w24w3vO2gLVfr/rLZg9HM8oG6oa/3sCAeuSgmMrmnFW3TalbCBNU/M
ZxI1nLC+0NEOFSYnFN2K+Zci+Fl+GfwF0A8quTQLDBJf542KFh/wz5/1UdAUIuTX
OoXOpIhOSCfKrI/13LZeBFXcannjC+scBDEL9OtQi7w4xbDcAoQYEQuCbnlr79c1
36ypdVKV6U15Iml/Ngyd+Dk6pjXKzgKvr1KEI5vxlaE/16GaPF6tZ9JUr+6681uD
H451rEoxPCuOUOdKvsjf3Gd6hFh5ojEureLHz+NTpK7W91BrWgCeQNOdI/pp4OZz
Q7SLVC1j2bZNWBVoGzhbadjPCYf+nXiCCEqMqovdTwzdeRS7oIWeW2GOGcISDUsF
tKJ+dkiYOjqC/hOzmSS0Ag8tuwiBtVBrkipF7uX3GZMFJ+aR/j4bOyfLfubaPLHd
nd6TwjNYAreLpSCqpLcsuj0GGr713CM/Wp/6ggdA/zI4yXVbkptvbGDxPzJg/wFX
flPaI+sKLbQQOEwu9jFhqv9PVdqqSu+qPsAnDXySa94K46u8mTLf9BVvlZCjtLzA
7Dcnn64ZKW1O2JQU/3a4DQeMYSCzMHX/OjYXD53hCm65wpRRBj08tAvYcf6llZPt
xnnkTYe41SOeHmV5Uej3aX2d4XhlmIOEjiqjZAS2x23Mpw3o2VniCBOernvhuS3K
1mLQdu7FhWvuujD8ZjUYu8bRohOB56yHwvcERyNMYwfrzG3vcnacFA327HCM2CYV
oaiPmjXtwIXR1uVyWyBBIc+pE2jRTVhnPQowcU8KEA6WPh7HK6BdPu96+5ELzDCP
wHVjbDXIWkgwa0gtbx4A2MPhDa5IvUaL5nvZvHs268WR8MfnhqPNGTQ1pcJHekdm
AZ5gV3RACGPla5W3pD364SY0Aj2dn6WGKLkdsPN1nygdGHiK2OAr/z9ICbY8loLx
Qzs2/2Yw5EPPbAQ/vOs3b/6SQxXSe7bZHnskFcMkqqWFFcUboo0HXFRsMOitb/qE
RcMNnoWroukIPkUk3jib7Qv1zY4QQGY2HhaHgzVMKmgKXHu0vWtpxnvMy2gDlXhd
gRhh51mC1TEb1kCoPCwTLTRJF3B+6g/XkIfXzY3sJC8b8hSugC13iC3zrFl1ewhB
yYReAO8vZPhgbf4s0JFLJQHBzA0gTd2E/hTeu1V+UUp0yFRffZDjIpaHFDoBqoQi
Tu6Y5/OkTZVE1RupAzaOSZUff9+ClD3iHDK2hdp80AIjg4B43NWFFUcC37V47dNS
MALSqX2w2g6pvgw366UXDneZlw8+/CmXurHjjeEnRMha92KQmChy67IWxIYCsgum
l6SHo19CfXk67+6CFJEij7mjDpelDOQDFPuy+7CpFybe1j7lcGIo7iTCVQGETcTu
ljDYJEuwZxEVF+OXel4mzUZ6xbQpRYQdXpSg+zKJ52U+RWJRLNLYV0jEN6fk/2TD
8oIln3gZ4Ogvboj/0cOOg5MOfT/5UXpsUZjm0JypY/2RlskVYwq94un0Rv4w1l9j
62PsbVKj64gb23WbUoZFuqw5dz6DsHMnWvJAMNpW22JE+462MOFqFVEduhp2sukg
tyo3GlUjLSasZQsH8New0ZpVJhviJLXMhCPV+FUtms/INbxeWjRz47RAgixuvHrS
g+xOgwPYemjuMSq+dwXIzduQKlx5t/+HolYHicxbItJRTNn2FCg3yZpm0XPInhCt
bD1ybiNBGQRyZ+xjIRxJE8NIQMG7wcuedfsnvjlQ0lNPyAqIVK1Iw5XoWYbVo/AX
ki47U1SaWKjgYU/nijKJXkS528nxowIVBoMEcXsiGA4hjh6ZYuUsm6mj8RWiKCNp
Rdu7nFrfPHrRDnOdnclCun2g8LfbmSlq0ulkf44dw26uxbHGvgthQX9GYaOY7I2V
oSxvni7oFX/cOrc1W8auPY7d96P8LP8WczAIo4HAdTNzxIWWMLcrD6Bp4aE2zTQk
MPjwVegmcTkwTosH6D4BO7P6ivW7OgFIXD0F/jq+2k6zZZg3TtwYF4JjExG5xh0r
Fz7I5RWnLj6g7bX5Xcye+sMnn8L0XgN/fm3XH9HrMPK6y7nno/XVPnbrP3HmK3Ql
1Ig7rNY8+nPV8u/vnVCmWVLe1pb2E94LSYY4/8t+EtMNqFs6+XcLduGM/Ngapmoq
i5zA+omr0jGvHiM+83U3/Mgqgkas5oXFrYfvfKi/PeSfyMWbWVM7Tgh/CeQ4Kbb4
FjLC+VFUZTZ8pskA7HX6Gp2zSAnytOIoixuqKNo4K90f7y76VCfw9Wih80kaPiiE
LcgJM3Rm9BBRxkt9ZVu2YBLJcKim7ckbogdcFoOx9K+/waAcoTTFamon/AXDOwCo
9yUcXe44BJGLojzqo9TUBo5DmKUJQzJmEqsafLKqjjFamx8mmPaKxyuOP1wQ4gqQ
sWO+Ag/96BFjnKnAOXCSumUEoYjM7e388W91VwSfK2IdSjLVftjzzKetCF931HNB
ik5YV6MDqTQNKDi2r54q2VG/SUL0qRKGcSMP4FbFPy+AsQ+RnacepQZ6REWAHSBq
oym8Hd6tT9GYnjsF2tIGClBrTnYmVBd9nmXE4vwQSUDGRi+hl0Z2ZjNXCSg60n+4
b31PFPjKylLpGxJWQBJzSB321DeBK/IwAjLdi1hrid1g44ZjlB/2Jixiy3z/VhVZ
UYZR5Yeu6+yhiDcAcPZiwMFRNcVr31jFShDWXLtm6iq1NIHGpN5mCGjihC2oC8Ja
T/mjGp61+ZGvtxt3UI/9qSLnDMxgpPvk7oCm9IRzzo/s6s3Om6NZi0qRSiFm/oBK
b5uOaOTOEQXcbIsjovFG+P+Z6y+xBg/W9wgxSsTIpF0bHfk6VX/Wx1m9PriyRF0b
0KCSAl3cGlwp/lnn9MVnlRcTkjmy3vnM0/5eN4mbhtzqW8eNbk30ff5+TQm69F+3
8dBCgEUmWcwZ7zMGKODrfniMfCeX4OkZJr925J9Gd08+3VKBZ4AzfWiwdMMnb1hB
U+durCPL+JQK6rEfkQOZvG0V2Wz9zC6pcFl0kaaiLj2tlklpSisvRs1pfVLyQ0CN
1weAUs2kwkBLkodMwuVGLgSfODxrv9FXFHQF/08dk9aMusG2Y69aK9Xs0pUb40oY
j38CW01AwrM5EMF3pEqDXXCLCJra/nfMaPwQLCWwsb7i0WtsujwomZWFPNj8O7mq
aKkKFwyIKyL2tWjGOHSP+djEcjVQI+7fO4m2HYZatT5seu2WC8w5iVlC+FQ/d81C
6sabClTbClAkfeNv6ht1LSqYPtQNKTKVdpbts2I7QGTgt+bvzFPn36v+MgptCDtd
ak4FrWarimKvZu09zNBu2qpUnPVwxHs+Git2lYpZErZFLlUlwScL/PWuDFwljaO+
J4XGhp4Iqq03WnCeoGDDZI1TTdLb46guPDnJR0iovJIPrE9j/ehZxkIfKMq6SHdv
EvOjZ5qY/zp5yxmXYbnY5Y5G6dSLrEzx+Hi6UnClGG+zUB3gO2+3UbphbpY0s+SB
KHH+gKMe2ONisIm0kcnXJECvO7us9rXU78QVpuv/IwK0ExsbGpflFWFqpCISyreH
qi6P2Df/D+8aWXa9sGuKYdiYLGPPYQ+/2hNJPzWrKw5n6gQy27bdrXRTd9GTgJeC
AKqImhEil+9y0yNJGTJa4rjFh1Zw7uSV+y+5TM8oxhMkOUkjEqvF+r6k/tKBp/sD
Pdf5fn13PY9O5L8vDjmb3cwT0HpwP1763e9fqy2M+sthwUk0II+dgwRF74Y8+Ehd
THoeFSDcPAHGB4iOjF1QvwUfAPszcJwqiSsbas2uk5PMhsax2ct+b1tu6vt8Wxwm
2prDrMEelFC96hiFkzqbIfPLREdQD7pPeFaTr/LFGtjXfRwpKVIioaezkxp+5kV9
1uVWNv4UlGWXUorsHGDud6X1T2sxVot2iIVsKJjSnTGkGySpUCtVvAcKnTz/P0sF
LG9EWFWWEC5pjyjDAJZqhICqWLx25k1YMnf8+ceoWXpgKONjlBth8CI28a6lawqC
5HFElHphkOgrD4dOAjfatzDMC/GHJrpWzd6WCBIWZJX6QDi+jzcLA1KykxIMnzeV
zq6ISd9oldRBgD8+uRMFurjGbzS8UfmplnOZz76iQieVIztFqpRFlIfyCS+LZsDL
higRecQe1vWYuFS1MvZh6GZMvEVw8PqDBX0r6gU+cIkTW2DD2bbilfoRvG1nauO9
2Ds0stUZz1lQ6DqSfU5N8xzehY7kOiti70++soH6o+l0qTddgsvegEOvVDuHJ9vk
D6Wqx2fDvV4byI3k473JbqEUoQHxGidNhSd29TlHSI5pzHBOpbvMrRzaBjO4Uf72
BSyxZFsNhiWV15QK6Q/vmS+w7q3YXGHcZElaJgDqaMzJSnyA7ZJPdwNOlveglg/M
DEcc+pkB1Hmw2cwrSo8x0ZB4uGptqPHhZIrWDAV84+eqHTAkLNiJenQdpjP+p8O6
dTJqInFWfEpBlOZyO+OtH3RXKlr1/McPMd4oZ6V5esUXIMSUhWlRoYcaMWFt/gcO
YIomBnugpaOnXX0VgxwWTqooQhaGL9i8NqQNmn33IVGM+R0YhGxZSX/lSpJB0zyA
GoXYtHvAWJLkD8CiBKPD3PXPRYf2zKq5PSjf0ZmwhWR6twyfTlcpNxU1RoEebaI2
Zh7h4pt1ZH+KCJZFZ/vZr6q8D1BC7pBTLPGNjzwiMPFJhrwQaJIa87oF8EDyTDFu
P5Q9OJq6F0Y9vZzcoBYSZ5Iwznx7DH10VufWzqigB47t826++VjMmtaCTrmjglw/
RVGTCt7fVGZGWSNoA5fA3MaV2vh7xsHyzCxaiEhNyKdgU5XF3wvorxNJ391So0mK
N6mY7pd+WFJaIphdv+c+39I9Ia/aNryBHlNyaAQTORDnVpQnf3i+dkLEKDn+DQSm
849HGnHna46xildaewtVIu3qUp970mDFjH8vkzLbJv5sOD+Mw7OXOXY0KOLm9Nkr
RS9kpTethSyGaaRhmYrnm/ZnhO1N1tBVWDLhabdL0hAFAS4++l9qnnOP7lhQx/z+
YrInWVUCUQnESjwPIklOTMUuOcf48mvmTEGoa1A/yL/MC1d4/1OAx4Jo2Gg5pTRl
YQ1j66CEn/azaPJ0il0/rUDYZyTLHF0PFRpuGVa4527Gk1vHfd/RgeuaRL27AZhl
awc0xhlUj8tdu/BAeMJ3tKIYs5wA+QuGQmftC2fhu+UfOvmGdsVC5DG9Am5FdLfK
F54fuv7NEPgLQNrvv9EiEniYrLt6TJYaG1lISY59AC8EOu+h2EYTPLkyjVchwTbE
kYHdHboAKp8JUjoSZYDOAdgrAw7lDxKOKFnL1ON0xYjb6d+amn0ZTJ1RK6m/bsK+
SNiLi9N91WhHqFx7+v2k27ed9Y6m9dheFEg30iK8dNAy7iTWXzeXTT72BuVRtFVz
zmjvhJNgfAtQCNA/t0+jU1uQ7vFyIAzkHsCl545LwmjJdAHiZrWZ39WGLtYja041
t93/2FUbqYDdxym3PPXmTDu4Gp0llYD2SprY7iw9tO6T+csZr/NmmII7AIOcwcao
8kJ0IgpuowH9XQ+e/ON+SE0XCrW8omqhsl7TWOxrHRaWEcCqjK91qFLFK8KNjTyl
aI5dHWyY3s5hfKbV3C+AIEYxm5feAaTPbJuVKfHAK4Wrwar9m5ZrbCzv895FyYFb
ZyDO6UJmh/nf+TEWIvJKozXY0IzOGnmJulAEIcgpTxDmgOsLjGDw7QlOmMjHGuCv
FGytbeCMyQA38OjOs2g8dpBZnb0Rt2rRIi+BH10octMepYIkwkVRuhG35msVTOyq
Uahq2eZ2dBqG/VYqPKrBH5OpN4i3PAMAv/PLtQ12BeuOdkbTAPrOmUr+V5NpktXZ
yqMqOAS6gePO/HPJxD+9wb4O5WVveJz2pkQkVHj6qii5niELHoqQd3CTZeE4kg0U
ldF+YrcRN+fmL0nk4luV9zxmsAdma8wRDbOaUCyxabdGUj4u6Sr4NC83Zz5DnrI6
7Rex+tkhnX1803VCo2m6BgoH7DKiK1CYg1+V348Yxp1+jof3wl5GAeHJ573WRc/5
Wf73tzZMBilx3PRUbl5eQZ1RJVAPHwxQ/vWjv5Mv37Tl4bVOo143tyAD9J4+0itc
B+7m/6aRwJtRVdcr57ZjSB6VL34x20nbLFModK7FHHzrstydtIQpBaxwU98WZcDp
jkekTrPk53ND22w1dnYfoZqSIAhwQBmjdGghKkMIH3DQLTwqhz2cEuvhCov0nl7I
0tOqDsv2EgNiCbgrGMf5TzBY3NI4lBM/nZ9glJ9dRFsUtZ1KFMk7SMBRzGSEYT43
znXbX77R31XPCqxdPy/4wbBMayWLMEmqLziv7DF1xltHZyEY58C8SZUNQdpwpBbG
ymDlLrHCFw/OADlAP6BR4sYusBroZHYHATlDJVYyr01NKCpppMkGXCMRAEAojgxg
EODhm6e6q68bQNdwtGyXsNkDeYUXb8T84nVxnuZ/4FRut8LMVRDtaOSOSPgP491I
zHdOzoLNKfLOwR8G63u9FoM2hEQtdIxVg+taB6XZx3fZo2dxLWP/blfCNo0z+XkY
OL/R6N463HCeQ0a6qkwEoQbL4uqNiHxcFzFdCFWyW1VTbkN2kef59wbSQUHcBaKJ
yA+kwKSMvUIWDjRW3qrtGj6wMQ8njpdMHNONosFU3kzkmnLnaEnjC/IgS14wZ+GT
dwyuRS65uEUZDOLZMRBg9IQ34pXawARlFar7BeiogDGsQiftHoN2iJy3uctzPp7c
rUylmYmHPwAs3hrZ9NdIGWxkLGtBIr07lXKBGOPsIA8rcYGe8LrNdMg88yj7KHD7
e8AD/A7tul4i63oYJv1dD0xNL+qm8MDaK9CyniiUITgG7FQwtbo9++cZNBskAs1L
3xIN14XHDnmMpAnyA09xl9NYuumh9qJ4BQelb1jdKjFDB1w11us/2GZbhGK/OEsx
+Ii4qSnIKI5W2bl3R9V0rYTKGGHLRjLEUvVPPfPAi4stWI0Yq9JEhrcDHyK+HUXk
Zw421s5di5q1q5qe5KsfxnmKru9ehR+NK4jSigFOYBGNkPiXpKQZDwYcW4Aj3rHr
co/WCTyfHX6jFn8/mxUdCsp/3OtitEF1QixylLDWZp2Hceb5lC0ZPl3UT1Aitufp
cHgjxU+mpLcxRjNaBlZb6xHszTSG6LNOYmAxMIdfEUrcLe3ULzLon1etZeupwm4A
BANU8ZDLyqBe+RCNwJpl3kbNPdOMzo8jI6tqvinnvpkEvJhMhDkUzOSKjktMe1bw
aVyuFsjrQXki0gKfgB8ea06A5C1W4MfxOkzBYVWqWJPbrnAGi4C556RD4Dw0E03o
hmEpKslgV3TvUejYeD473GEgmKUkw6pxk4RRyST30aHsZjcOEnyMhzF0SAy84/99
vI9qZfMZZ2lPh6FYiwxtoxSnJ2ul6SUYOeHi7jx3vtgDqfLABZQj8p9LPghpXTOq
/mrCmsjoN67OUMvowDDS6r8eETowERaGa5wveT0byL+ft7XubevAbu/8ZoIP48x6
6bhSmAMTayadUqJcWjIpUaKnqvCM800AwC1aO27C55/8V8MYjjHvjpjvsSlKmQ75
+B8RS69/+w1F13DzY9tFW/OQOagWqZqw8qxmOEHYp/dPh/x7cEWqSmG0G1XE0V4I
sl2JCvrldIITIfpjhYE/0peoQqOHzZTIxN6+AAoQIdLDTsHJN/xQvuZcgP7WBTXZ
QEyZy41gUtb5vWn5UaMlNzJavgVaipHf11lKZ1SSyJxxI9dFQsnirxUVNoIJ5OHx
JJbXxDWAqPkCzsFqr2u/ezdnjtaxeVq06iM9V0nui2NdRrHM8j67HSGlhThV8Uij
IeOmt3BoyVkuA6scSbhDzvPZyzvGQkfd42PTSdRV2M6v7oCWnsUrIhh/aIJN2yq3
7YeYD/7PJ8Mo2aV4LcJiPcywpwQA5Vc7JyVnwFeVq/oIjba3HeWQfVolJuY703VW
vYDfAldWptsX0sp+0hWbE0b2BQ/2T+yQgyLE3Dc/73qizcSuDgqMIri0ceJNBWKm
17Rt9OjerdwyXKD+aplEtLY4q6fEJ988+nzCmbtIgVErFsKjIJYgxYEvV8JiNgrJ
9rwHsdPUM4pmEbmKtpA/4ylV+Qq4JgUEtCWDjoolpoykD7K1D6FPrnRWriiytDUk
R80D+U+/XzuOBmfVDp/rML8uUudAjuqGmn0FI8VwN/cZDvbEcK4rpsV/iyl6Fy7U
/NtxQH6f8s7OMOVc5vGJ4/D3+vDTeFhzc1ShGd4SdtR/Q2eSiToYZKzrVvMamcGX
8904MDhgl5mYCnS0Xc82OYvQ9u/y2I6FveI2wXAoqIlvPeLlEaBcmuT95gQIrIsS
k3Rj30JeCuYFRmVMXoRyRym2IZytrOmR30VZ3ecs7Trl7J5qqNd/7rOmxsp4grLn
GqZ8rmmQ2DxrMlTYZDHgGBYhPe25NVpHA0if/AYSyGt9u2PJAeScjQNoLDkbBpcr
lxG8cJpt4MA56zqL2b/scKk+xKfPWABd44gCFvSejnhTHzq7/mlcM3qk+o52xpin
5cXvCF2Ymt2szS5SNo8BMtt/P+FGf9c/+qneVd7ko6jEk6tKOusucjTpPUquCoGp
VjFda+8rb+vmGvdIiZuZXw8lJ2++3BqyahDhMXYBfcMikLGyWNW/AHwNQUfjBzAq
uiQcYp+E6gwAiYbEhBqT0HBh17O8sij7qAJRTtGurjudntTwhuCztR9a2j5xdJCc
UjpajQvVczx7ZqFQ2Bt66/MqTGe+d6HwnxXme+Vp2xht2cSGVCBcrx5HprDVxOES
h9RLTIoWcrGIcpFg/D/kFQchJKkjsMeunD7MyrF4VnuKlYM8ChV/49aSx4RmoLBr
iFMtwLmyejo2xZ+mGhWAuKWhFnRpVmXbyr0wutzpK7UvdSCNLZ6//0G6IMI0hetW
rUBKAKA7iyB6sMUlBhqgvCASdDvKU2sMKcRRjyEzlLFzM9DHhAbKdUSGIdhAPWDT
dGllPpCbV1n4ifgRsd9s7qPs6KUlQz3zDr71MpXdB7w4qaa4pCIt9yHZwlztRv87
a1v/+nHdVEvadLoELakq4LvGnBjva9jMChKWh7sggKUrJQB8+TtBgr+zUFNZpFdV
QbO49W6n+R6EpAsn++vdMA/sggX0DQ71kwde+d780VWiZGyjO8xNXQKIh3E76yft
aBrhvB+p0m1SUK/UOLpy/Z6fWOX9+BiVMRqy6pOtdGnC3uH+u3Lwukwo01XtOFRe
/6CoTs4fH4HaBAwk6qYNYyb6Iei7TGAnR5vqRJ9O07q1eDi/wNndJrfAv99G/kwb
zYJ8HUH88KL6vCHCRyJw478iNIHOhdkyBJUMF6hy3MWoxDzbG+YzTBVqlhvBH1ef
0lqGC7KjxabudBMG5FMy3ZGWfqQh9KqgkCx1S90BFYstO3DiVAsw0qaaZdjYAm0W
Iqv+JX5J8/xYTGP9ZQGxc3BaXg5GQsVaMpPQn9fMtIgCuffImFUr44mghkyLtDmx
Ihbw/9qdjwEyG2bvRG1+kzlB3g1lH1MlJXnsdLPdref9D8SLc1kobtuvzscxBuQC
EgNxl0jpppontXr1Lzwut3kLmKsI0jR/w0wc8cds1gcalUBsgMkubrNC750/PNSK
cjNpLLi5hE3ynnaGTMs+4OZL5/X/kMjszEdjzmS3/ecznEygqhBLlKKX6pRq7vko
y0gjzXSUTWb2s6lnxgtr1gw86lUFKby49RWEefWBbgTdyL/3LExcN+0GzJz/NLnT
d6gxdZqqKxayItopivEDbJgDj5Q5e9fcdsyfdyYyas4yPNa3FtFYBZRdbwKcPkFa
tTs4M4HAlCB9fqoDruLTJjOpo76MShphgUITNVnbKoIKWD0DPGd6mNLqD3aoVyhB
WPRHyPIDGMPlW/V/0FpyXJ9FWDi6gco0T4UsJgwY2XObpWYUAIn0Tz23bHreaAC4
zoXYZw43pt2Tjs1j9KjBbFH3khDy5vaAK4iDVW5GQUVt+zeTKM6Z/Nx+hmKnuScw
CJOwj6JyVTXm3JIoKB0qjlPlWYPJqKSg3kL94fDxhqXBhLrcbys/cAlfRzTl5j4J
uOm5t1tGYBr2eYiaF3620GORUlUqqLN/t+q1gd1MZOtebaIoDtARnY4EnVs32c8a
93+D0npjiAurZ6sGecUVflrZti5o60zyUaLMrRxhvrxUcidbMviJRL4E/kHFKUxv
A7SOxUvinS/QQZLpA4M3BAv1z96Uy9j9hoVQo2HAb1ufL5CU8UBycmPf7WyI2uBt
tpeUEDCjfSF0pSGmEvk3MwafjKUPb0aK2S3z/6ZrIjWrWK31hDCSOVXFISNlm27t
wqp8kvvFFCeoL+3cKsk2D2VT5+Q4GG1Juvbsb+a+Zm813cNQj8+Gxyq0tSYxooPc
qpF5kjpzXiXYo0mn/oBH5auwxGKZIL/Tq26aZCVW6W4S878PSiSTgqxdvNzEX35/
8/0wl+7IlW9KsR7HV7Qj3IeRrzODz8VPFOt102EExOzr7PLxhugx8xGbdm0nSMQ0
ySRnp2CiSoM5mEgqYIxGVvg+vKRZCkuJA7NtU2j744nZrsc139W0DVtbSnIjxLO4
asTBrEiriuWSiXtQp/6178L6H5gopowN4Deyh7PfAvBVWwOUKT+i58fGzoLVuTQ2
/LqSHzR9Za18lGIKO53oNqwh29BURp1SqupsShrryjKuoGHbKKEN9EpsMTP1Efzv
SqJYNlctQjYTHalHe2634TgnhatYmDMyxmaq8TtZ0ma6ZvRWmEcsqdWBZX3wQWlE
EgFLNvvMZWN1PBxqD6/LFgRK6c7r/6Ak0sWG0Y9lV8FhwvFD1CxZfxmUR24RMfj9
7UM93oUWOXtR0/4DfaXD1tMIUhh+m3f433rLdCJ73J/t5SqjZTpFtWFC41tYE9yF
+9dtLp9AoEMec1oFBD5nB/BtZryzyEX02N+2hTKUZFOg99ho6KDyWS2ZTXWzqmi6
rIoQ9iSIrz215Q84bjJ41ajwtCRN4M1dlTR56bBwt6ipdRLKnn1SJn87QYUjhhX2
vtTd4gFypghAj0ikDdJHaLfGFJX5K3WVmxDK3h+eAMcmYpjlZbuy8M/gPAIdE+Fu
bzNQYBeow3ZcAy7jLNkMYBt7MWRblcaZ8c5PfWhii8BnvOsYGan4yCYrVKZk8dx3
Iq2h6VMRbctGXfA+xrQhz5yFlyyHrcRl2OC5Xj7J9mhwBlrzPGWrw7jNvzn9U2ed
iw46Zl1Rr6higAJPvHrA0JFjhu2qpKIX8AB+8PAPv/7spH4ckozamVkpg0DIjaaC
3AJtBApQsJqYiml4PQ3bed+C0iwxFa+Azm0zI50yTA8BSqMVAdtzb1w//K/Idalp
rzrgW3dCm+h8ZpLIIKJEECN3Bu6b2AskK95aqe0I2hTi5T1x7ySGTSOy7HqYbkJZ
0nstaq7Wl+3bSd5kvyXLyNbJdAw09cztjXy7VJhGBcu65GaNcunNYvR8nuSapkRu
exr/Ub/LuB8+RnOsfOyV6DdL4gufWH0q2p733pkkOFPFFc25es/FJn7JKxV2UBWh
t8fU9aOuTddOqVY7n5CorzWTI5Od1e5NLM4n/hNLPidX7aatbrSevLfiinGhYf3g
KsYJ9zcTp27hFWgb65E/k1SO/oTllN2xMTF5kQ/3zTZuJ18ChtDpp5DEcT+6DCdC
cul4IpQcqM4NAdLBolRRC8RzSiltoQZeHvDrD7niUCVDqzwZbHptu63sKkwsVdkG
nTcE1p3daQBsjSoKH26R9bgNaPTtPJJAABUNLBBrgwyqVh9Uo86I3lNo2GbjCfaN
oSRm1op6e0ncm0BvX0mAq+6+d48puKdWNBNskzmQ8WHfefmwtcgv86osvaDFDwX4
Bm+FCuTyMGDp0qSv6VJzT77LvZ9Og173F4AUbNATjdFfccv/gE5vCWJzfw7gHBC1
bUBOgqOj1jrERtvPbk0KydoErAyt1RlNm/+YR0susy9bDWLr5vYAjnw3nYjSP/IG
OJzrz+ZhSyzOEmpjR7R0p/cPh/ctwgM4V3OvrDwZNzM0TUhlUXkkE+a2ejlSL8Xz
uRtJ1AMSAlDVCCZjrsOqERLoAWOoWSsLIF9JfCgPzruFgPB1tdzMqvjyDt2cKQxU
wbJprVuwGoRUXrFYqvrrWwOK41fOBmgkbYopan6E2HnPyvMdJtNTHq7xlcdUa+9w
mPfXG3FrHBjnc+XGqZmPYOkJ4ZyqfSDnBi7Kfxk5kzica+qrkRvcui/5rHEL0zbM
fdHKN6kkjmciombY/dnq9qJgB+wpGhr+OuXqHHDJus+ZEQQ28q1W228E69o51QPl
gTitLvwH5ynj3uBNjLpbv73Nawk/QT84WRWA5G3Qru5qCGvrtmQlqBRT8fmTqrJ+
Jn+K8MdlpVS1b/PdFbizsxwHjfAEKFOa7Vdk6KVawpnpO7geMTXL2+5Rk9YhSv/J
w3fAk3kp0Nzub3HpJSmT0N8masSfaFhklYD6QiwDm50k3rgcw1jiK/8EUoQjtfR2
lYnTODoMi/ZU/9p8u7Yq/yHyoPUOb5+rcBKF0QmC/pkpg5gB1n+seOMf8Kg08ftL
Zdw6bh+O/V/as2DQFzvG+ZxClMTW8HCj2kjl2CyXTjiH31IZfaDm+kEeBFCyDoCG
8l56qOIyGhBYLvtO43Iey0gokmSVKNqGTozE5iti3qe61NErWAy9ZaYq1P5qodKo
oo5SdXJ79QNabaUJxcS30baq68LGa2anWCFjr25JxZSeK/uWbM0+QvTPafstjBiZ
wCmSrdUwpxbiJIa6p1z0bxJDHEqJ66JHMqt2HHQJIQ1kVruEIno6F7NO9emoeEz+
JJYDsOcI6Pfq/bDJXpqFuznv6PwhHBTVSRrLmYEcSbk9TCdCQLILty2jbIBJjrev
+z2lzF9Kf78nrqreUgJwji3SSgQ5WWVoAnRAp7cHB4rNpgZo2gQAbZzuzws52tos
e+0/rh3QggO8+GOuvncIzaFX5GjBSyw8O6ST5N6+lRe10yJrSaHBPqfXAt81x+bd
q7sUD9pgYQciUhATrH/A3HG18WDNMHg1zZTTejeLJFEAWi6ntZo/3+NjAvXQlW0x
XU4TAfMPMH0kYPhxqSMOng8/T8kt72xVGZCb74hCgLMiW82XvPiMYLiQk/p5Rr9/
Qd1iG6tMbT2DCFVRDwRvJQz68zW2OyE0NxNrYUhU/G93PVg0VMgAKuCDq/z/uTbq
a0W2TkFyQcaXolOyiOberaZ/MgFTnU082AeHqS3EsjKFliTV1ddlV0329108moYn
qTyctj6XDPy3h2U0kUUk6t0cYPyJv8gqI95eQdW0CzBqbXS7AUqTNbBaRZwE7zsK
hsz8gjuC2EhzoSSKIpuJ3Ms3Yhs1UyDXsqYXFZlJwnY+1yKCXf8DIMUVAOOfW28f
4Sbusa23VVWdds8p6qH7+GaNDpkDp30C68DwAwCr3CFxzMaxCMNtmfY7u2CwyRBJ
hyvvK/5C/Md//0UiSCzsjqpLVwFx/QX1Q8g8F8cZ7UrvdfI4fNQKlE8x6ghiiZai
DY/ui4gPgMwBiHzzh791Bnx8ImB9adEAMBJg4gKREKdyAWo+6OxO260T6CsLjGzs
hEiMuH6QxmHcSF9pVjH/h6A9nMq2BPvu38zzHh+MNAiV8ljXcm6vEhPY3AtSBxv3
Y1yPpApVf58rkC+eIBuzGuQfVNQMMxhFwHhUS51kGD98TPXxwvPM5QvyYIe/Y46a
L0cYrG07yMovX9M6O/6UZw2vKGwp/6t5bePujqMXQO3+Tz5l27NGkIWSBzU2Dl+f
gzL40GSSjr0U1zDZ84m6zQrtbsRRQDy6blRupbYXA443PJXXxzJlmNjs+TwkPKvZ
qOEGXsCMGrwWR7fSO0gzOnLVBeMngZCqrKuEtcV0z7Y4D21Xo+fCF76DL0k4Qrf/
zI003T1Pdc9u/qPYTw6tGrcqEbbM4n5/BD3PSRuihhtbGeBHIZSK4iHkicTfKNjE
/MtygOCc2E0/Rn438PQMtZoYQ4jp+NmIUKAn1flDk7828KDedFs+e3xJveQEunTE
mB/2Phuz+2M9NsA+KQTZ2RHDlgQsBh8xvLgFgXKW44L7yqAE78A2+jin0TXvL7cp
9e8Q/EJpZB+8UROaecGI8J8aOszcV3T/WxFCKjO4aEuIMtVAwUjXtvUVRwIeTeTJ
5Xiuaubz53DXl9zWa4LvRRRMWx1WYGHInB4VCOBZKzJ0MvDG/Z1kHJLoThfSOo7P
EHQOSbRp+XdPEUfvRpIa22NcN81XIzM1l9SzYoLOEUVsCB2T/AsAZ3wbVSDXVSfY
by7gFiWpm4Dv5sK/JVXtwjlySg/b3ngvzCR7Ulqk43yiIQbgy2jiZImCUZNrFpWO
UPML8EC1N24ItQVsum3q0N8yo/npKVMaDg6WYGiKwclL/dj70pjuMMinmkL4IwaS
FRDOW1ilFlWvr+8HI+PgpXM3wD13fYBCzy5CLF/8KeTPJmZM+7QwjzC8nr2yOe6b
DIlk0FIYqbBAg3vpujHunQqMDGdzWhsbjYSrtNsl4zeflXGXEbeF91R9p2XMxfuA
SZEttzgXCXNmWIP+IcEZK0aoDA9Ew+9XcIpXi822aoZnrImSw8WjArG7taHtMHJh
tBL2wZfeXaNUHHi5jXGXWJxZqsr/HG5MlqZVPQCOYeItmOIRgKaKN7z2KZ1hgOv0
v8tLcFQDvEDCEj1DciePzf5g/2srVmUIbyFfxPPqvHfJKvi+7FfXEky1gUbAHvRF
JFvj/UBAJo+qFuovgbHjx/lBAdOI6i9ZG1ON1K23wvD8rPjvrpR5/vjBNeDBdTLl
H0rSQqdpyV/K6H6lNkrTrJp6MPIGLn66k8oidLCOJk6bpVZ+VJVUhjVAFCIp4gpv
h+Sz6y0E48gwWCNlHvdvGWvaQ37H/vZRi78FDOcfpie/shcFX+CUypGoqa624xtO
omRdg9836XBVpfVe3tcNRafmmH/TcHLDL1jk6e1u3RYmBmvxjT50N+B/8oJu7hKU
59Qh3WqM3vrNGTr8+rEYzlY6dkWwEdPYgP/gtfHzJXmrQ90ZO39jKjtKllkq8Ku6
2KDxCwD3BfbwadGuuRkkFIZvcterJBRHcDhASHLozOnPBRIcttQYJpMANTUnj7VB
D/jTfcTIzvsSKnugK6NU9AYCPDOJr1KT08dOFGQQLkhzD8p6o6bjlE73ojZFhPqa
tSmcYRIIoZ8Tpzxl4dpt+glArA3aw6AqcodTh6EqlctaXSs1G4wPzl4SjhgIa6k2
g0uzx1Dcaj39IQTSB7b4xkrn0yOrTV4hRut4/XFDWswkNvInIQDzNitZGULxviX7
Z55MIC5t8yiMCn0LuYPPWNbVwsdkhHfDtuBTeEuaDx4ECcfjaXC8hv7fslES37kt
m9MbmefbtZIZ+YTGTvcFmrxbjjeh4eXIGWjbBLv1cNfIDEwQLog2eBnQa9OiKWX4
VLuMtLGHOC76J0sqYu0P4mZXVfiyihp8yt0If3U22rIWf1gJy5SVawRLcRW4Xx+H
Xu7cU5QyfvNrh+9GXffGIgnjEDe6xeGUryjfAXd4/vP3XUSGR57u4iYCsu1tupvQ
vXpRolverB6UyvJTL5AlSGZS74vhcKvJSkzuqWbxCTIBh8m7YqHqaPAm73IRb9wC
tUpj2fIWet7FZuyiHsZXPgiuoJhvOzech2CY1miYZXTzgofJnK0RueU/SrDu8G8B
vdR8s7nUWJiWz5QwrmFsfb6HDWygUxHRtt0O2jePNZ/RJrJdSmApTiWVt2DO9uos
yv+dt3GUeNIQDNhZdGLMZG6+wjfy8L+ohHKwVBMgu3ZpUvTA9JruPKNT73gdYZDK
UtG/5E3dypMOjCvD44Sc9IowD4rmVIgmwn0tbn0HY8bEvcBdJtB3uJl/p/6zemw/
pegkXJnbxMx5D7C88Ed0TOsUBnq6V0eP7pU3muB8sqQxa8El6ybQJRreJPIgymuw
ufQPEoXVXZpTjkdMJ3yDLXthMpWMBgxqPq9g09NZpA3STXTvO8Ey2jvGItmdY2iH
+AWpC7PFP+F04tjaYYRzNka8s25lyIc6CmlYPoFJCeMke75XvQ/1n4jClNChPjHL
Hs98l5dxTtL7O/8xlENGZsJyAx0DiIyfnGjsxt4TagbjBhF/ECTE5Pen4GCpmM0e
LFnyoH0p4q66Hk1NVu4FxRHhnVtWxohCvSeQgMhFGXylgtXZ/CzxwT14X9LFnspq
JjMs88JXdM+pnbCvjkFFf/V1OXHK8m8wV9R1bwIO+b+tYplpxIqCxBwZ2qZcFRVf
yZBLCf9IuwGSus8HjPMrRIUCQHC1nC4WSxo1rIEPrmShEAaLXilzQ2ZjoPXz6fYu
tei3J83Husgq+0pF5J8a9x5BqZ6iZUgGtko4C8X3knq/0LyfyHwOHz8LI/wSH6mm
6jvJY6D2oG1PI7pg6qtWOMkJl4vg6c734agMk5Ba8i2PRmUHoinVpjCpWZuiVa43
3gW6lY7XxQ4yQzMBESLAFoGnsypP7YPDVVpbpSwLPoHEremFasJ/9Qa+6Cry6ipV
yY6bdhlkrANixEcVou6mKdKI/qOEVzq0M6y153HWiMig1PgPayuoAaBbhboW8saq
wnBmKBBeMjH2a5WLKWDsqAymHkTfJ8HQ3HYwiOKpnmE8mPRfRkfsVTB7T5WMzxOb
rkj9+NYSbxf1O93aD3MRgSGU2MNH+11ZekOv9tbeEREqL4+kRVBB17ioQBoTSraZ
Z2zFHoKH9ZLvhd/1Fa7FzBFUA4qHfJjfvr+gM46e0c1Jm1s4+iS0JV6l0pDpQdch
iuVoKbqqo0WlgHEVwjtNxKqXG4tAJeQn6j8f8adDjBA55JgibvAsTVifI462OMzS
6+Hbph9OUmLk+APZLOJY39rUKAqyyHlNza/LheXglddkLNULE5CZGsP+oJdmoPAa
DboG0mr562wUFpfjF6q0Dcof+M3HAh/ZgHb8A/6syKiiEiXe+/sN99HGXiqTDuBU
IWnGiW4dlNkddNWzvreNspKDAVfaJvC/BkzK0tEaCEF69wpWgKkPmgNpWgMjRlve
YMTDU5d8xiudgNkdkpzqAW+wdHxVlEC1WsYMM1NztaTw0h/hMItDi5BGY6K5aBpJ
XDNtfoJbautCQI354o2zwzbwjKHwLiSLjyGkL4lcIk3OlktI5xb0I6y2xR2ifgfu
m0aimKCB+2ABw3bmm3RHzReIWSLnwKL5hfhx+rexlO0EC/S78PY15rb7FqeC3Dml
8YzwcxrQulxdknRqUCBeSOU1knCs/j8sv0jotoATJ5ISmGrL2LH4fgoqOPk6aSIh
kO+Kj+jh7/rhWT7uGTIdfl01NkiSv7Pbhu+/OWHe93Ck8U8/ftly2vUiTSBtutre
fy8rpsUvjVv9xjLkZzgWQh+jU2LICv7EryaYEZF1ibSq5HyBLgZghfnc9PedPZ6u
njJ+s7nYcNtp8XdbIiOYJTpEjiIKtf0HTr4R9NFDCTNO6vKu0+VshRYSK4zgBT+j
MEAnMo5wKnw44hFPTQT5qKLsFl7wwFWQF3gRDGL0dpCliBYveS1EYuaSGqpYWkUX
cpbPN+/EMvK47Bo8x5o3peUzU0mGEEoM7m78UJrWmkyeqyp1EtTtEuldymQm+nDK
TQtcsLxRjrz25V59pyI5AS+TRGqCefx+MMISonBz5cwjrKRNbwRRMpn1J/QQQmqy
BsCnbXgHoCk1SHn/iGay1hfZMaSvB/6GRfeba12dnSsp7l2Et+5gD1KfSQoDlX5z
bCxKn6LkRzsAyE8PkovKNcOG3qNM/Q9h+zHop20A+YEeHiNq3aVfQXT2CF25W3D9
Wh9GNil+94wSTiZ0dLMsfHkCD/eRvmUjyTA6jN3VnwhE+xMdm63DlAIxlSrsdUxw
bgFyWZmTrwyKqZxxVKU+QD63MhI9u0LXs6Q0OGHc/TJh158Z3jSPCFBiexRMURmP
QfhmBldWxFvcG5ME5MVyHvxh7jaLR5BtSQr9Awy3nVlvQvBLNlKQjOaZuffSE+oZ
L7hvulPz8Tctpu0x4/FG8H9nP2nw6u4OsScnmIDh6Qt+J46UpTQxN9NlRf4/pddI
/o/cfBdQcBe71nCLLOqr4yREoiHsfUGOtjlJvNRotRHpeOqGehBdA+GQjSU1RZHI
D0aND65uoXCXmJiFSGkXrapN2IDUOD6LGoZCSw71gDbKqcylgjNUCNe/ZciJL4yt
CCeO+Vdtrf5DlDC6XGi50B+QvPQYV7CVktRRh/4EOGD4CnL1evMQw6dBn2Eh0/JV
sHpeuAJySnkJDJ66NBpri0FriDUSo5AvnV+XVyE7iL7HGVG6caDcT2E+GMUyISgy
kBN7WDuifvnZFOpOcI1gcNqgJOKcsNt2OullJkza3T5rUYUqt2fDYFCGqRX30rg7
G6Xvnp4uEv57nH4q0FmGP5XxZLtjqXIEttKv3O6SBzOwPiEb86wHiOJsWkKvuttX
PQ/hiGlU0abNTzrdXZHLMXcceZb87zlbDVs6zu0uAYA8ne/ImkGqAQiCdF3SvZ8R
JM2QPgU4vqbsRvBCNhmGQ4Oq0hoWzW/whK/hzL+uNJrbezZOPtIv48gXkK0ZbmPY
U8Ueyr0bj6YLvcgapf2M8dmNto2WMLPJCBgavxio/LFosjweNNj/6Ig6toC5ilGM
O1BdCNzR/zotC27swyMG/eoVthO+UfOaZ8OkYGoO+fg57ybeOqMX2952JZ1jPJdu
bqdWDe2Lh4xS/C+OZLepbXySKK8kZzpIALcFgbVbBNtHKw1xsAXSI9eGnwFS+KVZ
YE7KutZGR/lPe0pJdG13gTuaTjoJpPImtAkERWYrUG+j5WTZZYJ6xcLTRX2sqoHE
ixODvwvhfvSnaixITrWkDW9uNKH8WpcG5pCKASGiAiP77brK0aNRLZIuptiYyYu0
mFv0nsGCsAqjW/dymiuzDpTLaHZagTMOVusPYQCQfQdVauE/LaWJvkhgKQltcfT3
lWAad7L/41BEdOE4GI7BeWBJAAzrL3H0Fwr04MiprrmxyEZeqG7m/xfvXIe7sMXT
IG8zIPDAccZuBK1RMxCYIEzD2jD7zCNPpv+YqaxvNOLoAScy60Hc44TlyJOjqCRd
mz8e86GXli1qocWh26ViatfW8y/jNsdnLwypCRjj0O7sfPQMolvUyXV9uBdVgAaa
z4UVmQ6HM1SGDBHpLD8Zjwas7Zg7n/DiRsgwIAyRYyw5LkMKxN2/GWdRj05GHqUq
LDXxqnDSQn+QAPONP4ViS/b6qT4zVhhTdx5KK3BNHHmDR889omOpR4vtyMHLFhhw
yTDYQoIgomgT34jsAfVob16aOdFaufOSnFVGxXdg/tudtttSgbO4QQEHwJzMAsom
Aj7bSc5w9KIUCEha6rNWZ6G/CEluj/biVDX0wPlQ4/cS5SBb937p4prEXneAcCaZ
PD+x/S6rZMjZFUe41SsjurFRit1uIxvg3vG9Nm3LLKnoFMPd0FKDOABVgHuDvpIx
NA77ka6dDy+h/YE80X8N63ILFFzXven2svStiygO+vYClqeaA46fMJ6mtUc8uTjZ
KibErXqj1mS/kM5LuK4fpdnRzuGLR853wIjhVwJtgH8OP20Ez9lyLPt9pytjyGN0
AJoHnsCIfBFwO3RLCW3JqhJQOkztQfYDKEMlf3UVrPspp98jh8TKquUi5stqw7Mh
/OUTdoGoqyfBDXvV2qijdR5cRbuV/fuKUnIgRhPi0mMFSuPUKtvA7aPEbPNr48tH
cNQHIC2HKEEpcMLT4yf8xHymfMSnogPyX9pqnfHPqrDHMp1itgP+ezyLrKe8f8yG
EGjk9YSkWWJ4gEpPyG4XYNkuuxYhvkugEpH7gwatu4MdPynr+gjB9jU0ctxz3ebl
7wWAkHDikCRXEG/vXgz4OAUVoyj1GLSjyVbdqUxXCcEf8bg/+KK503JdnJOW1Xs7
AMraVJOw72JcIMP3eldk9U1shGcNwPDybqH1JqKz3uQrWXZ23Y8dHE4MpFvJ7U+S
XPr56GB5aprwnxQnb69pABmC5bt5WKarPLu+BqEHgnonnEFqK3+XMNo3cKJHYFZp
YhO7pwuTtargi/2pY493gDskwBB+vTxX2trded1bQGXryxChxjJP12aJCBnrjaaP
NxMfbkESKADxuoVLe9WxKLhrDCSSYUAvoi83/Gtyg3qteqiVw0mSjlnSzzeR1WRA
Q8Sjl3WJfEJKiEyHhnMAKJzmQWM2aDDcgpUHapYhUfnTQ9nkfOzHxfxIpnphmCb4
T7fNjDw7XEqcxK5/IVPm51MYhwEISycU3g+HC8q3V5YAQ7ZFYEmw48Y+eIi+v5sG
Eb1v5/fqAWLkedEjPsb+XZGqaWSoepExmaqRk2vBcTY5Os0+6rmZo36DF/VcABr2
NKPhAkslRyqZAeK72Mh81oSpLfWCIik77t6ifgA4ujXq+rKvfA++RMgatdcef/FS
fDwU7Yd/H4FM++O2mvOo1d/nebrb317fGVP7MUjWytNTpRgss5u03m4cBEe31nAs
s53RyhkHQmYpF1O0UePOEboftBVTB/Ej2vFvyGLQ7IBtzQouFZwqF1f9bMM5jxLt
XDdUAJUxizPGYGRbjhv0G/bG23YkFGb5JqoKLOk+dpgmmq8JWByKJUG9S5LRcZPI
VCTiDUbItZBsRvh9MHUVStlv6yxz98t4ST4Z2PNoJaK55pZ3CwJQtpfZuMRyu6AZ
RQGxGZBJSpiNPeC0OkAYEH0GRsme1Pc5tj9j9xmmRR0agZedG8sQBXH5JV3kE1L8
EocbAqkRRwMhJabt8GdPisa3AK/8KP9C+rGuW1I/ANqG0Jbay+3z/02cdsMmpATY
fj1B/agjdm5PBxVJyyjKdro1m9qoQa72qCB1ntjY52T2ru7KNlTR4IFt6SApMoN5
rA4m+HpTz9cPeuaGQ7YCKfc/FJRKOHlk0ZhvVgzTy8CwRYxW8pqfjFt9YhVjBFB1
T2tpiSAxz3MQGvPuadHJvSV7ypnIUOysUqYDFDX0WgjB4ss7Z3oPBvwokIgCFiyo
+GQqC+JClFgfaLCk4q4q2uXbiZeAsqpd3GNLv68TOgd829aFgKAc2e5WpGa9UBUP
jgjoQaHEvkF0m/5LH+fhoIN4BaaumNtmvl/lXIc09z0uXyJqKGKeHYDj1V2+TvOs
isOxU9JkOJaex+Y5xFBoOXLzbuxbUG9ewgAuLDO646MOnMC3l+rWGv8Yulbe7Rfo
xql8Au84dIcbWwsca+JHWErcUkEjCDGH+Q4VgI47TbyzZAfmXPpFbG0EY7bsX69G
Yzc1JUqBiVC/qxt7oQBRUBj2hbHWfAS8EgCXww5rARP9OS8yXtUlXEfeGDMcB/kb
S1OzN05fv47uQG63VTIfIQMlyji2MvzC1H7pn/A3lLzTQ4vTqenS0iKU50n1KPoN
YcETCOc1VqQQF/CdCaJ5nSehh+KW4d2azFKKxIIQqXot/o/ar3EKw4/oNzKuIZFJ
VKCGgD0HACRIvWhR+uHvN1R0q3euihz2Dz30Vbh9JGwDZOkF0YLPEddmH8lhck3G
RVtYPcgLhQCq6EHA9Pe+an6foNnLYPXWu7fWjDpOAcf5ZrfAZE0M5F25NI+E7Myk
nm4e7nPohn4ItyFRuhXFupOb8J+Gaem7zm7uMQE3DxSitMmtlSCXPoImubeyut5t
0LdmKCI5PI3VEE3TV426ef54graAIrUbHmx/4ezlPb0YHHRo/i+VkQ5NrmYr/v0a
Cg8ANyVUAWUEdE9/tLPKdrjXQn6BgZP3v9/ONa/WFp6Z7GenUiBZ7JN3YKx0W3fD
LNKSwgFjakLQdfHl/0V2Qu5yBxWukw6Uf6UL1nE+FGuOSHdITeeIcLCa0NqEWvQR
qOf+qeX0aMyP2r/G5dblTmySRUr4QXWeWJ0WcJC/tCfoNzBMNoMrvjfdBd5sPLLc
DgE2L6ku1TnUGZCD1/lEGJhT6mOd9/t1Aa7V6dB4fS4Ve7wf82zpS1mZ2mHXDdLq
oSsNEJIH9uHG4DAcytmmM9/FqANzKNbaKTN+3KD1ebExhUvHCDdxMtjOTEjQXIpy
sHsncFoNnGVn74krcSSr3IC45MNTMG34Zw9RgwPz5zaPI3S3+2nmgSG9dvaDnB55
EnuE4V4SK/TL+XEzQhnY7hx63hlerAepCMmMxYyZ8URjgDAQtH/NtFrs2l9WZF1z
RUq4qSIm7RfWfUz4mj6bLWMLykJs5gYe7PEewV9+zrKSwhjsp6bqLHX1aiQixhbM
Q9pnxgS40MjX1naoRwxwUdzS+wFp2IAWQfebBYk8szHDaf4zzoOdbdPfH2M6R2tO
kMgDKg5U1XpsmZwlygr8nOio+JY0LD+LihfkZwT8LZyo6a29tON+1s3njQ+KcVjD
zEv62PI+JNzDKUFRz31I9M4EniRI+U0Ngy4SlHNaHqU+zPAPO3x7/51MUt1PGLbc
1u0lZAv/13ivDXk6I4Vc9TuCiNwXnaxw3fjfBbfIKJJcpmv1kQLehhFjI4vDiKXC
Fb3lxLJy8FwDNJOgTJWEQMC233Jr4ATLRTjSVQukRcKjVuCcuQv92R+P+jhoR+U3
lVevUh8iGG/TUBMKX9J5n+TT3A8O2VrW0lTzgAfHmW654A6TYoI9X0OXirNmhMFL
iKPuGpx30QfbMFfnUi4XFFQZi8Zv6Rzpw5QEgGX6ekR/kvQUdRFYKsA7JnHq/amw
0fQrnzzdNkFyXmav6nU6rwTIWs/m73HYC6qcQFBSgGIeDakNJFoHcpZpBj62nkpl
J3W/R32RvdmMGkCIbOMgxtMyfQRYoTzydzXsHUDYbvqBY3dDXQZ5NaGNSmibkkr5
IrhvPSFk6TgY8u35MoMdl5qRcNrJQrdyC5VI5p897nkk57iJuDn6mht3cesAuuGt
snbyG7RIItNoqtOLyGgpuoRfk9ntPZeW0Dki2FZb+jOZhXYMFYUBCa0tnsIEmTNE
dClr4GSwDAMHl0XWhzj1h+ElVaa4XuFVxgPJoEgx6T7ouNEmQGlEN47JPSQ1hU1B
7gvVOrubZrfBTkucR9hiQEyhVoRlUOpAPmBarVKZsmEKqnr1QAzbWuFJsY0/8A7f
n/PeLaYnLmqGUtHj2+jc72cGQ+5tjnrKn9U8qhGm9DhaGGgwXLey2nW5wJDMvZQO
N+LD1IDqFo4uDDqd9V52AneG4TVo1CLug+HWPI2ONv5NpKJq+3GAMQGeQ0jc/QPq
vMOGT5wZ/+e0QEveQfpkEFdq24+VGeUkXsyqOyfwuXhtD3wLNh2Dlf2Dl2fYu1Gp
fY0HP45tyBqF6RTkqh9H+GMC3vCSi5prtFpNYPQIACFBS8WeUHiiY0GdmrElE8gL
ePdkslf3q4/cR8HQ21MKN28fS2U2avbmZK/uV/qiDQ0B1WXQbv6pmsGfpcbienfI
mhKIpTs3Oa4fVaD0mMTktEvdOgB93aLibXEOYSlUjkOs3dvTkizihHd1hWLeBe53
t9MoAch0Q6qPnrfypGMKSNZDAZQgbX3anwzXMSpCqxZSgnaEXfWT6EOvU10Yw3Fq
yg7OtX7O+NWSgMdvp9AlZ7wvgBmkSf/64yRUTDberY477yVVyBPWQv8XrBtw7Wnw
7p1oJUc9bFq1S7aguDO/kt2ysMs1OBJVyLp/FOg2isMW6cgyNK6OnBAm+hrgGCHi
ZuW4xrb3MAj8pX9z98jOF/qWt3nEiwBaETXRYAPw7wd+/OuZ3tIvJ6IcJhYZLVlm
IWBP95kIB9UfkkQ/Orjhnv+e3E7hvZ4k/jru+bF1WZblZLkvCh45p4GeUQh8LCaJ
yrjhFVC+rrj3uHvNF+HVX6zVQ6LTTB+kfxDhoAJs3TSF6A6ZGWby/ksVPmI2ctBT
42xElud1k/J5G4xIOC3x324kNcxdwXY/dtJN1iQ+3FxvKzPZAvSryXFp1yin69xd
kwXOHB/q9gvgXtdlAGPORXNG+DQiJ/oetXTihl9AK5+p8KHSV27hx+XEegvoEZnq
2wysFBtcLq0C4hqiIzKSm/xGIA4SHnJcusUbK4yfIFUcPjIll1lMEw8qFJSJeDY2
yv7EQfPvA9Gv8zagCGMd9F86OMvhfdTv0V/Znyml/op63q6Rne2EtyWsbqguJF2y
FhPV1X7PrYJ/yPJDQEktzVmYqmMPNjRMdcGAVZZEKc38tjh4qOTIA6i9NbH+jaEH
vDcJz9jHgFqwBfT+KA665q+/fHZVmTryQ1DifLYaio+6MZSuuBvU/v04ww61z7EG
2n188nirBUASBBYRqyAp6AMET5UsrwxY1Ke/eXD4fsfscEsWxGB1k8O5VX0O3Po9
R2J/L/viR20xYKpOmwyEl7sIwe405sxVFrOKzYqGOQdaTFVzEAd/osI8NmvYsCy1
ODqrX0uhfwUuKZ9VKuX6cfNVqMAeWHGCq8M0CfjIhay3Ja3anTviyT4uHDI5na0e
5ULNTj0iFCBpA3iEwMcWB+3u/vCayJttMcAjHTB58tpxOj3ppqFdogKlKiLT8Id+
JXta66nghZKEI7FkZIGTQ8RSC02ohAEx1mgkdg12B2Hrc8xgpsDWLxDH4PdXQHvI
cqDJMud/e06OQT/04S3DTObT95Hbl3FnI55lzcMWDOJEwhITffFdJ7ABcJMKzQg6
+KvGXOqzB+Qik6hcqylfd72i7oC/UDmmnu7uSCKITpbHJ2bpSfHMgPbzYnt0Rd6Q
n7lodjdm6l9N8KmZHLc4r1hqHS31O8k2ENf8/RNGlviW+U5idgNvp3ehKubYkRwS
GpkDoSf8GNjkSMUrkz9QVHegBHohCTqP33rtQba1yp2Dkv4bOnFb6BBlvTXr9S82
KYJxlQSPRgFCEcDDuDziB+gzh1hOrrzfX3Kqpl0GzvzZayPaTYZy2GtvsSO9PVKb
WWxOh12/By+0fbgLMyY+m/CxOP+at3UxzfI8qkt7C/lrS/2SIa7Q8rWVmvK+700V
YcUTT566PJgiPWNbn/yqon1pE6BL6Stx+raEr88i1jToME5MFfO6af6brwZ07SQ+
nwz4l6cggJLWHW48PrtNqcvO6FRUray+l8eBsZ//ztNBmpenvlla3BVwywsZ9v8A
LpJWMt9Tl9C2BkQ2o11eTRTIauIYI2J0+X4tBxjGf7/dBq2DniHTE9Its2XaGctl
+L8VHNxRB7e9CGKz5OdCp+MzAZ0uiDVHA53X5OTEKVdFsE8NvLiHdX7IucPzbkmj
QwEooh8OjH+6NZzbNEXBgIBaYekNtBbGGX7aI3izx396aHvkYnvS/3M+65sUhOCL
7zwCGdYvRwO4cAAaVJswxxicBBbjeQhFRaw6HknqLua3Nr4TiXScj/QO4Tt1yK1W
/MVFSX1XrEYrVXUoQ9XnzrG9FuRaOp8TmP476KEXSp0mj2YkV5BM3X++eNdEOEWY
OFt/ICVY75eSxR3paImVtKXLPScTrmcj8GMLbVR/EE2rUfYBvRm3qOXs+fIKvzA3
Fze2tFs9AoaALK+wN+4uFtMrYWZ8iJLmTvuKV6k1Wx/WNY4lJrnIHSf24NPaOzHC
c2WkwHn+3xsyQc2mk09gIlSKp2eHZynDr6Ge6HRn64nGCC086FaaMt7H7XFbKv5l
rHbHlEEni+sPVQGnuEJevcrAy3CVRUoveoVGzlMx3tGi4cN72ite+w//g3FWFGFc
YCK9DJa1FnvcgvhPxT4nD2Vr4w9PYLX7++9kyRhiYSy40Yqgbum/MmQ1h4NT6pWj
oIfniOU9YQbaNB1Ph2K4QaJVBwBz/5z28nlylNxdzJ50Z5Thh8qaN2Web8LovEHq
4cFhfTNMhUiG9UVs/HWfI42lJEzBolH6N5lzacFGF1MRrEeO+7EHr3q6p30OB58y
j6IZRnDu+XlWr3AIjjTHf0zyV1svfCWp0jy2Vvx/a6uH+Ve5fRCmr7VP8v9e+ml9
lb8F7LKhik2iVI+8590nR7SH9EEIYg8t2v9wYShEz6ruB++AVv3u0JwqwThFkwas
291odBBMBymPLSUvTDvU+mJe+IMACgP1etqpKXUWoDrJTlvIpywjSyimfSZCKIjh
zRKAGdILgmIlQzTSxr0OWYGicWaXhLq3aFHPLY2A6lKoJCZWIdJneQ+lK3YgSbQ9
xuUq9E/wwI82PPKITrg0O/QRRNi4wbj+fCUTayBNW1mFJKl8wr4uJ82GzrFvTsMV
cmQcFu2ZHRfg4YPkkFoN0AQ2FshgPcotSwWHXSKDuQwrFyHxWsW9daB0TDJpuZoe
AL+vZlMXKehBMhSyuItyhLbf9RRAFLSdpENWnHZzzS/PvDo9SWnV3b8BcFXr16/e
m5mnOVJ0xispWvZibIh0R6T/HoetdMVwnAhei8bPH0aQzDvEgEB4EV4Ru3FbwywZ
clJduhRfoTYNA9a8fNuJ2HBA3SafmNqbzzVoiy2sxb2M54V7VfwrPry8Ngp9ktZe
aGGIP+K2hIHNcWZupasCovDPIS2HBu/Aa/kVLrkB8Etg6WBZviKaFdJnJ/n+Bdlx
KJp2JwhD9TVKIi+cG4G5cJ800BGEyTL40ctJqviys7R2yp3BHCKJxGwTbFtdyFV0
yO7xsGLu0B0RvLi1A9Qa3x+a+vnr/1iZlzUSIeat7KiaQSqa6B07OxCcbaCT6OBt
WeansT2T+eDiEmD9A864JruDsmote6w6eLu/StTvFIvHec++dS6BrsHAOjh5Yb46
3KOnLzfQi2FBqXv9l8ybu8+Jx6mxlf1AiDUnVRNQZAmtO1enDpxw4Q33MAp+zORT
7Gs7kuEdLvKt39gFV8YP4lW7E47C1QPkjiyqkteptfcjPx32g8Wq4yllem6BHHir
HPj8vMEifE+hxn5WrRqq7qrUKO73y5YOOpAtdB/zYvH3qhtqika+UuzO6F4YaBpd
J4VU3Gd5IauvV/Y4yiDKVts4B6SI0xLxpsiwBYILEcMpORK4OchjOjVSco7ApfIy
A+8liQrqweAqdFEiRkTp4UilWh2ii/HJ3DrtddtfBYdjFNpf7k84jnVdL9l7OMzT
owJxOdUJd9VjPxJf+mzNLOtXzwcp1AHR18fTDGIG4FgQdMh1ALJs6Kx+EzPBQTQR
uM4GEiVRTDwQd5ClkcEyrTsvzp1gdJXsjxIWUeRCr8qyndTqoRmrLCyKM5arZ4n4
qQSq8DnHqRethjy2tiRsl8kB6n7CwG8rAIqEU12v0+kh1FpI4gtFsg40cJ9OpadB
ToQTM0ccQQ9UALKQV5xM4/yLvaeG/jL3AfPuOKY5Cm5u749DeO+PO8JoqyZXMkBi
P4k0mP8+DhM440LTvaMLAnKc1wjggNY69Aho09VZjIwan5nJWvOpSWB0T+q72sM6
HJ4RJZ01jBfBT+6hIqRroJVOsqpmOMqukAjZScwIzCf3srBUddXplUi5TtKlM1du
CKpmMNM5p4ez3dMcxU8HnBBJAcH3VVG/jHUpuGK8RJPWJxzyINO3QpXHBgCqXYr/
qQJL/Bmao8zxB+jq9Ux4p55RN9QV/bm+Bt9FN//+wAJjQ4ps9ZMR0HfkjWOtacyl
qo1HF04qX/lakXapNu/E+yW+nj4Gb1pKL/sa2vGxhpwl+4X6YxzQElvn6JOBIA+6
6oinciGZaDn1TUA+N6xrXh1GPosDvGhrEnaavl+cm6PGUETSHVCs0FjXw+oW3pcI
X7i0FGZ57UqgnrwhwtmZHz5QUerZAfnPWMCICrEUQy5JIcq95wWKJF0Ft/Oisj3q
sZ6biRaK8bzR68bpNd9XoFXq8xvwTlqOkZH655dxFXfH6qH7pVqqIJ8n3MgCG+sT
2SRZtSDB97r5DBESKImVxOp2ZEu9pMP5bGSVtQGyk9qKJX+HWyklx/ypeXwPHJEL
idyengH6KcVgaujMNhCBT88kCgekbD6YAhcNe8z5Nh2nxjTmL6fjKGBsy0LZcfSO
9KOu2pmm6t3Ob4knh7Jkkr/VsSdG07X7GlGsI06sObaxY7iIi7G+iHL/B8AT3RbY
jHT2FWeet1GFXf+KXhSBGMdlvrClnxVOR3YZ0SFJPF1kenINu4hhrWEBP4lfI27t
CLKg0s3ESQyXmXn2lq7DDrI0Rq40dH+E2LMWxRni1FDyxBHz0RBx+hL9HjHzVHV2
pA/WxLjjj/zRjhOXMMpl/pHjl60Bl3EATQlSBUFJHcK1sfZC9rmH3BeYAk2KM68a
4QFcuPgZTvWExbD05wJE9yR0o/QeAezwJj9toMz1ICjmFKD0aGrSIHnG/8KPZMgl
JhWmx39e4PNtNc8ex1di+FvRldG5IwjjNrtgmuA4Fe6/qLrh3RvS/LVX5I48ffRV
eYSIlOfwGHAhrm/uOX3LoYiYlKx31IcloPNTdHghS5d/2J/cW1C3PF8Dn6tMG+95
EU8456vLJ4qjqsB2KiErJA/GIdqUzhdQcS8eGDqnNn22LR8gM6dU2y0qbR6+AdGj
kGv673PrClztELJHKmB/gy9U2piWmwSLLJ7Q0JMz2Z0k5HWApSFhLVO7/x6KGk/3
7uvPU5yepxTtaV9mUYEN9TXkSqFUOUEYFij6HU0SVrrOphu8Oq5qW+iFCRZ/zENO
in1lxhsNhS5msENiPVoigRfn5/SKHbrQLaZPxLGaa3bcJONygy9DAuQq/bwETAby
meXfYymSvuUidhoMuFNTm1jiOlhg8XoRH70m4A7DpUxhNSBqX/m4xxu93fCCW41I
gcPok6aoYo/K1f5+P3E2V+1PAbZMYbqUzZ6GxPnYzqb7GfUPc8DmYpQz4npYdgkM
7JMl+ZSnAZB4hOz1PBTU+OfN/smHPYVuzICMCC3jVPEIFi19IyrphuOQNZPgDgU+
BS8zLrCSF2zbRNwBwH7YGmtHha1p1SvdR8h7aAk9rzwFC/6jgOBbaBnDLsIadggC
Zn8Rt0+s8DX6VtSKerFzr4Dcx7y0UfaW0uXV1M16SDj5k7eJskIgXXaQOk2WVFL3
7MRAmAwd3ON4V4t6wr5eLrrPxCqqHjSS6r4ZdCY1iRd3Hqc+I73k6JsLHGAsg7zD
GgeanCdLmUoEUz5g+ayQtrb3+vk9LVufKIuYtBJGb3RuuRDa4tfj3cJPhDNalLc4
OCURw1H67lVKTflbuXIWDhiAZe+D0zISCVoTab1u4L60eTH2b6hn9Q60tOWLyviX
Ni1WaPkMYACUdJvv/hh07O9U+KDEiQ7j+5Q8FCzbFQzY3Wdtf9/PrNCvobgswihR
7c6o5DerUuq7YQ0lSd8QzCyRgzEPNzbDUq1vaJtdkrnIMjvaFB7cM+J42kEgExQS
xM6MzofIucai3RHRZlIfWaZPU0VX0hFP/Ptr+jnQ/1qHdviXblBB0XULkfgSFfxP
qEK/8l39OE5i5Ozv/czFBQgoFHYILFL8GxP69jlGwgfo5ZPjDPTsvgUaifxqxwvW
nzLTx8VrXexgl82cVglLGP5SwQ1ZK51KMRQKMe5iaphqDOYEY94tY59wh4Pq195u
LZaBW4zP78UKQL19s+/VjVBmdJA/bjwjTMLoRt8CW/bWsTGGT3PQT1PGaDRxrBLn
aniwHnuW7UuF15T55r1c174hZ1zlLLNpe0LoPJEN64+e7UPfajmV1OCz4U9iiiMC
+ergeUXvmQGciFguIU5drruxRJ3kI5GYaSxGaYo54nM21aypEBbH6mb7OnOoUlka
vVyLfvIH4kY1vwz25tXToJoG7KdLmYEEratLcel6LOrdK+QiQdgHOB2Es12En2si
u/nSjZ7Xz2WG3wtMFBB05unfNAf3MEJsjudif9gVxLsojJQP6/U4H0zsuH2JS0aj
vq0MmfUnqS5rgNaUInmsxBe6Gd46fHOIHpqvKdoyYD303EcNCObbKUq85mU54Jex
i5BSdv2Us9MsYVgvmI+ox8D7JueWSKiAiylcI8wSX6STQWhy+vUcqPWW4+olfVGb
Eh/UpQ+39YMH5Jt5/3w9SzQnnjcRmPTv4SruN836ZxURx+hP8Li3zoB6MzeqYZUt
plO9lIufxBDiSgzpd5AAG+aj61nAdywlvXwuxqkgGV5pV22cmNRdHdXmxniU9Gmh
Jqr/CTYVKdgii16Msv/azdd+gdBeKkcqVR/+YCCW5SIAFCfF5iESDXL44PRxE/p0
o5dMKQUIIadxesjRglgiBrXb3fFYmeqpex9B0H1b+mrD1EBvWdL8DNysEVb9nS+x
2gF4hfR1KF6egc2m5rCPF9l9zOXxe4n14NQvA/7cHD9hYt6TT0cjtaocCT5VnrLx
dkt7TsT93MQCGBwiX9IQLKXT2y72aFp1/J2zguiX0TII9icXU/nkDil2bO9b1vEa
+X+E+ag9eGg+11xccegcRynSTgV/lhSFUL8AiCFQmfLhzr7aZ95Q3kgtoh6zXQi3
wGFEZC7Ne8CO2OttnIC8VSElN76sNCvVk6+mI3uNljAJoSS2+fC2Tkt4nk9pMRy5
MAYqJn/7KCH9UFren18Zl6CkOgTbKhWNfNkevshtt94GkhvHjmJm7QJ12TCgp32z
8DxfXAmHiqUcnoezzBLclGUwjZJwjrtBb8OOA7mn90+6KYrUVV5KVc2ewxEeBlJ7
C2rD48FUAut5etmRH/5KLS7NIeN6I+W+glklIQLE/EV3JQryT9Z5Nqyfe6nT13hL
Ctg/A+2uRG296VAwRpSfGkNMQWEpJ3m0mi4e4/MXH6/kD/2h1jsRLGhEAJqle6w9
vabsNNI+LMBnBxylEL8LPjAydQSHRm0Y5+RnV1FIyw8aQVYRdO5/KTu0KkKSF7YW
pLZm4ON1pQA7nQNMBloNNpRvqGkXWADtbmLspcMuUVNN/PBvuCdmsHe8yn9dXjDa
Fp/vMdEni8BKGa4MZ8pil9AEcZnGLcEQ7nso3hyMjI6EVPovY0ABX9Bc7pglu9gP
zxs3jEfE8lGqiQAwWtsXSU0536H2m3aGL26zY0opDbg2wKErJN/qVaoCOnLwEVqk
La61Lsafv8DW/rjlkJSYrtcKIS+IeVW7lIJ1pnKKOUI0LKVXHL7J8JJ+uj73CEmG
sgaViJspou5WgLXfXTM4AlWe0OcTsoweYS4kyOrKUinG66kPdg1V+mjtw3CCskUf
QBJ3OgfnNLasf0X8wu7Yvb7ZCN7ts4FhV1kPD3PPGUfqOwkWP7nWQ2Sipbepwnr0
3j6HJ7NzLUcvxQNBTkV+MWspt1bJQZYrZohcqi3sL7iiSMjk7f1oj4Jv7ENvloM8
9yHCRqMRKVpFG6xK/svNR6Ngi/ShOVdvgQcy2tAC7N41Fb+3ZtGRA335p65W/VIA
U1vl0Ssmayc1SM3ZMc9C/LDzgUM1WE8hwCyI4zrh5OvHAs2Y90KD1Dmkks+sCsmg
8s8GoO4j0XZwdfesZ9ZucaWzeB/jHoRzpZlsJ8y83ZpdPyTWmvGv4tT4QTy4FtMZ
PRrS+Mweu6YqMDdfqzzXI6uVrnj05e6j3ZRgNgAWreN9nCHjC5Gj/hkARove13Zy
PpyZ3cCnEk0ZvPT/ba9Vn28x3nBO9/Oo8sNhQCRdiHV96T5IhNORR4OvIKhfk+Uk
nPMmZh+GL0tswnhzseVOIj8SxopVOzw1mjN62Au/Nukh7ae4dQt1kFDgVa9QIc2R
PpfJASPoKs335OFGDq0Ogl6tIMzDv0acjLp8KMV1zKlKOhaZm7NtbhccLpqJpCSC
nqKrexhz1q/Yi9hORHT/qbXGfeCEPfBecjCB5h9z88QJNsUnHUtLmNmY1OzE4R+4
lPIUCq7W935YEwqECEYzPVBG3pvRLrsecoWoZhHimJMe2OQtgO7YnfSXIPl/5SoO
datj+sMfkPZEz+6OT1DBg7oCCF/9atYIZGEYD278S1sZqlNm4zFRVKWHgrTmX5Xu
+QUPA75B5SJVyCMmamrpJ9yK8vtf5iNv4pYWUFJqCcvc8HMCzFYHFP/EewGGhYwO
A625sa3HelPl97cgCZmhv0b2iw5/SZz+7oPa/zdh588Tuo2PqGkUT5ziT0EIVNXC
YAPBwFwq6NzIujjzF/+XMwHxRDCj80BL6yAr8cYpfSbyYcWNGECZPg8ZZ3WcJ/PC
p3kXVSAjIZWCmp5o5eQzH2+qjKMEmjLYvqqmtLlYvciPPwl1OJJrqAwysXFfusEy
lGpO0OCh6C6mar5cPk9w/B0/P15rrgJKJCHdSINAKUC+fygL9MoW+G3UDd/LKCe+
O2omjkpPQqTDpA9BdcdRqdt5qwEpt44ehXBtDeq1cOYpU4RXIu9ddZfinvMetzFm
EOVtJmhl3HUY6azhr+lHK8ff1aOIx5cG3I/jPw8MnpYykUj2WrpxBhMLbm0JiIHM
otweuEQwSfwrgO3WqjFcHvJFCvioj9C2pLSrPR/kUdDrILAd0MGNdpgG+MuW/vwm
RCEedZC8fq6koUKMfBQh8IA0Xoyf5jA80S//PPxHtsh2yk3HcXb2PlqEUJovJIuO
1DvsoZT1P2688QAcpdk8gQjwqXh36SKelNzMcxT2ATHPZMOru2MwwSN7exKJa051
znQ8adb/U4ynce/Ot/s2SOSteAYOsyQDTXN6lb/5apj0EbXQwyDYhjOcxZkw3v72
jpiUyIEpGu+S4/HAOJX+woBnqc5naRnlE2PbstrDnvgniCLCa1TCFjp9OwGGcY/z
cFYZRamsRqjvKv+Y/X9fqdqbUMIewg/hYiSfxLugiVkJtseLu4PC+5VIMYxzsZ8K
NA8T0VEMNHgo2sWaejii9D+Ga/n2HPTzOa4o/I2VnNCDtIAwhnC+3hqiyvTAbTkn
RF/FsIu0gsZSCLudITa/gVMK9bmzGivRnZvyd9Je5NY5L/81ROs9G6RTkbzoJ/NB
HP0C5EPGFzeGjqPmmBz24h3nxVTEwHKORuXEny2V/1o2PXawKEP4gMBagK1gMkFG
qjaHWlvvpr4QJjKJ1NnT3jBEStv5ucCCvYSL7tT0CJAZc8KdYlR457T3tE2wGQIV
nv7sWBh/mBLqQTDix1oJzTSXGR0avRJHd2k7+rPObNHPcg0UDKiaeyAAUM50QOkZ
HuTp7/AUe5qLKP9FgFI3eSFh0daNJBqQGcgHekumbBEDLXUh/vqOxI7j7DLj57+H
4Ol0Axxkg3vC09m7dcsw/hjKfdHVtivQ2dH+k1t0crI65gbq4kkIeBlLmLJeDfIt
nAMRxpRRqCJh+w1MDsMQmj5061Z8E2fey40C7KiOM86U3m/T9mFchIKWndHIRrPa
9rhV4iWP7/z0n0/tcCWATqoGXYJ5Xn+QD23cvG3W9zRN4f1Kbf2M/AstcRjnr4We
em4sGsFxAIi4AFE0Z8sDFrUkE1YY83Uimn/xmYPDJ0WMDMNoN8FzldTcxGjYFcox
pZEaazTTRehARjDuhgqHXYkwooRlutdZIDAwpYw7PYIixtrBSLA3/mCEu+VVjy1G
e4+jq9Eu9YJfdI9CIgrYl9+EKDZmY0bxfOoRhfRl5F7Tp2BehyzW/NIfYT5VhTe8
g755lMNAZ/G/Tl2PwZaPC3z1vNEyc8llpce31hFlfzdrZ5I1QaOeJYeX9/4J5L9m
tLU5N9++nLzaoDyVNKQ8VZ4ogqnQk1CadSpu1+9bok5iMIojVZ83K5xRihKk5O9X
QTaXtpG5toEYOSjx6EuXKkHOqPiL0GJcxxfx6KMimKbw+0wob1XHZ5RP3Rnd2HNa
f6eJLF5Pt8BUarNefOy1U/jA5G4iAS5LuMNyB1WljOkniriAbVM74cJ6v4tSTG76
+L3BFOyy5sSW6nSNCWrVmRJ/OneFeM1LE/MMo2bX8npUK3EHMWBQZ2GC/2o5xrNi
xBqy/B2YsfrU+sopCmNSsZYSJt0yieYdvr40lecrqnExQjugtlwglHtts+8UsByB
C/VMpz2pXg5Z846R+MDcEmo00K3GIXlD3GI0XxGVcGjVulUNP0icggLs0R5qFg4O
yk4Rd0fdI4yWHokgAOxkjXI6/w3CHrG789zAF0zWKgQvJVV4JE6a9BGWXfngdE6+
NC8ieFANjCzEk9YeQtPc6UYqIDSbe/tnb98yZY8CTWUGQXkSFEhRSPTt/KVw7B32
4GN7QUgcVtwT/p5qA7FHpWxgM7/NNHr1Sw8yAgvsuRqjApOpx0cdvok8Zl77nyIg
8njHdTx0A3uwFrwUQc+YbfO9YRU3Ww4RBma2E3Ct1k22zJHQSdMzDd9LaWA8UwrW
tzaNwLCTNERTch5mxbXv1vTcE7L6bOrqWJYxuWqqX+Yo5326pFV5W2LNCQGtl8Vw
orVY66gPSi7M8sLq1eH1Zou/v/1TzymfcW7UEgjVST0dmGisdY6ZO8BC+4CCh/lY
H8IBH5c2gNbzspb2kZ4tezOkrBGcUKwRHOpBsiSr3lcrD+MXalg3BDhZalKqKQBk
qJJjsO0i2seBvAp75o9fH9NWGK6FYHIUnzDeGqJrpgYJauaPh7kXMuHP0MFkk19D
U7hgrTqmgAtTMdI09em3zotsgbj3Xxhnp1gSbib7m0Z1FnV9qqpM4UlKb2PMcAZB
+/tNeR8lf5cill+zI4vVDih2F67yb3A626TM1mTUrIo+r9VwhQsWuR+R9a1hCdJO
bsRdfI5VQWOtFjydYH+KhkaW54xv2SaY5Z63sRHIWoKtFMQhNoekligGLNNrCjYN
xa036BTm6Mc1kdUninLrccZz1FMqX/MJGfoAMpu/4TDeo2TF3hL/6hMM9X3/Pr27
I0hGI0eoxkaqurR98fNl39SAcBs4PbHBDGxCGoMIC1MpZpkENX+VYKzhziaVd3ct
1SgCcvgmp2fsl/+wMeNgfsU/5T+9t55gABhpwU7P208m3u00zWK/zh2dwXemRLIc
EMNGMxKl8yb5Xfjg+CfU0UeVbVuFfB7bv0rq9WTfTnH64fTEUOc2/m04n211SE7D
lTbqXDV0OGHZwJ0jtHMOwtOPJyiHeUydWHS72fvqbO101luC89FjNK3YFfXFKqtw
aiaa2rbKR5gASTkBaiOmnpVn/O7yCQdmsPGZ/GjXXERk1W0oB8M5N2kLIxDG0zhL
HADUwTqbPBeh8iE77ZxHLIDxH8v1obycWjv0FS1M+VPoqZL4QEmPh4i+95JRnj9v
qeck5+6pnth5IRGqbz0Kdf0kAlkdzAz6z+POV6EI45p+/gVLs15zUbxlbKklMLui
yIYpEqYUtwAeCLRfeLqo6kT24+GCaq5vcVw3FwTAmW7gG36W7Pmd7H6bnfaI09kt
sHdGn1NlEO1vYjwzxFduI9D/G7SVBkO4wVlripqdxBEPL147ul2BOfEUVS/YTSnG
W4GIMk/W5TTYmrOFjiKnnetqpXmbl6Hpf/QqEIUyqQgEZ8zfheG6gnw9Du902gyf
33mzUmNH9bqXoUm1+AdJyWXdDqlltIOQuso8c2l28cEDEzwXqGPboqkZsoB0jTZ8
tj1iSOx2ksX9vEC7+jApFPjE1jwXRgLXBILCN8/6C/qmzGpzAfymDdK/NZYdbmgV
zDJVetxq9NdOGW06nlBOD4SdCs7gFbJfTJu0GbJmAldBbHT9BljkTvoEPpNiYpvl
PBem/LGLL4iVexN02YVXgf0MpHExXn/y7TDQDZhLnR+dZSZDLOvBB0ypRjMX8qIV
WT6OxG3cZL0WxkGKSmH83wSmjtSSrPl8sDbJxK47LdnppjpXuc8Wr9Np+lf5wJUM
RxJwq/L/OxaJJc4rv261dHKX0zhRHoTdMPxpgKRZfuhQJKIvM6wU3+ZVP+R9Jv23
SHgNgFQZvMZl7XCYncnW/WEZxH807Rh77OObYLaIBhR2zwENoVDnTNt0jotA2yb3
KRG4g1r7wIdJspfohZjcRmpg20/QhxCAMNJ6mh8We7Ost3XbZ2JTcBZmpIpVkjLy
nf0K7jLhwcMCwYUCW97gw+rrQFhpToMDLAvV0Q9wRS+f/CyG749w6uBnWOPK0jXL
LCybtpyDPYHk+Ruuj5a2KDd3VTWxtrKi7yN6qwBvl/KOiCSSctTZe2lLx5NAqyql
k+ho359ghtIwEZJaHVE0BZPCi+OnWnX1ISzXXXuU1ICChDUUW1VH+erCmiVkCTXU
6PP8ZwRp2peoeADyc3pLbeqdDvm0uuvM0qwRkq9gm3imYnCVRPsKgFbDePoXzYp8
xgKaGW9DakqcssMKGUpNlBr4O8aSaikiu84DqqeoZEynlOozjCbUtiMO0tGrsl2x
h/6rvDdL5AqvIlBeHmz5j/qFAM1MSYwKtDf/CCl3iJEhxLMZMyC48tzTedDAWmBy
nIiKIleIp6VMnNU84pNDrZaF8MX1c9aSbXp8cOmHRjyTgIP8FfWpoGfiQSMoKtjW
NxcTJBorNSDMgXzMFT/1P7O6Y8L9elYPFnsLONRA4C+YJx7l0ja800FKt0XHt/ab
EnWCXvWTn5BQQ9KBWaI1wmESuAwQ5EpzGwx+NPD066oRuSuacXFbb17PmyDNuL0W
kwsSFs0y6ZCdsJzV78F39unecHzqiw8+3QznRHIdpemB4Lk7KFLQkiyL5bM40gBD
FdyKjvZ/RU/DKjCw9MzvCLv/5bXmt+bNDqTWLkXxyN66fzcWyRLrdka8YBp05Edm
MxfrG6fQVlaCZJLmlMRv25vSPmh6aHFmfDTlS8GDFAMra+JdHe8JfD31SMlzq/Hx
7AQ/x4H3suy8dmGVsKhFdamysXkv+ByswzaxeoHSq0J1MEol3FobQ99Wws/Td6g0
l1TfagjTcUn/0PIK5t6q3KCixZ9yHj8RX5yOxyvlo0SbAyoMIg46FET4PrQFI8JQ
2wMYaFi26CInOcRjpV1wPuV1vIHNXK9GStHNh7XBXb9AE1Sui8ptrKgljoFQNyHp
vWu8+FosLpauNeFRGgFdzNQwTqzWkiW7UNHEELGTtJRQ/RbdtlaMsk+/Eu2M1dr8
jJcHpZlMkJYSUKRvH4DqI/O0XBODjpFxxWPZS173RUP82b0yr/erQxnQDkQt+YnC
39BnQePihDyQ514OwBB7NBLeG3UNnz/1uPaEAcbRHgEDdkXSzRYGLSOvbxpFxUg3
jNnIbcEplrRFbiw0lwvv+XqpjRx5G96VAxAWKo2Afn7E5igXoiwybDA1hlYN6cX9
PLOVv0Nfm6Jz30vpAQ6PNfXUH0es7YqzW0qkknGRQ+KDPT4+Za5pAZJwg7ijL9lQ
paGNRULTsnS5AGN4/Q32orXxhxX8fVQrifFqA+meFC9pVs/JG1w/2g2FpLsO8ArD
D3448XSGL78Co8lCq/v5kzdxN+vGlQpBc2VNUjyKzybA3+clcAzJgKPfgAzZaGEF
eGZ+aCVMIUPPP1mwaemhX3m9ZCgyCOhWjiVFlnnlO/XaEVR2Y7rgtVRlPaKr2JXE
CLrIZXZnYd3qlAzb1ZqGGE7KadiT1PeL/G7DDtrh5fSGYmUKIRhvSSwAejjvxXUZ
rVCHaeF7n23X83Mst+r+GvkooKq/kjG9WvbEpQsodfzybJ9LZaNSnAoNo+Sq/k9j
ZtRaNfXeSmT4pxFwA1VxoXLVMvAt4hOi/5ZZE4MKj7S3hgXfiDhb97l4DplssSig
CMHhm2a8TP+UMsvjDEsOGmzrfRvDqb9fsk3tt4R/mygK77jQZmbqtYEqFmOFDKJs
qsUS2tDNGY4z3eCfHszp0iiHktQuAGqOr8Wng1obrFAIvY2npm0CZcwrgMWh1CVl
2k6tQWC4UkJkVO62M9mb2UhFzfELELqAqmZJBwipqS1RCE9E0/y6YOMuanDP/qgj
kwxZ1GMGiWH+wLxY4ahWCxnK/zV7HiHjOUzBoc6dZ5kUyYvOkzar7Q+fj1dnN0Ra
gNOf1WPXhCFyMdbujQXP69I7WW8r2QN6b3Mfgdyv/iWf466NTZw3ob7a5JvNdCxZ
ixETKmS73j9hZcfqMmk7NkPBZGT57SAHztxioqDEGQkE3FYgykSeZqdlbQHGaVi8
Cu9rXD9ECXWF5E/LYBPbW1cIUDjC+6j2wAnUFolI4p/qJTFtfBThnlccfGgc/SXD
7LRhLgDoCqI1VChZerE353BMdyd0l9/YR53V37L9YskNQDbzgyESjZHHBE7ACdyq
X0mzuLpXbJ39EV5T7bSLuIFS/UxHJPcGZOHgQvN3VVjXvGXeV0u4YBJLRhPogS6F
yv1yH3n4suagL3X0F/+SRc4uz3O2SAb7qYjjTDX/o0h3jfJ7I73vMl3bhWUqN8Lf
ifuS9wJqMOE6fNnbMVOOvRqvAGDRDRL3oRmRYKPWvfFNJNQKcrrdJuHV9NTOaiRt
U8MQUXr0I329RwDqKz9hhbC16E/bSMO0AupmwlkRnCCwh5UD/+v3Zy5l1PYgx3w1
LIWPcnv4zjNkKxYaJ5Xfhd20m4wTvo1TkDSzQ2OzIlVIEPf7Yks9T9AX/EWgF5f8
rFJBqRcOjnAAdnE/vXL/2Z9dvjYliPVpMnfQPR7CkCghwGMNvtVe6FPXTbODIq5J
5+Twz4RbPTnIsVMAAeZ0buMHlpFND4MnsbFNgUKmWzLMJ0ZguJSa5n8YhH7jMHsD
F4vqutwur3ggQFFwt2/sEsjzkA520cj6hUBOpcJMwQNq8+Bs50+aXqKbjWcApX3w
g3vPuSF/PP96TQmGrhksXoTzwrVwCoCztNaUINtYGPWFbixhZ2y5KxwrhTr98m87
v4fEbGmP1NkQjcHylD6DuPHVpXWqXYuyx3wObdY+x9TQuzA8KxNwqmH4y4Fl4sey
NJWEz68bFHc47jW9zJivsGvt8a66IQH/viAgiMuXtHcSmfSaU0W+fItUiqThQoAy
DEa0t++vuz+vT312jazllbTp1nVQiBr9DeNHfNkN95MqCsR+YmdPbOwDywdEpqZ7
kXCKw5zXWhmpTKoX/jMWmnZmdS7cKI4I8SZCXTMRTlNoz/FxjjVI15JyBiSsEqjK
YsfiGs+cryrxHCAUa9Viirsk0YmN6zF6T5t1rX1AdHxokeL49NW2X84yMSayH7yM
sqH1Ih4gJGmTwLclDmWUIsexk15P7zCSaRS8yZENqG5RMOTsDIj1KGpVsvqv646o
64IuIyPjifKt6Md5X4SVHFIb61E43wkm+d7NpVToQ1sZWsDsG9xMjZ9tvb6DLreP
t8znkqT26vv6TGqwtaIXwI/vJSwLHu31uC5W0TVb+GTBTHopovcaXbVwfZ7P4zuE
AB/aIndjUFqD2klT2NzYNQ8hf6zec1FfON5lkf/394tz7zBDMZp031XxAIUopk/2
rdbDpn4mHsB4VvRRjtcAmC/gufjcDXIl/8WhNKSQIigRJQRoKFiFj1dFxSXu8U61
npqyRvabGDR07veq8p7zJercYA40K24gL+1ShaCHgay0yw2vq38cJPRsYyovq72g
fxDwDDdbejl4KBsDbL9WXGT6YWe6WEwKeO6BQFwHs5lcNTd7yT875fG1SYu1DK09
9LJm10WuMi1rVgfdbKqfSukvHkF+/njjYNhQNE2DRLJmqdSiOng5EM9zA0NnrAZK
XE0KqjuXv4z4zKWmYYhgfGjwpZhV9nbR99cFN2+TH4RyL86vMwoUNmPXx7NMFDYl
ueNGqKORRNZ6Xm9HuJPUmtnh+BTxU9wViifHSxbpbaPhCPVI/aDkOMK+xYTn6M7Z
hgLf4W/EgEWD+2O1MS/9wrL3udTCxU4gLu59J7+etD5BX9TJAT+E6fflHe+oNphS
daNbLobqTGBT09TahMYg+8f1pu0mAp5H3ytyfYGUB6fpXSHCijj05AGzw7PHT2Fb
e4itoX3/1qBvH9vHEjX7/xNcaLowq6EIlhdVR0FCdHSV9KCb+9eqou/FhIKKDNBv
wmd0KqtBI9xSuVhId8gX3c7hy0RXbXfd5x9KHdJouPWYXtieapfr/fiewTsls6NV
d8ewvtJBQK918NfyMOHm5Tl3yl/0ftdmWSWy32XakoIqiAzUtBOXF5VCzrkj7tsR
Bone/uYPFOkyeaP8pPTW3Xh8Mnid5ZoE547qFIWu0jbIaAgwKnXFHxohP4P4NkCh
IbstfMzegV0BeQIXTHf5SLKYHBLCCZ+VUYiD9ycOLwDf0xZc+n8tL9xqJqCOXRaF
CLPtOTWn49dnXaUrCleFP8Qezrf/+ymgEHYmz+VtAenXwp9JrAZWUW2zQAgewBH4
QJCJaFHBFVaeChkm1SaXSQsvwXrz07oOzryR1zLso+8suGYV9M86irv8E6WhVqaw
YKK4L0YO97KAIMPWmp5z0JXi22A08MwbVJWCGXO5K/XzNvpndOVxtzq93OY7PnQC
+C/LRQKal6EhnFJKwkVNJZ8Ebq6ZwsgKG3UrtVm8fpKfwYw672wlKfiDD19zMEUj
Eg17Evn6cahhjo1E4EKqGDyY1quCjoDx+J77OFczasCuIfwUrHxJ1KJzCOZ3FDRf
vDWJ5KB78Crc7I3QM50C8ycI3DtymcZ6LQdlCbVB/7JQEmS1yEnPKMLjUcRH9vSR
m2kiqjOm2DYCbbVOpYY3DSCaBe/0Rnri3RZ3RpjxS3GUDvmyGmuZTpDAUaQvssnk
pp5GLMwmFQwKQ3c7xoIrMyQA96a0Jx8sPHbQKJEGhiALAhEATZgyBF4YQDcsuef7
Tm+xQJ0P3R3DoCqppmSwxik70Ah+AUQvQaeZ9cnpZKSQAehJ04eTKuUHYzfGlJX8
HsoCo60328YHWyN9Lcv/+wOIGvhD4S54u+4YWGkO9T1U4D3rI54M3NwQ7ELuf+4S
Sv3GIzFx6am7cBOU/A+wt0NAyRd8A20XkNcVq0PUH9wSxKDLGscRJMe8JDj+tcUI
qARwXa4Wd7+QvAOY5G9jdwm5v7FCq7NglzT3LtofPQg/RJIoLZ8bexLkHXci6YBn
gzLIW97q9UH+s6HsBnsCidgxZY0wbGLMG+Lhu2472CecI2ltHy4+EIBZMQKz4NNT
l6fe5kQEcCTnCKt0Wkcw9TrfdDWBbR4EHl3x+vfV16CxBF4VPqe/voJc6STYj9qu
IDePdvWiA2Uq+D9q/HRIIUFH3Q3nTTqQtj3mMFBW2hxc71MIazEXOYm/2oVLjrBT
SVMz+nDBsL36xRioxrgQh1k/LW9uiyGwKpvtas+hNy9hBvqIXE0KkCfZoxl5xjqV
uK0z5YlmFz2ANecyk8I6nNrH8y0wcXUORZOuOQsGfedxrrTu3ILK2qGgtoQsYKyd
rhl8o1K70DTM9BTi/5V7PS1c0oYbvzTKm1ll6f6ojg3reFqpnoIssfwLG8svhd+G
we765zdWKAt7Z8whFcqcWrCub7RyA4pY4XAM7Vv10yzj9c/36ikpLLRqMSYDXJqx
bEB5n4NMbgk1VcIsMcCwTKakgMYIPbUCnfHkZP8+EoC1gv1NabBdIBmJp0hICGx3
w14jhhbGBMfvAJvs9HLO7x3SsyZi9FVw7pBMk8IU2i2eyn/TMaPQqIgUXbBTFFKu
1dCCjB823xD3qRZumBxr+VzC0ZK86FvkPXnuve965wJDtNe4+p8hcp48bM2Utix7
t3rU/dTAhW9hZXW9FupalfGPbAgdTs2m6lqUnnfLolGK7D0kdJ1yf1K6ywWAX/m/
HDPk4+G7XGIvSyZjgbB7kqaQkQmNgIyLlwWZKoD7Y6e0IhvWXPyA/aahtnj+o91r
GaZYOyAX5NtMLJ7BIm22X5b4A2srJw8QHKBpgUF5EHbU4Ifw+l0PrmCzpsVkjqKE
69XcEMNDlgA7RX7oHA2MHlr3F/SeuicKHxqX7pM4vr+y1fN695a09kmv7ks29WR9
ISPAhl1GRw6mL4J5UNa1ZPa36E6hjlikh5jlEBY1g8XnmydBTTVrJlq7nB5h9j4w
j5Az6JG3iRwVcvzyPeH6CTSzON9XpAw1pyLkrCM+6Z8BDjhmR0TNMX/gGtbM2T1K
/9XnLCgPC6wRv3ZdOOWpe1bajT3HNnNSs3L5GUN6p+7a22Pl5Tw+hYpjEgjXRFwu
vxwlOl0VJ2zJSzW063BfSN38Ej7eL5p+nDBQMmC/iX4=
`protect end_protected
