-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
BRm3WJpSRSdcLL51Ws6stI9iHwjXpNgn8jfqYANT0J1fW7hWJlMAwWdN5ifIuyTr
y8gr09gcqSBgcxWTQ80xANDlJ9FKLJ3lrXs1mYkjiaPFKWvZbLjWcgFIkV727M+f
QUTiM3DPeZ6kzBO4xXuHqn9VzCz9KxrMh5weqKlIhK9qFv9oNu4UIg==
--pragma protect end_key_block
--pragma protect digest_block
PBDlxaFqFadWguqMaEU4L1d9xy8=
--pragma protect end_digest_block
--pragma protect data_block
wxJlmlIe2VBXZ7RDb4tHFGXNESUEwYrtmceMxX6utCVwe2dImbFVm0pB6R84eOrz
oW4fsG4aTnBd0W7Y0SqoK+zuPQ1bjWBd7xhxj9ABK5qi7Gb7wM4UjSxIAHgn5Cp/
9BeWJ6zYkfft2bqP7y2XAUr+CDwFyvm/npdUVm6K0nRsyrCdS1Jc9FDuPlLslHTl
DV6DTPhY17+rvuDet6Vhr3CqhO8F8mzh5KQvOyNKa8TSqv5ut8KZQs+Gg3FIW4NU
D01DN1rUuOcJpkYTb824gw4V3EirDU6Gtb2N0cJfIdvYxHiXiXy0y+z76iFGNzOs
GKqW1M6trp0MDWky70pVl+FLIRkzB/AO2WCpBoQ0vIYTfRJnFbETBmmQDEFAKuOY
kQBprERAbFRt6fIZsvnW5010w5Tby34n47/TojNGHhG1G8xTojKdkEBecF8B7Y9r
nvXcnq51M45x2f29M5cS3QqGFFJjSfd9rD+SwsYLiJDlfYbWpU0x6rNvDT12Ogwx
MhNCHJuq5RQQyV+mWINmABY577VH4dtUekHu4/XbgbpfwNm5uDlDfklH8J2+iV7O
N0oXauXSc+SgIdgeREoMSlpTVdL/304HbKj1y4pQPBxS8C0CB2uqo/4Vzg8mcZSy
PKq1e6RxO/7DUoy50MqmGyO1Btb+VG7YmDC/K/uuumGOjklVfJFsr+KjL6We6abo
HDkBRJt3PdZ6+oVRnU6gLStS7q+m2zm1AYEin5B3otYwKkIIEEuVdeSQS0dA7upv
lS+7unxigeoG6meUfkREzzDHZUmB5oTJkfVjRwk5h/Kp3WrGNSVmiMZRiNhe6QIA
ZAzZw4jPjTjPsQHAbgEyZmtjWeCgDuLFnJkqUqiKX6X4CEqSzGxaDDlg34Wb6KaN
vS9mzQbT0biJDTzRh1g0Uw/XihJw45DrSSLKi5H7k3K/TmsqhLBF98zWYMHonK/8
hdRYnrpVoYhH0LtY9KIZg7QQeuizWmpzbTfRZ8ocgO5u0uWDYTuZod+eq6FMRil6
lhtWUKlwmE5OtASj2zn6dX3s/8nTtnkRFTJGQjzXw1z0jFFLq0mf46sRSdh7VsJs
BjSjG+21VDIXwoYnn2Z2dK1O3q3jJW2alNJ9u1eBDilb3gxXWgdJp0B6i4f/MqNO
zOoXxKFBjm/iB1hhhmj0zBVYcXsir0AJxF17rTTZjyV1b5EafHu11O8saeTGD2t0
mzS66VK8BicAOLE6plzF5pf+XgKjHyGhbImezdW0kGeDw/da1pqnPXXK9XSk8u/M
VBeqXuttoP1DxXpi50jDCTxK4JkDtBbQ6ouYhyEMETG3HuL8IIN8nWTK62P+fBFi
7pdDsNwe5A5Ppgri/AFWVaTnbKWJKchDS3knaqA81C5ZtFdwrAYoaWZ5LFeK1+Ud
D5psokiUN3y7HSpjNqnXF8YQ5TXDI5058TbmRKwVSaoUmLKx8Ag7nLvj0hbHK9DL
yDHmvaAzWD14ZnCrA+7COZ+rKtuDsgc8wkjkaXbiTR/6WeTkbwQmYYaJdMiES2IP
ova8kibyU3TAJMZXe07MZDjGZqhAMEq95+AVBaY74OueanI2j3aMnHpLgvXFEflr
pN44t/RbvIXCpAu6HtRl4LxtlFdak8KFcVX0+ArYrXSGDqaLngTq3J6fzaMXZ2i9
bZPtQ845GkvFLClF18nIecOFB9yVo5+aUunDAwAmq2ArDCy2au+dcFWwjcEDukwO
wd68f4EWNdguEDymIhI8VqUzoKJTjJYf24jFC1dKj//2z0AMnWO+Y4vCDizmh5c2
4CoFOrNly6icbUhtVu/571PvN5tRP20l92KMr0C2mOkyDk5liyrF9MegC9XmrpAP
e+Ud7bZvQMV1RGy0RmP27Yhn7Wk15hl2Y+spQlAQBfNSMLMqXjy4lyezUrkbq1hH
l1eBP8Z5HS/MoyhR4K3dFKy6ZkEoACOmtlPiVxL9zBFmxDGELn31hL/liDGbJTty
EM8tchwGaU1SViqZzHD+qMPeVT3a7aD0LZBAheS78GwJxtfK51HUmPAWYLO60qe4
OEANrCsozfLepcwFePAhDuNUQjMjiIYnrRZh+zLMc5lYVm/qezXl8v9yrXav5dAg
+Jsh6Rice6Zds4cejBUT6GE8opzjLzn+jMuX8MjqJD1N8/egMilCOx1nTR/tDPDI
iqQWISUG7Uu7nnfACTBQCsJKRwnGS0Ptru5Y/s+5qsJ/D8T/c33pD3LAI5in9nBr
EAftR2TIKT+prq4krt+YTHbcJzMUaeeOAx6lATmNftCQc/eJbgOHbpFE0uco+SfE
/qcBsPOTH+dqATCG6OAvqJbPo8buLti/w16OFGlBMZI+q6E9piymhBFLqaf/wWuj
wd4eaxsXp9xejj0ON8GwhYmlvBYnFlU8XpqaDwxZTizRq6S3pA05DnGfaWwaaQe1
xIDB0NsTNCZ59mCq5BHm7fAOHuGGBtpX8bLGqoya0wz6nYcd/N2+AWpWPQ91f6qL
B6TRFELbrlQHb8WtlPrlNgKsNyqaXAsGhjEScs4ktNpvllbCRucxThw4Rluay3j+
2Z985FVneNEvsYQoRn+brnLz9RhpzN+YNzFH2icMgO2yQlFFDojgIaXmIHBzyrm6
yAzFNwOeNTIOJs/jY3Z4tmSw72pmc3dxCFiHjzFMVEA9oIA2CsP5AO3Gczb3+WPi
NBuKxdD7SjW7rIYIzGypYM7BlB4Ahr4nyy+fOgZi9SRdPvc9g4+MRaM38P9cZPmk
3KW4ZcA04R15rOOvGf9tjCqY8aPFH/1sLQiDq8YEcW9iVfwVzhdYZOd3PvVa578L
8nMcJVskIfPHkaBJjSO2RNICP0CfxHPs7IFAkdZCQf2v9JkYR5lE0dKeoIQgLdyu
vOVa6HJ1yMmzJy/HW1p7/6L/wElqCjr4ULknH9ZVrce167VjcT9UCZjK0a9DFYM3
srgKgb2caOzX0bML2fY8EZEhkmHhpqrhBE6Nn6YJs2BCVEDbEotd6fljSNMjYv1j
7UoR5fh4iXdLU5ESBEhPrliA0s3O5uOntOA64wg/YpUM8mD+BopqGbGF+J8HECu6
wkUKlC2Lo/CvqwfDGnY1SLvPbE/ibMBRSylDofN16bB5NBP935Jh4UEqnyfwu62z
QCntq38JTGPAr/xGYlavosJkjLXWfqjcPvPOrrTQwKHOgUDLjTgbKP7BZwZSftb5
1au1chkxY8RZbBLbIpXqZw1/5hedZesTBvPFJOj0HJGIa/nPJCCNcCXLkERkm90R
S9kmhm+E1M+dbSSBer2iZZzXnVRPz1wv9z5XV4g3LXAaMLnEcw0S0KvqOUf3Zw8M
XDmJM959F0m/YZpkanBv+7MIvv60XjPnFULd4HktmXgy7UqOk+pOv9gfuMn5ftc7
IQGVDFsjfOs2ZNjKTnI6PduYiTzMLdXar+bguPf0Gf5TMH5LHdv+vJmSk0Uyrv8A
DGZB26CBqAJldGSNp9cb0+2FD38f1HKNh6RAwu1vEegENu6jXm38kPYUX0/XLmYr
tkNIHuohfYkgtNqW5JHVcgwj1sDPJeBU06Eoz2rkAYxXjGVUZGzqwIOMEWA6kVvH
S+k/89n3Nf+pQXwZJ78y+xpoai6uP7GxmG6EIfx+W4iPyCR6Ngh8Gc+8uOn/we69
jrv05f+odypx0Tyj1nklLkoHvQiM3qG0rjAmQWq/qImDVT+bgEsaGYTgxcy9rHid
BXJaiyJMRW9oOitZeuK3lfHj22XvT6NdRY+Fv+VQZlCVM1MLdbVeFoWjTTp+z+jt
M5oedv5yM5iI9UFT5PL72oJn7lmqIXjj2VQSPaJFNorzCoVhzf38c2zMl5TIHJU4
EGJujGaEVciHI+52ZAc/Ovxq56Io+BsokFh1y+C6KsNjeV0JCff8ylIyJd0Evbwn
pHK11AMTsL8cbtekbhLEXPLbVraTgTJBMYFrSH0+YRjtSdBg+fLUrWLxOb4uI+eb
dZ5Sy2TglECwh5we8GPOd0TefE860+MgXndGt2n+wTetW0hhmhr0DEQWMLlnAu6j
pM+w+QPqifCRwSva+Z7fPCseosj9J3yhcdcIjIXd7cblAeC+rfmTj34Izr2bOmEh
eeGgcv3A6NZ2QRATxvCeAie63MVL9oq40BCn61r8ovijUqa9Rej4ex79G2SXaasg
ojavamJaLbLT4eneAvtbUkjPe+3vGr+jm0aprrwbftyYhkOKul48n+rsoMJvvEUj
20088c6BljZVGEJSWXCwoZJmiEb8e1h36kmcsWyKYGuKAAQU118gBY+NnjwyIBy7
8HDtKOsLfGiHAc951+WXXr60RF0lAY49YSR8KAAPxUEtV2vMH6OpUYOn/R6zto8s
6VCl4MVg87E8La2ocuTFsR3DjYDwHZ8fQRQj8Kb7AvMS+N8zkrvj2UfHoLx+PrFJ
2S10dAOv2oH8WnkrsBYDlJ7K9KxqB2WCgkxqlo5oLdmdVNSfMOndOb4vO6YEhN01
dm/oOFiH7lRNzHjYMXTDSZrjkDPimNdLlFC8OdypwcGDhQ14ZtC/xrvmSxJsZPrj
nyepWvySvZvb7KbZ/IHSdj6opwQ14tIk0156Nyqi3UcFIW0f0rMhEmHBMEnwvkdv
/GBQlvcUQkuJeo+Nl4xAPPQ4DJDKctI6qmYN8p6/g8fF2EtJv3kez8pMI1VR029f
h2Ad+NK1WOKvbE5S6CtdqC3RaTPTvjkxsZIutwv7Ip/uu67LZ+o/yboHlB8PUbwx
f0kt/cCjrzzaSPDGO1fxtGTP881Q5BH2TofYJ0t2rW4HhKW7RbZWewhohwjj/Yv4
snVksCoV2FGBg5eodrVjEbIEhPn4dWvNIGUQ4REwGxjyCKtXdycxlvcH/0C19cfV
9axZRYfo7Xd0MA9MrZ89uao4ynKyv/WWamb/FNoJ8PUDuFW7k/cuTIAEHEwQcus9
IZPQ+lV6Wrbj4GFpEB4TrAJO1zY4aEmLmEkUEX3d50scTDFjRVDEvafaJ7RBs7k1
4VKh39mjuN+wkiPNRQSdDvaMiARSXxhLxz88BxUWuK+HwaQn3PRaSQZlwzB3UVI6
3A2fTRS/vgZ/cUWUiY8Xvk6m+zBZ70k7Kwdw1JbvuhiARYUEYfzY9VrqUIFyDcvH
zG9Dc2WH9hZHDEDbzO59jqXLriuHYIrckp05526NB9WTZuoU4CAse8PM7/D5v44O
ZGP9DeuIa41gmJ6jZLSBr68DgM0yb9QAUgDDBGWO52H9DLfJKTLtKGkiqoZrPcL2
IIvCKxcFbKmd4X9MCUEC6b0h2oNDCE+NAst8Gs3NxYyKveAFoc4xT7T0IAT3t5OH
rGNcVUgx4KWmAIOEFr6v2/C6lfEU5vq4hpOMnkGRWVA3UANgwdYMXt/0dhCDSokw
F/RUecBgYFQ4i1+8+4bRLjlce1yxsptZzdEWOC+aYv8vNRplO5vIX4Am/76tf1Kd
8YMIZ/W15V3LkqoDxHdyH/pCTBwHJKCGaCTRWjyZ+1o4DKRS3iIcwdvsFKeIMgEJ
oRn6Fq2l6FsQPNYJWWJ3/C+UURGhZ0aS0qNf+sETrr5sdyMN7TFU0hzsYqeS/ywG
cDqA+k/aSTOFkEwFsa8VSFfuJbHnfRwJHxBHc8U9UfBLFeR3/Xg6alw6gYvdTcHy
Zj1h5qw0VNguTbrOAl28APxNHrZetPkxRzQJhgeiGWPzuQ9NqK0ivLiTOP/wxVZE
GVfEEwpmdHAah53U0pSn0xItdgs3TfAKlLBvRJsVXzSY1ilYxD5dO8DeW/qvrN1o
u8P5G52M8XS983MW/PG/yRn8PEYmKlh/g1WL6v/Yg2bAH3+iD3CMcP8684AZp5W7
wfKxNFfyoi92dWp+VA6yM6SaYYTbMTxtPxgxkDw6KqRbDFbFDoJ+dI/ksgyAbkzj
LnJwEq/8SsURulHYARbyyT5GF16XFUZofDQ9j7Z1lgyj7LHITq8No2ZSpOcZOLOK
S/JL53fVV7PCrDMspljNra5ycdndlBX7DvPS8HeQB+mJs9lX1UUu0C6trpuAeM+A
VHWQVb22bngLnEAxALk+Lj/2nr6N9WcmTk01tB6y6THy08Lam4MVujP1RzLn5HZ0
F3y/BIwCSiqz5Rl0VW8n+3xy257JI5GkP2bHdbi+TSa2uuHAEq4L1y01hg4tLyE4
/swSEdKroAByUYJIQopAe75EuUfdhi0qmqVpaA/ZH+/6I5BIj/XJgg1YNSXz7Uwt
SJ8jeBetMucBPp6/G3rp++q2uSKxE7dpUcgybgnyVYd4+9UMr6OC1BTYCQSek4Sp
pbiloOqjZy+kDnBGDkolK4MyEtX5RaLnzIR9A9cFh1hSoW0Ve5jCn3Wm9pGogPYC
O+JV745MJ1CZV4sAbvi7Agiv72bwXHCxsgXIkjeJw1UtSGikq1GB6S6Hhma73Jv2
jHMuDLERv7GFD2F4z3grhwgS6580c8clspmW7gqRsS14RbFlrrBT/uWugTkEE7fs
vcEQVOnsmBBVLBkCDuMFXB/vCLX+mfN0L9w7eViuFMKD2Dt7LLoCw4wlm8s+kBLi
QmkLQ/TtMahzxOaTmw8hWZy73kw2XaEOIR01mld3Qt86Xvtyzx7czSIHhvke/YjH
NZScxio0coNQe/8prQhpfEioN6vExo/tDevLM9I8VEMYmycsWs6b+qhgHf8JccsO
rR8HDvXsd13wyK29W65bKK8GJmXeUSrDW8GtdqcbmCkaiiez0XjwBRFz3YSJeM6P
p+asA4AEB4cH8lVdpnQvOv239pkDOXK6MrDvE9jPHncwdFZV9JTALJ9xcvHJnZ3S
XBmz6SIrQV8+BY/+ZOpdfRYucCNvQaJSvQvsaxXesHsikxNOZOnwCNyz+i48sgEB
VItnUP4RU1Yl1VoZgkTZTJCFZLKzQxxhPU9mWmd9DlhvTHrNOheHrE8JYFCYZ1Xx
a07LznO1LQVH84K3HzqliRFFddPTFrW0Qts1Khc3nZbbEn8tBcOb2cUkbfLdAn6k
CHFGR+bzHuF8LmlK4j59d3SlqOjnHaUJ1shNpFl+IhGpI11DBqIacYg8UWVISx2y
U3QuUMezLY+WSO5T6byGftpvi5i5DHk8VM0bcMS249RXl553l9r5sWTEBdTre1u5
EtpzCA/HxicsOIhtX43vg+TGXYcVpzryTWwihqsJQbaf0aticMIfs1nIhPLEEedP
OL81cq3E887Mb0nZ1S4qYQL3lWh23pwFHBbsPbsQ+Db+YukMnE/aK71LruF4YK8x
X3VaD2+4G2H8M/iKlV1Diaj0BSwFCzx50uUpsSUnFPaEGslJQyV49biwYLX/HjQV
FgU+x01PbDJwmW4JRRPWbgR7n/znpkHbBdctldVnHCtqvQDkt18LauSTqnNQR9pb
wKSvkUZgLRK18fY2xcgpB1XtWLlB9/ZEXxsoo8zZBYN9ROz3tgbu32MARJlyzDvX
wmmC2Zgbkhm44LrJ9WirDwYQkhf+4J01UZGumZscIvi5rD/deQdyG9pkPsRP0VmK
v5TVN4NcQvsj6aCLw59f1K/qm6vKIdfDmn0qFeaona5An7s2CGgFgm/U2KJNuHM2
paVFyomdH+Icrb3m5Yv+FAfVgyHcoCBW341efq+TKXRO9fNMffrV3/tlCxQ0qi6A
5gL596SV3zjIlU7awrmueUpWX6jWv9jhHASeUL0QJ/EohJwlEf3FK+8Ay7gTmyVJ
KWlE90JEgoZPlXH8CePj6/BAXmfpQboiB0xEodseWzPH6RwSV4zCnb+bbxC/b842
t1eFDZj/xhXnSHLZJQeWmBLnoRAq+TBgGTAm1I7S+24b59O9phvN8I40fq2Gesq3
KAV52IJyG27Uoxnk5Rr8ydUGSbzMHVn0tKtUhlh/7TH019LKGMvpgU6njgHJBw8g
2dgCOtxIPqjhJfYnKHPaoZoAldJH9Gewg7ZtmhMnOfW1Gsqkr/pieb1aDLGrLXed
8NeC6VIjMg58O7WZ7Va12FtZUpFVSDBN1Wm36/s0Fj9NPbXvXpSZdVvH93ov80hc
VkoQWPHGxWwHHJVkWfCqR91eCehjmrcw89xi/Eb/A6eaBujNDf2YhEzQHiAoDxTD
Y9LvujefAfjCR+TGICzLUTvSNR/Uo/YgukVO4hza+bjPzn+7OEDWcvhgpp1VxP38
5F52brtghWau5PKOACYfOOr9Ymg0Pe6iqg5MaNbB3F3Qxw/ZLbcAxVHdYZ86yAYR
YJMTc/E+vLScpSzCpone8q7//4LYa6EBksTkRw/lHMze67CjG3r56Sgrfv0XuGsq
OjpQlgPCAD6Cq36JTpp7Ef5eCdHIWVP+MU0Nn3v+CXH0COg/njUVfZ3xP5S+h03A
D7V7N+7JgnEiE4xM2uMEmuzUx2kv1yr0XVmudp9gCO7R4FJB0luUI8yAMPPYoAc7
x1B0iiOFgah1DeBLGKaHHqFpXP/K6TcY2fhjKFqvWC1ULTxW4XpJil/7DbNl84p7
fb70JTXRr/ohIl0ywhHYu3g+AJhm9s704U2oyARAdX5AiIhuSBL2wBiQxxbtT4zD
HVdXRfn1UIBfzc3UHtZVITbJYFsIbg0hpaYvtYwuduqspXpB7xkRI6bBXliVots2
3tZozmyCjBDqmrse8JHgDqcgM3lHDKX1zGj21dR7UL0LfMEUVe64XR5GU/cWacO1
8BjIE8j3ZO87zePFM4gqAhOM4i8noCddWMdnKujkwBYnqHr1N6CxBu9emc1HBYwS
Qp/DZbxD4gAltxW8uwFBOzNe3mrQiXEPz9ziIZ8n7l8s7JcLJtEEaWwey0ImWabn
2Cg1yfFfTZvR1finO3IiqUhgpHrkU0pZ6O+xfLx0X1KS+Np5Gnk5zTXff+aAbU2a
pN3axK4ufdA7vcjeLSSNfL/Ur2MHYFcmAGh1HJjSPojAMOtYfJ2wFq32HMgH8gr+
UjgkQ9x7I+yvDc0rxB3YCzpZNP3dkXFWN/diIUmN/XQ7davGXF6WNEOtb5jRKbWS
FoC9l5mZXdjbwBEBiAUYCpP4TxgSz7gJCyXce8V2ltfWIdUZqWZsdDpaJClgC3od
/OCwnIcdDXuFDYXDllaDs/F9SXEItwZCbfZvjISKbw9TP9oColZ+dCswk6mzssGo
4HtiHsoY3aoghi/9jwl2GAWmD2b90ZB3IVzW43favxm9BW8lSMQdI7bl1z1hIERO
ch0B0nqTy6tNY4u5q59eSvJTubnlKoaWURESbWfzYsw5PkMaZSKrCj8dDjr7cNhg
DPEE9fietfNCpao/XVdADOQalEQ5GSpkxgK2tU214F7pUlV4CFw4HO5yy1DlRelS
xhrGlf17Vg2BXNtNKFL9xKhWS7SWKQhH/exu+a0Vu4ZUcgoCRVJvL86xj346/sBI
fn6negGfdRe5Mqz81IWeA7lCE+BbZ1Z9xOZXfKAeZ/j6HwHzosgk8lmJdGuf7EWq
Zvhcnj4rC1c2NGIrfzhelswr9xZV3Yshe8nzRKxUnvD++Ogw0+usGs2GyZbpI+l+
yKyAwdU1ioAStfq6+jb5zKx9AagSKsCR253u8udGDuJn8dYViBCHZhDQX7EQ8a0R
BLJZCeVvUCo7YxDnCFmfNN8/tHOFnip6Hn7I2o6XFJOirsSaNdRqjnQMLexTQGSd
UTBo+MePal/dWCoBYRCQU14V3iIuviwbJimVYSM3yRjEstmc7L6sLKmg5TMiA6x5
B6VtVOALM/6N3a5zNGgB/f1sCVi/6Ck9oVzFRh/22GhPmRda+2vGCe5I1C1w8i/q
3kRNNm6kB5Vz+pAIOHz2bYRdCIy0e3bhCGze7bZ+vpDqc7KPHJMRkilblp09fdLf
A52pLMOdJfCe21POYcxYBffnTpCrAIrzWFoG4BgFygcmB+oTX+2ljgUjpaK5WkxU
syqUbcRq9GF77l0IvDp9/dqFrtpJGsDl3Mk/F5jXoAvtkJpp9xsop1uZ3J55tGUq
1dlAudrkSBAxfKJRryOfBVz4wiFif7ibbKYq3vyNMQNMu9TIqOk0oR4myIEz9OWb
kXLKvAjGEkX/I4cgCqDU3OvJqcxOihDSDiSmvZDHA9yPF+pSDAePKMqM8bJWt8Ol
jrWCYV5jk4cQ9FvOTLehmj3KQTXGZrBp6JU4LuR1YIckj+cOO1iNENZoMdfXRYiq
ZuJrnktBCE42/cef3T5cO9PcyhJx/L+m47f3zQx0S4oqpZ4nVpzLhqDbtW7XEDLN
RgCHMAWJUz6F18X/BluN6Kuc5GdND3MAi0LCsZzCy7HAHFf3htAnURQqqeod5pUj
pmcAOwhyj38+/34bPPmwmRz1JiGmedblRUhHtTPhgDvStnVNvLDSNaMGR5nNg+Gf
ys0TN7R3cBZk5RDZoh5SP9ifpAZ6gtlZRiiJYjpGkYjLT4+X1+Pd2qn3UXfisZ8b
rDN6sBqQqSirCY+eg7ZUmbRl88jLzAFxnTWWBB/F185R1AMcX88X3FWvPyBi9b1D
D6NDhC2mGqmE0B7+2tFdURuJcvzIqa7jh42aBnczuzGwX47j90DamGxTgGJ5ViQU
AxQQlbAqlOvpCxw2+oVfoRLKZkvelWZneKkoHXAqayL/xL2ECQxq8olpHjfaBLJw
ie73bD0CXmUw1yJpZo0XrKsQzag9v7KhnWOicKmbR3iYlolckf3s8fA4AAnlUVHC
AkN/8xO41aQ//lf8LMq8rVwDDBGRbWY3+wrMdS8om2Z70/Tkynos3kSfx+bQ/EhQ
13Mk1rC+5xmGVpBlrf2H0dUCXn2nGQzGm3Qh4sc12Ws8zexGY2brm3bn9z70S7Ky
7nh7b36TntBLk2N4LNGS24m4MO1dtkCja4poydXdC9lHf+mCm0Z0P/u5DZm8bxZu
8qs7IlfR3wzJ3e4c5tAV/mN8WJhn9r8f+WdG8mNfAN4tPLYprBpSz5q8WpnM8qJg
+NSIWVIi8EA5/wp+lh33fX7FLCDEkonLrBrxLAb7Fvu3W9WFQ/eN8fZNfIP0ro9d
q+Qnrwt9OT+jIcbwIk/UXOCiQcomWXaPs9kkArzk/PjHhz8lHvEhQY8AAeR4ARFJ
3fRxuR3pFzdEYwxjEJF8yWvwi1LDo6jkqx4IKRzaUQsQe9zlibDA6/QEdwg/XuZz
ZomzMQnbEQP3GlAsc+ekrtedNI38WXxCQCYqoTnMYAE5KrqiJeLjjofD39CYmOxg
siw+XwD3PXU1gYwWSp/OOquE6sDOVQcgaMZ3vSidftHFqAdU84Cjd1hvnifuC18g
oG/4dSVvKkH6uuCMp+IIRO4rzpLOQde6TXRDsQcAqCH85C+Kv3b8S6IZfEtMPD3D
rafVrdIB5K/mDpf93mJB6NIz21d7pp0C8OA9G5W8jFapT51f5S13eib8MIsUsSZC
g+iNEHZd0wxIjTRwh/T9suONutvbc484HhynFto0IZBs+U7eBUNJ4NJrdQZdWg8f
5wQ0Y/RA/QRazBQ+ml5k1cPXxBD+evabrpdId5NUSEXTmfLBiP7WoJ1182wNFuKY
70RdUtNkXT0B6XBEezvpNZFy9PdsDBsXcY13B01iSIK88PWohxq/9uUKkSSuZGW/
ppFxXzo6LJK3TMiyYs8Nq2W1VdMzQjXOgJFkGno86w3LQjw7P31zqbmBXmgt9Z7n
bX2WbUjgXPlGe2nmEzFygH+GvRARLZAvVAFEpRnyfAemzcQoQb1LPPs0nOsfJuqY
Df121VqXCk/z72GXX3bZSvlPwQ5hN4JZvosyboPbrethaUPoPuYoat4b3KNIfcnn
Jyy+qOE5QzasiqjApmhhgnczqbslDpmFg7Z7+xNvQvojmKd3xjWp5NJIImepjfOM
o9t2PaUeZoFyzDRkPf6s++2yjEECPp80zcs7YWU+3mJvDfbDbeYevpaHUWrB8qW7
tXM3dy4k+7TvrYwHIhFnX+zrBFBhHmV7h3acS6FRHZgYHt+AR6d4hOhYlOGfwnVp
LkgfYo1kM148ReweAF+N0JeTEMUDM8gng4vOUR60kfArVw/hmKlA9CHa+PbzCoXo
JLyMN6VOyYLCmPObqGYWRA+qU8k/uSnuwP7X70sRMF9hW4OeQ4IfR5f09ZgJZyU6
6DDiZxQuJBO/J+FXuLaEXXXqlwfasmRftsHPYfuftAqRMVCf9hsdGsXLxXgBKpiW
U7e4M3nzsaKgqLIv0l2eh5Ndoe+O3oda9X7cBGnX4M0W51rMoLGtPGmo945bLGRd
Aen1OuGnwTpFF7FlNqZb+cOXvrEDx77Sh/xphUC/cmHLlutP7y2tHFDmLQrbFept
MqdraIFvYipjDdkgSUVkLbz9WPjS+8BVm12/SAh7o4ic7/J4rJiBChI2W6saH16T
81elydcdsAgj98DBtK9jYsJ5oFTJAfyvx6aLpCX5IchUWfVBzExlgOiS4oTVaHTY
wVVJ4lsjA4NEHPSVrwQ/AVjWLxym5SGEiMmoa5K5HtVU/56+tnG2b9RZCMsLGqye
CFf6c9JrKdKlxKimFlkkqqkq9wEKvNAW4latfbIciRY1kWjUXzaEMFb1BzUZPnJ7
DPmHxwDELD5B/6FplQkDgTAXqQTVtW1QG7wELhsMHjMRoEwaUcuzUs7e4ZTrwBGf
yIADhmz+qfIV7sAqfNrkZm0sJ97uYxIa8F75ojePzXAKm2QXHh2ITUbtUI2evcg9
KOH0L/gRHxRutbqAd4EBQm/JKPXw2NSNbDVzpvMEeaRmDdaLViqh0EAH5330ueVs
/60ASGrP4GHTddt04RKk5EVtXv/137TtWs902eOP28HGA4+GfvB5YkYOQ6z9hxAE
xi0x3dTq/dhJBQ8PBy7oyQeTTJTIMtXFyzqwKTnqlwR3UyUQgxO0Q9GsDRbDd5pF
Yrtf1gUPmKgot2V0aG1azl4BQe2nZ+enYV7m7bFAQaQYsB/2lwj75Gaxqrm8hs8o
GlHXLuRYNP34qFO686QXMSkVTZUQzM+iMya1iFwjF6PPBRAAGZS3jAazYLEbaKD5
O4s6RmkDI3xiYzVDp8dmtcrPTEDAiMxpNOmphUo/8+xgOBKhC+0hSk+G2mZW0D8z
pX/HQlUXAEkNJB2zcKEDJWs09aQhlpqcJznAbNZmFkIA+vzv0pgyD0RNjOlm1Ux/
cKlwBhn6IFo6UyWd2MPnre9nDsFtvwqNxGR1J5JrJEijnjgd2okx/maeBLW1nJam
FUv0qZmif6br/NfZtv8t7YQ2CY+NobjEvGEKW5bZ23cxK8aH88fB8H5h9JsDfTAF
PF3DDgPithbhVwMDQGYMTbdsnGNPFvo8KDiJfN0G3ZcIQRhYYVx/71nu3AvuxeRn
3WOL0CeXlTGC6/QW0ut6DYJXs3bEZd7CALPBYqjO+37zjzqde/VhqHBcu4Cxnh5c
76MMdJ53FKB9mzawtzbFU8Ob5bbUCanqlACV3FT0UInuL6zCroth7EH8tSlLngMH
uLWhkjmv5uunw0Ccuh0RjZtVMqghUdVDGJfELE+LusyAi4GsZLVXLqAqXernKXpl
KE4o+vy57/r9qwfr4bQhRcBuW6d8Twrj8/QQBXrYDhnpAUuFc6HCpznJW/Qk9Wa7
ChvoXivsAWseqSdpgcBuNEbmvmxHBOMbk0N/j9yL6KDe4/1KTPmjcb7LHnWH+sXn
TQSHB5BK9hwV1FkOHSi++FVrHchDfnU6uAde69k5t9c292Bwqx8dBVOAF92EdSp9
ojRO2S8ykEyj3m5BCS+pEFomPht0ZRIlwhkyOYFG8Z06oclDVYGJm5WEXDVOncSr
26/TBBvlbpXLkisGSb+SuEpDk5JMZMnqJlKWZEdDSH0SJWGyh9k4wdVkpMqDWdOs
vO8WQiiNgYGhmkSyUPaimwP2zy/dkMdWFeDEmFQRlJvfEW3y2yOZfBjLzX0XK0jl
MSg6//Z4Qp4DH1z9OMBfSljmoS62lDE5j4fdA262/DTrzv7nJMn0cr7NomTAjSqz
fmzbSMOnRMWCgVMZ9vpbYR28IehNHUGPmpMesD4Oavk5ZnIs6TtJQQlBUM8fs9I6
NMN84B56oF0GmjGZhBffS7yxLcbb6+BE70j7ILumBO5qjcVpbbRIc0xupPiadYsc
q41G4RJ7jFm9E4J6yKS5qgMHTtdtBVm1Jk+CYzsLCUiFFSuCX2BnWZq73Z9Mu2vx
AbdatyDBYObTFsWmt5dunbTqJSr85ko3yQhZ/ib4DY6rUFQBEx6KctbsTJ5VwPQ9
Y2qz+uAPy00/z95KxxytEEQTWGN/krF8u2NInK3RV6fUxkvU3B/2zgTaiiOD/fic
iipQ1vgCpjA+P7u6DT0eRQBfjZiid08ueeN7dMRQ2ik8gck492Aaqwsb/5jLhrBB
oYIiJOZNyWsS080jd9s1/ZrmcUnV7pxzK8OAAY/Q1svUT6+sISAKj2QIoANQOfm+
RcXnCnc/zIaR0NqMg7cjDe8nQ/9UuWhaNfLX9/BZ+FUcA3zxa5N2q+dnEU7rRTNG
Dl8ORQrJ0dijXYzGhkqdo6/wJFtX/6M6ZYLLOpPyslvcvAdwuIxBewnhq5UJ1nEb
pb3dW/weB6nhhKQz1SZv9rsb1kzsVM7qeEDNXeVsw1tRGScyyRWZ6Z4PkPTC1r8/
/CpM2FAh9s6qYa7AM2YWQu04DozHoNSYuwxJZszkqa/+NbBSkkCj0GV4h4HPZ/g9
tWX7+2TPxNjzXJTBebZHICxQgta58MwvhDqKJPSCxc7CcWQNzh6J0w06GkxplLGE
drJfr8x8nHK/ZwLAgKHxunqT0rgVQLdHUFQ1PwA8DhKrN4yR4lXkC6gIXP29zwU6
RnUMDpkbGo0KPFlG94n7pojrNHBu8wK5pHDkchThcimAeLJMsJ1zsPkwphhKq0X7
vjbGYav3J7cvJXU+RWHEy1H4fhdbLIJ3saUk9KnLhPBacl6lyghN7ma4ImDFNplD
U4WoektwYiYcnss1DJi/yxwrB8rvyuTpL6H7RNUMwA5kiVndUWG/qYhvtN2FrIGT
IozNa6vo5QIML9DxQL3d2KQsvYhVfTOHd/lLUn4N6EU4eNDpRhUH7y4esPubNXWT
9Ej5d9XikeZIxW5FCxeYDDKMjeuHHyUvcDNVsUHi61m/zlsrnDjSsc57TKvf98r5
H+xTgI9yEgMumPnzWFzjRRUd8QOLIb96xfpxacmFW+jVyxyxyAJEEu+mUPYEp1hz
xzjZTqvawkF6EWhW8nBgfEBEWGpTCY+Naq8oNPxrGYY2f2M292j2TuY+dcHO218W
/F5UOPvO8KbLhp48VOotu709ssC6LgHrm0zvUT9SfqxA7DXTzzD4KYm5Jxu9G0AR
nBEWhjO/6F4nauS5jY0SDBd7ZGFFzv8AMEYsctawz0qZ9u5oVRsPHpTzISf+tWu3
PeNWYZ80umvru2bxerpFjiP9C+IlT9UjdmuAgfhgU+BKQSqeJEgT/vmJRIMZfUEj
7KSVpI4I+69T39HWJ4YaYPisH8AfHfsjLtrGv6h5hkZZa3BcDluzI0aqXW0w7O/K
592ZD5ozjnI0MBWlBZOtgsfUyuFZv2RakOkSIO+UOrHC7vGSw8niEKDlq8XRb3Lr
2cHhQ5sHcJCKJpgJrnwPUX1ch5BLNDMt0MB80RbjFXY0iECNCLeh6TLkreHW86RF
x6I3qy+i0QYsffU9OwkUUgEdjx1keUsWz0vbdPJ5M/FH6Cyd6kxJoYL9tpEqHz1n
tTZwJkGgjv2BPIPIzOzo1POCPticwhPHzqE9m8PfyIlf/Ncvm8a9DmcfQJ5afmIf
lP2n/UAILOjMsP8dXQPP1xACDFz7Zu0D7ZmBAvUTnemdApqZA51awUjG8fWlAALw
zJLtF+nPMI6d9KEs5keVrUacm1gA+EzMEsqNXZEv9KUVpbRTAB2mRuzVCihS5ENo
bKUpdtU6lwalJOSfLzKqNDgDTgXWt0KbJEQdRxEwkuxRsMDdJ7vWRVgH8pAEgaIS
2D3EePBhcwUDrzGq03+k6jSzFOcEEmTqILGglr/L6Rrn0WCXuTIsmC/FlxHPzQN/
KKYYf1hIsjpaxhNUF3QaiPc4a5NoL60oGogU+ODcYF6gJnP5+LtK7QkCiIhoRbcI
xXuKPfoEjXq/ASqcCTeShE/BfR594GiKq7nnhNV7CaWxQUenHyMbTADjxY2+v8a4
AdZVknbNPCT2PMUvYkvPnMuJx/BbNpA0/tb8mpVU/AUsuFpG1zZiJTrpaW0oFKVs
Kv6TBPA7nOFw1B1Ym403mwWqYicm3/ZMY1tby3F3Lkt8JAfpasUkB37FZkDjFedy
ZAAE8/Mz5IW30pbxLG5rL7sQB4jeb4mTL7GkjCh0Ihau980g4LOLMJ6CA1vo5Dqt
AQ/x/rz2cQytQmC0689ZIjzpFmqMx7wywnNFHuSPA8IMnlYQdjuUhIloHDzopZcB
30nYmO4F78eJq0nTtNjvYsgRVEXwh0B+N7c+mjk8DkIFNk/kICrIMJ3VV9obmh+0
TNQoF2CSKXl8C2+4AlVO6fAucZx7md56h3j4njhZDiGw8SIRwBpnTRDEcUtqTMbB
Cw3XH3MyizsS7sXswXeVmDS8Lhi+GPS9jjHFYBB73mQc2m9IixOt11GTZn6udDrC
jOjUQp+XAr526XjUK5SNPRFLjYt2pAS2qyN/f9W4aPzwf/+LcFFJXwMZ2LaLx8yn
fCzUY4NQuv17IDW5jD62KtCw3O8SqmiHdxMuWQw+CQqj3TbheWkZg8jkHDmanqBQ
00/NeGU7eZ+cyxQA8y5/zN7CmmdVrpQUZvQ0oKLrQYt49X8mhC3/SxTCI34ESrdW
V39cSWTsTCXZZvWN9xz6gVVVldhXlT+VRunArb7FbRhSq2fAdp3GLxaapAkQ28bG
+rl1SJ8Q8pm+7lWBBO5R3pwwSGAUy+mWJytcGH9GDTlii+ctYV+KKVmpVL9knQ6j
dW04e3vk356QPXjutkXA+ru9gSA5HQr7nq8fygz1l66yBMLYDzoS8VdXoFATZjiy
IQw5Qsqlv/xbwaRDRuFkyCHNFRKWuOxdJBpNGwqAJwf/nuhbXamAmcf9OEjzyhct
0tshvwrYabr3IGufiYbKFjD6wZce104ScQyNUWr4sqZOznEvvDheYepUCUj8gL32
Wp38xEiz+kMUW5/euJDijDwqaKbjHo4TaasHremXyzjCt5TcCWnNl6nYqb5YdXqO
4QxefAwD8YFY0W5DwWJ0pd/hqPk0Ydy91ORegjf6zidxEjaTJHbpeaJTa2zYKvk0
WfWpobRPXn1JiQg3SW/YvMTev3/vZjWgleWoIwjVmQOW3F/XVJifGuDgI7GuXxUn
FNlZyDem1LAWCWFlgeUlzAIkT93QMjLXRBYCSB62qK264xxmQeEECo58rrlWykET
HYGyCE0HIjEjUntMlgHha3A+RjOuIr22EcEkWf1wnSeuhSEyvTVISbbBsLSzeVXt
4nGltOmlg84t7xCk15zrOd+VMOd5dy792Kw5w8c3ej9NtOn11D1PsbjEUNBz1TEi
VZZGgFursfOVGUe62metdTTcAirvaUSVfy0FdkqYd8HlCiHzJSx2EeU3XMBBcnrA
Rs/JSHDuRgvFB+zrHLOuU0A+Ypns7Molf2w0gLU5/KZCgKCiHvbFi28Y6NE6N2GJ
QSf8CYcRAI8hPSqG4giMuthQH7ru36ihIcSWvQqqAQoEwXbPpiFYYOxtB1Y6F2C1
jG+sc9QU/4ouYMH/XcT295uvn++TardZ4dqKdPxAPvLnsIbaGk9YaTgVdLReDlYk
9h641bGkU7MvT3bLXpKt5I0t5Wr2nDojKbWHC1D/LoXVuDZkjuRLZIToYu/3g0HK
THHFcjjTf/QCK++VDotUyfiDzsGmLHIYmbprL4d22miUisAAppf1zoDfhMaOAplE
MRT4wiUv21lNbakN4al6xoE+pUypPUXgiO6G+4joYARwbKJCNTegCVcry7pOn5kX
DPtXS6zzSgwjsQ10Cav92OC08+NKDTcFEBcmUYt9a71daogfhatGExGlV4xHR+Yn
bLnD2rgMO7aaC4VOFBmSDuofCxZEwxd4jLEmvIWk7DUhT/tgu6joXpPzuiglIink
6JLQZZtRKSJ2buP3VQZ0KThyMc37P5pUxgTHKDWCUzk2EsrVRR5AvGQBf3Kr6Kxc
Jyucx9Cq8KNCZpgtqgdMOaZQhGIf0oMWLUUQiX8stMlyYz9AxkfqoJ2+CwqyJfTu
hFr4O2XhbF621yBZowVEfnJgwFWHW3x9PQGfBufmC1aYURxli2PfVq8KgsH7b7qm
qej0p7sKtywIdjIWHUddiOXhVHyAxKfNwvXdNvO+n7W15vUjilt4XuELNWXg8DzI
vgtfDIGt0ZSPUVNZej3Vhk++/vpu0BagONbEfJC0LEITtirBeDwvuTdHC0eLQKPU
6+Z3APgMTz4UNuP1JZcr1wVOldxZ9sYNkdAoIgT8owG65altAsMpUDe3vj0wkcCO
LH/fJs1nO0OVhoKCBG0lmw++P12NPC9PCsS3EDuYF3g0ykACL+YGG6huQTwumsvg
bEZUbNfq+BKqOdv2bxGe8DmO+nvvlFJ4fuRVTWD4nzHd2UAV7dqB4TYs+Qx6zWPN
V4Vyzd6zEoMoleZhBS2EdfLiLAKaNRuJAH9No76r406DPvOTthJsjcmd9Q3hK2Vt
SOqwTaxNTkhqPz9z8xFZFuKg3mtNeixgwa6Wh/BXeYAA9S0mo/4dSwKQM+46CWu2
vyTKy+VDDz1SYBBW8AvPcqs5UhZHtwBk7K9XTh7XVf7+QzG4GQS5cNOGGrRgVhyR
rmX7tt45L873HWBuM33s/UtIYpioqiDgCUfSmKopTTcTGthxMWyXbON1/872lQfi
mGJG9bZEuOengNiYKz2IUKrXTllKowRF6z/5NkBm6EcEfyYZtDCoMTWiYXncCHnv
pix+Y7+33Ep5BZUqX/Yt93Z0gQf5N5R8GzV8ae3aMKSClJB3jnTsBU8Bx+0t+BU/
XWy/UyYMIgFI4MKKtUK20F/D2Mt+0H0S6q/pjL55Xk5pNor2Y90UZYr+BU1k3Lmw
x8hTwx8MvKkjAg2tu2Hkxu6hf7YKUCxkFocBm7FkJvmziEK8MoH1JJjoim3y9gyA
cS465Q7QgFJeoYlPqwYSdvOJtJ6U6iEMWSJ6qNZ3ei/WsOKcvK1A/FiN4NhdfJfJ
Yz8C1OQJGA/xvgO4DeAesIFpJVK/MhIh2kM2puBUXaN7s2V+ggf8WaYXNZvccbvl
+zBcplQ8zgOX+eqVNWabM/hCSvmcubosfi3VJ6UKFjCbpFGABap70HlpyHppUEgA
CsFT+xfEKdavj3oIcjHMyOnnwUTLRwHUI24fLoJigjco3+8TzYHqwoG/T6lWGgZ9
S8sjq5FLWz+fS/d0kUlaB2sXHRKBT8OHdeRW+xwrlQVTXOORrZauC5BZnEVzhQDo
5bpOJ5TVuaABb3nX8ZRriu8ttZWF1AlnpHc5jj39RAjO39h3ZAH3mADHOdLPUo4P
Yx+ch/fd6AYCkNnW4hxxr8LXcssVatbtMvTKOlpCD9hx4/EqrZidEDPsRLY4cTMW
yMQwlyWmPi9i93ZayghSqFk0/M0dyNAACOCoggWGo0B16+b0s5lXzHBwbfsmSrt9
N6sRQELEoRlfD2+DTYaUKatG/YFQIMownrOovEZg3rZdqiX9f1JqgBwX3DTRbpyA
vt+OzuyMFfqXf6tic8FHo/ISvGZfH/d9FHItEDrSeWgTFBuTbsJB9nk++Y22wKiR
HOuuEf9Y3QkDJ1NQdmRLu+nm9dyP2Ihay+nTFKz6WYmULaIXpRe0bYTGyJIZhCF0
km7hbp6yOUps3bOdx4vQ1mpRq4tKOI5bAv/QmAFbtZX4GPXaR4xglkIuLqfCE7Ms
bey4Oir8ELTkxdh83+j56btZ9jsc9dMNAAO1RehXESMSXgGWncop+Mvw0s5mpuPA
Qr6JKwdHKIkfW2vfBCkPJuzz/Do99PxBPh9XZPtHVlsk01pldsE+YuCMZRuCPU7T
5LBXBRtbNLJI+xxh5BR6gti+1gq0vgvIv5paxqsMjm/gh6FzygG3awVCk944krRf
CXu9fdM9WgaXdBCH/KDSV8uCx+9J1u5H9HKedUTAqRoesfy0eOLut/mH4C+Q4iMi
sBUyy1l2Pf9Y2qFr2r5p+fYEqnuYsRC4I+wyZUUKaer42KLUk2IrDeT+IvkfcZH0
bOQ4lIpmTy6bFijnFQEIc2K3/JzNbp+AnmiTiXlmMZrRTugw+QeyDk33Gw/ao/Y7
Yfblsa36EV0vw30GHOVLVtzO7iUv+085y5ViZ0A15aO3eKMAAGRkkkphvPkR+J1c
snVoJ/TCx3YQFoYCiy7C8JkMjHjPfZhRllsZRaBkW5vzkoG1/roUNvDuZpufcJuW
gsNhn8vcYBo+gA+HbU/FkTTuJ4V0uXA5hNRit1A8g1nzZT3nBZlxt72tf6hotI4X
oTTz2dbCmj4CiLdNa9fjkEywpwqihkLfZs5aK2B5Pr9R+VZkPeZSj4TygZH/CUFj
DXvXedJYZ3FT7YOZOoJfaEBgAonI5jAUuNY3MyPAXikkghATGDH8c+taeKt590XB
gbfFr4SV8A5BLbDhl4jyPIlWnReVcwKD+ExTFgs21Cp2jp8iriUgpFK4+KaUIQVw
K7VC+0C6vzOsCRV9w0At+gy2xlCu04eDO1DNo5Q6Nphl6lyBX5Xas8L0ysmghqTK
hfLzzN0IlWMAcBEsVSk96VlhTrJSLuGynLvG72Dp4O47k47UMs20qrMg4grICXvQ
O14Qj5DyNfmdfVcfJBEgoi1fQ6gj/rfdJn/BGtOhMVq+XKhhSY7MQea8NGSmgw8R
IQ3PC5I5rh+KMaVWnlCJzWAB9vzpyB0GLzMkIM0wfqGVRn/rKZ5gkegVqt0a6N9R
tXkUO4lIjEc/jE1twr3C2nvuMUutwaabh+maxC54YwrmfienFY35aeyvK9TszGpC
j2Pn/am38vY2erC70QHtQV7Xv7oAQG9wOiYn8tsb1P51xBuhmMqxfPIzuTj7dhW/
E55MsQy9h+EVgx8cWMQBomzJ3c9EubI1ttRNKe5DaH3uK5NSjglk/Kcs8zLnRm7e
MJ9tguenHqKCKNZ0SIVMyWZtcQ6XknrYtkE+MGIK6EtuetCiv5tczNyfy1uXGGY+
QIoPuhKjyI+sVrFbGZBDP2YyPq5FzXB2bFGo3oAJj8fwkWeC/8+i7ThEtGWB9eSc
Jv07AIwQM0PbghLnj4/Q17xwi6TDCPUqSnqEt8lTaC/TtTYH30ZDlkBy3vGuJAHL
o53752fpYfSSq+w+gZUCISYkr30Xz5zsAR7DJpW9ty1kniEM3nDteXtcK3bee0tI
QHPcxbzjXObPGK0O1FtxtNoOMEMSUhAVvUV46+gkR9rfOqbHxlO1I9e0cXYKUzre
uDFtRjL9i1mJyI5QCxbk40L2AYX2raIc7GzqW6qJTRjLNeoBjEFsKTrsctiDqwll
wv7i+PktLJ86X6IY/lRtCXGPpwFfeH3aaqzqhyg/s8CWCJ9+PYGnu+0gMqSdyCtM
KaxkgOnLRPeo6LNdB/hcnVfOfQs6v/olfn2r4WwBpUXAjgam6nubAuPvG7XZISEH
ffQAzRU4zqEn0txd+MyWvpJPZKfiu4EXETdm17rKEmC+4ISaC6r2JcF5SDsok5mR
lg4wYCFJ1CnrILhb5am+6q6wW1+xzdnKfiRJytO1BhisYs4jGi/vU1G0lDiwpaKk
E9h3lhZJe+LCIcgjcSYPl9RunjbyRnmmduYKRCpBeEQ9a8vtQ7DbDydH6035APx/
JF8dlxPNmv3MK0YNhjQD5uqOJm1Igb4ShU/8bYMdys7XQXilRiX9D/Y0ATfJgs/h
UAzw9e+nq4kY6LHlkxsKbDv1L7MnjF89qDFKTsqZjO108tIxxlqvLLFNtGdhffsA
ROmymObLwyDnnIpycs0O0m2ntdLPDgLB5k7w7Y2KK0YCozVtra7XaPdeX+vKW69u
c03xiA+U0rB/4klkl7gsDwBSu7zprKqLWWiZBo6ndL1RCaSqNhqVPIi2aouYSM7y
OpxqVajITbFneZOnAj2fH62IqNes8YYO+8YlgtuptnpWBT9xYrM/zAWD8bJIBlgc
MPDq9xzYcbkogZwl2u3LSgRcDjLQcp4M6oRXTgjAwEIXvqq8pZhyNZ612TmypVJR
tpRS+UrIUHRdxhG2PXIhroQFkUvTSo2+Z4Te4fx2SY7YGO3Q9WKImLVt+4jDBm7u
s9rltHX8ZQiE+r+EQA0pvMEHC3WhHRVMe67fjaWnL8GcyAvxTH7Z13Vl69uaqtsj
IgyNqpNTOR7JTPq/TeEwF4HR14clFLlU2NnJ++s5qWr1fZlN6D7Vgads/KNo9f5V
i0CaUuO2xBR2ANk0eOi5kuEqcLy9oSqiojPgy55umMQjY67QMxqaysy2KHDNaGMr
zIPnuT3E3sdjXNhtf1iItYo3A5JDhVSUQfB0k34E1IdcwJljGdY3oi3HCYWhboAT
CKWxvTPe2l/Cdil6usT/euEfJvzGHgUY3HhiJtvfS52DDUni2J+EhfPtflRqEwPP
w/I0z4UqH5tI1R/AjZNObv5MmLtGqUtjD3MVfTxNVYNAPXm4ZRxok3q0SPPiIyM0
X23ZDBzxGENp8US/uZZHXjUxzend+zY3JgRMZSYcY2S7qJEr5uJ3bM1YVH7A4eBR
gzCwQ24a2lic461MBcDkKt+W9i1+ZHPG2aC3iJgJQ4YavNl3c7btsg7yq+rgTj9r
zjEwSUjSsu2TJ40dNlSK2wbl2AIEJSE0IEuGM9w0w3JdBZMz4AvWhRIpOuWC363U
QBOHC18A/MIe2oiy3YWGO7eyaVDQDpVYZq+F754gRjhn5DFAwZHteVXqolvC9zwc
bMUQkVqoWG+lKZt7UCAyKd9w4sJizsJOaCR0SgYvrKpTntxSchvENckfObFtxT5C
D2EuPc7i6TAspR0asft3pQGHh9EYAMlcfO7gLwoR+NpgAt9OR3Vswn0uskA0Aq70
7do9pzf9cuXNcWwpnlTyLhoOtshw0e8gw30ipvTpdgnU8pf2SdDLnNxMEPrFzRsh
FHGHK50zsqJK4zn6DqPSdAZf9C0DT/Q+ubT/4OsrOoy6FUEMapWfm8w3Ovjp0/by
tsKHXvyGp5EHcSCQiNGZdvuerRL3OujfBRPJWlwy5YsE7Vm3Ba5Ii3trhsTahLnl
ipSOZ5sYdZTUZpj/GgOlrPENgfSXFXXIYNdNx5uiGftHTEuTVI0Q2khFRAOvi+NM
AZbQJHDaiaMn3bq5XOAgSBwngM6l4yTcJTwhgwHSTcVYR68LycuShIsav9MG7HOr
D5TQATQJ8dYIzyBEBi8/kEy4J8GUUGFSxt2uK8aJl+8uib3JJsSyrHMYTQO5bV0F
+dD65T36xsVtpiNYF4byz5lPFSCZXoJ7rO0uoKYWFvUBqkTVDANEah4y4EIU+eAo
3GkTM+gG/ppFMbrcdqMkYZKWlAr01YHLtv1AlC3cVpRkhG/3LOUTrKiQvFY1Byqq
5MTOgdGaTnjkTCXqTfGWgM9fwkwu7FaLKZmpL2Jg3DVlQwG/yX42ytqh06YitXY0
gYriiX6CTFGO+BqpzwOM+Pxl3YLqz9ppg1C2zqz/ooXDpGhusiwALANhvrGLJqwH
Vl3hO9J0cnZIImOf7l7WO9BZEEKm12KWDMF2+tQBsxx9yE9zGZyvwCHMoI3Id8jh
azryaKVTAGZPARF5q92YF1y66cGvbxQ8VxsYRpJ5bFMB17Mfx+DIciByX4uRT0u4
11IFTaly1LafJvB8vBsXhuBiT7XOt4AvFRLhgGMMVzCobf9wlw2cgBMRnQ+yr1Ak
BM+7CmRhKqgLKFBSV0+QjKAS48QhXviGe9uxM09ub78UoUqBgjshv9SPfplFNxFT
vTmo0i6lc82ECQ61rnnX0FLZFfoI5RG5moyOEZdTn+/f74Bp974Rw4eevmB6t3JU
U2u2EpC8/lYr2r4ai8l6kgF+1comipKhoN85d0BZWLGJPsiLllPQLzz6jwVEddvn
vdw+MGdTl7ayD4eDC6QT7W48qwrIxZAPppOL/rrrFp0H3DvmdTHCbhg9T8/eRqCD
99r9RvTuWPhsQAmBu9wrQ1tHn1eUl2EHpIoSjIfW7LhBzK3QW1PK2ArqTEi/e95L
LYqHalAXJXhIEmO8djbr9akrMFXmzVctrSkCTt/ObfLFju9Wtkl5y9/Ztqo3Cldp
bQZqRLMQa70N78UNstgo2g1V7BOg7XFKvabaHOEIJTvIO9DD8MXzv/bN15z+zRn7
oW1BzlRV2rKxpMWCmvMwkw/XX0TzgwvS8I56tHggnkmbusP9nikkueAwa0dOKN6H
T6mnKGrBZOXeftoY4SF0tM2VqMxgAmb3W9coBHuCTdIwrk8BPw5MBcUIjF9A4anE
Zmne/TWrNlfRtC30TnugtyD/F7roVcIKBulx/McJnWgEWU/jvgBII+0iutWVHR03
X3BBp8IxifeXJ+cJGqWoRzu5i0325qx7vFQwbf1hFjkeZWK+M/RlPj4Yt1cN/6Wg
ctgaVFUzM6OkqwrBHP7M8cSuF2vLEpnJbCJsgSDB3tZgBUKqi9+aAut057fQeVaz
vFbqDVm/Lj0de/x/X837v/7HfIfGtR+1G22OvWbstX80PirJiyjPGnWWV0R+TIQG
Y8agY4NSKhj4QfZRJT92UUGDfiWqIzxCkvSOTF/GIbXUOkcFIjceZ3FUdQEcBXJA
hUQvlzZX/xBZwYlXrTdVGJnjXtx2FbhNWQI1jp10SzrxtwIwItF0Y4dlx4vdTJZ8
PYX2sbtLTdGNPV/FlPsNtU7OeuWhGqs5BAhu2vXkk7kPFGvgE8ZLtQggpGszjyR+
IpyUDs/q6+pqzcfP9k8cv3S9gWnFj+1079OQggtM9AFsKWN2DOIzEIezsjhKVQ+/
e94vddy3DIeelRHf6e9+EaSVMqPQ7WCO7d60svF6x3v9pZh46r5uQjNxIkqg6QHi
APU+XKI8fWj22JLFIADWI7PfvjxSnNsjmLnlN9HuJoIOFLoiVututxGi5kIjk1Fh
5qU9ibK6kZaFCPLshypuws222zSyhvk1SmzvBnQIJl1AiSxBCczKyMKFQhYbs/G4
oefYImkmw/msqLcFunTAttRi63va1fJ3VuEib/8nnyu7Gvrk6Ex3CAdWqdOvzk/4
Qyh2KQpODDxwCENuvtlV7+4YAPB0R2Qp5Uu4J+Wtx4fuOkLstHQHqwSHDngOJvHq
BZE8KEi6EcG+BZ15XhHCPsiM5XJ3S2ekIEMKUW2OniRdSovnDdpKuuBhABv2Wcxf
ngvTjSm+H80emCAy+Rk/KOpTpwYvuNEYbFPaAzPXyK97WP7or8M5pdKR3ck2m//k
n8+slBVosOA0v4FNXUpORuAvUWqYm6OCKUi5iKyhSmo+eND8Z2l4he9uM88DnP1h
bG0q+bpMoIn9YtRHOMjqjnK6JtRFZTiA7l04YLpoqPrxgZsbG/UD8P476V8azeyA
aYWTQLxgA7gYUTrYiwilvlXtXkKpn33B40vKwwAu1xYYt3wMVDdAyLveBX/zSUoC
kfBYYk0yfcssLrvi+NAjSGQtNVVIXvS0wFCYT/npYr9oKlon+PgGlytW31r6Z7Qo
Q1iGqShc8mNavCuWlw0paD+clwrQPBOlV0bQ2+fcLKBirBD/rmtnyrJEL9C8db/d
3AqiCNmj92L3B4jZkitO72XQ5le2LImaGlwz4HJiJ99GsETquUecU/j+8aTS5y5V
/wEFzvjN+C6W0WntHnV3JFT1hvylt2S73rwtFcHxInV5B6Gg0V8vEGTJWghbtxcV
yXPyw0nW4DG25KVCvuosVa9jMbhP+GGN3iTexGCWhOd0bOf/zaBo3PfJe/kCMech
5hY9IYXnob/mJ/yn+SWyVbuclRbQ9wemrvOajq4+8PaWs+no7cBzTLrLmareqTyy
YtcVNX5hjdx8n/ILS12AfKUhfSYh4Vygfu2KtTDx6vWwC374TmjNzy7Zx/fFeun8
0j8iYdKwUamXDRuUFEtB+1lqMatA89socMVIp+NTpDzDZn3USHfEcAUGDh7thXfC
YddhIS1I1YwmgDuL22s16bvyH3iEGW0E3e+DmoAikev2CMQngha3Ho7WbcJJ8zlk
hlaPGwPcpY/I1tt7+sigiAcMBPw1l/Wx8qhKW6QyXr7ig6v4xRyi7unQn8MhSNel
n8Xp6VV5LQPw8YBVlTQfo8lGxEXDKESFK2v+1lEDBzJFOH0kFXGQx+9wQwU+kExe
zdgLnYeQ7x95k1iksrKJJfQli0lSOQdrYy3uGBPbAgMfJ0p502B6o44apyyjuFvs
9w1Atd4jqbGrHzTmgnh+FZBY4/vKMKuLmqIE7ka4OeVp4rTrdWno3vAhnyiuxQDw
a13QY8rWnQHNUQgtbquN3XIc+CQMvQXcX/yHFhVf+205qf7KclTwr5QmbVxpREOL
nngEiZrZNaXOApQH8WqETsM45TGseZyiPdhHmrmfKp4pF8WyxxAPfRwU1TYOEK3q
lm3hBoYkBx9QZN4E759yMPi0svgDYUoNW2lbnmoAmGLdXu9gen76Rvt1aFn7x2av
43Btk7iEIK6KrMsQRZCwE2nwGK9deWKZzN6vWhM2uBKpW1fdPo6z/NUbeHQlhji5
TQpOCVRq3hSaIizEQJnrZUpkytC/bXmiUPnBRW5DBwiM7oCi9M9m/Anu7cSZPdlu
EQ3KmWhLIkAPvy5XyW3WxE873lkLLV+3C3FNnl4DabWMcN9HjdJnVqhQ17QOGYbM
4DABsJAjI/+wsAYkX2uE8hjCAXVkzz9JScTxeS3Vt4XZuYd49CpzKRol7xZuVZEI
4j/Frzc9vYBTiPjZt5g83tfeCoTb54bClP6bAbHRIS6KFjPsJMthE5pIzvVu1R02
KaVPYaytX5jUsUU/SpFCTjpEJuhiZMXG3QRwFX/4ATTtyvyjO1Xc2rZZqJEk78X9
fzTi2ZnHw3bkGFnnOsAvYpjWBU31nJP9vMQG5rffuyVKwtnwsP4zubONJKQa2tJk
04Lyq++nMnskn8wjTxu+o++SyQsMwesy5uhaorLjvVb1hdItpoWJTxmpPCTEeKmB
WtpxkGIzJB3DDrkSAE/cNoJvrhP57Az9tSIqHQ2Y+VBG31uVhfjzem1dQx7KKSzX
tvkJP9V7KUQvGjSRCTh7Z0fWa6whothOHXnFtzIoYr8Bbi/msS7CGjJB6NZ1Oani
tr6o0Zu1S2XxIuyqDOVoXZUflBG2ygpNZEaCQDtk8p+UNgfxXuGjtkBBzPsh1ZXh
auDqE67RLfLGxt3nF/nbshqgvV79RqE9/kZg2r8xkHEhDTkDln5AGnNjIIpcEkuA
6HKSCd49T6CgYxOfvD3WlSRwnNY9K1Gt3TTWGIcUdau49RK5ko46wWTA3+s/MoCD
tvgTFfCW0bKPi9cmRDe9QGPJAvqGVqUtdKWmSwDWpMGuolP+0QO6NVla1Xb04tRG
txXAfzxX4AfaMFZqJHse7/VV9Oef9jOoClxmz+q8oUnCw7bB+wIjUxeTrzXxgnln
26uiA7mQOdxlO5T3ovm/z9Q9gP7v9NkefmWYiSSvx6CON3zAvg56eN6b9gu4r4as
rrIu0lF1/Yp6DJXjuFcolYNI1aWJpllz8nlUyuqoOZfz2dUIAO+uUvHu/b3Zn7fq
Lex1lRNfCjFs5NXhvr8CAXUWG/kgONqNGZCpRp7jhDr26FJmp1OFR37Ll2sZGW8T
foeydHt8dB21pBZ4FKRQeelUjKzoGsjm0//gySiAKacBQMWoZ8pS5POs6o4JCBS4
Rv10MC/9XDxK5F0uAK3oU8QgAEizTeoQ8vlKQXfCXUyNP2oMo8iKviQLtX8Xw4VE
8KeAUy4LRFJn5O6ED5jf3jiqL8ukyg9kALZAbLUvWO7GYjXV3t70GbEwYn2udDa1
cX/swqa9bzywqS6jTrgnm4tAatnb3YgWYZw59KiYcn5CgZjuMoMibfJmsRx+zIoQ
xjxUuNN+6TTb8452oanvRI7IQpuk1n1srVe7FMH6OCnxk8T78q39ktfWNVmEifVO
Edh6msZdpPx1NxG7KkhjjHN3BvaPvRf04lZpqV4YaU6s3Z1RKODZFP+MGBh/4StB
ZxA6r2i0VHQRicO5etquQamxgh/6XK3gZ9jXgVOvsdxX3PSZtCyUKsICiRt2ZH8P
PzZHwNt2ZPM9p5O8U0tbLZtKnx+XFqHk4efBFVy1Y/N+wOsOuZUjP4hewxDMDSEQ
oRoJKxVY+mJ4l8p63MmXu4w443W/IAP5oPEgeW0BHE0MwJADk/WpKDCQ6yXOIOPR
naq5w8RJ+6JyYHULOMq0TAMX7ksrGP9uVOYctKCanEcmbSd7Dtpth2na7eknuq/s
CbOi+mP3QC6wiweeoGXpxGuNOb8RsLCnmVnWZU6r18a4fGGRvczqaCcxjblXWJMy
iXz6/8fYkAuHp8Gy7bPzKhLzQehtfT1FYEPZk+BmdsHhJ9O3Zwn/KvRP821MSJBS
mEpgNt5T3GHdldNfjlS4SkH5GGNXEaTInSje/p52F2vOfdig7LWa+QZ6EPhz0gRt
av4kKt8GTWac1Dl3H/uGL5Zhynzvh9p/mcWE3k1ZBP9dvtCT0E2/e3QPktlVKIYs
dTJtsHKNjtw4fKaqCpAWsVgkyCIgZQmSI9hctD0v+zmzutRt/5ktgjCLUWRXayFc
WNaTLaAn88bNM2cpsXwMt5faRzj3cjBKop75Evw8CwUMyaf7uDNnYccvOB3qOTls
M6+10+LtFG3xQP92VyA6YH1ZNTiwOlBC8ogUX4KML7HGlKstTHcym7Bq07nz+XTu
NPQPGZ0R+FZmnSZMzUWZ2GYif1iE2yeUd0QSOHyKr7RQSCHT3tIHaLES5Jfz6AYw
HfqtjwbEWmzhmQbSX6pYwVkxlOZaL5PVGlvh1M9w2XqBd0u1iY+6qxKQ74zUkKa6
Dcr/3321A+jgT3pQj0gRFyp7bykiy3CLA0uN2lWOX918O0s6aTECBCVvSZtidLhY
03oPhSJuKBQyDwLp6Yuzgv4978LrB0KMeNYRvHi13JVjDmHxvGk7UeiGZUGQ0CyV
BkKSeZ3g21YfA7vnOO29hEA0/wtKARHQXUQ59UEyVUETFxkEQkuI+tkRGvOR5yOQ
Vk9gcnqiL0aVyukjzOZQrDOVVBdaW8MVSl7rDl7VWl4svRBAgm8i81OWdT3cFY6S
aI8/fzJwwuTspRtVqIqaMvMTiXnRG9BtJs7czuLy/NzABY+5xkOSZrQs5srv+C3C
ycNWRnzoOHtpcN6oU1K/YngxpfFBNmurPY0p6DgKbl+GKwJ1rXsxRqTTTaEZj5Na
O3ku8hbfI8BV4d2LtiNE9NNdoz4yI72Y8wPrOk+f0CIvc4WxVKoOqZYfY/AoYFuP
kwy0fxo1PXUKj/kbgLbFk0ct8Oq0fzfNPpcoBRnmFclQdGuBjajhayZ+aVtkeArm
J1vnbwThTYvf4asL5snbd+9rxDNRSxh21V1tjaCArIuG0F0hZLXaCfiZOSZC7fEa
ZG9umOLnaR/KVizQrl54yfj+qJmgAuIlHVFCMI83jW6a28Lo/u4Ud1lnhCV8Gnq8
eZZ23EkgRZQ+mwQ8OqLIOp6sONtTQkTaYdd4SjpZCzh2fcYN6Em/X7A+POlJ+cAR
UzAkZAU8gqMLa5trkiuGWj0Y9vhA3WNLjTdtpkMPH7I7Ucn0TgyO+pTvsOOp9Isq
HswOJzsExkpmEutLpv9xVwvnIbS1sOV1Z+hnWCgsyUpAk/XvZbZh2I5VRlB0XM0n
eIy+wNEE86WMQxORxTMoPtGtbkG80cGIFwIMo8+f/bq0OR0ClxGKYGWBtccEcyZe
VBeNLTHG/aHW5+/saSWSekPKfowJ+1XxfzzkauXepZbc4HijLGvm/rITIkO1PIAW
PyNyP8rTO3dMsLMJhVKEb0kIwdo5gHN1yBAyY6q2drAEgpOEdVx8NZ1sbKWLOLEr
gv0hnWMYgwARr1lPyLBQ0bCN3pY2vPSsBGBmaNWOSCGnQvQ43mKzlUfGWh+kxg7o
PY8uiPEcN1KFxQzzOVyYchl6WvY1HS8bMMNmbVa4pwMp9sqC+dkO3LIOkB0XW6FQ
/NhKv9lVw+CeRdkXD/0c6VguEz41HbVHROlw/zFZ+z8SbT3KlTDwOZEUqbmSMB2T
kD0U5emLEAKux2RI9W0SuVXU7zYNoC9/wRaqBvYNmXV6P2TrsTKxM/aZqOIkH1Uy
kkWFKS04FN9Ewiy6LScqMRB3W0LXjToCkuJR7kCAc7vrCHv6bKRHFVR+LT5uI4un
oIrKo1eYgRt9Eu3aAleX56FXWe1vrjtT0al4rTGLeSf8jvS8onwsut6YJodofiuO
UT3/wNVXZu/PQRrj0AnM7Itu2z8GBocwrufGG0I77NVZp3+uPcV6QWOn2Lezu4Sl
P+YQkygQ4Cawv3SmQspy7mOQ6z0S5n8B5EovJj4zayVzjIOvi2Ix1BbdLrtAXeZC
T7L7PwnmhJw17Eo//F739zx9C9zsbuleZU0OKnq9Z/gBMdOjURhkkNzX0osEap4d
8HoRW68Dg1lwlX7dqi28Zi3Qqlc8ZN+7R4rtRaKputU3NkqOqzIhJI8QvGs/0shy
KKan9j2eO3Y1cG5Kob0XhfBxNgwrhROWoQd+9VH5GKn+qq68zOY0j/w2XEi1atdP
mB/nbmWPbaWdi1yH+/muMbrFQHI0kEkDiAHTpP/IdIv1wMU7HtmKvB3CriEiG2/j
TOh902TOQdBvoeRKKCtfxhCS+q7n6uF24PzCd8JuwAvKDoz2u0q2nC7Cp/hlBZRc
03qoAaSqghz9fz75rFT/bHlkJR/AoLa4q7Gxx0qtZCAcWBt9TYeaRAx7Ab5av7mk
iu4YuK0l5dSe49H0qwLaBUpjptLTAzk4tegV9boQMm95gc7nPyLXDOBJDKNNxQkD
ZwlntSj5Ix/S6vfmMBP3B0EHjlpFdJrzxNEL5Mu4vvk2tyNZU3IkAuPynRVLBq5I
tgSCDlr1aO1mfMrfmQ26YCjT49DqL7URnBHnHpKrTdMvrJowzFisW3hTxi7r6qnu
Cfp3q7nnfMoj86w/NypykXp5xlhyQLwgUDyXZ69wr4hZbigS26YBV9iCtJbMXOAs
u6TfyoGps0p/u8XYzILqXtipqHHxpP13eRGgZxzMnh4VZlNk3R5lH4mGPDjzONQq
e0HeFT8iw+2wZuUHsS9W8psYfL9hqgste+Y7MFanvv7BJmCt2ETKtNVX/PnwpiLd
ibhhqIfMnagmre7PyX8NuLrIP45x6k/zwJefxtoCPeCH+dR1RffSretvhXPChgbc
0RV741+fiZxLtdXH67bNdLSs+cLl1oDuylS1plXov/Uk3bilzfiX54Xptb4jJZ2A
Px0vH8HI0e8p4K28Q91eTSJ1ZREr6/9VtKQq81LRTR6NIeziXbkHxKlKuPtPouRo
sp+dBrsNYZmoIzzfh4cjkUO5401eyHXCXLOC1Vzjr81rIKno83bF6BYGk+sgA5tx
R8hYBJKj615eqhhQNyTU+WDGNIown+DvGKLC15jhAqHlppRJ4gLlt5eWrkDSDtu+
L8JAsWlbVFuyf/XJeF3tXPRUOVqH24CNxTWivTBR01KxTEb7PXywgEVo+EcFHnwp
TuS81kuvcSPR1ZS4BRs9DvSaknJieMirIf42hrjMXI0MruIMXM2F7fKyQ5qdiEpa
pdbKJOqUes0wj/cqlFtIkUoRpqNljmGOzjbz9V1aha/8O3VbqhF1Z2pYDbtt3hvV
IE0OrRYYGhWn/j3cB9tKhwFP+dFITBQcQowKjC5HdL16X5DZ/teoEpD6axf6wbQr
ihztn9fceBabcOKCBD3FnRx5ZScl2kygRTrxiyVBe8SwCmRAhPpbCsn89/O9CRZ0
l7atFjia+8Mpx0cvikGyF/2jkpIFI4xtayN8ubsutPhwRCfXc3zXW8pirUnA8cWZ
WHs1RBC3xw8EoTn+M3e0l/Xq0ftJIrtttzAViAS3K8goNdjO89KlO6rjDRLVtqOs
4eq8cpIgjnFZAdBnVDDHKa+WrxSq2DBJp897zuadJRaavLApdY2M36byPcYusGxz
G7QZQeUYx7AZ0AHfamHmpkfhp7K+A5Hbk0TMqzn9Hw8PjLDVBYuBRVNxdyUITTVX
WzBCrqIHL1Ss6m/YSCRDFZC//j7AEqArK0ZQNeqowJxgiIScbLALAXicDKMUddEA
+o+3gzb3+8TJK1TcgSLsEpy53AovR8KAT+DZP/E4qGLGKioy5Cbhy4X3uv4DNr0m
xAGMkWpHsEZpaNNICIeOEqC+M7mmE5WtV9SNw1ejV+Ljk0oSKGTf7hNsjyu/y288
n206a2SmxMtObi5ise/ZlLJscpK/0n+SGHdYosb257F1sllUSFFGCTW3j2fsP5Gr
ko/MTpLAyO0N5B2Upei05UzPzSxnp9ieLUL/5sMAcpq7goaZcRVzU0xzeR1Ygi2y
Dw0cnyLY9CTkA1kGWbjQBDJZgrXlEHR2K7yBjF8KoXlCNT2mxNuYm0XbqwbwCs2z
/Y3ZcG3vMC3bw/KQBflMyhT8Mj0PaPoyzEJSYKPmj0Av4MgbJitvCvhIdWWoYS+R
taIW+oxbZJhmrBOE0ur40//Z7h0pxhB3eUcuIBUxq5tNxaM8wwuk+0CZbzL0Qb5b
6Kl/EaRtyKjJ4+f9ZI9ghSuHbZfVkdA1GIIEnDwWJt7vUsY1eSy1V1Cw/D4pLcrj
KyB2e3XTgIl404Qry0IZxgeW0/+5sHqYdrC6w4adBc8CRzO3Kg0dqZajIAwWkLTX
dsY0BrpJs5d4tcITs+Mce+vi8R3WyU9n+H6k4dyF1D8ndpDWYGruZ6znDDKF4+TB
lJ5ILcs5SIYAn7k+PswuuB8vblYxc4sibslh+3Ws0L5anTjYRRDSC0J5zUxUS45v
qP/dL706jPSjP5HL1tjMA6/VZMk0BD3XflJ271rRRwCmmuBZTTYHJZaclBh9i6+c
w4NrlnDHDeAkx8yONVOfX88pCiQlY47XsDGQnx91W3dhNdiww5MEQg37OhRlKvsi
81y90V3rVnOt1HzOD3kxH5hEEaLi3TSYNP/eQ+Ve0i2Lg/G61U9UKndpafjVxsTp
wugEJO9CepZ9AgsO8JrRSotsg21mH6fqggygmZ1oGqcLRR82W/HfJXKE9nkf6Hqh
6DeuNplb5EHDc3eXpgzxIIb4dlM3RVLv8V5d3U8JRwOkUVgozTEqu3UwYnpptt7p
P6hcHS1e7aP1Zuc1YFItg6o8eMwXN3y0q0crnzcpAqhpruS04s1hBSoJ4WIRubDN
h3gE4E5MxgMIuMVAUIIIa4mhDP/kNe+6QZwVTyVL5PfYiQBuEaFJqcgwXNKV9/KV
qVmppO+fGm4rn+iOfnGnwUNSQhUpgyW0X5caYtgC/EZ8Qp+hiDAfqD4Vs8DfTZY2
EmMS8dUX/RtsNH/pP1SAKF6dM4pdu4avbMrflGzll35Fj4nujHtVaDx0vUrdQODD
gwHbIIY6sNwtvDlCujeGdn99VF3EvFdOQLjADSYHx0ZFL1zVJZbeKEwx17G5cDlp
ce6fsZfkiXT58wla695NYjiXj0oyF7zypcqBPMSKBWBXzkg6zVTXF+CPZDmBdi/m
H3FcAUD2ASiGYwcZ4hKh8leOw3GQ9LHAKNzR/XUJztROqZFC5HqEyhoRx0U/N8ix
p8LX6gTK50D1sCyVLP7WU/7uWcyKb3aFD36QOAicgii2R+nscdzUm4Ba116lpdof
UUJbCaWyHgh9BUn6O9xJ0mE8WVy8jbJdkIeo6Cw1iAYC/eHBv6Peii/tdJfzN+zP
mym9f++Mr11SrEjNqS/eQ/2cyWeTRIKIvFcGko+YS3tuIul0Xj35qsCpPKvWpkOB
yxfEWeZcVZPKsHRIPmRMlWogQJf7E/x4f/grwbUFegPV/eAs0t4XHAYh9JRG3Kg6
FYBf7JxviCP6+FN2b94BQgC3T+OoRd3VH1BSp+prGIZnrLvL5L2ICc0dl1bo0Wti
vD9SSAWZRV27L5HInLuyolqdq16+5cbc7bnPsJev1QbsetQaCRrXYplyTFkEZerB
qNBXm4Wztr2uCEkc/H3g0F/NkzaS4hHdHYCQld57aF9W7cv9q6X+FfqbONLk3eH3
nXYMTVo0cQoeZ5qbC4ihHiogZgbyplChdIjx+UQi4QS1tXDwEpd92lyCk6Nu+2hh
HUzA5yI8LJylBw/r/Djub99RjGSViu7Z/tBIOvQqZ4F8dhXasfoJHcPNOw/mR64A
80l0KzwB3BAv9Y3ZAIStPD8FWCGRiCoSfEHsvMqChw+vAJ5+3c5mdrabpTTWyRWf
fxgpCIC0kFANj4Y9IcrNEZiLAvB4EP2P+mCOQ8QerFNA8AEo/CWJLB38CFwJuj4i
usILoL6rg/mFWWRXLcAb0P2DJndqSo6/2+poQgmW+oYQMwooVVN8Sd20lywbn0Si
U14AnmhMMViPSv9n544juP5C6c9FHchFYgShGpA8UiY7JZgsLuSq4niJlQNOJXDt
ZZWSE+Eq7Wbim6MJjxUv5M1QSbWJh1o8rOTs2iwrAJkVnApnawYrXG6w9gaM/t6R
vE1bECK/+lvlWDdVwWOIQT9qgttKjQKQZBShzmNwe3uYCkeHYOqya5ZwrCorSjq+
38r9TQBrITmLLUaEDHwTTvWzKYjpGMB4N4ViCTPgZqxoY8UymLaF47Q5UuIACJBr
JVilMeP3s4lbtEpeTTplGOJg2LzgU8s6DCZb2F2NQ41yddsHyP2ZT+5srarBRPkU
UqWVZ3nTgTanDbBn60vgKkljsb+Yc+eC7E0q1IvWAr7qmiFl7b7APIzJM5dzX39g
tiHYOX6fov4Oh3GPFF/nX/eNLcZlPo4c1b+QLW/5SGiJO226JOiY6rzqTUJQMXFE
CXsKO4lfc7A0bD/fLKV7VHooPa9rm4WYDqYyqdSwDvGBr8ubYcvFnb7KeEbxmhAF
Hi28uJ2L6fFn8ja6QDJDsDx6GNhT8q37kOabMhCa8t6Kou4JcwxhALShqJI9vcOG
RzGut/jmhnf8PeU6Vv+ECcYmHf5mJGJpAmqeQhWGL4EhwJUhH5cyJ3Xd6i3tBqYi
wZ3x6u1h3qXMoNPbzHYMh6AJrLnX5cS/gKTqw3LCoezQmqnnmezEzO/67WsY0TNf
z5GEpa05sgBlz8GMe1PWUPx7m5bg+IryfH2cbWfcx3apy2CaaTScOueB8AvL3XHN
tBV7tmBF0BobiAlJvfdTxKdKKqaeFl3fD7ZRfqdj5mM6YGjEs+CcNm5SgBZ/MpYi
AHsWZKkzNTyOQs5zmcx+6IRWwtsdw2Za0Ypexzp5KMhseS4A5DZaqtFdrw00/Nqa
zKktrZ2WYFGS6TCFw3jb6BeeIQP8chg1HRyp9vYVj15b0UYcSKjlSu7aM51KuGM/
2uFGTNoQ/XBqMaik3RoQrwwojzhZnoDGUDFXlLBVs+l5bo8lwGUIGFblXKzSDOFo
BXri0A5wFWJd8XIAj2R1efGd68Ft46ZeiaFC3rTgWJNzk1XoSh02xxZiIQ8G5kaH
cMPbWghX9g0xfXk/bq57bQFXycQR2LWje/ADcJACRi6/GJ1HAFGsvPn86rcDqkno
Buz0RucXxEMEyvxM6XLrsVAgPJQWHCSrX39UHxjzTMd3CvU50EZNvwg5g8I7rNhJ
ap9DdLnUV52ZFlEA3dGH5olhMfWWMi3WHfzapat7IV4GXhzcRsJv12e0adOOetVx
1x/oKF//T8QHN3dp87yUKl9lQbeqU90AEfPfgAaFcCjr7wNnSMW4fyddpAs32CYf
EugyTw7WKjhR5kbYPNPBWfSbAb9i9x0uknlfwWX74IhslWNZrWn1Da6JBi8cUPC4
7oMDJ4tZticFacFRJGYGz3egTjJ0rwNlfkk9fVrdUUwokHhcNYdiZRyzsYxaTcy2
YWc8XNe+vCf9TB2ulrj+A77AmugHvu2u2/EJ47CMbXecfD2FTmu7ThLdhle+Hq7E
arGwVpkES1rtg/4GUhinxbdmQRxKBYaVkfWlhkhp2K7geGtNHnqBVXPJ5yUyYRKU
SPxakNk2bzK42FqGNkUy1nqpkmsM9qI970RsyO1MOeYF0o0XYbjEa3IOFbf3cAat
k1AfvFz2ykF9AK8LKE7+EQjPx9E+fYB9d9uILzugsFX9d8MIWLj8nfpxAfIMrrbU
r8XSIhWqate20yQFOSZZ1km6gI28sNmjX9WBSzC6BJZgBV5cfNUzBzm6ADrLo+s9
uQZ7XcvkV8xvnMw3a4s1WGAGfcoUpRT3VZie+2o1ggZkpZZZA2yn0NTHHE14wJta
PwPGaCS08wqBCnfEDShY5UX0xlH4StGKdwXTgRkIQYz10cDjn2TfJdqPqurbNrQc
UTis0ZqS8slsrlzPMcXcvxEJ2k7JLiqhnnFSVeTUJlLOxZEwcMbDpoBJVQKUf479
1l9pgBjNHl0X/Mq6Dy9Xj0ayIf9KrjkBqmSZ4zzl8349o//wgjN1wx+ZZxDTRyzz
XL3Q9bLEmw5MVVF3rfyOOxwBmAk/KvpEB5Xqm+KBxCdfZwojLL/SSlkKREQoNd4r
pfOIcTo7viTMyPvb3WMo+ZdR2y5gZBuvaGcFTpK29aw4N7O6srntEGU22bSPq5e1
q6iQH5uM9jDpAPcjtlPxKbx8+d3Sy8+5HFC8bStuZ38YVOf6TUBRHwAGz8Dp9LQ7
3MPP2yjpNU3uDd9/3+2FBWiZG5waRjg+1xQD+aSbr/G9ntrnIgK67QIgM/376BR/
gja90edfRwCnaPcCA1RvbJlcYBfRfI0/tQwOsZYZSa6A5gHIh838tlPCJWp8PlbV
cw8VfppN0ik1AhGC+rDFsyIlA5dnI3cW5QGRiAqXqzVTY8DMprED2nA8rqy07XAs
C/93puniuVXYF52Nd+hQ7k46IOoB5j/jI4GVzFxhZpfg0POZOE4o2gjvjVzPsOaP
GxfCs1AEryThP0UrpLouFJt7Ha7Cjsj0JUqfhJvzqesVsf0v1lC+fUKBy9V9axY2
f5GChdJMstZgk19hWYFLDFRBmE8ogfLZC/ZDEZZdqXMwKM4zvn9ux9ggz9lPlhjl
O8WHYFJpuBNpOCbH49tfQ8NEz93vrVE5fQVr0YAPcPSF18qW2LKlyGtTcXFgCfi+
+bCygjbwGEgjfuZYS0/ob0hRaM+26HIyHuO6DZ0E1myGfAxd4cgm1dM+GabMlD5W
ve9UIEyCWptMrxlyFXmrc508xeS2Fm62gK0z2EgixW5cLhPwaSZ+Ugzkvs/fRQXF
rOzSst2KVNFVACbge39deq36rW5WyJqm5UDAr1e2/Fkb1r+ZFIg5t7doSmumaxew
v61OmFxQ2ic5t4WOKB2CxSoxg2wkr1QjRIFG7lO3X7r9cCmidlzvJbEIMX0ElTdB
raDsP3nthRwoaM94quV/pg==
--pragma protect end_data_block
--pragma protect digest_block
zUnvRXv7lQF+xlf0XRz/gA3pvic=
--pragma protect end_digest_block
--pragma protect end_protected
