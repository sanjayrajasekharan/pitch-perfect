-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
AxWC3c/XpSGKY+gzN2FqqRrTdfL9GOcj1Hn2emvYfEWKkqyvS+pgydydvyD1DfAG
lRSkZPLPRyxHM11+euj34hpRW3vd7EJcVOy8pO+58S0VrxMeDU7zBiAf1sHw3WiC
Ohdv8I++M8RAe73QPn6euGcfnAvVswWVZPuWNny2nb8hW1of5uhRkg==
--pragma protect end_key_block
--pragma protect digest_block
YtrgR3cy6lqqQmy3B7h6CLVFRgg=
--pragma protect end_digest_block
--pragma protect data_block
MnBMh9XKHAyVRIyzk+IpRRHXwrvAaS2PuLVRFKjjSEY1U/DP96eixfyI25ciTCiH
GLjUiTTKrD/VNXm+fcL6Ph+GXDLrJ9KhAO5LI0sWecBur6u4mllGfar6DY75X2VB
aJ3nuJF39aqKc3bdT5ozSZB3Brhqz9h1SxtUB8Qn+E57QM+a1qpbbieZ4Rj6Dtc8
uJuLeCZg3Nwo3P8Z++hXXHmi0SlEXM9LnmqAzd8E0eMKq94qirIeIIA39c9+0I7x
dHQc65DJIyqv8HXHrLlxbfc2ZSOXbFila9G9J0XxXuT5CW6LI3McpZCb7EX2qChN
9vfrOiNxgyLC4pV23zHi/cktJ+GsccD/QcbBXDtRUi9/d7tcbruuajCHs38aVMjf
o//SNQ9Dm7yHztp3NhFGX/NZFAF6UxCijhp8BNjE7LGPnxlxjv3zvEdmPREWFYYe
s8MO8iS1iCAitb9/vlEN7h+KUlArBqwsUlCjVfDmt2IaeuW7blujKhEY5+cmQuSc
STE9OxlGNDQdK9tIdr7PLmyXthTffMPuPZpopLO6/USQPbBsbF0+yleXCTwjYzHI
GLfPqgrYtmlW40VqcxZ7q2rAkGQjIP4MqR3X0gYD2AW7LgYpjlHT5jsQT2mnTyPE
HmQqz9YRnE99W0nrFP3A4Z51f/jDMB4bsNCs7ewJLYpda7MiiQkWwvcMMu4h+lFC
8b0N4Yyilwdl6tgyqT0umLZ4hur3p7xehH8Cge6mO844492fUNsXGJAhLM8iNo27
LhnDmuAmlI9Cr0gXtyM2E6I9D6jqphIIdOUaX14fvvvdez+s8uAtRAQdHJbhNQPH
AHGrVJQqwhEoAnp2DKw/IHm7LhbzM6QsfG+HuNhLuYtfDAje1qxxK54q06DsT6Mn
BJMP7VcQmNP1uE0Bx72KJy48mMN0gRz/AGZQKFlgx/toFY5RWwhsGYQMWMHxCCbH
joe3jmmGlcyzwmydsjXDwDYJRn5sbnnWLjE9EtecxssZ/Ic5LBM980qZHbWsp0BJ
lP9EsCSE9LT7TFle4ZocpWxKzyKP7DDspmARF3bdgsHU9qAU1BCziD3woCaaeomm
IlfAiDRv3yWljXjFWQ3N3GusJ8RIEb+G38gXRGZiAQh+vcq192sdVRoyqPPVvWI+
qt/U0qpMeciRB0TKVPYl7tAAXDpc+cUcEJEGgSti8pxUmNQJoLpADepZ7Gi2GGbP
MTxEGTdM4dHLS5LR2jEKU0PRiZJ70iAFYhx8s5OrAOq1+C28olhk7s2Dnm0KCHM7
ecV3NM69Rg7fEG0f/CMayvTvlCeEL9l+J5asN5vi22ftFphDsleSzd5FqILHwGou
rlgtmZEZkUg0neTirUTZzHLVEv/Coe8zsNksdkhK8uSAyLcrVcr3X3VFc8mQFU5I
uCdAWeHRFeYLHB01IWpqM+gDvdbAiZ/QCe9CIHkfc+yvJ+EFKN+bAAAm/zCI7QLm
zDMdBPTT0PZ3hONXayeTGRgPLI38P7AJ+los4L7d9WQSBh10Mq19IuCyw4tpV3BY
7+c4ndL/ygVVjzbvYcqBImnPWwPw9DErW75u4JUHbirlN4mQZNw1+gnaLga0FW2n
xpKUGa2Un/xbqPUe/2Wny0WiPsZucNkRLKEMbiNkvrOJ6mUOOfcy/coLBhAO30Bm
g1/WyxPH1s/hdlGhwKOre3PUidjdnYWf9JYDyvy6Q/+3y0WiawMvv+0X1HNGHWi7
5liW4kRzPi2aUlCZjDmTz7Um2OkAkgjlvdn6M++Afe2eyu+l2OMW/o3GwK5/DkP8
7aYfmEsWwqzqf+W/Le6u+J1fdUCWFGxoJtaotRiXnYS21pCchbZp4eWLP3pVdgtm
Sdtz0j3m46sxGfOvuGOHHAZRY3hmw/g3lLfuZFvueHVm38f3As3Y6Ejt5y9tXphZ
X/g9dg24Th17qP/RPvNlWNwDF49mnoNkEta4VOrERIJidJzvscHLwaZI+zh02Uto
zha0Fix4kDJfjxMBH6tJmsdXUMY/bAZEskSBCN2PCCBL/Qo66ubziGFu5KaR2cki
wxbLtNg0Z6JK3B7P+oS+nUSKR68qZ8wpRctjHGkMitQmmxJMCY5+t2gl6Io49TXG
pVY8esHqtGjqek+I/LuZP/XIXN8n0HoPzkcVKypRhF6W4LtKpLkhOn6xY3Ae8Nlw
rhLypgMHlqTHYtl2otQF00OemkitZ5j1yXDmyZV1hBNzOCPkE2WB+kG14x2mPGzc
IfayBNLNfUbFP3/A78o7yZIMnqftunRvfUUsau7Wi1sowW5eYGk0+UL9L+HAXShD
Yb5ltTB0v6srLpChOSWkew1YvBIetMZJ3XqKNYiSilNa6pAKpJMeOSPeW5k0xW3X
WC+xQDZXmL7jHUoNXLqRDRqenFg2RgupFtKKxVwVq2AnXTAnu2RsiYF7SDMxkjBB
8zg6SWfORsjxi1yVQ0F3A2Om7cbTRmvwhoyW3tbziOJ0X2erAeCmsYM/Epz8bUUw
3YtQZAOTgeiB4MSn6b5mK1DoLb3XwzNvMJFDkoLsWextHTGk7WXByu3KEpx5Y6Iu
8oBA47VRzfL0adQniW1UY8O07Xlo+NWDBavJP7TW/1/pn3YADrbnase5CzV4sUA8
CQodVEm9m8r+Ff4tyQ2ikPZpo6beASCmrgsyAczz7FeIhPwwlk7JCIKk+P1n1ZOV
mMrt6AOqXR7yrW1Je3iMVZbiKJuN7kd1CHKVniNpt6gdkTCkXfVQL0rBZwFYVD6f
S40ugYyMmP6+xjxjbgL820YCPxcyTu7wGyHLW7nZX10SviZQYuQzXgS/tP4J78Y/
m0KGp84LKfzSQjP+AlDO3HWwCdofCAizTEdi0fg5bvmnQw/ka7cJoDXMMGPLzfJO
jFSGrDc+RHwEgQPcxQgFYyziQgxvrjpeF0yXXPjocTI7syoTuFMvriBhFTuthHMh
+5DgkDsbwlKeC1RHfNt+KIVLR93gN9S8yfQXthiFs7pG7EhOioDW8jHBvWHTGBNS
p2H5fu397SEeWJMbB7vP4Gzte0DwY56wvoImVkuL9o1RYSdgI8sbAKv8p+SCZQs8
Gs0YdEAg5HTnBHeZc06CqKxUSuDJQD4prlxahVtIYZrSRJ/NraTyWZdH5eD8HMxn
zI+0WGqwQexe1AOc6X5E3lWhDFWjBH00W9/IRHZNwzpJp/RbUjLDdpshJpRkMnyl
Z5X1zLfbnvKtuToBMl7aMZUheWIWNN6TlV06s19tLRqSsReoZ4+nMB/G1OiMlUx/
AWHI0Idqwom4GwWW666imDjjX1T4kPk9J0d8FdZqiF/MRzB/DCQy7Su53uQO6dOF
LirhTUr+YG2WVlVv7A9rouObFSTgJD54WxZKUhWeylCgNGnBiAJvcy3I0NcXSv8V
36WvnDeG/apIk6mlW0qDV0LgEk2N+DkbTugU89q43cd767/kH58urmzEr6XeJxPh
ryjFH4HHeH4NXmKK+sfW/k+A0BJGrMXgY4vLF+MbzHEAOs8R5hAHv4ThvI95aolt
Zxvm2mTFIaVD+xuSrIW/vOKJYhYD+cAJ2Gi207aSDpfo5PWND3Zqz7yGssFWvhJT
fwyK25fbwbS34lqPbMqMhUlO3GcP03ynmob7wbI4k2ABarl/gFgbZDrH0UPpM4CU
4VTmA4+v5M5zPAfaVFL8OXJacve1vnzG53AjfLZXMeDPJ9iy8B0yVyzlq4D2FzgN
Ic2DuirfraLVNuJZLS7BZQayu89gBWd3h0FUxyJidZfPWUa6Pb6iD9pNfYHYxwAO
yVnVHdjZu2hufjabPCjuNmRKovMP9HP+y81APc3QVJZJneOiPxjwxJ9xlfn6AkKV
MuXneg/7u/O4U+MzaJXU0aSCLcZYYk135WeUJ6vBoB5RwYgL3gmfpGXYc29JMhIK
18wu72ZZPEUuF2VbjTtZRB7Y+0dijaZsSPdhm0IU3VNhQLcfmMPk72LHcHVRNvcg
wQZ3/hTLMM0p278GSduaequ4n0tEsUxz2SWGTySGaYqhH2FBoev/ks9O+CxfhJ5j
wz+ex1JmJvRs+843rDt4la3i9mbJURiAP7f0nx0YqWtDVXFXByE4AtXorPhpCEaq
ZrZjgGapRKbdbAPy3Ff3M2oJPAQlBTXHrK2QEFFFZaIkBTBotTnvqd7dJEkvMv1H
qnLuSAH/E0yYKvnZ8BvNWHr0Q4dA9D41UJdLlRR4/LnASzQ4xG0IezpSEtD5i3LR
iR0CP3ya6jB2SQcgBCk/TOlAC/brDYb3Q5PTRSQ7PdjcbMA71DkKSnRn5TqxZwSz
cZaL6XmVcmX33/BYpo3TSdO7wHbkFTMoHEhKNVL13u/O000WM5y6TP1BLJym/JNo
M+1hkCnALZqbE++hGnS69CHL22zB1Np9+nhKglhBZxtPvICHEP7VFmZwZx4lU1fW
ah9yIbNTGjyyvq+Fueypy8qTDZkPptD4WYBCgjHDQrw5x7GsA50kC4Ug1D8Ioo01
kLoe6AbzF+JZpRf5SMMYpTHRV1sP8H8ubQMttJpB3aCGAIAJbQdTqTBE3of1CFk5
pDbrtrlrcovW0Oa6GB7wFSoNNIBIOVCKVkQnPJhuNTUUMd6z2Wk2Ds+uWHCW/PWE
9c87+z8noHUdLCmN33VKCv3mdFj+J3tPsY6VRY0JyaUiq/pYO9pMo8ZiIIJO5E9Q
WtIYChoXl0UOyX6Dv/jyVKP1zR+IRsAUsrVfFUC1HUeNVf638jMebXFmg8DL9UcO
D4U0XxXUOx03WouRSHeFSAbxRnYcghBI1KTWy3p6wokICY+6ywCrh7Gluvlvic8H
vEF8h1pZUj8j5XLf6FSSIYhJh4rxsqT9r46Y/bs8WwSuuU2WowjRNaEMr+pXcRch
evpIxwfU0Np3CQwDh8lfee7k5XyMLsMxO1i/9r38JDZWziDPtKv2GSj6uVFnCjVm
JQPazbP2u+xBOqLDniQK6yaI/85H/woySDKqv+N6N9RMqV/EMtE3800OaNGzsl7Y
LYeMhgxvGa+SVWj09UopsbVrP7b3dGudsDEOtQXQrkaAgDl7efjGXXXF5aK+ihTM
3WI0unHMkOkCcTGF55Ve9MUhczkzr/dd7W4ehSZRHTdfB84JYqcvqsBr+DFNWuCe
1ep4XaWTO6CnPUwYdJi9fvVZ8fp+g2DAnv1czb/taLRAaclEvJFJ/uvcmYnPaLw0
sMlqkRTTxg9Ag8sZsVfIXz+tOeOcw03jMyZ3UQvmtYP/qMxB47HOvGS+YMEFj74E
/mgbwYnG8u3T9+fDlg2zw2Ean0eaCYKyPE3HtBV50n4U+giFHFxl7gnDd9MypyTr
vUKtApgECtaVrXRMOQjJq3D7JRKjvMcgFcm4/eZ122OcdHU1VOenfAFky9AT//NI
3GyNqDgJx9R5A0sCUYZ3AWXAneUHbK4KJ/kXQZ7Mh2dSS3tDMt2wSD6xmWvWT/og
gYTFQVFXjIYJvE6ulEk03jOZL9bareXrSQ5oZKmOZHJtStLpM+CJB283GctXGAIl
Ndm/0ksCl7lDvl6GhhZFF3kuXwXbjy1g+mn8OlvYMdMor/3g15xU/LbqveIrMdiX
UbZjFAOtnok51ozbz0gSl57pY2yMcW5LAlUxWs2i8ctJE+70W/CzBO1GjcEBi1sB
pD4N3hlL+sNbvmyVnSGtkwUWQp/gXEFRl1rlpviIFshDReahFn8Kw4ZUYac4831z
Zs6yhDQ2U+F2aRWNSfgRwfV0aKwQt6a6IyZtLhcPkZihnpCcpa44mJl4UyIWzmee
7l4+Y0jD46RgPz1VgyRoiMYQk40S0CjuBUf7rS8xSyLBNUyZGSpJf+31y8gRWGDy
v+sILET6vaER5DQeYJLWBlIsrpKouprqozr9qpcSAOMHRIC2vWP3qxLaRwGBgvrj
igBnq95blZyTcQ6sQIZaGn0P0sJ97CYxR7bIEl8MQRBBU6iCa+hrmUrHjY4KkOzE
2IlQggwU/R+d0NHOLwa8FAaUDAnz7akkijbvlf1IK8/VLCCpjPZXfOWT/EMiqSfC
o7grlXh3mLgdysx7DKwBr6h8B7sBsb8/FHi+bH4VelB5aGi2hcAheknxj7Vdo8kq
Khm67mafW1SFATamDFQw2DycZid6sFLs2HfVEZStAifYTmf+E+XySi2SFfGUOmIE
VEcR8eBqYndR6sb5Wqd5owJRRAHE5jeZTdA8aqVcAMNvYOZEWIx4oUYsMi2+vN9r
KC07PJtmZzud2atvAbFiZQ65nR/FsTq/dzNuwQBx9ZyiewAb9nwFJdyUQnqNtiDE
vni1AtwR00jTEEvvXuWlAYVG/Pz8YrmGe9DoNdhke5TOUsA+rWPHamAH2EM6wZWu
vjq2bWwaBWgG7vre9yoJlpzMJNQt+OswHr8hbZxUTPRabCjHQDLahEWGnzrMw38G
3I2BOd6SEeoXHIlQuVsXa0osRwerhsMnD5rIgK9F7OsgUibg6iEVo1r3DDCXdKSl
kiZIPrQaEx3SegjOmZE9ibffZLB9lDaldGmO4ZkoOTt2uKzqDvYBZ1vI5yV9Bu87
cJUioHrhaeOyQ+gzoa0qfdkF1nn5SEXbYFA3NqMFFW9/urMedQF7/XUcBp+VQXrs
wJqdks7SypCnTHK/MkRqgGKcNSXakBrSxsh1HGEwKsCKEA2uFQ8Wt2Vf+xL0I7Nf
d4YHTb6R3Zj8hTBx6cYwzARuAtinDxnTye+kiRQr/ihqK54u7hIJgby7D8e9H14J
1mBXiVfCofMQ3ItB0QGoljDnEQVVWk8mW9xQbaYf2E1j6q0Uy90J4Y93sDzdMMnv
hq/ccFK6twFWACWgL4jmSriNrP4k/YhC2XBiR+Jiq3A2LrhY3cQJ5v8NspH0AmHC
vxNnA67Nh5yZ5QAlsToqjlUV1DdcUVTt/IMUFpGnubEI9d6DLhvBe7cv5A5b7F0I
7C1ApFKQhQY1aKRdxZepb/DBuqNHUAoIICs6IBh/mkDYyfsUG0GwqauXlXooDJce
iv2FZMoY1STRkhLVyTpksboJOi2uykHftf2cx4uKMCxeedq6mQCySHzhsAgU7pre
yPUda5c9BSj3D2enVnBhfBrZxi6kDKyZ9MWMwz3mCChqpJoIeaEqj3WxIedoK3iU
vP5y40DxUA50eNWaRfiPI6r/9Y79hOa8IGQxMICzGEmdqBUbee5SMQl4f9k/ZO3v
zH8jkzF0PJGhKtmb66mqxp3ZWDY83fmIpBV7Qy1fX+Y7owOFJHgPfLDX+x+eIAAr
jIfmXZms/Q9y96V+lZsdatCXqyqdSgzrJH9+b5/ZRWVr/7AUKN5IbISWmu92t8X7
KLNN42Zue2iz9gDjvVl8sLvT5sLWivnMXVcQoJiFvJ8yDG+85Hl+n8p3EzbIsnzr
ddNqQBADPcrq6IeolEZwKrGDarphdbPDm8Ym1cOcqlz2sav63dFI/aNBMVXwZcIe
UURUp3MNLcebiZNcbrZfSQqNCwGvlmX5YhIrbuBq8ed0NNMyVGe47qQ+guwiA+db
Sr6FdisIOf5xhZX0xVewwLtg9ajcGeto0siYSGLo4gBBL7pC1MO6vgqbWTfoqN3C
xByOaI3RiC2bP2aXxwSWIaXh1X58WuUn9TtuKRnTQzWrcCfaH+buuGkyH+1NdEfq
u1BTyZykie96KzoTbXRlot2I4aa/f+7K51xntRMwXIla7x3r9hfui8BYPfuSTOMc
LyQo3YzKQSU9vh9X6k1VP13m7y1OwWSVOQJwQta/QbQBGDurTOL/xrMQ9EXOAL1A
ozu37FZDBD/dGXZzCinZMlMAOaOcYNEqrw0rOrBDmfCKO2xsaTmGTHKy5cn7HknE
8ItrF5+HC2TM7qOV8+L8/uACqomDz2VICUHUTwdTDD0ZaxwPne6/aNjeq0gA9P4j
yFS4qiZU3O/WB9k1Gh4Cnuwyzz3WvncOplY5rqUW7IJZdNf+0231TKZ9f20Ldp98
GKa7zagcnSxNbI0BJaW9lz8oIQJ1uYdxCRO/cKjJUwgKIVtZ1XdGU0kpP5+JBpLp
eJJ7PgI+eKQePAKciI+1vMKoOdiT7wMPEb9MnFXV6ESvDsSjINrBbV2QScnbYZyU
0XMrTn8kxV2pWHt14frk76H5hnLHTX7fcGkZ1dUyAiDjKYCehkKlNY9rbq/4CMSG
Xru/JVK9QuIwX/BKwJbz+ooRUcU/1hhwGEMOzCf/6cNzbIRI530b+b9SGU5zMfPJ
pPWjJN4zfD3NTkgZ0/HNEBr2FEB9SFK5aBSR3WJ3GWxpndEYedEXyuTXX8vxcq1a
DnP6AysK13YCzWGdf04oADwf4u/bopk6u9XS9NMrjaIqDgEFygQw8bnu2hdI/nDW
rwrGRL7tylwjUqYTtI9S+/z/OfTJi6xAhAWUWpYe6hP1uoyak1mA6ZFNZeFtMhRa
hHsGMOBAEnusNm0cjuTNmQKS5rSSqTCNZOHuJfTGGtr8a2Z0Gle1pOEDFSUIQRXl
+zfjO+czfo2aX3vp4fOjGYgkK1tTPIasZsZp155PuQ08r7CF9QbtX8gnVa6cDErG
FiyB5nK+LAqjiuxHVDtP9oDBSt7MyrTspoQ071Hkt8ChZyT00vr22yTZ2HliOPmW
/DRv2TeBWybTqAUOtTNy+PqxZpMlsVxTvSkRFw2ArmNyVxnzqhTMtSoVMLTqJSU5
qL4OKtfwKuIJ66220pvsAVV1mCRT5tE5X03bxG1EvD6x+g8M2Oo7NKVx194imDhj
wvOZbY8uPS7LI2VUfmJlJSUhqy5t6gv3fRALoJ6aBywJuljWmGd5hsOMSyhrJW2j
wSrgPZFeXIB1K/PJlRJe724U33md6jxaSk6xQGJATfQzEaYuC9kRPR4C1WkLGmI9
to7uVZfXa8UGwTI8JKtZnNCMAKjLl2uz0bZQFUEWkbRhs0nsXrnTnu2aiiOh1WOP
L2XKoraMjiz8+Md6+flBVj7HoKWawVjaRYH61EKk2vhKT0IYWTe3Az31VeEmMLbx
Z8jEoYRRgP0Pmuq90aOT7xN11gyFezLCsujKkh4s5OUYfGfuFxM5BqG+ivmefjBb
LFc8pmkTbutE/ihFYkYwgrru2M4Er3lO9oEdSt3ju22QUdxKxxsTAho7XzI+Gpyg
sDXZxlDXkIf6/jUlwz56L2K/rGJgm2p0FfSAcBpmaj/oq9hY6OlkzXW+mbzoCOn0
uAfg7oo38BgPAs4jklJ9PSGVh6Qlb1YoTB4eSAIJanGUum77O92yanQFDyxyFrNf
PwQpFH5RcqApJuv6BuEL2x+UwZIIBSn55+Blti0fN3B8NAssRXDo3+wg57hJZUpv
/CKpYDXWogKYR4DQzPiqhg486lkpiZQQjE+qgdmDt8K/ddlcTFjoU20PQGwnqoeK
ndTyzjCbWbgRYB11PCVxf05O5u5TKOcJOAy+9ATPTrcSq9Kza8yIiUFIBCLrVIUB
yXhyJWZKgsdavB7Zfg4PZKlpSKnsgbOIPv8SxaU8MAmTVQe+6u/xmLsGUWEyHYuN
KMVKWzpMQrnIyO3VcnsDGRdTqO2M4sZhVejsma/OTP9xQQmLRfeDEV2b4ihf2u04
fFlC2eaR0F07H8zETwZ8/vltefgx5Po9e2UWwiX+9qvGBSOKj6nvuqcMQbYjoCE/
e4wyhhCS7beHl/BHzAERQEoyVt2hwWt4znj6W2aJIZDKuuc6ucDvlw4IPIqtAWRe
hu8gzqemaqCbEoNBsod3QhYJhV4+G8SJdvHO2iLRPnf7MYDbjBtWbupDiYb3WDM9
V6Qzak6cbDjN4ByVwBiQ/+2BWQW7JgWpR/jY+pGJdy8zX04AFTSs8mR6OjJpNjRg
WdfkXgypWoKYlb0KQXSac6uE7aGu1DIliz+RPDpBRl8btd45XKQ6aeHcQ1EK9ehi
HmmHxn3esvmZbcIiNHuEwKaFDrIkJ44xn3HZPPnbGucoFYgCfr+YN0ArBCAbHmtD
/krIzTbBv+Ag3uh2/y3W/HIFoIVt7YwHmbofIYEM1dyeKnojUvpy4su4b18FoZBp
2C932WzAJJq+vqcMxa/gGcsy3uvzbWMuv0msNMwhWxwmKt01vT2oYmJgKEFe4h69
y5h1dgDOTh5WsJH/OkI3WnBjOnTxru/1m4Nclur1/KaTNhVmndegOX4TO8yID3JB
sjwlWVdMth8bXeziS0KsSIctLB1mwyTcxu524gUMt/9BO0uA+xKyqVcrQN23zWqf
OB8KPuO03t7DrzoTbc5up8mVz0GG6ceNd5FnoeSfO/mK9jUZLs8citcO7cfXQ4qe
lFNGe47re16AGbZwWJwOEzkqKGUlevzcDn3Y9Pn4E7/9kLtlj0jFECm7ICuaDoJ+
igBhuy9CMgU99lHunr3HuKHrEYfBKepT6Sa2gWg77tQBOL2pPrbzLXmw6deBo8O4
9I9LMOqCiJHYt52qlLq07Svjn9zE0+/D3dchKhrQhFV2oWrQW2tal2pfm+dxsECR
JB8Iz8JlQhSBrYA6wQ6pW8l4t6ifpgua8uNvzmKm8CJ8AxQdBkgzHNJrc3BhFRqV
6UpsRGNKxSN/bLIRqQlDGsvqSjiEzuy/aY6Gcr0gIFnDnD1GvBTdQ9xojqQgpqQJ
ci7JnN4na8rie+eE58IS7j4X7zjQB3txVOmZBFa6/0Qm9wvHR+IPoQRwYJXL3leK
gFuqaJ6BTQDDwJAzDZsYXd/mbFzZFCW3gbSpVfEIRtrsz6p9aSR+6dUjkaWkBD3G
umjS9OOSaQRRNhY2/k2wwgyHabUvzh0AYgO0UrBUQLESTDNz7lHA/eADvwc/yGMP
Pl+v/XWB0K2PGTLwwbgH4p1W7uvZp67ArumKa9pybxB2uDYQky/Lym9a4tzuyDyH
6dYLz9spEBVtZgT77T5Ag9NWMQDID6af5w/7RG7Wr5pCuXerjvhTZtI+PGQPhEM7
OXZsnaPRGSBOYj0VtN0JFsotXxpcCwmJ5TKkCzADtQ1mwYfBj7BuIO2NI+afQK9c
JlYHg9BPUHR20Apv3C/Rj+WPa1j8cVlYUMAXsyuVsPDLmT39UuI3y7LbKsh+zAuB
I9tVn8vzKgZqSvZT/OpPT4OhBnx7tr+68n23ZGMxSOLuwGUckosmsXk3WTEYK/vv
8WJnas/pPLVg7Ay5TUAufPBEt/uBxcZL2JaDtpqKdUuQpuqbq0TPQkuMsNIblwaj
o6JcYkmLShoj4wLN1jAVS72EaUwiFaPwgCC7jzM7XbgZruKfAgE8/SABs90JXkp7
zBajrhFDp6vFUF5DuXvR0t1WXjRdytD9TFBjefTty4hKT/wcfjhbz5mVuPz2f2Tu
aLUGVK5/K1YIefzXxciPiffqKaVhLYZzUi9DF1STIr+6nk9BPYS4bjt6ivSp7Hdd
UgRWdBMtxtvLahznXXrZFPATZrG6cEu1yfZgireiPffG0NG1ME+ALkdsp+7OGtEm
FWnib13MMpnzIqlqaw0C+ONdOMPdIhbipLq21OJECK4WRCZP7Sc4r+KX4oELNByZ
9ln07iwhU9Xd7v34dDQWue9VyFfR+iYjenVE2X0igY+N4KUwb3iTs0JCxdq70TG2
W0tMqJmPdpacemuiivnLKBL+SERxp6q/0gKdEYW28qzIvKnpBop0QQfyTcYmTcx7
C0iko4XM6H/v3Kw/+l8C8go6VOL2dxTvNthvSK7uzbvCFQKMZQOENE+/QpwWGwYL
VK1Mcm4em8ZnNMxDokCJZljiM48hGcvvN0PYr+Fa76Y+8kqQZbluReRZD9C8V6KP
j1Sw4WUQ2aBcilcexOQqkrM2MmzZS2640SWG0sVJ8iW4K/KNyh5qkCSqSVGk554y
PH/C2znM1V6dI0anktDXPxtaWI+x50jsa/e/X7hdwGfnpvExLawCKB9aqPDYUpR3
OAAaYI2ubIA7O9+m756kFeIvVgQB5lb1/Y0YO5HjZGx5cQOoamPZ0YsCw17TRMn7
REN9qQdh0SuaJ00r2tMgHg1L99363+Jw6bVEIAjaNv7fD37SDBUgjiSle+JA88Is
osgl3j0XKgOlLLjMCgXESrrmX4VJZ+8KXTLlaeP7YM0cvPtLqXsAfRqeOCJUGkSm
kzohMzzYMKpBz1SL4gTH+C/CbEJzlV0x9JH78FntCDWGWhF82RBtdK0/ai1g9utt
EfsGGA+LljqnhFakABogKemrbyU8UTRvBU1B/R0DP2G562qrquUUbvoNxICIfLnL
mbkWfdHerR//+tY5u+HU5jG0M6G1oBebrBMLJJP1wuB2b5/G1+aqj6Z+Ztyipap1
43wceIAK93A83Fob3krtLIUQyGXsXPm6ifsLEcITCxS/I0lEf1aeYcmSDFU70zue
AslaeNMqHvKxpF66S1PxRqZSVtHnnZgBWrjbUpD3Wbmxph4KwhhrgQJOOC3FS6HR
HuyBcbXSBwuhPMGEOcNBK11fQE08XusSGaqGR5yEot5uJjJR0QkBT/ZE8NOGcb9E
B8L/b1kIv+Hn+3B2WkfjFRU8/IYrSE45dSdsqDob4OC0VVLCDgXPDOJe15JEysuo
Cg6owA4NSOqmDWb+3+QkmXwpfr8Z3X47Gkx4vKBCeQJXhdG368PEth0G0QTmhGHQ
KTnqzve1PuO1utY7Pq8rDDBR4CXovs8tIgf30fCTSVGwipRyE0wL1qBZCPcAHU3+
hjzgagcyP7rCyKOvIwswDph8VETFTYcRYQueBIOhNSz/ObQYPsS8MP3HxuYdcd0X
U2lv29kDDoRFHHTk2cX9NOkQFl46xZt8KRULRNa+AWOqC7rla6n9GLRm0jrNQ3WH
2XD/NrNk5MHk4TGlG/kxxBq8ji0+RxJPfjZh0/GrEVuws94n9NLSzyTNV/BGILAH
Hl/yvYtLUxwQhB9BFgO6LWJOaeWAea5UT2SJG/Ni5ZaNwcq/Lwlfj6obbJFhUsac
skIjjX5orEtoyp/50GqaRCC1fWUGU/M8B9uWthqIjJzb6nkH6ADIRKCxxFk977an
AVNvFTsFNWKXDzQGrnwnEikyz6E7mXhis6ItDu4KMZjeCJUkprFe8OSBi4qJL1z+
1ziMKb09qbBPipj/8SKGADfKrU0oCFrZymDX0dWtNp6dMqtDxuHmlsxqbo2kg3Iw
RmkN1PnNbiQjJtUS3QAu0zhygjBQuU5BJD9LerGxmT7w8izaSzGMTiWx3zzNhmf4
AWP7J7EOJT3q4rBvTauEdpkGYOb4Zxi+IS7bQZ4fyUcAaWBQ22unkRKDVe//ju2o
TjR6wFL6R7auYDXdNvYTqD8dXsqYaW9r06/TFM7ntrgVk03JhlzKF4KqCveTC4vw
FDRTISYAxIj7AZ2pDish9NGJx5AjsiwSstOZiLazY3xzNR74PaPGubVvoxo7i6Pi
WBgR7xLgoqD9u69xYQ8NoQM4K8UMflPl/NDI3n4eeq856ULOfW/fsgEA3Xy7hZbv
dDFQvUwFMpuBr5yR9nUCpZcpZ93DPWws4DrVdvEaYqalLVNK50VLf7LWJ4uzN4nC
cXUwUK5fzJxh9JW3/DO+VDMQTP/pj9KOLFDuFSaKsCKUQ1z1KNHGOqLqWAPQCiCK
BC4vSbZQ7HctLiTc/JCbWWWJ2TfmgcByMGTk/LPwuAax2JJVdIninjTwXB9AMQ7z
3z/Mq9mpVwbG9YfokYXYCj4CIZn+i8eXLgbFwtJBKE3LkGpdD7hAjcIszDNqUXBp
y55qCnV04UPLUHxOFtAD1pdYQskVajzkfBgZaHnzhuFUW51k4MmvR9ew975dFPKv
4VZJ6lju/kIQYIhmA9JbaTHCqMDfJkfJkyDmLbZ+4vILorhPhCFf+hr9Mqb4Zkzd
2fEyaEUi5Q6gw2CWXvJW/niBtQr+fYf3dalrbgTuin7a26arRVIJydAjzINIBHNi
SHtmuqOlpExkamAEc5ebKZr+djpGEFsXKeBnCJ3H0uB1tqzWMRJYuV9zqWN/Q30L
ci+hTMF6L6QKPgnxMUXlzr589Ly5m/iUAD8uDm7FEMtWmoQoElkccMxMcE0CKbgv
zJY3xqLs2iJaQ2lbbxUU2bYVV+jvAQ2QHaT2X5N6eoHpJ27Fw57xm6yaYrQcHYz5
8qErJND+Us58pQLdOWK1NgEYY5vZ1pP5etVRdwpNzPnTgGIqzrT61xjmjQS86L8D
6iMSGN4AxpJTiid/xQbH2ILo6PJms20trrn3HVXY3ODMycSCMLngVl/vVahQ5m+C
WWsZ8J8g01MIl9g6hDesh/UVeIcRtQPCUsvn6feTPywLnRDYKcrXxElqE3xLIVBU
t+iGX5N42EhYniGqgkjWs7VwVKnqpvqUKn7w0wCk6j6kJYUqOSUXVLfaFYb5Tfmp
yxk/erPmNFKtSqc9iA1b63E8fzon6dTfpk9Gu2uyPcmWX5TkaAoWefvSF5/tcGnr
t2kpRCo6zokSqo/CrwhgLHWq3x5hNzE+7DtTcafBVapK6X9g+RV/TRaP9nmDCZUS
UoazxpFmGougDT/4CpL7ltXy5l6vu+vA2xOO2jiYW5KHcAxK9YT7CSdv7VRXKhj3
6QbyWUFX9B2k6rTmtSQc8bLu2WfWF5LxVaKvUXOtdM155x6SPRPU++aRVxwc2dHn
Yfa1Fv25FmQ1VBjQziwKYP7AvA0XRVY8K3p376qOnCMWwxVNbTz67kKHINciZyfQ
w2ggYqIxvFae5cSsO/l9o1HkI6djArITsexGgwk7ObGQQGry3brbx/3C+HLJr+Wa
/+OPj4SJOJQEfBucum04B86kpKa/Q1jno1UiQY0Pji+8LUr6WCl7l8bLGXf2P/Ox
yQIU7IMCI8jmLrYG3HkM8EZYnQesTLrtxM29XNFI1faFbX6CD9Y3LFqvA4F8TVN6
HFhGbberjS4ECw+kV0cbQ6MNOWctDTjMoZnaICy3Eqxg+uyagv/Pzwi7IAU1BBce
WZafhpq0hs3DUSqzgrV7HDASYn0TD/agiONdQtaIT4waMalZdYvXv8dpck8WR/zf
esRyLtRmT2cpmV5mMLtDo8DNzmk2mV2qkaJ8FNYUDfA8mm05/fdF9UAwGrnCnDYU
21gcwKu4I0UeGsHY0sLEmnNi53izQUoz8fP8qmJbbJEmZYS1NCcCFLnuTgu5y/UP
mXCQGvp4uDz6BgZGMrTgjPctomxWFMqNjrYv+6LfT2sSwsQGPBj3nRysU4KWpbvr
LzzHt+WoIsTU8ItrZL6dtY7oBClmoRfPilW5oZ1G9nF6HzpcQ/Gb7mIcwbE9As4V
ldw81SW467yzzfyypXYk0TzVoEE1ROz9IFFh03YteQHO+BCINAanCD9bg78TUFXk
oKAwP38TFMbRNxDwyD6sZ4M/dJj9cYvdGTLiTiCbYp/YNjxsXcisRYEPI61cjbkU
m/uijrIIhELh7UcqyhHbWQzUfgvOhbWrLMFmqOQuQrIecgf21EyCk+GWWWVGkRdF
T5qxect67os7jf0b3PPgi7RHJodL5/fuCy5r27q0WQuO1vSyhGMTkOLJjKL/1tOU
2F1+VNFYs6qTRUkvUpa7xnXGXDXmYepk7jy1mMv9WF5TTCsme+bIR6MsitVSzsSQ
upVJqjgw42o0YlSZvlB4DI/67R7sOh5dLPGStmqJODyaY5Y6WykL0gFxtyA42qVi
yOgOA8OpKG/IYr5Bz3c4j+GlSfwpBEGTvoshnc58ZTMkBlSRb5nywZLiE2Y1G06w
eCBS4GdZnoozUdja0JudPBzst/NfjKkCB9BXj6bz9t1Wzh1dlHp7yiYPi4NhiXNy
XInLpp+3BuwPnWtZblLa4hsJAdOhN5Vq+Di1cU9XYNpiD19+kysAod02Yr88NHOg
e502FQynlaTd0eNe7ARZDvVeaXHZVEtoi6S8v9xcyriXhfV1dTzLjAVRW9ls05x4
3IS4CpnIZ17oGR7OFp/gcGrvFvZ733DV+N+4cwDTFujR26VkLGS1wVptFahBN1dd
QQ67HdWEZhdyUuDXIRlApBkEI3rs8HOH35Fs1qEO3PY+axHQ8mSC/8aknB5eouaj
5wF+AldfblcL4THdCEXNFQH0k/zzAypVaxACy/K9n6SvLeH147usVh0tsWyy2ktc
wDwvyOLzgyrJ7j0wS36YHQtsnos/cFj1BvtmG5ME1QLVj6ONl72Rd9G1Kv8BpE+N
MR77e9fDwnMKtViB1/28R0KWkwMqChsWjgZ0+INlsznkD/2fuUDJtfq7CmOnbwyr
mF4BRbT+YevW6tlc+kwV/248jb/xOdb3bj3GyHYLl30p4gbAOL71VYV34LeBnvc3
x3ZvK4viu+mXojXbjXhJfrMbC6Fetv2ysTWaVPwMBhmWmIzAMF1KymWoXRWiz777
eQdNLFzuoRD+o3wbX79DIFoTxc8jmeNt2Gr9V9OMpfbByZolyUkQf9U6oVddAHUT
CtpGiIgbo7qIEFNqvEzmaPGq3g7KZt16GqIl1BuTRPegDClj+3kke0FRx0uPI1fv
tiMhd3AcFpzAnmwT/wqNBfnctXCBjCIFQRvzdYMF71ocMYqho0nNeUvpTMdMWPj4

--pragma protect end_data_block
--pragma protect digest_block
WuYvVJyI4qpr2DlKpLeP0IcFoxA=
--pragma protect end_digest_block
--pragma protect end_protected
