��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki1h=nb[p��dM8�H���]�ҳ�A�z0��.�"p�q��yp��#/�K��� �ܽ��F'4)�V�,�Ҍ hM����;��hs��j��+w�*�V�j�';w����`&���`J��M���v8���0��_�Eawq��,�,j`�P1��[}	�z��>S�u�J~���u|?_�,�C�O�	a^�u2}��/b&�x�fSwɏE$//��]��&7tiNƘv�4m;/�PoNwx J�=�\*$d������C�Ȉ�>�#� )v1�s�v�=p��?��)��	�п�����^p;7Lć�kh��t0�A�|�g�z��HJ���(Қ9�V��L��5��Դ�L����B��S��X� �b-k��йS�,�r�!�N�^�(���I՜��6�r7G5�H$t	�ЖC��W���0��a �)��L�$ºƄ�Qe�k���ke�S@Z�p��w�?��ĥ�4��&D����?y�>y�4��WE�A��E{T�!��&���v^��@Y��Q����=����y�ՙM����rS��|��1Z�RL�\�C+���j]*]fN~�����*3����B�S�m�w�H�]��yHZ��1m�4�%'�E�*��^�qj����
z @�-���\.�ı72�>q)�wH�~G��xYtq�� ߶��^�KYCbڱ b�JL0��c��Q��l=��%�)'k�nP�5�(Vc���/�&���O��*�(e����Ė� }��)�/��^P������K��h������z�l*T�ӂ�KIU�PVm�tp��e-W���w��Q��?���TT�Uԃ�=�C�`u�������e駐�������l��d@�YM4�`�'�pi�[��v���ȭ^�^����ngX:��F�v��|��e�a#{���Ze��m���ը[Hq~ H��SY�Gp\E��f�4_�8�G�<џ��Z�]���&��pؚOG0�U��̣��E�rܙ��R�����$<;�:�kE����?#vp�kzIh�5�&��rGNy4hq�b�8൏����E�ct��
��Q��iy\aߞw�J�"<��o�j�������x��������?���&���Ij$?oz�}�
j]~��F�j:�� -U�q ��~L(�~z*~����x��B������1�Zq���>�B+�]�,F�]�c�1u��=�u�|�Z��C)P� 6�H=d�2��)%�Bhm`��3i�ʺs�s4~a���bT��iSgz�[��-��e���_o8�����p���:u���W�n�N�X��+	uܘ�8�"�X"w�O�W�-�p�p�ƪI8�dXm�=C]Jíj�Yf���h1 �q+ƽf.��qb��>>��A���|�O�V(9�4;�%k�Nݿ�~��n��s�X}<�����zH">�ǣѴܶ�l�V�>rk Z�RL��ݮ�c�d ~���;�v��Rj�v��X�f�{/O�Ƃ�_��Z�!(=�\OJV��T;`��!ky�)7d�-��[�G�z�Z16+z�D;����6Y��v��x�^N��i�R�ѿ�*2YPҗ��d��(�q�HxccgkcS��f��suX���v7�j2����w���tWK~f����hL@	&�������T_�M��,{7�5����TdD�����8`��� j��+v;��1�"�CY�x�B�}��kc+��ѡ�<��Eǌ*&�	<��(Pt.$�sȷaYJ��l����"Hb�s�״[,�h�o�Z�s�n,��"��O�ݻ���~CK9���7b��f>uB_�e3_R_�.%W������ί�����Tލ_�?	�n���%|��}u�CG�{3*�E<$�HX\�F���S<kR%	�E�LƏ�*�����4F��Ux/w��#0U�	�G!Ĭ��O��*N0�i�!:��b��y�zs��lSܳo�&(������S�f�Ҷ7Ư)J*%�*�����N��ܻؠ�sW
ն�W5X'��tKw:A��ݴ��$�B'E?dزB@���XG��,ua�g�따��.y�-�^ ���n"~�Yq��+���.�h���L���m__�^��h�PY%<NT9:����J��[�(/����auH���!A���9�Wj��5��ɀܙI%�������0U���f��c#vn�?�v�����\ו��H{��^\;ꤝ1��S�c���-�.�|����W�N�����.��o�.!��/ȑ] }�6��]���^����1�-��`g,�nN�Fԕg�V�P|U��W�(|�z�t�03�� �$d;�py	�9sǫ�@���4c6�6�	��-|t��7�����
a�&H�	ЅJ+�W8�Q���k|��D��Z�e��bp��EH�}����M�$Y^<3��X
����ц�ޖ�J���5'dZ�c��2���/�OP�:d\��M*N]��mZ� vr�D0S\b��]N{nil�}�o���D�F\Wc�\Ǳ��J���3�������Q���$�Ǔe�h@�K� @��ĝ��MEbD?�ם�aXL<�6v�碐T06�9�J9x�Y�f{H(��~��Ga�P�2��E��v�l GS���I�`���qƠ�μ�1~��ޚ���O�z�1�5Є��C!w�o�Lt��m��q�[q�����~����2��W�9�Ū	��Q�p�Y�l[���I6(�i�ͦ��W�˱��3�Y�;����w�j�?��L0	d7i�Y�_/�k�.	`ʑ�.���faU�_�{��ЋiJc!����[�H�ڈg�*L�s��|j�:�����,4��5��.�h� �������'�{ă���=��@��du�W�Q�7�53�	����3梚໖۹&R�^��[�LANu��nI��p?�u<��s��8Ę����� d%T�c��,r!���/7�L8Y��$i_ BA6�O=*����/8��M`��4�F��lF�4��5�^�t�������VF�K����te|K۵�!2��^l�l|o��4�=���r�=���tÇ�t Kyz����O���k���ߪU�+���X�wri@� G�����X.D��^v|"a���"�H��u�2vN4ڿ9`�����bs:{�������ᕱ��C�Ó�4v��N��gD��zʷ0��K����肄�1�`lغ����|�9�2��� <�VO��a���N�䒤ʨ��tz Gp���NsǦ��^�30q�7쒦�^&�h\�c=7oQ&$8��3�-4ǐ:h�B�X�:����H�:a��* l\s��ˀ�<$�4?�˝���ނ/���O�����`�T��Q�}{R�3ڕ�������j潿��T�b=w�z��o��[�(��8�vDKfGu�m$���7[���n�.Nv��hI�5���ga��iU���!G�^�SNt�Mm/�x+��I������Vp3�C��M��B�~��2� [Lk�i��
����x�rr�mJ-�1]�8�$ݿ_�Hq�.�v_f�}��7$���.��9}�ʮ�Q�>�@Z�/o����ɢ��ZxO.��D5�2u�J�$̽� ������;��Չ]�ڊQ��Jnr%���j�PƼϾ�&X0�!y�#�F_o �pci�O��P61����.k>G��Ba)���"t�ii�As��Jt�%0�q�,݃#�o�|N��?r��hQR�Ƭ�eZ����CE8_!l���W)�k�iM����,��I���Ks08Q� �� ZlG��핞;,��%Iaqq�`m.s���heH9G�^,gQ��s��,�g�BW!�(���_�k_�����^�&�v	�&���K�K+Ȓ#�fX0�T�j�t>�������c���{p1�
| -�:����Y'��{�|�^������g,��9kE-/-ϛQm%�ޟm�Wbs�u 2�
u�P���#�eY͆V�:%����c		����T�%��W����C���'4����С�̕Dx�
����w��qNg�Q�C�ڂ�2�ܸ��r������p��(~3~���@# �[e�	]��R�9��/PF�E��A�':�`���,a�����|��:����x���(��Њ�� 3rA�!ç�*�To��mrmѴ�>�x�a�\=Q6���#y��Z��u$B����f"'�J���)JJZ!���}
��[/�uEt�;s��k��<b�d�y�c�aU�q��9hq�H8�Z�mP�&m�Ww�f[
���>Rz�z	�L~��gR�^��yӖS���^���5
8�q��u�e!�aɛd���+���9���$����8@mz�p��Qv)F�p8�zԠI���PT}@�%�B�� ӱ�\�:~�Ӿ�2*�5�q�ˤӇ��zq?������eLw�� =�J��2W�T���Sx2��M�o <=A�<8B�g�>uWf$�S5w�B��P�]�f�ؼ�}�v44`�Utv=ǍB�� Y�3�k�]�m��� ����4R)�{����h��J*i��i^O��y�)6�v�d�1�=J�xܲ��w�� ]�"=��ap�+��a��T�^���2��T�1���ivbŸ"@�eb.��17#�2T��.�)b����[81��1��7 q�N̠ih���P�'u����=MmE��Q��Z#8q��4�)�x�4����o�Q���ZomY�Y��!��T�ӛ���-l�<~8f-$�7�EJ��%ϝ��=ء��m	&h��D~�68%�šg��0-f�.�s���]��%{�/zԚM��z}.j��^VU��D5��f�_T�S�)>	D(���m��T��r�8�f���e�1@���Y����$p\�k�6��A(�YX�[zy��m��`!D_z蠆C��["��	�m4T�p�ۥut2apV�}5��b������	�n�3�Jk'|�)
�&�3�"�!Q_Cn�a����fQ�(k���͆���x���O�;�h��WCaښ0U^� eS�&M��m��0��RR�T���0퍟�mKSp��5&��p�C�,���~�A�|	=Vwe�8ƶ)�%
�����D*����?�Fp��S�7{�F�7C�j��E(�~0I���A����Z)�7�S)XC6M�e�Ӑ��#؄������N/+���>
�f�h�Rz7�/p#��jIM�]G?'���E��Ő�J$�g����ECyst�BxG�CT�}���=��brnb߳�S�7M�s�銟���;�58;|����v�����+���h�cR����(F��5f��_����Q�Y*��b��{aeG���~�\�q���]j�%�گ�y˄Ѽk s}�����E9͵��rLqZ>����|�f��E�]�#���*�u ��襈7�Y��װ>ݽ��U�V�Fį_/�|7�C.��B��<���8�]nm"M��5�~�M��T�	:��L%r7pv�r4�sK��5U�>���3)�5'�����"~"]�f���:�n���eP8�),:����"��s=>C��}�2�[��I*�_�������F�̖��Ej=�^�9��\�����}��=����sK���|�I ~uK x!�ajL��Q��,a<r�8�ʙ�k����-#n��\)g�j�l ��-0],��-m/�:���-k�+�|��œ�5�eG-�|�x�([�uOԳUy[��Á
�����6j�w�	���L�1x#a�L%x�PY���5�L�)}�� HP�wȡlcgQ�� 2���zW3*A���������hr-��JP"�Y�Z7E������_#H�C��3��ƝZ��k�3�Yx�&���׺��`"YfE�Vq����".����N���?x�N	��I�P�����
"9h{R��k�����h��!b�l�0'S��ܰ@���[�'n�q�ȏT�Rq�&���l���w�W�L������� Kh�!�y���u��]��z���ט7��Tj���JyV�[�oG�m�n�+��sN?�x8�>��$: ���?gB3���m+���W��2���3��}Č��V����KL���_�#��,@��7//g�گ��(d�yB�F�<Yi-,Y�c�e_"�_�!��3�j��ׯM�`���=�tu#�v�2��S�ׅ�&��4�<����je;H6CR*�^u���D����hޢro6���q�Hũ�*�݄aoڮ��@��m���[��
J�w���"�e�Q���*
�2K��5�4`����2w�m�ft�V��11�~����L;f������<���#�q��zr�7t� ��!��_WN�&Ķ��Ji������ `v@��7f�Mj���s���3�ا�AqF���	���q���4
�rON�A[��QflW��K�k��BSe�SI���crL<��qNd:y�k����s�����s4T׃�#��!�Y�H�_)��mЉP;�g=��JU/�5?���4xP�g�v�~x2^o��`ۛ;.w,��Q ��t�}l�c4� y���APuVOXAt&ꐙ		�8��m�z�����?$���Pص��-����� 7:�9�^|�w��R�;��t<θa��J��h�Ni�[�?�-����� �W٩-D7�E�����|�8"o������c噔�C������u�i8�d�biA(�o3���+K�s���2K;p�)�o��; ���ܾG�5����?�����Vڝ�.V'�@%�rʕ��uH9N~���VI \�d�(��ʧ��
�\3��B ���6��5=�L����.�ҭ�.��L�q��b(@ʽ���4x�ά�uP:>7^g�i��%����#���V�x�!���?�(-�>�B������
])p�.��i�	ڌ���E��YD����L}ǈ��N"R~1�RW�t�ݽ�[���ˠ�}DX͟��K�%
��tz�ԕ��3�	L����h�.�X�g�#.n��A_6�f��k��*����3�B5$����OӍ8~u��VQ��p���-�8s�� ��7��(�oi{^ᛩ�n&���E�}�������c��h�*����n)~��!M*X���$v��~s2u��=T�ұGQ���i|!&Rho�u�i���W�9[�N|��� ���A��:�[{��}Q���Ϧ�����\6#���䷘bt ���tm����˦���X18JY$}B���+1���2��v�S��j����-���cp�j\|O�hBF$�%J0�ur}�'9%�y��O.^�f5{����G��%��m�Y����bx��;2S�1a6���pQ��=���/J���/"�M�}�ݖͮ/��
���t(й��S�Bߢ��*k^k?"��+|��aclk7�R�f�*�j-�;Ĵ�/��\�vY�w���_r:P"�t��Df��գ3�6�(&.�%'���+6���+S�Hj3�
�$&���y�|���a�;��y����?�h��|���ۓ6���_�`���|3���9E�#G�A�b��o
�h�2�lK��R��/�-tV�-���y�So<Br/@6��FV|QSr@�&���h��v$���]����u!�V��4�J�gd41����[�p����R<DO�@[���N��LD�'F'Dm�S��3�@ ��8�W��-�<W,T�3�B�������8~�Bђ���Y�k
/#�2}���W��dE�����V6+ڊn-�g�LCҲ��ʞZ�B]��L�R ��I�˾|G�Sg��'dz��<hIM)� D<�3ɹ��#mR!4]��`u(N� s�����a>�UEh9>A@;��mBkf��L_�P��&7n��AT��9@�ƛ^��Gv��<�X�+%q�V��j�_���5Vd��M����a���QO���k�H<P�%����_��a�
�"�w�}��(SV�l���%V4;a�_��cƿ��BCz����N@D���H�Vॖ:?�g��B��;A��N��\ֱ��.`j�E���I��_��d��)�_oR���U2f�|G�uR�ģ�D���o��A���h�b���)Bl,� \�!׀���.`8�.��@(c*s3#�W�?.�<U[�up�%ԍ&U��qsH躃�ɳs�{j�4��萫��z�$}+VAX;Vi�)et%��-?�4��Qfh����tű�v���Sv�gqLżI�N���ؖJk�~;rp��m*�,��BvF��ĝ,���fݫ���w�?IM�DO����?�������1��9�5�G1�����/D+W�|k�0�;1��~��*��N�6��I,ҧ�6���09���.�a�#"��ј��WF��Y�Vf��b��M�heN�s{P& �0kd?y\���4�	D��qQ�U�G��������R��H�qs �G���!�e��Ek���r ]�;4H{�Ybo�˙Lp��r��~��D�F�=2�L<���.���������
���Z�%���:d��t74�k+n/��z��G���A'_���¡� bt
�K3#�.���(*{��[��a��2c��X��3	��HjӶ{
ٶ�mD�||�0�.p��.w������>\�U �2_
�u���^�t�L�޺���~��&>r�+߸Z��_���l|��+Ɠ�t��b�����fl�MLm�Ja̡|��=�ԙ�1
���i���Y%`/�9uZړ��貭��v*��+�ĞX?5��:�}82$�`����o�F�&r����f� #J��g��x��OB
�ّ�\�s��6	� %��ѝ@K�xgE�7�E[�0;ɋw�_#<���S{0��/��XDa���q�	�ǋ\�圮��:J��9�qR�/�N��y�R�O���.ԅ�q8{��ADȡ��	��L;R<$�m�?I�;c��r}[�Ҹrr���bo�(�G����<C��pg�Rjn�������Q]W7�JmL��BT���O��	>gí��٘�4b�ȡ�uZ�f��
���W�o��W(�P���-׏�6���2��ui�%v�O@�Ce�vb��`,| SD#P�����������o i��{���7�`
����9M�iv*������4��J����	�9�/�s�׌\�����\5�3�Go�W���Zʰ�{��>�!I%ؽe�C"���M �*��f�}��T��3�d%��n������56;�QوAI�,+6�Ԩ���Ѐ�=��'�
�a9��:��]�#������w��;`�Z�k�$�O$���|��KVυ�S[�-�� 2���u���T��U[S�l����9����g�흩/э��0���<F��Q��]vȐ����v�{8K�h�I7�/4�D��%nָ��>�r�-��;�(c�ޞ�H�3y5(n�4u�D-)�����ϪC��s:�Ǭ��%�!^E�щО�R��AW� K�#�sH���Ȓj\���g��_��O��=�5dᐗ�a~,�E��6�ȸw IoP����;��9��7bw��M�^������B��B'�>�e�ǐ��<��D���K�3 ~N�_T2��B!,[y�؉�U�/�˛�@��6���N����.[%�E����2^�'�(1%(����6�9�S�������P�@��� J�:�	Y�]�	���~�Y���7t���U���K�}��Ň�]��;�^�r@��ʰʨU��i�ꕱd'!͍A��mz���q�xT�A�tS#��d��M�V�X��l��K�|X?,�9�H 	'��GJm��EtE���!���|VX��.�1O�l�j�����z�7�����K�|�i'"QUd�VP��*�/�k�ꩂ�U롛7܍�'ֻJ�*mWc�X�;z1@�@���^��q��#�ZG��i��i�/��*9T�0нF�C5�UnS�z���|P���\r�u`�*A����nK��R�~��`�qin�3� �PT�w��A�!_��jz=QH�VJ�������Oos%%#��$I�<r�+��!W�yfjnXJ<P�u��/}��r����xA6՚�4��<�_!.�1�m%�M?o�]:����(MTj���Ě�g��S��Y�O�eF��}d��Q�Wկ^l���fͽ	���L��_��T:4��y5�,����'��<�"?}?�����nYu��Z�Pwo?�j��4�&ڋ��sB+ީ&�/j��R�瀱�@�Y$��3�G!KJG�b��H�����6$��#���%�y�����'Ju_k�i��F�d�@�"(*�q������t�h�'ϡ]�,L0k���.���hTi�&\WH$�V�Os9m�6�aW����N���