-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
OYwKOZwZp3U3MPYRvJPdvoySfXfgXGyDWFFXkT9Nsv8G1O9u6kPVl/nfVix5sGWe
lN1yoaAGV9l9zVH1bD+yvxDHiWWmqfR55pd/KfxWQ/nHg/z+eXa9CwJ0+S7wQ6zN
JzItXlfPIgUeOje3cLD3nZyyh2bLzAZDFuUMHnA9t8o=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 23374)

`protect DATA_BLOCK
7zTAf6yAgPgsnh6QlXrtOmbxzbjWgxEFWzqZa7eM3tdaBe2zYB96gsrOSV/jVXXR
+APYQC73HSeLjlT5jP/aLywwmjnGIj/VIW0TU4GUQZxdCivC2jCPzUMBRTKmDGXS
Bu6AftL0R1jRK9fyemodYHNJ06lcwuU83t91axAdKkRSWOBwG3iVqqi9So6dHaEV
s5yddD8mjbREoc+sj2v44671z3ncsc/wBtTG36jJOPltDic5S3fztFlHD+DS7jak
kTv4ogY7spNBzJ2BHqntL07llVKC5GgWAqv9cq6oz9wYu5DzmhdyObhXjgLzC6B7
w2mSthDTN0cznsM1CC3dv7ETUJGX+yetZ0BHKN5sKmyQ9mjk2oODW6GqFC6jV2Fk
xcX6c+nanNT6DV7K0cBI718bnChf/iPyrKyuqrnHobvLKWnY9ZJXp2STQnOTamvY
nMuOJJrJHIuejiinrYPGE216tQxCx143G5UVIXOBFmt2r6k5qIXP5/TvQXTrhVTU
WgfdgRPg8NhcYZSDAcdZC8jkgMrqbJSkrTHTo1ONaR5J6jBJBKJtc3YlG1uGPbE8
vY/BbjTFyQy4ryi4XIyxpk85j0CDMEJrBTDryIETQYuW5QUjSfz48igEcbeuBcfP
+KwFt+6kyPUwSC4uaMJTmXXz7aC8KOFOWO23GXiCY4z3ndGw/byYse3cre9yag74
HHfxhp+s9+dJsOLvRnHKLmkiwz1UEHW6Dh1OWEnPgD+TyosLpoBRJrfHXKqYKiW7
oEsf9/WVM3sm/zmUbxvszkXqO3EXzXxQ8YD29VErQUZ+BUKu8ukN5eF3TtEM1inQ
P/X6OKFZZumA+vwHpLAK8/6ISwhShpRu2bZ2wJc7eAM87CQr6YG6csip6w5nfQun
EGpcNkx0ktzW9Z7yNNaSdgT8tNUVTlF+8WJJBcZTocY845OYpWxliyEYHdjmsGPD
gPTdVUy4qc8IUI/axdZRSxqCkMnldimHVhCMw6NK3S8WXTV9PqHnk4wpht2jQu9l
E2KGGScn06T20neCBErMiYFxlkeeJ16X9BHPQ1oLczXFnzcNkux8pMN4jNgQhY3O
qvs86L/ALTcS1lls0vdd8ytzpmq5upJ8muHAPF7JJZXVpKfyFkWWmF4eJV+NyPsD
11t4h0SxhIGkBg/yRCM99wW9mc/Bo/H3mHb/TxRhQg2aQCOurINLsRojCbZWPM5V
A/M8mOYmUC0MctP3/XNrsGzx5FjP0vSleENTepsqFbqwvviXefvhst5LR3P1atIx
DVBNVJH3ajsAYMcgukGcfgpDa72PpNBin0gAB4/gihb6OYjw1UrMfqS1VbEUFG+f
ugRZmsFga8CvW9D5jKiFBGB+k5AX6SGEC+eZpmDxbvAR8QzQb7Xfqf/NlQTPRfE2
J3/QcO1Xv0MQrz0YMCfxCNmHLrix7R/WF0C1c3Q6Hi7or//ku4Y+tfs/vNz8wBcw
knLHjgRs+bdTRzP1J0VG6jzBaPfcQxdwiekOdUkTnVYmHiHtfHC5qZURhK1R6pVv
cHdDg8VoWoa3HNxqyjgt3M9Ve1ylELUIChljfY5xfnpTL9esZFTtPT5cW3GNJFNM
BeUPR4kvZ/TcqucuHf3bkqkEJHpoeIjqHWwApQTzM6MTRYuYbMRZO1B6T1PfRACB
4XbfHRiyvN+oOcW2M0DbLYf2dAMfNEnU4xllBWpBb5U6ektIXfCtwgZMVPvVug1L
o5DghZisiGZxZAsg2xCDdZ3Gb2JxX66r70KTOLQqltaV4m531ZksGeqVRt/9l7Al
Tg87q+hCZnDJ6LbYlXSMGpc2+ap6mrsj0S8O8hi3QyY/MHIKdRajbJ4q7KV/5NlO
uJpjFv/a3JOhkSh/Dz6Jq2c9PiUpB1jpQMTTtIEFAPqbiTYkbSt/dWYgWF/A7jUb
yCE9DYLuA4PxnGOtIlNDQ3kgEtozSlZsU5m4NFjrwdTvNG5NtZ/Kf4Ntyugf77CJ
AfxBYuk0ORcuWJINNupeYN2UbdZBhQPhy3bLSgKCVNwIGpIQfddj+MeDtUSHVijC
MBdxavT90Zmw2iFjnYn8eNZCVw36PaeyojkgpLpo1S20s92BNYOmkyVIsqfN3OKm
s99sL9dFJQrSGZXsj5yC+be7zXho+BqIQKKIEv3SVMebF6V9zFZcUXQ7x6clYZsn
mBlm+FgCwg1Sfh5AYX/XiU6jGO7HHkYa3Lb9InIKRi0lYWeX2T9jT71wVFRhRN2z
dgnBUBAXHeY2tCXvN7gXB11+oa+IZcBFxIJYFbgdCzwcf5DzPe4X6v2zbHKGu0zc
V2Yp2u0O9dr8V4GLSGgj7N7n11cKm5KvvRUmg7L5r6JIoWRvFK2GSXZHUhWo8U71
o8fQdBIeubc/w6HpbxwIUNtL1a4hd+CLdOtvY6RVM+XD8gxVggk5EjFujqAeQcas
sPSLuhxarMbfrqOwZhBzywTyaeN2s0ny8gjW6YpP11+FWB7zslyhZe1TuJWINVf2
LbT0KYDQHNqECQPhXHUjamR4gg/kHIVcZDWmMCnq2R+aDYfcGuTWbnyO52iLLeGF
nsMZ+Ir+6W0VH0ut7nNPZ43RU9Syj/YVDMIXwfMG5cIO47xuU6573ur2fetW6ETS
TBjf+riC6NPhGPn37iYLt5749QpTzTgGHtbdYmZgR/59K2zr3XgKTxs6jaPeOK1U
ME+fOCD7/1xE25Pz5GRd/MfeyJPWK2gH4uJF0AAyj7v1ZUEpywqYk2BgY86oTaK2
d5JbxZz/dSbqGD/TCTM4nNALh5Rj7+qMG+KCOgp1G9KcZmVMC7gWSgS8RGbkrZjk
znnwLGYu6wZN9TyKeZ7Vgk58u+Gt5eSmJbEnk7AWu24SJMvMWIbPw9Nc/nfHAHM8
YnYwWOy2RTQV1HC5WR+zcQLzRWseiltraUZ22TtYMetyNZYA2X+eQE07/jCEx0ag
QHvcF6zF7/sMJz5C1PI97u+1V3BhORZbyGuL6wSB3FM66jNRG9wTl1CsxCQ0gPBU
URP9spLvVFmI/DhItUAVzZNRF4qDMHNxgQZU6bz7zVdz2JlHEwdjMysfuddrf5zw
wUxCiTZH2eFt4eFKbhFEVrfo5xSRfglP01PwtaGwOigefAnwQMkiwLpvIqWJPESt
6jAHRcwvCrohkjIXxewWacdA/QrRqT8lECbR5qHWxG1YlsHZI6Qyo7c0iby9HSE4
AouDYMzeofyTgMgLAU3seuNNMChxdxGkcEqr/wVqHlM9W7cmUT0jNN5HE9BtOJLd
OW4glvJAwMNr/SDJou+BlhToC5fCjnmnBZ63OSx9YKG+C9NH7/ubpzFp8kciiXox
ruwjBwTf0cHxSHaoRsWV6yBmPmGjoj2fWvWlE9B/r5sLk+bYrVbLWKxKtPL2hW7x
EtJ2QQaGK5VZGKJDplH9cGA5Z/Dg5tUdcz++Uei5cTzZlaFslO9PERYDwQvyhk4G
epqmIRo39UO+8VzW2sv+ATMc7WKvhUk6cHnteWk3rTfTZuZ4TICc+PlRO6PAe02y
HN1GlVsrTefmu7bOY868aDGjR8wvIsSKDppZCflY+hojMU4kdrsfiOVMLoqiuxDu
drETYkJvJ2XYDLvS+d20b24RglGgtVtIom7U/e8RloHAME+fy4lHiW4+P4WmrlyL
al2/10rIy0nSvIe9iRjjJD+CuC9TnsliEW8jaOyxw0a28furJoXjJg5XiGGdKdzU
VnPGXnBbyaHd4TzYkrowNshUnF6zWdgVhGaflQNWzP5xeTULb1VX//TPr+bYT4Mu
3ZMuW8ngQVvGG/ptjCQrWv+uJRVLQIQk/vWKjYDny6FdrRFz+gsQtcB+BAK9d6QF
xwjPKQ70LhYhGBWexQclawZ53ugsGsFRSdPJnXZGN6hB9RL31kmfzYlbkgXNmdF4
aROntjckJtu6w9/V60igsS1JakTeS+tiSKO1XdUYW2rk/+2FKm2rY2fFeUU0Y3hh
r2TPI6Wctdrf3YY1VOt15GuvljwX5KtdliSjdm3yizJeGRUO6/dCXKFLINVZmjlh
n87i8n6rtcMvZTvbVssAD3+ioAKkdee34ds3ftx/iL6LL0s8jYVrxf+Of28n0o/i
dBe8Is3rAJj2GoZef4F/2dpCDcYgxRxQy7uI5vYzSZ5g959kXZY/AjWkPpptvvmm
WWj6rMAyfqBZlc35Qr16qzBgNdgSYBfvIoLsYF9PpRe+6oHz2bUgnNkjd0uHr7NJ
2Aj0GY6v5KClL90ymIBUJH8PBtEQfKFysKtwdDRrLB9vnT4EJm8sLKo5yXI6K7GQ
Oc5te8dY60nLCA6yAN72J+VRI4GB4I7bV36oRzlmwVqb7ATjs6AN0bViBBejket1
wEBAPOzT6FMr/jwPMLPr/Xc/pXtP1hWwFmcW9kyF4jE9RkBf8TdRYSuTn2nDCoO4
34kDEGw2+BhDfl40uajAX47S2bKOMMyjJ+JxrBm7zRgXFg1koR6WBNxjNsxszTNU
5pJWHj4bv/l9agZ11adV+Z+TbL2QZJnWhmb78Dt2f5K78aB6ktOK6C0SzkF1A6zN
5OO8BVXEtTj3KBH1eDPFp3M8klqtyvH5C5S/8b3gSAn9/0xxx8D6gmGYxAzWGG/7
4uQRI9lfT8Sst2QGO4P88M2r5ynSbY99Irt71VZ7ESM8U12qAmG2z0R2jqszs2r3
doYhqNaDf+wHEbJ3OBLRQFkzICXxmn8VXfkrHNpZcnIC943TcFQIkmByvTJaGOwT
MAX1M8JgM5/Lfz/QqmLfwGDcpVoVMjMIf5XXy1VMN5Kge1CopEdxDOyTCV0X0SGC
fFcSWuC8ZSFeKk7n7+gIz4oMzBO6kXjwu/qRjWEzVnoOh1F/5zG7B5zwDHD3zh9w
CLNqnTHbKeB/a6ds3HKbTnb/SfA9VH+4wsDI43QzAOihCiDxK5d0aZXxvc85Hrz9
xReKJTgKm26kPZtHPuzY5yQTClyq0kEXLj2fR3PTEr0QLWCHVdImAmassK3ITT2p
TLoI7MJn9TsbrkyjP5IAvvEBLNsp4ZvX+9jOzqh2ua78+z1zNI76N5fD1m4DiOTE
0w+6zsGF99bmBdcImF0qzgJDGPzGKsOEMsf0dQoJYM1dWV54sa7J+7pDuLrcd+ky
uMcoSVLQGUX7KZo+00jiOAkG6xom+sUxeKBexI4IrdPTbz/3k62k+Bpct6jQ88lU
FPJ9uoyrcyouj+VD6TxwngH7XAs5PhLzwHke0/PDkRR8AiYppcS812hPwyv9J7iT
tfigzQsfinrU7IzRqxfDHzu/n8xpzxe2EKB8xHCOaYsi5oc22rGz0vIywarK3XUP
3T3OiOlktcXBOzvdSRnyuOaLELMokaUuUaon7GosaYjExG95qXaIgRDeoMzhhMGo
Y7CYwwldLKac3aMimZ7kxztA6CjOiNjFWBpcBrXdeDzEDGpjNJgc1IbayrXrk999
ULmK60X5x3FrLQ26L2YxoefC1K1paXpRJRtj9a0pa/6D71slGiEK6Mul2wu2uP0L
UhdChskYylkF/YJ3bh257g2zv0KUa/bjVE9S2QiLx1/Dme7ZcEYkavPMYeo73Hx3
amNlo3MARO5YOkoLRlRgarUCWmuD0/VRAyQ6rm7RDL+QDxICImf4kPlGgGDplqvE
ROjIAa4CxerNVnVUfryyap/PN4SyDPgwMn2cr5m/qo/Gxaq1C5509FTMa/iaJLAX
5W6JtYsRLT3ZOKIbEOCSh88sTP8nc4/8LrsKuPjrI0oP9tdpcctNX575Jy8rckZ5
aV5L4ueib6zzjGY8leqtVSpy76er4Dg621AjMdEy5pzJXMvqSrccDZNkvnAgT/XT
kzaHjMj0Kexc1YrT+RWPezz8kTcbRuv1qlWFI5FPvGR9WiJVBOvLb9of/QAwAawP
FBz+4+MyzBtcjAnlbibXFRhn87Y3AkPdeQbePCFWGJQwTryuTEj7ehEerTSsHMW4
V/6jbNrS0QQbikhZa1Wj04EgQg42iuYrDpVvF+MWcZQ98DEpwDIDWTcftpbtSZNC
svU1peB7GhGcPSya37nsgqzfDZMPg9g3F/pjdNdDvOZftY5GVwVSMoKeIykPbnkn
Uoe8BxD9Z+LllpVSLbI/IOLfefkRH8SF+2NwWXm4WQajx5rRL4x5hrw/Omt930gR
/qWcWgh386vBUNX77JnTxWYiuM+hhXcc8xhPhqw6dGwgKL0kZvdEG6fT4Xz1Aa3C
+8SXIXkAmPlJ+Cc1a9s9pV23UqwETTMvosoKD3sS30JJcz3d5Uhfyl0O3lkVpYNN
Lkq+H2D311sPjYH8+Lca+elyUkYVJavnommpMtV3kEuU68p6SfsdG0go7+nhAA8q
ckMerlCIAHvQHDsL9YeqBm54vVvTG53LVAAHiC31+yIFvwQ0u6pQFHW9Zk9p1Ty3
5JMGf3sKMhd+M0hq2jcgqAx2SCmJnzE7E1L+vjD0XVTpJJNF3erTnTZLCd1ZCp60
LFa1NWYU3MlOdb1+cv4wicF/OX3JvLi04P0OymZ7i5jHUXnHbTlk2vIAgNvycewS
LvU4ZsWrCYKKF1opAQIt4l0GPh4mnj5BiWm4qlPA2PGVBu33JUUvo7ZjB70oZ9yv
iNXkAvqo66vEJtOwtNL4Hrlvu7fKOLxlHA24MM3X1PxuVd0GD1A3mEYIYFmJEgRm
Hn+lES9uTF46aCBrl/Duge4FZ+NgndBwIpyz9gEw8ZBxuUywFR9qu7lod86pZ7KD
BnyQ++NpwdBEZK0ihIbnFodN/TSH8CnG0qXlZ7sQw9HfuGMNmatuzGZNMMcDeK1Q
1vsCxX1YKm1Gv3yJ7nNMefbZYzci4ufhgmIAF1QAD+SYY91WiKzeiafc8+YNdTIk
K0Oe2XG8PwE1jSLER5nTVLLUXHJtS9BpjnDRafRAuo39QV4NJKSp9Y70nG4Gkk8W
6OlL/ERnve6rD1QGbPRPCHlRsa+Qr+Q8x3AXRLm4Fs6wHrerZTn67W4793qjuFvE
VKYmV4+0LSKZjmrKdQU8wKJTtXvz/qotizmsmFIkLiM+RKSvYs1I3q9ArgeNv4m/
PRbx/FPtNDd3NveA+k+I4Tpc/+sSXEna8YN3dZtkoO2FtxrmuX6rNJFh9xBqPsR+
hrhd0gTCWKb5dfFnLBtMYRzyMoe9gcImB3SweD5C4roJhwylFsY6P7IA+UKqUD3k
1xL89zSP1PI0BLps7Q+xW0fudNeDdP8FJr5RSjRlYJSqKI1fBmytuG6csdvO8Csu
f+Xj2Bp4PuK+JxEgNQhJluo9C9p07ER0lswLPruZCC1c1KPXOaBDsDeZnoPWOQ+M
P0YaQ2W5TzrWT8a1ENP3djBSwhO9BQwJR5QiPc+jZEtjUUPHSFhFN2/OU/E+X8pE
LD2TveTqWhD9pQF6PMprIURic5KpZ65wWLh/+cOKbqBpf4ejUPmts36+5Y26NNV+
91W2FRuDpFBEHLNB52jkYubZZto9ePi1hMb1bnP+e1/SXzh3Rpte6+B71+w5jwhu
yG8YGKVwb1kX/1WdpPN6P+O5qUL+zskjTLqOOso0clgpcI+mybwP2hmSVyGRt27u
NACiXw5Nv/SI/ydAs/T041pmGTaLyjTM0fMm1E5LH5tBJALI710AQwUpTcDKDT7g
AW0PbpfZD4ErjYbQ81HkCfP32DjUXsxrE6grC7RXidRpJGBfrcIsP2BcjGV/sLHs
HOWMx69fuOL7H7WMokqiOBWl8TfBpgjI5fUjj4/NsAaPZ2NRq4+h3/ByNTjafVbL
xLR4szc88SkiDfRppUh8ctvkpOdsGpQagj8DLwX5/kROc+53dO+yo2uj22SMfUG8
cWsm5sy3pdJ6tdejf+rvkeVzPnUOLpIuKhikSZ9j6P3e2lRaq9xvUhSiec2q1rpg
CrCNkhHivAmwLpqK318DOptcOz7s3+qkxvr1M9ZPTA1xFIzxcgE+1q4qFaVaGnV2
aWGeTcZ7L37hM0cDlm5V5D+oMVCb3ByhXEBiVVrjC7QKX8P4srM/fp13xTJVlF8j
HITUZwxIcEGRgNVq7btWpLjRJmzjwvnxv6apiBMGA9OdY9o6Q2jCpXWb9I4VDJ4X
Tjj4R2jiNLTmlPmPDwYtZkgquXDCyiI2W6GtLH02Uf/k32uuJXo4g1Dka9TaU7wz
gTHDYWwXptaVIttNzW18Vj/kanj6SJ9/ojNhAsKjbs4W8Qq5ILJ9fmXN4aK2RRUN
JG7M6RSgyzL6/sa4GEMPkNUqd0JLzyTZX622oBeDvC80VtrIE18lIbJRto5v45VB
EIs4FwomVYoww89a11BF5TY/59yfJzcOn6IHTWp/LxG5iYZ/LzgWq1zANJ1g62pa
4+zB+4DeEgBoS6qcgJDS1hRvXZ9FOAQ9L39GFclhfxrOxuHQvrHTUThevgI0lYsd
ce8rIkzofjNZhu/3COOJU4uVpuyWAZex+eHJk76Lfiflk65oJ/s/UDITjEfEGpAx
YQ2JHKZV7pkTXUxCFidCvAdxTF1+bH2Qm1b51woka983cQESpHQmaCDkE87T2XXK
7yRaE7bPUqV+uORybIVHCXLfrLpypoumFxwXdLv04cl42CjfJ2Dzs+/RcwDehWF3
HcCAuxwC9atxHS67l0TwREOGy9vG8rTOJu8WPRP2aAaZeSOxLuo+OZ0RC/n9IaUO
wkfGv7NtSgarbMzOCfGVtXAsejIJao1UAXLjmsdROqpw2mWWiDds4PPRoOhyb7Xn
GHM+EbFXlXpFSfilsylqNKCHfnPu1MLZh/JJa3r3lzigcnhjPd6M/Yw251wEdp6n
rqcIzu8AC3/4dNayKVnX8dleJBZt7D8HdQmQpSv0cJIzkIOPSKZgQtV2/n03+fUy
eCKK/qAt/PnxVmi1spYlxR6H+EuUZrTXmZdVQTYFLInYZJgkEx/Xcrt1F9SAR7Er
oF5Ex5faQaf9he7e3fQRcr0NypKW0eyml2w1qjInljP27oKTij+hRVCbRhUqkGxE
NByjAR1RIUrZJHJmZD7BOGrVAa6Vx+Qpo4asQDCcRbJ0vL0+Qa3czUFLmmI7G34s
eYpjwiUMBoVnC+3q6I+2RZduUey22WdoKYuRJjUtw6DBXinyE2+I6fhpmEHwrSfF
80VfpBUjsXed5Kc6/524ZlTUjzuZfDnMSSwq3H1N4+TKKAcT6djYOvOL8jY3Zkm/
3f5z8KeD1YDMqxTcy9wrul0t9Cv1pKY97XrgbrRyGZLATMhu4LD4WVWA0R0P8aZI
a80gltGm8myO0lQtIWRTKTexLf1sII7EzFsD+ILT6JBDIM9dJgvDuef6iOCoUwLr
39tUsF2FEzRuIo64M9Bp4raTh9KjrNwnQfYUZrNNwqTfr7Et40v3DShihIF3kb6Z
dz9sxb3lRfn36EQ4tfLqn5MeFXNfN5BXn81dZfdi8f+1aC4s7YXZPl2Xqi2cF64m
q38KIhCTuGm0FLNl+wHw1jlLxNh+XQeznPXCDwH7KUn59wv6V4IB4YOL0eqvb2qF
Cj3+qL+AC3CG7b6koc+vUeVQ/jW3FSYWSOMLAc9qiwwTjaQhMc0edh7Vd8WrFzrA
Veiqiebqd+2wkT786l4bpWiiJLgTm4FcEu9pIiqAhHCxU052Frkcew1yQbkTptQQ
QPhC1rGfzI6vCWCfajsqj4eFCn1sDmEfEH12o+m3yfRIk9G9EMbMc9+Ji0DMcUb4
sBAGuaqTEoNaiiYNwmqy1/sDA1yBPFEyB3MaN8z5bj4ALXlEvMeTK/M3b5kTejrG
tn3EbJHx4ej5q4L3oJZTPck7c2udhYSFj6cMu9vIz4PFIh2Tj27eK165NQyI/CSR
JdBP4tRt9W/Qj/GzPlPE7qG64i4fnAbP+4Vyq4SJcmjozXF3b28GMOXIRaWihxtj
EmXkTjMKAJTYtKHMatCVP1pK57IETbjbzpu3a+tcSJVrhoEcVF4fFQaZMlwtT9OD
FvdyzdOl56D0etvlt5GV7gvDv5QFhrTBiUPLed3n97dtVT2kjMMqt/+rh1oVAK4F
SqxB7dKYWbZs580QPfmtpAEgp4nM/1eIZ6Oj5c5xyfpvdHpUhpSKbtVGR0bBdOj8
hBTWvOXSyb+56SCthog3F/UJooEOATOgepvlev5CkG8zJs2A+TQ4au565YqBVwrn
yGNtG/0Xk3DCGDYmIGH8Pvl9EBTGl0G0ogikUt6a6RRQp0MvoLVsfM8UNhLH/RnE
7HvzIxKlPYZ/lTOUzY4ZdrEhdRNe3ItRH67fsVzw46PEiQSsx7+x5Zyf9G8p0fj/
Stp3yfcEU5daVIcSqjtrwZ+a0FJ0qbzzKgx8cQw+YlhBmHFgHGe/g6gQ2JgnGitp
HAddp8twJCmMMy5tZR8Qn4I7N8mUFrmZwf/EJ+eQp1wdiX3VdtdxvSqrrhrXtcB8
bEYp59d5qGmtsPV7CTey3XlYWzAW0GBUY4c/2zIGd/0jSp+3LF/8wNjlgKI73KDL
PVLVSxoj8sJP75WJAqPEJoJ5pObFS22sr2NvZwWKyHehkmppV3VT4eo5ySzQVLn5
Hri0zpnDUuzZdaOi/ntFoiu2/YIFPntCRQMJXOR2acjnn7IXwOYTKzZcS1AaquXF
Tak/prJK0h/pDck1Jo3zf+x3ZeOmfO0HS3PWwi1LUqoF2vHuLq/TRNycluKAnZIv
yACi9fdPu9UnQxBBgdwpyD8OCiXiYYrN6a3hOwSIgLmQ72tCcODOzHF/ZmHvGGJU
orEni51MPgqTk/sLvusEZqwIzNhkoYLFozRyC0VDV26O1HRsWQaxJ5tH3z77ohni
bMJSehya+wfcH3xcrZA8mIkOVUPMaioaPp6Q8nJcSTseug1DkjIOpRaeQUePH5Sa
5uwShzn63w7wcCqzI9szxZLLQ1svgVU+mftLpBncoxaZkRKVG+leJ4pbwTJOytd0
BRjG8I80yph1WYvN1kyztjkhlhk8WhDK39alFVs4XZ2Aq7Coa4R8dcUIpgR6yHAD
HQiDR0XbhjEVbkH/QJdAI3qeLiMVqjLTjaQJQorLEr5VY7fDL5lLOa7xBs0gKgi6
QbtYC+VL53bIAjs+i00xq/3ADpT0v2SQkTxdB1nKlvRXsVogqUsRfaROrgZzE0Kc
KjHlAW2aRLp8re/HzDydEp626h/iajNnF9bikKbdcWbk/FQzLN6ugUV6xeCFF12p
SnRrr4/L1iOfa4ZFPJcmmWZl21A1i7lYYaBF9PHOQ2Y+K0PMoheR2DeXuslyx1m2
hyC1ZgFTSHiYzuZAc6u3U5XyiGsuBgdpXRawfXQyPDev+fIEoogrz9H9LKfFgAxZ
BYiuKGI8Hz1KdUiwFrTp+xVhDQHmqXIC6SZT97AGQSCyJxeXIv1rveGy3ch1sSfx
dJZtKncFkoXnXn4vYbruvy2t1aUmBWjtEhbqxw/ePVc4jgI6AhFFQF4An46xiRDx
Pi+iVN6ARMPSF0elPoDM+TM//LP7o3/+ATaSd9ZOzPdIIX/WeOt6EgUo3comkFIZ
eZ63vZlPEdeOqza69ghcL91Mdzzeqy6bS39Z1Dm7C+EAjAIDYwpRf9dODU1PGCCm
sKO8S9+QCWaJL+uj7ycksQvViM9O29npfqQvrlEZfy5zK4/+QDDBiFKk0gMAtqWO
QrWrpJgOW0fenaEQv+ybI4BnEKsm2WDM6kaKp3j+S0QbWuXH+owZH//Pb7s3SUZE
JqYbN1gvNPKmVcq2GYsCG/M1rm0OVdE/DWl70JP7sCZIh/ewFp8tn8L0vVcMSz2m
pNaMd/NMjjeZpKSRt1YlEUkjV9Ol8JLYUz/7dinhnfT4kv9vb8PGisinGn1tbZQv
s78XdC5MPT/Zl4q/DN6x/f3AJt4Y5jOhKkOfDn9BVgB9xfyChgtMtue/JvKTXWSj
b6dR18aoFbLKQ0JHnrYsD5b9e+4zb2iZfwo8QuKVYwPOzAWugQJ0WHnPmqYFnBa/
SSTwi+PyqsB0/FyNEXM0gGmmZVtxL2SGzeEV/PyTP04AqfDSJdPCqYGw9y/f7K/6
0bU98bjGb0ggrhmA7yQ733V4wDTCkz3IoBENR8na9nSfo+XRuZ8SahJg5tXyxvKV
BUuPGiupRSrMZrdRSjMq7gM7cGiylyRC1FDxQ/oWNuIfwPUbgCeZMQJFynj/k67O
R/396K+N04oNOg9hdjBR4f+YVMoFnbggmRBy/aGzyr/9m/X38qsvfLbYbczaB7a4
2Qcs74t04xZAaTGHvdAL1VGSk2kz5PWk1N3Sjow31jvjX2ETNxSqoriJz3BHVjmQ
Mt7t/w5elw9fkgOyxA6GkShQeYHnofjr4wGCdX3rgZvtJlcxvO6dk9D/2TLn47l5
ugaqn+34TIgUj9tA0hVksf0MYp+vrhTH0rQofsO15OcZmkIMYxAkfMhF8sS7V5+q
/yyTD3/cyNJ9al32S6JrvnMpqU42SnF1s1CdEY0n+vUK3pKWjUYwCjefS+YwwX+r
gKirfZYtv0ja7JtodhKUuQolY0bOJToZgEhWCqK2aBP1o1a45aZE/wSga9J6Sj6Y
TEvSdSwaEJFHPIYjEtUSCenhP90KRTHimwFG/8s6GxlefWSmQemouHORwJ4e7Ahp
q5ZV0anRI9hE1NvBYiPTimu3jdMYNRcVAyy6LrtJ4PHb5rJY/hiD0PdWHnzAOLWD
Yf+TaKDxkIE3yxdmaLY5Cr6njALGBTxLEeIV+ZxppCCeeosYNt52n0PwL+dq/25b
JdKtOGi1agXUfwEE1k71jI3E+VhsD/owX+TtxqB8qst5GN6XVJmHSvX1f9cAZyHg
cWc8C3Z9ITpBT2S66LMgqnt2g9wOeq+O3GQM89BvrD3mBWRHRhIXDXt3vs8skkOl
TeED+/uqVqOaAc9rb755tG3q0vNLouQL4CTEuJgNgEihj2dXMF8X+JXIsYTqB9bK
cOZItWwiRqHFaqb2E9FAcy1f8KTccgwKDmsqN6UDmRJTZsiI2ia/dPw1QviaG0eN
PgS1s2JXNABRUf7+bzGxk3irlWil76tYji3eQj+9TTR2mZepJKfBXfOSI8zx0yGr
PxkZW7xItCEDDKaAbgXM3c0xzMB9QBdz32yo46fCY+7vIoIBZf598Di7lpbIKU0v
TVjv1EVt8Y9JPqWOCuzQQB1AKsrg5oth/dyfScxmlk3UweyscMgRjH0ilgDTKzXY
0mxrAFnIidK3uNilk/BVFCyJpjyGgJJ3/m5eygNDK3F+Kjul+o+twviQk1cDsgPT
PsupNK9nD5ybnmEMwiyBOPCyXQyekpaZa6vQUoyeMorkwnxPnbIy8PBmgpmCY6k7
Ff0EG0ahAvKy1oVY2SSAYxNuJJCkb1flSxJeDz6XEEN5B431wgfkzGHdJWMvDTBi
ImzxErkAOPl2J9iCq2Ay+NjMtLl1zUxar1B2vQat1aHA7ckjTaYdzyiH3TdxG1o6
5AKDgYVICK0P28dYFQmwxfHP2SGlu6KS/Uu24NWoflwTAH/zIUVQSvpp8QLb6bVi
Nj9putn5oH0C5valtkxy6KiGuyI5uhu6gA1hx5V3XP1UBEAx9YUr8VE1kq6Mw8lj
1mikp9PxfN4SI4XivX7bww9m8T1GeucSepz8vvegGFcgJcQLOb5SNaxt/c8wHgdE
08Nq3sLFp4Y4c5OrFTj+T0z6tnyvaTTdywfLfLePGbytnwUs1hxwj/0TL15pWeMI
82LorcIRT6u3zp8yhoDsdz/JcTa2AsIzjpFr2lW45QXpxhES/c4HKI2M/8+G/8ZO
gZ51frJ1UbqeKzVVf/0yBjfVN5iPCuay1LkY5DXUrQaqYZM+xCHTc1D1E2aIckKr
yYtG/VIbFC1iGm5jnra3/QjOAJQlQYeX2SiXeDAIPhX8WswX9TvPdwW04dcZ6xmq
u6doMhna7vqT1jdWMcOILQ/HKCYwZ8VJ8zPk+iPgHtAnxsJslyF5MRcTnYb/+5Ln
nbsyjRrO7u/8Na826U5bwrJDLyPF40DYvAJf+FWWG6CXUJqDV9vvL5nakIshMRfT
jiqcGRRRYdR8qg1rND+zK6kKHKp2hvmxtZE1trw7WoTYnfFnvlWgcW95nD0PsLCR
P/tSFmkllABbeZvDZKCHZFNF8M3GN4qxGOIpqUudvqFRc5iWkH99iTFZoVmp8izD
L341FLEsxScA6vketAbz1m9aOLvHb0m+lpbal4nNL0hKnzgdYp2DhUuwVUqOsAcP
xoSNH/pgXasMcnDahz4GxaSm83bTXYfP5Q+4iw8enWeK6lXPDE3bjhGdNfagAcfq
mHjBsYC9JPEYklWcenF6uvcylWJtCgtPvai5CN+QryEeRpLx+3JGRcd8zlxBO1bO
f6D35F9Ms15v8JRAzSpoPou8rUOcJf6gn4LP4P5NsgHYuC/p5FdfMNgFmGS454sq
VSqrWq7Ch4tdSGJqx8SSlHa+Ga3C4hltti7lGymJF00rDoDkaHzcLiMNDJY/Dh6e
flhGjEQ2xoaP5NOqzxkwJy3pIFdcZgeBbk212wYJhtJRVEl9O+w4cd2YTHneRKN4
NXaCHD1EvDJ69pmm9keXrrvHLAYIAa0lgImGYxdrMpV7eS+Z4gRWB1Le2CRXtx8s
FoUhLsb1oBQSq6Ik2j95EozPqhKSDNyYjGXEcUJXKouYCu7P8UZ0oXV/OHEETKij
aMFFJiHL05N7+tqeAd9iHRfmL3HrO0Mxb2TFM06YYyt+YRsSuX55ETecrqGgrSxX
A1wBrFqsz8/eU3P3FLolgFnedggFrSWHxRUiOxGnCk5QApL4y9sI5aqp7+T3jPLw
AWE4+zQlgATCabVAs3lV+LyFi6+QQWXWCmojL9Gps0CkEQLdzRfFXqm3RcrTENiv
MFW7HwHEziEHeCTBgHdnHVJ/FTBs/premPbtLnDK0PInGYGOTftF16ZJOkuWz//P
xxDPZKB9hVBjzYxu691eFR5oZoHXmRc1uPobmahxoabxjssg81X/0HOaCjjnxbXt
2t+kz+1Uk7w2s4qlbz+YzYASv/lHZRX4SVmN8vx8g7FgDQMA2Ttq5A8wuQodoiPZ
eLbhIIdOBI1ANTtb5UySrzNeLIXYGrjlVwqNn1yBlxdM2LtMk56L/rGtCVey5QcW
vcVHaLw9Pn5HXs+/wY6QINq7W5ig5Abbu4KyLXay9uh+ap/pHH6kp0FK8nvwPmod
JgWbHy68+xv2om4q19jp9NRDFFHxks85rj35tJR4QP5qPlDEV96GJqBQKolJLEhG
TStnxJbkl536+pPMmGLOe+4Ora7uMJ0DCmS5fwHZf7hibqD7JzD+IUSZyOHuZTbf
rHLyzO3jAngabhcKFhEp5K/7jnJiSc1Y6lTpQRukCEik5B3pXPFDaF8tSUPUdfpe
rRVKoGCKjpx6Ay887jjYT7D8TTaDDuq5WLzMOCr6lcTAH2pFuBr/c0ybCxzclnZV
zdHKGeurZIn/IOcmg9RMXuEit/4f1X40mOQXRfEC8V+EW9zZeovr2QwTrLqy2jWC
xcNPRvZTwzTUTZXH4nhJHLC3SyNyacLALJ0aFJ4Pi6PCXgguosqZ3DxR5O6KEWhr
zMiwnzmAkRmdFMjx9JHGqlz/m5ljJuQyqY/bzKrWby8nkXQcxWfKR4in0PiTSd+7
Po3aEd/DSXsdCpH/eCxW/utGsEY+sKQArg+mnZWlFlwKY7QDy3dRLEbdC2KSJeWt
0/+hFa+ZIJLNDW5j2GOxtnYIL0H3gJFP0r8RrgeygMJcW1gSHl7Ui6NtECThoxmH
XuyQjOeBtspeMK4AMv3D1pAzHv/QeGgrOqHeNd+9MtvLbfsEa9GLp+XbBbJoYQ45
Db0cxF7n8omHaIdJSrlQ2krmrVVjCuyWLRCF3KifPW/AmtWqjE6uqyGek+CFoOqv
tToaXsZoucQbU1daoBQUDexAcdNEEs3dtW0pxHyFlytkBv8qBbxJdwFl9un7egtS
zmaYQ3URtVkCfwns0GKspAivLg8bm5hY3AzrfyFSL7Vj0FF8x/7qXGt7uO4PnwHV
4VBimg8DMw4hZEyrSoC5Sbm4OY0LbOqFbX5Gg/iuTpTl3obsM9mHQQ6Wpq1OShZA
8YuRvVQifuzHTTCKAWtDIoMkJ+nruoy+GVuXQcXskT/XYurrxMijvEBZVfJXs7Q0
zzMLmtYZyoQ3mjqrX7TF3FsxwpeIF0+JUKKS+/lU/MwBmmtwTcj6ro7aYQFfdjsI
I9xOo4QSTHQDiQ5Q6Bwt4iZOuhSFbL3oPmVKSC0373tcLGt4wgGHFYfj2ZDJrNQP
JY2ocz1otR78ZVIAOoqXWgH3vjRDzZSHSPkRSS9s2bDQl+CYKh4J0kOYjJKFfRyl
VhbNqoL9C9Cr7CsIWKmyTcEo8n1rNxZ0DnDproRBXqK110aN6cq6hkYDmMV6khWh
AMypXiWiBaL089NebkA4vfM1qYjzzgNAjYLIJFUvtWj6nY7qdSL5ZOoJQgpgBtad
wJ1XImJYf2HVOZucw6X2m+1uxFoqJTkxjMZ9uIVDb/yH78OM+wE85hCZrYEFZ2X/
cJPgzoSz3AcvtV7dlVVUgeRYRq59xk3dwdRW3KWNMW50YZob3PsOv2VIgadDgx9T
cN43T6P1QYRMBWg0koGQcLzwh62eRxWy7OBVRMzk5OuQB/2Ic2CYqZVs7A78BwWD
1vy6/V4eev38+PIQIwxmR529H4tGaIZW8q/A2euyKMRLe62yGuLM190LxYJDLxra
5Kzw3+OELxjMi4Gs7Z8aPAQf7uU6IKHBaEINTNEINavlHDqWqcMKkbk4TCEyEs9x
8dLL/OKBZX9iTV5hmdeSAV9fgZDmBu/FhFRmRcaUTuCWA+3PNMVa66HMZfsu+tn0
pkjzH9qSSFqpD+ir4x7520M2poZxAacRHK7pLgfRnmXPB3zDgkOHJmWohZxgIg3t
h1cgUJNZguLp7vwt1Glahbl5Fu09PLpk49dB5S39YxIqEmcgRotXyIxrPuNlalIX
7qYpda6Go+KlU0998VcXFAiUs2loYDmwEJMEHLyftvMqtdigs8PKcaF+N1DcD+R4
sw94AskIJVTKReu3NXw2+wK36sfYkZqc7skDZC+EAx2TaKzQNsBQqLbGobH9kLL4
JXo/KxPqwlFcA9UfozY1BpO/sxuh0SLftCNfP4vNvRDNx/yk9zHHbvtDhTMILvmw
u5EwUYR3hkfi6dpvJIxq9jYxpgOpvwyeL9ElAkGjOMX0tTCax+vp3h26IgMeaT1h
itim54j6ZgYDttN2meF3Ed4szHi9WbtMT5inCE69+rdfCjToMeEsQqWQe4BqrK65
VQWBlutsMMr/3307lE9AwcpmbpM1RHY+2Ft70fww2exME0Td1X6kyCFMOyyEgV/D
nKDmsZmXsN2uv1ri/fdkHKB6LSTHBQa5OUc2y+dNbP/7omTUKWIAj99eK6T9W175
ObN8ZXNeuQ/X1XWOXUOlyH0Nr7kITZU7cYtYPz0qjx6fD1JiyjBzYmOiY1c2b6+9
wGA/gkjbxKRX/NOSv9NIJH5rRS4sKXnQf9fvhawUh/gzq95fDtLuAGCM1lj4KvMW
s/xpQqlFwZV2xZgCjWba7kniX9mDLT4xHZ6y9LlzYPbONP77eT7z1FHzl9GMwLKy
2VQUaTVYbta83Xvo5pW2TYz7Qd6coolkBw5AAszq/K6SC/ayo0sjxuFJvw2SCLrD
KiwHe+wPO+XtS1oaNGI7H2q4mC5PO3cHxIL/xvK+ChgVHfxiyVarYru4pFHnpzk9
Ca3xK9n1fLyQmnuio4JA8eVucQwdNAPvDOoH8JfzQ9HYqxYxRAMzjbhToMrYZ9ju
qC8ef+UuXUtVYapAEcVPXrhIyCdrfCoEtmysiHzZs+zVxUIiONXnOfo4hpAsRgaM
LR26L4bVnzWboCcQLorG4w2OTOcEj0RF9k2UbBARnkt9QSo8an3c95CyZAQ2M2bh
X0quGEK2Hep89IqLFKHOJXmSr+Zgn0Zzqk9WQe5NcX+ijwqRAnSRHBumkRxGvNF4
y6s89YDZBIbj1FjxRvuPxaciLhNNzrdxHEaCJe6NUD9DePmlYeVIZL05zTBW/u3Z
G6Jb/HoNPlqC3PyVClw08xW6dQwsx/spNl5jI6U2c11mb9lLast1CGpxAUVFlc8o
4ySq2n7k2j8hFiBSZrnRaQ+p8Tr+B0iDjK+Pihmp3VyS8gImaCYksAj+0Z0DG8xG
dVGv55CO1U4iZROoLUGNERmloHgosdFiukV66uvPLG9yeJR2HjRneTVkTMV60/4G
lVArltz15ZYAvjrs7ChtlgK86wJNb97PyJtnFEubXf0ri8Z3N8SFX6nzlajnfFPP
3d6/LJeS7o4oNT3mZp/VRKYKGqC4ObVvvcmCjqFK+rI5MYdHSSZWI5nypx321hrw
7aNqvCHC3OckWEDjQAZ05wQZ5XT7VlkHNYbAMzw/EjLy3lFKv3qdCnpJDIgrFmEG
zLEJYOCNHjNKZPcYLEL4L999XGzEnmZkdWUibV3UBJrY7DDV1asWkX96rDYyd4g2
QatEFwdBLRybt03oVMHoAD/Cvrs+ZuvkXQKJiDSBeS7xiMzujiNIe0CmEOgzi4us
kRBhMVUDJQT9zV5hyr1ybGRAE0lk4uePwVgQOIm409pSY0V0wGDuzA8LuV9vMvOh
va3bWsFo5BCSCSZMg5/pU5gIl+m6dv5z4Dc1a2hSvTwiudVAEtZE1xHxo22Sbix9
B8QzDfte/Z2Q6pwsMp3UzUkxV/GQJ0x4GSmJFljkVWycxsYi7CTzqqPwgW69TiZK
jcIIpNT49O9zgNlaDmoB2qO5LR9KZFG3taIzk2X44XjLsHF4s7vmqdsI/gLVtKms
2T0N8Pu0jpIaWgfZNLO2HDaOpHSzi++P6RXqA10QlYUffVGd9hfltrI5iQIEgh6R
psvxIJBj/mq9AFaDgjzC5i+Yd/yoTly5dcNrCIpC4O89lOKDaPmuz4zBX+5eg32C
f3KWivI5De7xOqNuf8wfJD7iHmS6oMYauGmjt/A19A7hi+ilrrYal9ofLt9q3TwX
EjHAR353O41IxplEZC1yStJeEE7ts7ZZfarLDJ4QRHCfLpMBr+b6QB5ZOCg1Y7Nr
ToRIWnxdi+5RHFsc4SQXBfni1XnHtQZ/lQcU5YRJizKR1Lj3ggq4wwDGWtriEU0J
XFQTM4nmkzA+441/+vaM8RJD+aDGTVqmP+b5AZdWQPjRDusbF4FsDco8ZK+tadOh
uzxOVF0UVOFlmcWeUBDLVa9nWU8ontQ2syw1wZ8Z4GnuuQKlcGHla+GaoMnfCfKC
6Xjc+9lszpI98Z5TcHJjQ16MiptpC2ivZVtl/Y4I9PtErEHGK7W97xO6XpJu0ZLe
u3AZjmI726oKvVXWaNtq2XbC7kmLBM/jH24pm9XKRBDx58oGAU8WzZMjWcH9nTuH
u+xW7RXM/6Dfnn5GvFuu6y4Pcy9DuK5QwfWBIeLk0wIuaTCFC0zYLhdQyPjBTenF
EEi0YWcwTg7i8DKjEGLrrYsBtQ7A4hPI+U1E70RMC0bn5WLpOiQlMvI+bNkTFSFj
PbDwkFzE2E7JxcDU1hf2Iu92iEdWxLyjDgVYCMoWmllGLlraHy4YJUTr2vqg/bzK
boM5ghtBjXpAX1t6PMoz1murP/ReTeFH8z9rh7zfC3cUwAoFFTQZq1Xyd0OL4RNe
Pa64eyLyQVdZEckdK8m0AVP5kPj4BhtwxFtZ2JC4bwcWPltkfpV1K93W27KtBMon
AIu3A5BFUPD7yAQ4oaFO3+pcNHkx/LXLu7GzBuvhMxKqmtsg4u7/rQcPN0YKplRk
o98roRtArKH3iJb62CN98vb09W2o3KijiZoMIv1+nGMpByziavl8cH8YVUbkibtj
Q3R1/uP1amCkiTAn3QDVIoTd1C09ZjlVBx6k2wlRuKRgnvgQ0sjpvpEXdWEdBO84
zr/HLtPBNo7McTo97wTV19tdmnN+fj6v4aRerDRZaTgOZDn++Q0/PtNktrUfes0+
6rwnBQBwRZ7jXFGhhFlkpfoG0XZuKPDvNhbaQCTXe6oS3/5o+DP7DhttwOcPUwjl
vT0pYi6TwDXYHqU/ALlnj1ZvvsOQRIW/bXdMZlToz2ZEzmwQT17ANsFGV+PQbjkj
ztiZIRRLFljQNOVbmxlFn8BKeIuFtl0xDY5i93KIrJ3yK5n8UgdXcudtv5sbdvak
koqIAbKwIpx0AIZq3FtuDfevpEyN1QcXuK7AlgI1kqTQZtfq1Ik3i2f5xdBqIfWl
CYyX8d0cjuW6uYTzM74Xr0PJJawmXKyQC8ExNDBDVsYDrkINULe1DtiwKQY7dA24
y9iEVHW67Nc84fjtQ6/YMHDFzAlVH+ZK/8jse9mYr+ppKdAoi+SHRc/Uv6aTr6vd
Z0Uc4Pvk0dT7yz+/buamEX4ibN9xvrPV14M33W54Wprl4I3Ryg0aHEEi8YJVpOvI
hgCpE7lDS/ejFmFZVz+3wOaLMz/0vgBCHScMoPSWSFNe1dmsGVnl/9IBkRhZfrFo
TmQTVYaCgH5Oqeh6QZdq6XqX6C1zwLilXMyKOIxDFmqvdB1xfO9gwBIOdo19aDHL
u1cTklHNJc/0xvS8ClkYs9co/HvR9lq1eqhO8CG/Np74MbtPKQ4mi52+d/8/XkIy
BRCjfX5cNFxZ2LoOXTj/7j3VhuFDrWM2l1NcG+oXg3lIOpe+umpFolWU6Nd4Y2rb
5JTtWb/2zK+PVwIaTM1GhzwRYCZoHkpG5nhvC2ySPaob3WQmb7LgAYGKA8Y4TEeJ
XzBWzgpIX0rajCrnLMV990oJNPkKOLQRZgParep1IaD63Y+NH7V+lhwlrWIUhZXb
xVnszjFQc3ZEcMwnY1N/elWmte4rCImqvxxexQ1qoFGfiIEFATSMW7+/09PB620O
7DQ+QCT0aB0EYH707fDz3UV0ix9MVZxsjPXUWX8codZi+M3kTZFLpGsaG0h6GUdb
f2lohVRKaaxt1QsxipDWkSrBUOiewjX4E5DZLqTgPYIRAyEcetOBYhE6WECKAtsr
Z43xbEN4FhdSvBYrp+TtbaBXc31cPhToayC8bRCFZMFhXQoMSqZNyC4iZCLdUkSp
dZd8T05R7SYfhK9mHt2MWkucg6H8nxkhhd60chz/TCFTAwbMKOJPBjABgk6p6lSp
T6MdNyXR/65M75aDeIazBWnkEzsZ17VCdG5wuOpBZNAIlt3u0g4AWx0BbyHYSJ0m
2dxPPJEhK+yHjtzFNx/4clHmC8DseeoQAFS+uKLS7WnD1AJbK69XPkMdSeW6ORQF
NvuR3NDGFPPXwXoQxFrBTCpT+ihjGB8U8jtjPR9Rd62vgdi0zmbVahmvr37uJCA0
5tQyg8016M9Kdw1IdZ5pTPuozL63o4qSVApGFINWtrjjI2aJG+HHB97UBOLVGL1T
av1Z/wfc5QhmE/no+BZa5RxjuTHj/NjUMKBOQCViVoElX5GOSGLgfvE/MmruwM0r
hfvLMtvaoL5BM9b4NZRACji1WZOqU2RKMdZ9yhk5gZKGTSNx0iffdvHCnVfJs1Ug
Y3Gnn9BFFjSxHSxkextQfTSjm4+ZP56pPp8f13sTPOpqIAgCtpEMF9dKMSL+dj1S
C7fl2jDzSGtndfzqDcSeeMz/8Eov28bIgQ4Z1fvanJQ5np/jiFmejjKZ1D2wknY/
yltb9E72U2hO99x0HTShT6bnLXdWyIt7f4VOcPrRh56fIXZYNrab5e/+CMIP9gVQ
AGWsD9F4qIt3GPds/RZvQwzwWlEXNENNyBojpp4HD0hsGs9MMK9ivRGkYbHldYDE
ZTJlsXhh0mlZbPSDtkDT6iiXmyS1BK8mhoUmKxd6lT4KBKeREHQ2oz4ZEN7M/Fzu
MoSvD6XuCKVta5zCXEF5xoh9mvMkwEPw6oAOPGvNgt3ezqA1DVIsfi9O4KzLUEiB
RF852F2aqrqVbsbQMW0J9CwqQrvXWeA/sYSfHd+eOK2dNHimGDo47y6Egn2SV4gW
fAbSphTTobVQS4r7t+nO06xRtO1G/b/uliK57M4JoYjCPprHPyZvwqhEYeXohndk
CseR5oodjij/0q+IHUp+VAFyFXsR8OjCIqlf8gshHb+1TjsZhJ7nE2XSqd+51bap
92P7hAVY/FoC/5uv1szyfyI63AQo8E1C7/HwIcmcn5dGfcVGPNE76pxYRcXIz1uZ
UG/kvSYck3jrRtLZS88JeDoyeb1kLTRkRy2F+Vo/GgJR4w9T9LcY9drFmxSEttuS
jnxcbMOsy0Du7wNDwiovMEBhPn3hb6ZaZ7/Ale7H2NCLdtYJjTEBZi8Bxt3HtI8m
g1sOmoiBcxQwzFqMf6d6tgPInSgO9hUESeQGmC9g8BN7DQu+Z9/EHYuH/wGO+bNI
bgN7JNVuWFiUPTmAD0pxINNBgiedAKQo5IsBiSt4nGGr/XEfbzkETzv95jDhtMny
cFLrotvVKZ8nkRpdx27pqb453a7wkx4R5GUvKzHYtE0RBa/Fqn5COt5vX9QWkgEp
fG1lP80m+gSAdmGrLBNcQv0TjPg++gfxN1nbHqiL1RoZpgitLN8RRKImDPru5imn
3JY83A707674sdYpZ67hbpPEBN+XmwP+PRIgqpEee6hKPiLzI8U/L/jQD4t0vffQ
+XoReDbYyn+/+5Kdt6ZEbfEWwttEgp9mbVC4XAg++NCb5XrO+5wPdiQpr/FnrPnQ
ZpbkAkGEerz67Qk7Ucuu95Sp0WeItWb8SDQAh2+RE21fB74gibymIPMRBoX1fcxN
RLv/0lnDj1/1kS/LZr46dOZ8iDaqqy+HIFxFjJANHB1VjBwgqkPj04kbE6pQvHW8
zpO1LeWIXa2yiRvHZ9j/VH3BWdw4/R934iDkCE2yWXLbbfq8pwPe/IQ6fW2EqeAe
6yjlaqfN3o1XoaSPqV3qVMXW2P/+iRlm3XjQEE/20vhJjPvLnD3zcW6+l2l5Gpgz
kPlSulbgKRBC7FGgAGkMrrXxIP4wXx98fZj9meIzVAPzm7VyX3As7FdeR9hFeT5+
IdnrkZaYgXu+/N0V43KUKZrpN7yDAjSrseO7ZszOEct6mhQ9rHW23W4sivK6Nqfj
preSczXJluGzkhGA/8DhBkM9fu+8CjN6yUDaozmGKAmMMAJR2hi6MwnDlTjNzRCD
K3VV5mrXm5dWtx7+1GcGIvC+9VyLCntShMBkj31U2WDKi1K97Rr5DJZIpE24gzP4
5hU4RMnuaDtOCBmcIMwaFoLPeCVOr6ETBhRCdad1odEfvVDfGMc1vu9PQAUyyfan
DsVpdysqilM7qjRoiuHeDt3taaB2q0ylWdnGffiBas+G3PMLRpbJHK9KzDblJgqw
GrXG9mUdvB/ZT8Ay9psu3Bgz1J9OTXul/DoOrP9fubrQsSkLNUIoW5uRks4lg/G+
Lam9VnqkBK5roV1prDFXGXgkfCju8hWHyRzNS79mDC15iuQiOmkXj4nse/w96Bnn
V1i4RxiXRGpERcrGVf2k9VQfgJNuOna9TrrcTNDAPrHj6q8luu9hMgaWfKJHInPE
IXiqhizAiVR1sBTZf1Ps+VlwaCamLbfI/0t4Iwwz3gllGUtO4uAyasuWbJr9Cal9
nqDE2aDlSKq1G8v4jSKcJk9sq6ag+Q5IBPzefxnUp5Fxmcq3UYKGFCrp+t1niuW2
+5VooNdCagaQqcQGqbqUlj633j6IRItEC+HjiQIrZVWhGlHB/M7nqGagDAdk2irK
tW8zAwcmy8R8MGhp/jwBpUQgO1iA17Yg34zLOMvmk7hNHGRgBOX935ayiCVdzNb9
zP3z5t4avGnRrAGLNKFNIwnH1vI6GYFfTEc//XNPV+Fy+ZlZaCUCpkl59Kt2LFKh
+8SZ0lAouZ3w71oH8ce+QL+X53J8mpTzcTMiGbS6yPz2VQbRfONaxFbI8aXGYy0P
IGDQYAZ9ILhUSTjB8jave7IXUQRr01KvV66I15XlEsdr0/1pTZ6n7JiBANge6CAn
RCgI5W6utbZDFSsXwyWf/T+38tEuj4LVXGcIaMAJLcLdD8NJF+ORNLiWdLKpL+Ld
JU/qFyc/c6A8/9wwzgJPNoKrXq18dHbMb78zEuB6LQinPkN9nS1W2V6lxMfc88d2
NzKJaUEefzIGdyoBvd4R172QyEgZXvww4zcFjRqZ6yV+psrwDZorTnjl1oYNEGuf
vJYjWswL1mriKitbNFbksP998fySe1TYueQl3213YXMPSIKtUIR9vWeWmW0OKrEL
ECUQVpL+/HTSbKC+LErS0cSaQaJV/zIKb2b5YC+Of9EIGOoyq6qigsXOFmQcEaXT
p1twy9CWZ0qjnUG+Ow4imMq1wr7AgpWO4Gbe/r7JxlYCoNQRlhQW2hbaEiB6/hCu
05bmRJnaCZsV9jM8feb5A7dA0EajYdgXmaCjWhdwRNJJJ4+KMoeTf4TvV/omL1RG
eiuzvbGoRvssV0OXhyryFlgAmYenq7rz0nvrLuy4hy096fwTZtfqP2EmT24osuah
5HHEO+8wPWmj9TPQu3onvY9YmLC6gkQqlb2dgWn2ETuO6QCDumiqukaHMgSTlvmx
ZzS0+NCC02U1kyzVbKMt/1ps83pQpcQ8gkZiynnM+DPimwETHHwb3zqPvF7ekcre
RUlb8XxM05mq1ZheHQPkvVZcdCqncJdIXoyTUmsyYNUjMBuPlVMUebhTG3O9cB6v
5yQQ+EV1Qh+WKqMvWy9jl1cG7n8VN9TDngysa6d3vb2mxWbBh1Ctp2aOS573An49
vjTSbrua9VaiC6XoL8pfTplwsy0Q4HPmuW/REQ5lMNysZ0RBrnexLz4s/UX+Il64
ErXrDupkmKYiDXnxK2fS4Ppfk3MDehS5tlN7uyHXTdIUSZXk6Byo3k3dvqqH95Ga
sIpe39G+Jk5j6aRuijJZtG9K6pbh/Dvi8Zxqhdw52YVYP+kAMwprW33Lu0ZCfBAq
KMa8X5F8DEQSJ2XLDt+ZOkERJZvmbzy5vNWtoeAXRQ35qJ4meYdQylyvh9d+anI9
oc+LhRecQ6stbAB6/ztFW6Vd10FfiLspXOVKCjCM4R8/WIuh/crFpkQHY4QOSik3
QaOCG5ht7YWqROe7YWcschaJwVZ/O3EPeVFuEpGm2K6xlaXhVoM+Ew0L4kBq++HD
g+uBH8z9VJisvxuiKfanA3YlQvZ/YrHJ3+d9Z2LL/vW2rZT3j/MgLa3vagYpf6ck
fVjq1nRj1TIM8orOm9UamN1YqZRMQemTNulTQ7Ldoj/o1FqQjT9NCi0O/6JlnGwp
B7BH/g+eONq7o6KSncINOo1S+PjmRAam+jES3VPfiHqNGOS5O6GSn423IjX+SVO8
vtbVdWKLyfDRnc0T5T4XPCRfuSTMnL8QQR2p3NeWcJgvpQ7gJjcrYB1ZOgZZYyaY
HX2JrrLu17VzYMfxW2YIFpph9BWtZCouUFu8MAQQbBKjn3+YSmh4fnX7za+bc+L9
w3PKTKyMeusyTGmK82KZ4u/NtYwnjczTlDkNdbjd/ZU41Kiy8eA52N4/rSND1p+8
hljLqY0GQZV2B/Nn/6XhTE2ycHpO9tKl1AQbmtJaV39asB3WrToZ1ujXxzgSLMU3
zygV9L/n2zAf3vkR5GkjQIdBaJBESFLlSjPf0zg27VHKUTQOtt8lO59bnSKsqmjn
R8xjEjJs/YLLVSxGSghH1auHy7KU0NJKucPRYUAqsjULUHd8dvWEBCAMvMXXBXW7
7szBvIWhlW7Rg8eAhoDERCavJqwGmGbTbQ4YiyChpdYeuoWs2HNpoROte9198W52
9XNu7q6SpMsWiqSPqPqDdGt8fHkl2xGE5Ve5N446WIRI8oEcydVgKxctcXNJMCfZ
pQtnxAkfEJ3jW33bJlknGKeyoXQIOldDOQhTzQOsL7cJUcVZNMR4BJFvqqYv8oMy
BhxKn4AmFb49Vx4NIDxLbdFrp/IOqNVwfuRJJ5L0g40cFiV3Wt8JHQOKtRJAm/Cm
wMhpoVs/p/fUy+4s+5iaqCrOgLqhtesEwaD3BVown2njswJUn+KhjEKLueUnhfFZ
oTAn8BPOpud6X39Ro3xmyY1onf9qANvoYn/IBprWs4NiFnEQg0JN+pqww5/oStRX
auOCaGAmQB7EXAQlXielwEWoSZ3y+vHlcqMZBpSEkM0JQDetr5YM6sn76GmwvLpG
RmNcD3+Po+VSSO4vjjSeObzhkYqRXx/1iO+HVGxR7gr9bbwvQyh+Y5+lV5u2SJPG
b4mamqZTZMIy458JM0VizqrksYxl1fsCOtjHRHUG0KSeZHhwlUN0IBsi0kWG0p2W
d8ce4QrtnEd97dl7mkF9Nol59tnyMPmhOaa2ZTLKHpUqxODONPpTMH2uMiQswhV+
izqYX9QSGMXynOdCohuhZ5X81MSb9BF5GBROPUx9Iw087H2Ul3Zz4oJX5fKAitbJ
+AVZbtbjmrZpfdFasn5PgaNyR++Wpr5dKO2uOIV23BQ2I+tWG9+wO5kaLg95ct+9
Jhk4+mEm/5HG3Iolx1IZ8rPiNG7oy7KZTjLxXCqC/dSNKjSs6CYPGu9wupDV5bmJ
ck26lpxc8d3Z2E7X+LExtlXs/V9oHHNJUyWgnZCe0R5OixP9l4FYqextopP5EHpE
E7Wb7UqVegN+h7pTinY1MNy4l8eScnrMcnvxS0BzG3tXQzDKzPFs1aaerQ0I86G7
WGZ0EwAPEvY8QxrWwJhLrFd47s0qMTI+8dI1nq4z5H458QsAnLrWRXq2BK6XNLAP
ADAXS9YYIDDDL1ft2dmpd4mnP4X3DR2iR1NGmeUzFBNytQFoF7EBa1U4L1NEqOPw
KQHqu+dxngVEB4E8ltERi2VZekdX3Szlitg/gn/2FTX7yCEDPsyicMSmjreOpWkw
sMSPwQix+qLatCFlc7uDZoeOi/vkzHSi8KFiBCBJEeO0Fvt7SPqH6w2LJvfGYIlp
2Wm9PHaKW/vHapgDFD5TXQ1mbkphmDoYyvyqnzOlk6Z3uYetypJf3+fvBLdmyKRi
Q3f4KBo2yb8RzDa+mAXtAdkyKduKHNlzkEHTlmOTVDjB1jKJ/hlQf8TUWUkBUy/l
m6hyfQvPP90CiayKGg/7tlgIDq3LeXZCOfSbyrgZc1/Kd08q8Ovf/nbTpfCRDw+H
Rx48UI0qCKT3yD8xfO3woJfpiBUFxQ49rqeA1Hzo2oyvCLcf6wAuo5IrilubvXHq
KaQtUKtaEYG12AAkB6xad3+yumU5VqaaWaGlKWcxvazxrCKfw4q5qfPkfqTdz0Bb
Qc6mfgECaZOjJEI92Bxt1tIfXKZo0WEzYQrWrO1uDfDUBzhQFwuIGhnC93eLKB44
MxeDiaMJQkpDBpEbwq95EysW8rtNJFGQSDo4VDwMNH4fynZlxHBF4YOxEVnmPQTh
QHHsn8s2fxH/dY2sfSxIqK300Xmj1elMjWAjnR/qswLEqC7wZr9e08Fs6r82tDdf
BWHcVdW1FHKVFcMjjdXlwhjV9GLTvBhUmJT2i2q6D+Nz08yR2uqYhosusNUljzIv
1b69nYhsX4RB3Dhp2bzeF9+ezxAiPkbeYiu1o00PF3oH54fWucMM9SfC51O7ayf6
hAmE0d8tqLW1EgTqfL+dskiE4xSkcCpJdZcQvSkxgN7hufSb1Et53rFPlcVTYWIa
Te+uk2fjopKv5HcV2HnndVCRe+04SrI/pVpY69NHumr6DZVQC5Maym0covvlJlkF
P9RGZi0+Q6A88w8gXl1Y2YkygwpaXTFzmle6I3Y9OgWHIe9lbskR6BvTvYX0ly1D
L27Jz3YXVxaK+aeHanh2U5HkB/HQl01eg024oB3USHsrX2YGnIccYA2vB5cZhisc
feear1OJgvcRJ9say5MIismqjfkmp/2am3mSbxl4cdnzK9HaeUAXvbKsIShKf3bk
9g2AO7fyZ72I3fzdyH5ysXsHIPJTntsUyxY9G0GvnzHHb3KuRV04dZyNyzYfvmRI
MsykWR6abHDVyy7K9yQZAwgqUgHzYsiaFz1T06JC22nkv1ptZmeOBDXFwA9yG38p
w0k93HkN/qM1kQdffL1W+mwdV0hD2NdJeaysHSj8JOo6LfJ8uOrgQYCUhravasCX
XqRh/rtaQ0hlYam1zVOZTn5qtU1fFBIX7I9ErgzvvDr+Kh9IdneOODE/UY1eoN+Z
SMAajbi4NWtfnB1cwfc1jdIUZ+HGLALABIR0twbcCNe5vyHqz0tE+ZyErQYfbge3
sI1D+S3cXsw9sNC4QlG+djc9DiXtjdsNNjnZMtqyF7GnVtle6Kk/YR9S0PAvYPUV
7UMOfnzb09gwCBfChZniT27I78FQMIO96S2oIsjR6qRgW+utxUK62ky0cuottBj0
mPz3LDDxKpAvivs+emZnzAC/BzDBTJu/2zrIHU2n7R4D3Wg7Kajhwp7hCs2RtW6f
3g099g9jXxnOjSW0T7PqBuycOOCWuYLVmx9IFjG+LzyekjYnNfLiSB/wXuHhhfVM
3kPTBSVvbVeZDDR/s//Pn/VIuKxl2I0Bn+sBQuHnUhP+RcW1OjFqdWSeqCCy2lzb
pL4bAxFapYCWJG2kDqnIo7bMiAsPd7NZpgtgI2mhGQBk/+1F9jYt/DlP6oqT72o0
HLICsYrT+MLO88T9uxS4yEi2XDum/IQGkXpVGFEXdHxz1GxaQ44rS4FB+7G21fb9
Vth93vDuN7wkhq+SUsQKzFOdhuwLhwgLZ1Vv4G/HWIOySBHNzE9sxicsL+j0zkwV
p5ZV5ZNvD7YTQuPZ6DINy9Vgl+hkodhTZQ0oBX9kl8mKrUYeSy3Df40kxWObKDOf
Brp1pAyQsBQ95O7oANTY4n8e8z3hNkdFc+wN7u1X7bCSAD5DeLLFbU19sq9wkjLX
6RtEyKdXWSlli4I4bbcQUkf5cMcMXltJqRHTNUCskSy0QoY8M5UT/Y1sK+rFgcMZ
U1wStnh7nM6o4BzVRPQLOY0U85h9Ne1WyqqOwOcgsdvLp8khavfi+npq7raDUPt/
m1QuHHm9DE5z/A856CtI40/MRFSTWYgkUw+cbfJGSlDfrq39+R5sBBbXSiCmBtZQ
0/p+CbaUPsgT9cJQbwT96AfF6tf3TrWzhULWIh4RXVMmv8jNVCt2d02P/Q4XDs6P
4pckSWuYS4KLsq0qiwLF4Fm35BXShy2wsT9Z2MZ6aJrYwDMdfuL11AzwhfoCLjRQ
vPYDQgf67cvQweOqnbeJa7e3cQKqZyvoPPKEC9OmAifT9kuM8ubcnP8RpNsDqA2L
39eDueyiyf1eRjCUyJ9nFCUdaEPe7WSPfd8Kzoi5bYGuNEy6ohxRkH0RrO5qbztY
pnMh7Qa7d6logwmAhYkrsi+tdZDKXsLQEnjOKlbuvZ6dDUfDW7Cqd4j2/sydYrrE
aRcPV9bFBoEZba9Dit0ienKPslan5ApbFOMUaB17ZsAo2FJo4Z42fK0dr9GVFBP+
3Rg8i/jds40fCNDcT9bEolmNYngtnKJkcFOpzOdwDJt6ytPVJ9/wGKVbPdt5zqK0
v3N5gMjEghDcrKq3XYpimpqsKLJg5UbSOO6X0lZSb1TgOiySyp/1RxNjfFRIOHb0
zAIUHc9X6s1ReMJnULcmnd8/Q88fj9DWomURIi4pTwJmu3+tFZqETOYtFEMD/BqV
5QdU8FcyCEI0auDhkPv7LiyJaXsvZDJsytbRSJ+hfSvONuY7lTs4bVUNLyilr5rh
V1N4uG9WDSAw5rIWY3mPtfyfsPddm6yQQy19o1bUG5iRoiQahn1VMV2fTkxrB7o4
ozlw9fOTZQ8hdzt4eQ2O54GOcA8Snq4HxvqyTepVM9ozfXkdsqiyorxbVL7d8EqO
fuR1zzSSEPTaiUjwo8krskkcFQaiEf3wHEb0QubAoW8CEkGjL0MX1YgNy/DtPZWW
kyLzBy2B6li6ykgcfYSHRiz9dBJ+jdEG4gRjiWUF7CMxdSKorqSsMc/G3W8xfd0M
qgG4jHcyTvtiLtJmZQGvtuXZTTNVl3FpyzFm/tvcfls7Tv7YgPk+wRuwcrqxEv7h
V5k8yiucc+/8+yVSJ12P1ds4enW0D6s1e2hk29uRSbPxOI4DUdqzwUJsNaTKMnRm
6Zrqk9cod2YUsZJptnyb4avhqAohTfPGLb5zvxaQJWGeLY+YJkFDxaIa2wbuIWtf
OPc82I/xjmL4FCq2eaaQ/NPmrpm/XlP5gIs+8y5VHsnb7NBtk4FqwXkihcuZ6RwK
nIcnlgeW3H2gks7GvDBuIdEpEY41b3w5DuQN8Nr1zd0pwuZC/GhKrhOf5fyROGGl
CEszjMLIMlc4ja5otYiw8jM0z3uSPClm4/EsU7PZI3rJ+wUobUOfign62ocvrftB
+lelTe5+u8d9mSQCCoBoYn6oHZyV/2awRFMYqk9GZk9Lsxumx41M7UCV2Q/EsOh9
hiQQWukNBZwmHPr8MVUDo+EddOYe1QPjnofATk9r/wAiQC1a2f3jvvpLF39VOZ70
6fK2pJextzpOTa4x8/tbFhF4y5rkjx5yXtmUGyoKDa5yUp/T5nwHcw4I4Vy3OGjr
Z0BjuTtGGkh3Gt6xOAr7XYeNzY9GoWreUnyVn3hS+tYY2UhcWLHd7geuYIddya+N
f87eJNTe9BZ75TahK3xa3EFuEXIj/H0UYgV43C+PAQAOr8KfzHwWlJc49NfVo21/
xHHko7Om4i+WxkyEwysByM4KUwVUwvS7ZvCEJulhyy/x7AXkYOMIhTaqg33RTm6Q
CYerhc0AcGuB3cuSj+UXr35TVP4Tq1bQS8tefHh/TholZwvkRjwcAiLA1eYCujJe
K9XWWyURTVAOMyCosUZq74UI2OakYS0iTCPuqqf+L0kdi1QCODp1H8Fv38X65zxh
RYqx1ouJg4sJ5/5PmW9beR9qWyQxDCzOLkOf3opiZUa9WwmwKMHZ9pmGfovmyFiX
bB3148swbVio7sJzVYV1HUGZar9uWI8f5zvJXzCkeLcMQgKVwmLoM4vLwNeDIPev
aoVW6xCq7XsTJJJn5t72PNj1TMBIrr0mXd5ExcyIKdJ6+aElWl47ziAfPXjT2T83
K+oDxOuxxG62LwlMYADFXz+XIfoR32yiozhyN3cRGAV39Aq+PAEEAipN9TWV4QSv
Y4sJmVnHZW6d7nbZJJUJATZz9C7psi35dPjKalj5if2zCRPrOlE/932fsOe3otzw
lrNyKo16IBrDL6HoDRZOD3dBcFOqnFPcESl0N6y7PwOjJRZ3gwQsba8nabxntL7m
SPSje9TmAOrvd8nk85fVYWjuVxKbKJhW8VqfuDCusae2J55weFppVbI9hz7+deyF
AeqzPcAOO7MHPIXu5Srzsw==
`protect END_PROTECTED