��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki�N�z�-����	�a�t ܌Қ��1�׻����7�?t�D�Bp� E�b%�U�f�p�@�=l�����­c����OM��}��/W�B��x�D���A�'3*��
��z��F���Н��ս�~��/����v��Ra���a�ϖ���i:�V��1\Ӊcd�e�k"����9C'�a��bsK�bzN	���|z�P�i9\��&���u�|�d��j�Ǒ%����[�Y�����W��2��%��]"��x�A��VG���M�m��]��ã鹾���m*\g7%�1�h�ޗ���d�Tģ�����������!��J�eD3]�j�/aN5���q�|�$�l!�������d�#��Kh�&?�GM`!m ,#�sN����C�[7�!��O����{q��m����ε��,��4�۸,0l��>7����S��	f�o��(et��$X�D�{���۴P�G'�B�K��UiV���Mj�]�P��e�汪nP����Dr?��"�?�wqR=-=�Xdf�	H��	��S�aV���{iq'�G�Iˢ�G��<��� m\��NH_�%�?�xm���U�s���7:��F��d\�:ו�V�)�����W:��=�D���˱��{�a���	<�A�^Ӝ+o�G+��R�w�G�r�L]}��2�ϡ�f�#uW��[5E���[�a?#��GO�LL�Ir2}ˢ��cH�#m��;��O�+�fX(7:�4a	�"(xy���%,�$��T�d��4��)����Ɂ��;���A�uہ���}�%���P��/'��X�:�.��+u��Ϛ(Ք�����WF3�>U�e���M�P(M0�H���WWH	��ȩ�f{θ�l�1ypƵt��Fς��7Zm�ۋ�u#�3~K_Q��Bh&z�o�mo; .� ����/𴄖�#l���Jg3�L�}�"¾Br�{����P� a��h�9�0��H�Yc���%V�4sKQ/vS�%Jk0����,����{�~=nN�%j��g�+ 6D��ˎn�j"���;���v��8&��a9���TQDN�m�K{��N-pz-[��.p�r!l药�TK�L	�����X<P���(ek�s!�GP�I�,���!��$��1I� S����V(n,a��6����sg��e���n�7�BW��-�����i�e�Qˣ�#7:�)}��7��X{L�E�����mgR��.* U�M'�
^��8�>��G?z�VT���q�D�;"1�nִL����j���*��$�\[R�� \�1��n���ɞQu�PA,@r�.=�ok�\�(-dҤ����`�g���ejN϶4M�e�qBBSL�T�Į��0�M���2�[���$�_-m���h&Xp�5ޠ��V)��3���������S�uڨ�M*�Φ\�-۴jV�0]�A# ��Rz�I$����b��
C4���
��r係��!������O�p�q;��ᅿ	��p"�s{ ~��:nT���7Y�a9t��aYc�Z����Uӽ�b�سE?j�9�q�:P�|;���Ei;���_�,L�B�:��LU�ΆAd��Swy��G�����"YV췩䝳��	�	�2��b��C���6����F�n+�Zz�PռR���c��ЧJ�!��`�-�N�����2��� �-u]!��](�J�"'��B�f��)��TP@�lP�����,V��v�ׄe�ޠ���ǚ�5�t{y+����춯�]}�فOEC��#�L'��#�yb���K
J�W�e��w��T8�ms��]�����: ����� ������	M�#9ˈtu�Ӹ8M�U�G��I�'�{,�?B��:�0h�veW%�u�F�~��:�����3L��h�Q�) �gY"��+T������X� �4rFoX���D=q޶9
i¬�]��u�X�AW�e�����}9�g��$%o^ϥN�߳��"���y��Af���n�(�H����q�V@]��m�1��dG�WM�DvЉfp�j��߁Kj���,o��N��3��/�����K��
�u>��Fb�E�?��Vw��B��S��b�1+\��dP�� �c����	�fx�L����WZ�}��+s8��!P�A8��Z�u�7��$BxJ����<�b{m�t���ýfb��/6�N�F��[W�X>�n�֓���{�� m'������1Jχk%��5���}a��t\������}��k�bJ�"b�6��H7Ik�?qf�q����V�Hh��i=�E��]��M�X>�3*����AdӞS���qp��rGTaY��������)�ؑ
%;��z���y")�kZb_(�W�h�V%�Y����k��i֌b,�z�b�vjU3�{L��.\`�ml�����`��*z>)��J2�)4D,���㶄m$�X�e�˧	p�}����^e���n�w͖��m-ӳ&6q��r�Qrd{qC�s�;����6Z^`!:�&Z�̘�w�5��p�m�y��=�jI��6�;H���Ư�g���q�����U`�O�D��X�r��M�h��ɏ�8�#���Z�DdL�'�ASEk��ܠ�!-ײ�򠗸%�������/��7�o�Z�Y��h��񫋀���3-�g.���`��=����eY�~%I��E��0E#�ps���$�g^i5�;b�٬*}y���H7����|��A'��!���G��Ş\l�J�V2��	9	�p��X*$Bj�DQ�'PEe-�]ƽ�:>Ǯ���v��;�¥�!b�a���Kɿ&�x[��@O���*w�K�7v��l��>��Ts�6���30r8֟�;<�7������{~��qE�$%�*�72D���	A��d�պ�)�B=��Pz��5�'ك��)6��x�tGX���N� _�sS��#D�=X������C7�qH�ƈ�Y�3�������Z�v��F4F}������+��Pd�v3�������k*�TӠ��&���Q��t�fS�`�L���\�8��4Z�7�Ԙ�JD[��h��6qB��=P�@}i�4�3����� _RD^�]bb�Qq�a���!5Fڵ��
�
��z�y��ֱK ]��W�mbe&z!�뭤��ɦ�w��=��R�>��o�x���m�Gk�-r梬����趿�!6d��զ\ډߟ�޲56��.Ķ���ûy�K�]YK�浶m��:��i9o<�����KJ��:�;VlxbF���nQ�ʏ`�b���g�����i���ޕG�Ԫ1`�	���Vq_ڕ!���]%3�/���-�[z2SR�t��\7��i��jz���7��q�F	�=��W9�ZR�e��;]�%�zo�F4�C���������ś�J���Rc��8�������^�}�^A,��F;Ĝ���l�3|�1��#����j�@C����aτ�~�%�]�ig�
��)��7ωUN=!P�;TwXb�{�7���6�!� �~a�F69$r�u�PZ�~q�n./́J%�䒓��j��<��59n*.E��|��5��%G�n<1Cxx9��eQ��;��D��GV^��0>�_{x\��������W�o��)hN����31�po.>b|tva���m��Y{Ƽ>�����ny6m���B����,����k��p� -�0��u�QB��GߟڵJ{��7��K+��i�[7o5z({���;Nz��!�Wp}�����a၇�SO�p�R3@���rL��G����:�0[b����<��?�����fPJ����@�ܙ�֨��Г��ᨩ܍>ncO�g�2��Q�KR��PD1�Х�{P%���pMh�bj���U�O��O�Ś�zQ��J%$r�P��AF�@��Yۆ�"�UEݧ"J�� }@��`j��RY��f�!���b*_�@{��@�̼�|�	)�Q�6]k>���d_�S7�m���;�g�9ܷE�*� �T����U�ՌU��v��k���-�3ϵ�;^�}�9�j[NF��@��"�#no�n��[ǯ�U�X���	(�q<_��@46G؊|�����.ފ�ψ�˦&���W�� �p�t���C{gt�B��l��l�8��L�U��\�;��e���W�9��M��e\�3v�g�:+ݹ��(v/}��v�z�7��{���O��U��C�?-#������m>d��M8(&� f��':�Ê�<6���)}t�v��oeU�˂34����D�[�Y;S�_��\8��N��7������٦�Zd,��{�9����E����H���>��+POe���$��ߑF������0O��!t@z�9�D
����Ac$wb./0�j����,G<�u^n�}���pA��&�p�z \��V|�XU<q_��򜅬H�iڽ�u�̮���riU����k�P�M| ���T�V��yp7H�.�Z�@�VFle���1
��އM:e.g�`$1*��h��j��g�+��Lǚ��1�u�����\B�$�:T]����uMxiXS�����LU��I�.#%f8<V�O�_/��JA�wx���Ӑ����߬ēh*�jl��8?�I0�x�6R�c�ꭵ|�R���)x*A��0L�c�]�`��Ĕ�;R)krחD:�'1�H,*χ���'{4}dE6m�WRvW���@I�p.�U���x����ѷY��� b99���7���o��+��D���l�~S��^O��DЊ����`�4#�8�I���X ��]�W]G����y;a�r&�ln�f�WV����c��S��v��T�h���y���K~����y��o����������,p��ڙ7K�"��j��JS2W��6N����ӥW�,kw8O����b�[�ndg��9k(��缌5SlU�%Y-h}��FUgIh�{�٨E�:��%���U7Y���|�G��{�5zhNJ���)�6���$xu�ׂ>.��o1�6�W�w��I7˅��pF0��'���C�z�woU�>���ccΤ�tp6az�'�����|�7H���fPKQ�ao`pv#,��֭Ln���]Mu�1k�ET8-UՁ�xA�n�ii��f���x砃,���X��OZ�0yť�*X"oy�F'�>y�x��J��F���T��q�T����_�p^���T*�.s���Ф��r�(��w/i8�(�л�U:�Y��xOlZ���<�v�ر����rQ�$��-�
~k�@N.	�Ju4����wK�M�^)�(22��{���;�`3����c���/I���uՅ_�hsK�Ȗ̻��*�H\[��b��U���INdm�2�v����Dƈ�x!�=����{,&?"d16p�9���K0-�k�:��H�*�̌5=2⳨V�5w��i���E��[
k�Wz��]de�X�}��|ڏ2�0��s�SCUƚ8�9�dO�ؖT�G;���j/�hu�b_j?ew�?�H���fW�xkk��2�S�Uh�:q�PyԒi1�q��3.�����C���ʘ\{��"5;���-��+t^pv��st%%� J��5tMH��)3�^T!���'9���Z@�c��t�p5�����`��!����ak/��]�7��rk�e)<�2�����L���as�yNy�ܓ�P�9f�/<1����n�(P?�T=V(4#���&r���b���|�J���
5��MyFuĕ� $�I=����k��I�ݰ�n<s�0��Kc¾?hx�/�jq����%PVwyq#E�/������W�43�dڿ+fv�.�0�ޜ��3����t_��;�R��vG->S�>���9��@��K����Ú��@+�s냶�� ��n��k�w��*����mm�i6l}����E-�Ƈ�W�;�Z� ��<��s\?ƕ=_}|{ |^��\o���&���O�f�TLn[�U����E��8�6��xiWd�p�O�:ٍ�{�7�6�ο��	Թ.�Bb#X�vw��,��v���ry�#[c)�ΤȮ�Q�@y[���7E�=��
TϦ�-E�j0��_.r���-��sϒU��}^8R��b��|q=:�=��?2�i�zb�u��ϿJ%�?-�g;�<��]\�&>��z��ƽ�(�� �0gq˿0C�1%X�����0#�w��7�М�-D�#c"�AR�������˳/��T��(U[�0V5�Bt��'�V6č��W$��-}8v3�8�/� o�W{�|/|m�Q�Kx�X�Y,�G��:���	R�oYC���bL�d�4�����[ȩg�~t��=�l�P��.U�//-���z�e�M�\���DX{j�����'��k�(1�����CuI���mm�Uj��$���t��F}��a�ߓ�p{���7�/$�Vi�H�������	�"mک7�66��xc�E��Υ�#��e|�-�݋�}�ƿc�᫔,
���^���dK��7dM�/��>`	:z���`V�5<K�NMBֲ�c�(����<��s�{gѹ�n��$����H[��D���Inlv�Z�a�^U��p�r�M��C���0$şohjC[֬x�+���[�R�˺?�j��jU5�Qa��L��#��K�_�+��1f���k_�&ʔ�@ܦ�����s����߫
P��	�QӅu��9E��8��.�㛻~�w��_5ʑ�I&�(��FuǉWw۝~����vPv�q	ǻ��㲥�?��ـ*Fv��pG�uJ���-����?$O�?���j,UG��⨼���^���{�
3�3`WM�\�,���MQ���u��RF�� MQކ����sH���jӿ�����w��	����K@���}��x��4ڵ��j_�
7ں)zVDD��������@�O%�B�����^	Cy*.8��~����,'� ��U�1U��5ԯ��(؃�JP)�1���g����ݱ�R x���J�Y��i?"4*��k�u�Tc'�z�����*\=E�LPQ���aMh���@��4Y� ���7@��M��o,�pW��w.����,�� ��z͟��fPMV`�U��_,5�̀k�{4��tY@�d05q�2m��@ɓQє���F�'V������h9]�.>\���bI����^>�۠���>~�p�] ���^m!Źc>�_[[��Q�R��
`"� s���'��
ں��b�k��W�F�_5�!7���':x��;V�!x���?�/�3��jOr�lXK�H�ةDL�ϓU�,��eq�� �6[g���VZM!(B�D�B�kҶ��O�V�~2sqMN]��!B���/��'8ENs��S�x�N�⍍� ��t������%hq�BI������e<Ke+�����2�U7�|{�g�cՏW@�y�l���By�ɼ�2\sR����r�-R�z7X�1����⟚Ԏ�Y-�sCx�+'���sC�cnY�K�è��@`F�O+�����$3a�c�O��	�؈E*�S
�����n���[�)��}�xU���^KXz O~����;rP[G�{�nY`hueO��V�(���ں���O�_x�ݐ>�Ԗ(ob�z�p����_�x�݆�<Pź�Q>ߣ�ӆ��0�*qT%���B] ��������	~��YbQ#(��2�%� c�`<&'$(r�/�-&�:A��_P�=$`�3�bjRf?�J[��n�l��&�j��&}�B4wڶK�j�	+����rQۯ`.�{�'g{o�U��f''I]�?���[od���(�6���lR�=q�Hw�;B\�������Y��f��i$ܱ�#����A��Z1�Fۿ�a,�������ׯU肸-��S�ĺ��=l>��dj��0�B�*y-���!�5��/����I5��=)xra_��X��'�ʈ��9M]\��i-�&4am�����@;���~_�x�c�糢��*�r�/�����[.�﹉>q��"���ع�X�"�+�rИT���$q�'��6�SZR��<I��a�t�kOo�T�u��k�>��Ƀ�LF�������.ΐ���U2�!b�%.�
U��y&����"�@Ь�cnH���M����7���>�� |���(J4��@k�
��� �(�*P�n��o�i4�2�$x��T#� ��
�jH�R��$l���V���܋<F+���f��e2�Q�-�1�^"�Yb��Ӱ�J�������KH!���`�����3�BzC�u����6�b?�j��f�)����y2��,�����?v+�;I����G@�>��20� ��y�Q�X�-ۋRfO��L�TS��)���hL3��� L>GQG���΂�¿R����qq�q���?���[�Z�c�H[ݽ�#�~� ��ۡ}3p��Q,_����P�#�v���%&�]D
�)����m���͙֜��Q�.�?���d$==<7h�	�e�O0̶*��5��[�[�_���ᓘn�+CG��5j�k���@��诙�].e��p����I�C�bG �d�:�e�ɹE�D�8'<�H
9A;��ћ.�R��H�����h�;��M$Z�[�k��:�=2H*��mw����}�ŁH8���D\'>��H���}٭PD[!�Ȝ�]q�g�}��(��2�}r�\1ZU�o:����ko�*��*e�R$���۠�U���	����Ϫ�������D��V<��ɼ��(��d�ށx*��++Q��N��x�m�6������L�T��2O����x<̠ C���ҳY���_���i�}"�kZm x�У�]�~u��8�W��P�1+���D"o��F\�w��&�b��&�b��%0���i��J6��p%P���Cu;*rb	#���͍K���G�d�T�̛��R�n�k,:{"FU��E�a���Hcx��Wi�'�K2��ȴy�'ς�0�A� �&f��cdc[8HFkA�W8�z�e��td}ϱ|͘6���Q��ni�
z�->��%�D(Y8J^m�
� �5����D�K[�]�S��Z>�*���c��ūeW3ig�G��<��� ���������̹;��Fz���2�ú���eK��pt��󙌨2r��R�n�1���\MJy/� �&�R}T$
�d{F[��%w��5����|*`��{�'<�k�zj��W���?.�͋���]�}�*���D���:�#��lqq=������{V��������j���d�	�}����P�	�Ք���>�A_�)���l1�KqG�U�m�#Dw-wl��U�t�ѹϡ��4�l�cZ���Q��\�־�g�:���̒����#gW�]v�)��nDn:�y�z�J}vIs�w����&�pYIkE��tؗi<������jٰ8�?ϐ�{�F�O����Q��aNgx�ك���&�,�ܷ��Xk�AXu��	��Rh�{����#��2-���a(�N�����5.�0����#N���e%h�5�%��}�y���"\�����Fy}8f�m�Q�aO*sg���Ü�T�xb�#�ud�9��Y�/���4���1趚O��Ky�ج����U�
L(R����m@X�҆�� �R=e�O{01�-�"��|Ҍcv��{��;�~@��A�$���Q�~.���d��������1��cО�Ǉ��=s�F�4����!DzG(L�Sp�tS+��P�p�x&k�*ꨫ�yg��E"��&cǿ$�S�E)�;5�ՕA���?��c�?G�g����K T�1xm��w���>ﾳ���ɣ|�g���@��ډ���|w�*:A�!ש�`��D��v����B}|����ѭU�ӵ�ttq �&|���(㗿�n����
�o2/g�#Ƭ8�I��P��%^<d��a#yCɜ���7�K�1>��2k�wA�|5MK�_g�~3sH�53b�n9[�~v�9G�*��N��i�G�y�E��0�S�Q��_1�W�/�8�?Rӵuh��b��I\ATR��'[~��*T��x�1;����!q?�A�q��I�4"�!I�8h���?�_�Qq�(V�;$�d���Ќ�7�5��G"�:kC�N����9�7>Xm��3���%"��6>�B��X�<�����a>�R�5�Q�ˇWs�zx.<�љ}npC��UQ�<��/������W�-,y;��b�μ�W4躊�B/lz^L$�񂩖w��n�D��w�
ߞD��ޡS�$���D9��<e�`q~�O�����'z�LۍC� 0^M�v�BI���Y���T<���<��+�w �^���QB> �J)��>q�В\3{}�ZgD���7*����F��64��L���g�-8�Ӷd���%�3�u��mB��6iGr�w�a�Hc{Y������I�E�I{�pʊ��K��v�t��t�ҧs'܅Ƅ� ��QG��l��wG�|ǝ�g�m�Bxe1r4�)�R3�W�vc�������l�e$֬������5?K��J�x�<�M�+k�J�ߺQ�ٺ�R�̾y�fR��=��t�'���
�	�Z��Qڻz��sL�opr'�eq𯈡�[� �{B�Rm���C{V���{�ݠ�V�N˻��c�:$���aa�]����5'�Cb2� ���ʒ��q�=���_v2��eNr�]�¢<��(E�Q�R�X΀�æ�w}��z��]�ڡK �D	ݱ�t�Z(���D�$��I/P\�2R��~�o�S��P�H�A���%� ���{o�\���N��%�P�;^N���j{�Q�Ց87��-�$F�͕�]i���%�Y"�Vad1�������j�&�CUS��[<��Ǫ�R��e��J��#�������p��)�����J�=�>�xn���ztA?D*.�/g*�J�d�yHW�HVM\��t���V����2��ơx��9�<�iGop-����.�F���� �V'Nd�=I)���}���M,s*~@�����������x�B��uh�vN�����Z�l����{*"l*�:M(6=z�s�%�U���'wX��1��Af�y�|)U�jx�zqTBr$`Sa��X�$2sHzp=��L1�.i13^�yWn*���1q^���5�݇��@+��#��7{�S��?)4)�������M�+0�{5��+H2�# �WP�ܶ�tI8͖�:���m�B�|�'`^��caC�{�"���#0=&��RE> CB	������8{�e�չ^�~��֙�&���].���Jn�7h�jU�o�R����K�c��K��K� ���� ˵�;.�O�mf_A���qF�,d�h�����%n3R*�us�#�}�	�y��f��wwX1�#V�K���!�y~޿	�g�v�����1��;�9�x1�BVn�"�b��v[��w ��=GJS7Y*H�q�B�[�������1�&ґ��>1v\(W���=���3Kha��~�2�k�=�Z�7q	�����	�/�F�-�4tĒZ��Dɦ������a�2��I�f�I�@��P��l�^a�fV��E��R��y�kj1�Zq�$-MF���R�U̘o�"�\.�ZQ��YR�v�����v�)*/,UͿx}�?
������%�Z�'����J���!�~wGD�ϋrO�Zq)��lk�y�R?o�bRo�fX=���A�Z]��y�9��PH��[w3�I��^_%�QH�t7 �'hW:	����Jyq*6��Bt��w&s7�!�D�u��d�:�g��
"ϱ�?��1�,\�W�ăl�(�0�g�Q�kJ��"9(o �%%��w��g&���Ae�4^�c����Ȯ��3��ׁw��Uqs�2�Ř�犯2&��J�$�k��1�H*��h�G�:�=�`'`&L��1h�����X=����/�!u��8�E%�_��y=\��I�n�e��쑶?c���]���V�'�-�� �ťG�B%~��yh}�p��!�l'��!2�࿲���G��a���HG���%ɚ>ϕ	.ּ�R�~��V:m�������_w�
�A���]�6\ޥ(�A�L��eA�Uc���/�,�0n+����,���-����cGWߎ�oU����<7UR�2�w��p1�3F���$E&_4�ɶe�Nn"�y�}�|��:7����j%.�к?��2��e������P0�7�M�1�J�V������y�����?�����,#��+u�b1�5o�d�����N����� ��H���9*���Es��8o���ˇl�%����t�8+��܃�����ӝ���΀K���W��F�O���V�3f�Y�U�:�Ξ���cE�BZ�/�Zz!
=�u__�v���b����hH�[�wq���=P^����-�'�#�d��*�9\7�?�աNF��N��]�pԚ��Fu�{#D��Y��"����~�>��DG06p��/��۫mHJM�̀)P�[���p�WH�"u�B�s��O�X��t�"w�|�qcY���5uTu�8j���Fd��y�+�#�y��Jkb�+QX>��S�k`��s���&�����,>��k���7��!Z�K�s�����v�1*�"�ȷ��j��H�F
e�7�K?�A3���ޙ�-�C�ꧩ���K����$Xx&�8_z��B���j�l�Z���͸ɇP�S�Fik�,���I���*����*o��#��� �켪�S�ktKI(��u�ǻx�׀�4��󃮺?�$b&�h�g�iK��I?���ve}��[��Y _�bHoQp�Wį���寊6�'4�R���TՅ�k��7e��򉬖�A�8qr�Dw]~�N�*��K�,�ŋ\z)���v�������ѐ��?�s�r�L7�;B�C��:%��QޑS�(�t��p2�3���l���[�_�"�:5L#4�:����0,:G�P?,閧tϸI��<38�����~��F�#��1� �_z,��q�r��y�M�d����51xAq�'��h}dbs̶����0�ȍW��*���g#
]WG�"����Q��.��F���s9�`������o�-Z�eӍ�t@f��_�'C_�j޻��*���n1��Vmc��#cr�8Gm��]�ja`P�]�Ι�Aoq8���{7��jh���u����Her���60j�Eі��\�wQ"[���.><�7j����2������&N�"�7=�D���\�C43G��@�P�8^��/�Ђ:�u�'��
���b<P�k`�j}>w�Tׅ�,v��c'�aU;^�#��+=�xĀ;�� c�^��6�,pAi�Z9�E��xe��H�"Yj7 @�f��6קN�����<67���a���O?�ڟ�畈EC�<fI�S�u�"�	��~ݖ��_�`3	��޷�>��WQ�/+��a�{���'l��3�<����=��yMM:��Q���w��&���(�o���L$�P0Z�����M4FS-��J韾��~��h8FJ"�jZCܚ���L�:���;�H�0v���:�o�p_��a_-�?"i;n7��*����Cu�RI]�-����o́;�T��6&��?I-�}hd:!�LYl��E![}�+��+�mBA�=8�"f#�>��!QLh���	�����qz̆���6O��$�sfJ���NE��6��Yc�6�BfQ��{E�G�m���(��2��|�����؁zx,����1��9�vJΜ��F0��J����s�������@����v��b��b(��/�/��>�{;��x��'~� ~\N�D !Br�'u��S�����T�Q�c9:b��h�J�9�,��F���<���v������n�'�q� ���ṁ�E�9�D�oQ���tB��o|�o� 6��_B�ϊ�	���t��n�/�d���[V�f~~[W��<�g�1 |�҇ap��Oa��h^���8ʢ��W������0��ʛr���WLݜ�!"���)����rߋ�Waa�ߖ��ی��{�l� �����oW�c�jE>:�[�7Q#��ú�I����#�������y`L��3@+ݲ�V�?7�o��bR�{)r�kQNz�	�%NՒbH��2��A����g ��.��3ɜލ��Φ�8x��r���܃�J���#�S�9�Ï����P���uH��/��P��J#���a�ˀ6�2z�ǃ�ӧ��!���S0y���a4z��䕽�{3� 5��辽�M���0����x�G�3D��c����c���x�c�nU��q�d?��^�3�[�׫��k����Ƴw��e�s��n��U�K��i�d��?~ 6��Y4IW���͛�Rh�����N�¸�Z������Px�fY�G�b)8�C?Π��Ӥ;�y�A�+71�BՂ�ae����������"N�_^������
r��3�h�D+^Sn����t��Jb�8����䓫;����pS���Y����H��U�����5�w� �uƀ0.�xy��Լ�t� D6*�|��&= �z���XY���'khbN����z�({�����7\�<>�R�j���Y9��~�h���5Q�#_�$Ŝ�j\���e�e��8-����?��8�ꎘ�M#"��?�a����y
�/-M �AĆџ읡X#1��tVN��z=~�F�Xi���~�?^)� ;,�xE�P���	�$���'P4�5��8�S5��gk:x��ZƸdEr4Z��?Ȇ����T�Ek�������mΗ	XeCq��@��Di�	%��8��q<U��i���槕a�<'A�Ѭ���B��y�3la9���@��F\7.�	n=��;�PI�h���$��
/Yc	�z!Oѣ��sf������8
�nT�����~��k���mpM��(���Zc�7��mp3RT݃)��-	kt�W�ʊ󾰎�?��\��Q�]dQI����� I`�?9(q�u�]a_3��J���8�K��<�:��eD�N��2|*�!���1��Vju���0"��r���oэ��b�
���mZ�1o%"7ֈE�tH���7��6R�=r_�k6?]��[t����o�ɖ��F���{x*����W=�q�xVN+g~m)T�{���SM�ץ�RX���!0��*<����4��y�A7u��o��I�r��z�_bBLp����ޫp�g�SԲ{9U�Ӈ�R�!Q�m��,b�\I�W����1����D��V�K�$\�.�
�S�r:�!�K*���\�Rd��tR�_|J"HJ��qoP:�8���>��N<��
f�r�^~4À� ��e~��a���V�MG�d����P���CxS��'9�����;�F��$2����]G��7fCN�Ϫ"��.��LYg��0K���q<�FcXgxA'0!�|W��B*eB}���X�+_�grɖ�)`{C���Ll�A�n9��:�-���Hl��'�x��ڋ_$�*���a�k֎ѳ�}��{��{��m^)`�\A=���@�u�@�~]�!�z���(6�xD���]O���[��Q��n��>G� �S��B1v�!\���+ۘn.U
7M�H:�����˛d�����Q7r)8r�'�P��E��,�ͺGb��uI�ƚlȠx�B�p2��;����t���"�O�FV��$_�o����$MQ ���.�N��I��f��j�{k���{)�L��	
�8�>g @L�"J���9�z*�����y9닲�"雫9�#嬙�:��Ѥ��cN��n7�������+;m��c�A�Twi_6�"x�z��q����4.D��L�k"E�9�ε���`��i�XR�z�]�>nlfYHĶ�58Jڹ�)���$�)��3��e9�\�>��%�IQt��im����duxv>��=���6�r�'}��4x�ק��2t�h�Q�^E�����>����%�5��:g�d݆6Y��e���ew?�z��?��L�=T��Ԉ�#d��L/DG��$D��q �"��=U=���K�������O��<�a��{4�*^�B�>����C��9�ں	{G��ڻt�|K#����Y��'�t�ޤ�V��f�Q8)5����O:l]_6wa-�}��6��=.�<�5ކkOIQ���[�?�;{����6��G�X����a;����?"�I:H�}��c)(���
V0p�5q��~;H�������!�p�z�*�x�_�9�Iά9 g
�7f��'A���dQ�����t��X��`O�^t	�x�����1��L�"��2�z���~YJJ|&�#�@�r:�ޢ�,���UV���hyh�{�p�v���݂f=,�6aC��Q�U<g/뎤���V����hL<ĳ�r$���6e��bL�4r�?���+�@�$;$}�S!�Y���?��6�OҌKҒ� � ��ɐ�ܶ�X���cA~D ^@����[����s��3M>�p��bI�R/r��W7L�t�����nuWo���x2���1��|k�b��X�軬@	"�aB�?Ƨ�@���P���f��)�����Ž\p��k�bNAo�E���e�{�`�-�qQ��Z�g;z���/ŸN�ߤ)8��I��,�.h~�a��=y�8�q_�T���fx�%����r��UH>n��7�<k��.�]!D��������f|ٶy����-�_B��`'�iҽ;q�4��]C��~�Ƭ�j��o�.���ZnN��m�%+-��O���8�qAz��5'����e�E�(3�8�:� �p�<��Kl����}3����.j�B���)|��>aH?���`ۡBO
�B���K��Z�6l�u���!�x�!�۽"�ԃ�W$<��JI��d��ͪ�+�����Hv�7�HR��N�����Dxjus�'(X	�$��/cM�{��/�����.����,�,�C�im�K����K�ڞ�^B�O�1z��PD��ɑ�D#�,��+#���H��/�E����Y�P�����KM�$��[;ֽP�R��*���������E���*w�����}t`t�6���
eT��4 ���Re#��w+�r°P��#i�;ʤp�:*�M������w��#y>��#=�3�`�y�h��O����ի����]��;�1��l����n�p�P%��5���mW���g�@�������3R�uV�j��G��LD)��^�R���?��� �Zo��T�J+B��Z�x<uc���y�h�OW�֭f���R'/�Ra�� ��:����Z�~�4l�� tX��ش���9ܭ���"��Q�Lm��)�ax���ȠΈ��M����ꀏ��R�taKpĸ�>=G���.e:���ƙM_�2��35^2�	�I�rqyj8W�gW�r��J�6�[��w��̶����L�?��tL�����m�$⇊{�z�}�_�T1vu�������|c��A�WZɺliL�����;�Y��d@��V�@�zA�H����h§������hS����Þ�4���6�@�n@�״w�lYO���u�� 7Wm\��[$TxQ�q�
��<�(S5���ڏ�c<c�)8D8~�|,>[i1�ͣdpdv���1t���)����X��i"��t��{3;�!���-�(v��'�9��f�`+43�����B��8?���?�������U�3�c��c�ZO��l�%pH:4)�]�y좱q��J�)r��Be(E�;�<j��J��G��:�΃�^��w��a�BG���YS���x_�*$��^Rb�s�_O؞��8;|([#�ȯ�RuSɘ�Z����Lgy9y.�C��Q��8�<�8"&G���|5������̰��7	*S~�8�qD���:��O��[ӷ�W$#�|4��_&#7� �O�)�~q�D���Q�ʇ&��VY�~ĉӯdO�7^M��������Hቈ&R��L�)SY���6��d�m �����6�Rl��L�y���M�K�H�{S�ƃ�`�Dv�U��K�BL9�֐ӑ���9_�$Ue�	Y-�p�nƤ�$�/����Сxc�z4�F�-�t8@X��}N��|f�#K�k
�m�Z���XlT�C@f��"3��XT���N�,�֭�S�Ju3�y��Dɳ��2�' ,�ν�=~�yuT��^`��O��������p
���'n~p��m2X�]�����V�~��8��hQ\�p]�eY�z�����ב�W�m���5�����O>AZ��f�N���ʿ��}y /�:���t��U�l���&b�T���
�c��MP�6�ǉ�x�[��?@��I���x�;w�^���5� \����Я�n��{����)|�3?�){-��Z,y��)rN�}9NW����M$���{z5���</�-7���%�~�R����Q}�͓�}����ʍ8_wz���Y]�X�Û���G,Kh'[ �i�Kq��&,:c����H�v�B��SK2�5����"��<eX�*�k�� �zk ���	�ӯ�d(�i/�c L|��0���P�� �D��ݰP�����X����~�pv`9b��A[�~G@ܬQ�[�L�W�Ѵ?xD`�1�b�w���^���@׾,��ضD�IH(ɥ���6g��X��i��.̎�fE����C�6�0^ч#v�[l;��!�
�k>إ���O�C.g�Ε�ȅL�k}/u�?)M�uI5��o"��h�Mh��+�_��]x]�6S�V5_�«N���/��9o���Z5s�D�u��IuAjZ�5N��������{y\Ti 1gw#st\t;�>�j��fôA��h�9������X�J%D���&T�k��� �r25����"~�䷍�O�"e����CD8��Bɥ�����W�B��=RG����P��ϲS�
��i�!����?�B&�n�JGC#~�S�v����߃�9}�ɶ��)|���`�[�To�^OD�`�m8Ӝ/DYu�k5������ͷH�&G]�γ(zĮ��&���v�7�`����JdW���"�H%pe����W/�����2�t�K���Yx�
ʬ�Sv p^��>+�u�E�:�}�t$u*�a�TMP�)�jj'�2��4��e�#��Yq͘�������o���f�X�g"B�O�\ڷ�8���z�\�)�0��@r�<����/�&���5�X�tv�Q{��FR�:UC��K}�s|��.��i�����VZ��p�)�q��#x5B�� %:c�0�D�ݺ{%�g�/}�^�Fv��}��G#rC\/��������Ơ��ڊGd1��%H��	py=�a�Y�����jA|-9Wd_�yT: &Ob��<�jϝ�u���Ϫ��cld-99Y��7#�P�����-���@�/�H���v��e����A�lɗO�Glt�ؕS�ȟ�Fn�U#v�8S�Ho-]�r�����f�Ć8���ϔ_FN!r~��}Yw�Kr*���t^S�9���ǣ�����=�;�|p�7��-[rڼ�A�q�*	4���©�@pzOg8�I��g~E�����IW�KV��h7z��F��O4{cC�b�#����>�Mo�K�R�z�v�?�������k�W���-k&f����c����"eLLf�"�dXO �,� ���m�r׋�� ��x�؃9J���p�Q��&�e"ƣY�#�\�R�[�5<��UQ�}������S���l��	�B+�bB芤S�ą������V5�jWG��8\"���)K�{)l��NݮG�'SXs�Ω��q�湥��*�G���}*G]�2��x �z����S�o	5�D�N��Ę��M_�&�N�g$���^ s�>��P�r��?zw+@��٘$�&<����l0_��Z׶��V�25ԩ�x�ً�Ӟy�ƝZl�Q����@:�\�q�� &?=먹/t�\�����o�޳f�j�^5��̟�	Z[Ori�y����+-���1�`�a����e�+8��r�#�wyd}jAyj��+ky��6;�/�;�Z+�b���uJ?���7L���^�jx�T�O��t$��w;��"��N���_7�]�\D7���G�I�s<2�",�,�]���a$�4db�deR���	 C�����A��ک\�kx�Tl�*^�� ������H`�؅�/p�i9	%_������?q������el 
�*o�܊~)#�fDUS��}>
�cſ� [�:�ydɾ���BmC�A�)D�6���t7�ߨ����q3�:y}��=U��9�~���x���Os��lN/���m
��W��	�����Qء�t8.���K���Q�W��A����������4�#�S��LV%��5��4ܵ����1yJ�2�B-�:6'��Ј��m0�wPť׻M�ݿKO!�d��;��V��^�8��*��VzBL� ^�¨./���T�)��Cm��|5���G�E8��|@GX&_��tN[���+xb#G���1ߜO|ا��,ᐸ1�t0��x���!C0)�W���}.Y�Z�9=�ħ�fK	�z��"P���e�e(�	����1�nI���RH5jm�i	��G�kV���VƧ���"����ta����h7�n�ꡗ*�����I\ xp��qiO&iK�m�s�
�s��6 ��/0����7Hk$���o�8�5
�͙Ld_@�� ��_�H�H����@b"`m��}��|��{S�2;�� yC�c�z��������撵>�P�D�.A����aihï�����r?�XA��7�'1���_�g�J�C�K@��<��"�c��'! r����I�t�w#��/�
�W��˽	\¸��B����&{iW5�\��(#�-wI��m�mHC��T�#-�Ou�|�fMt6h�4�I�nl���W����K܊%�a:#��]:x�0ǍW�B�l���7�U�Q0�r�n5�I��&O&v�cj�yߐ�C
7����+���7��̼N�S�3������J�%1��:���E7�x*�j>��lt��s�GI�o��3�7��<T�=6�<�L�JG}�M�w*�cj�QE1������h�3_�$j�՗�0;���ϕ<�kM�Y|#߲�`{ߐ�����
Ć�C�����`��>W+��.n���b