-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Otb3Bp58z/HA8A81X//lQdT3Eh1si+sckv1UDWjTvrOcBpr2Xh/iJH00nrm6fjsE
2UsIVgImgH6r/cFiZ9rFlxiuzjTfprP+cUFDlZzHUSm+X7HS3I3DDjsRHa+v0x4S
dZGBpeZALPmBtVWxAT9hkiPZ2Fhu2vn9PUVYCv0y/Z8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6336)
`protect data_block
mgw25dcKj2bjqC/psIPUxEs5gaoque/TlX0Efh58zosrE9t5rbNofzlbCg+Es/2E
FnTDUtTHyO+nE5XlJoVtcTj/oRDE7B70zQ4wBWAw1MAZT7OqVW0ZGPeIVam0T82L
SsWlGLrOjYWehtOAymUa9CFVLTZ96TU320P/bher07lNf8MJbgcWCk31Wo2iJUOA
EAHFR4kQaWkBZ3l7Dpe3JJdUphN197695ciSQJ3Aev6JUyIuiBhHish7krx2GzK3
ci4fraBRpV/t2DxavPS2/8LLOtxan4AUtyrtBsHbP3lX7eJx7BtgI2LwUo6oTZGl
QWhLIiRNQ9h4hJ0nRMF4vzxOzbCCKWXsMxNLifq8W8bxf3gjaSnT3K+aq1eRBXRH
CDiH+nfHaGDz7RxcgvzVHxGkeCAPMTxf0wU7eFDzFLBAhjgZ+dCgHSv79XzoGtTF
hdZC26B3Oys3g9GFRO4C5KknfRCXo3Ey9Gyrj7aZPj6DIl9NkPdPTEhCt6N+ki+g
br4+sn+/9AHKOUa1T3j2cDSOWQcYzQtafmmDIM19HuFg9ug8stym2wNVpwxhY/kL
++qoJFLq1fYODwVKW73pKJW7icr3fhq4lQAzJu829ytEBpiBf1rxeEeqzgQEIQyG
j6/ym+R4FdOMckWWpUD8yuVLpfWKhPPJLbkwM+82CbK+9JYIh29/YAMwm6zTfyT+
is27WYWweyfPq9k0GHk4ejUxLETph3zIhK2S5kIlDvIbiFIHMspPy35v+BxIFtnk
aXrepf3voYG6ayx+yjDUT3Cvx7YPLygA4hIAD1JVsGuXl5+sXrggspGRftRbo3tw
DNPfQS16KK2Cd0J9s/w4Q/lwHzaf+zBRoTzXsX1vRwQnmao66FzvwC2gyRmkSEoN
lNFzki9aq6zDZK/klQgPfttfl/H/SXTzROqEzkmsJTmCX0lrQ4jk4tkwapmdXORv
QPWNIElr420tKFK7SiLb+Y4LLAp+m/z6eN3F6SQ4g0abPNrzlrBoHLPTPxujRJNf
CUY7YGvvCmUA+92Cl8glUqU5ZNS9U3Pnpd4/yeoSCk1I+Kz12T+imuM1B0WdC3qb
qvD0xzZ8rgCN7fcacHPjAYzS0Sl6nVe9dEl5MFWVgXwjqaKJ4z5EOqBCgEYTg/q6
FebRDA5TJt7XFDK2usSJv8D3gv+tYybh561DipiQ5RYETl+4gbLgDpgKj+2XJAfs
6dhwyvNW8zoEjGRFbYc/XUzyGBrB52gyu0tmj/jTSJQUn+7nSuZStoXSJgWj+3I9
g5g7NCO0BLBFJ6RsHKsX+c60EPitRXMZxXiMQnaQRmIYLL8ThHKsFGOvylEyD9KJ
tMdJUTs71wu2z0QOXoImb2Yj2RjVb7wGmQ4RkmNuO+SIKSinlb3+M5Jm4X48wu1p
DkXDFYPILIaU3DoHdv2ZnPFxHUZ1GGLQj0cJTB3YVA1dgKVv7JdmyU7Z4PH2unez
28Z5DPQb21l1CLhiweYhBxw6iWogXAK+dQq6LZOjHr0CJL4CE7yUiFen/FcvEXAJ
op5IPm9RdLuKe3d9kCvb1zfR0hD82l/aenrbgRt5n1Ep893Jq1dRp5HoLMjGekZ8
W8LVVBqs8bJFG4MB1XQqH/cpfukaMeWdHsUScK7POy7eFZtWlJQ/vd1PRSQ8Ft1W
dDGWU2yphv41Tkr1Vl3Zz6s2ont4quVNMb6Nr1blZJp3vNuB9SbHf/dpo8HVG+Qw
cb3GpFqBdi3t+mSTNx2lmIXsVnttnoOcoPMWwVef/KDFFQKL1KuCZ7VnqyLa0Bfb
y3PZxtl8Pn2YtLHQSFn4qdyqqn72ufbvw3l/vnZ2Fv0M1K8ytUBpU5lrGVM9l9EQ
494DshbRy1DFyJjpeUkODpxodxy6GVm3vc/RwCHN+Q4ikwzVS4Udg9N6frfwCy7R
fPBPhSyULaq4EpLWb7pfdhnXj9rEwgl6OTOaUOwsn4jsuIulAlTv3ogcQ3wNYdGW
KAdrkEMwGvWSbiIAA23TE1g0RSVaXbocdlpSfaRtyq4wBgnBWHW+I/PzwgKGv+x4
GAebmGPVRqJRrRupQSxQYHqLYoCLrc2Zd+/caDjzSzWB5MpOKpwepxzWjn8ChjKA
ls6i18UUChpwpM51RJJit7xAztWqBBvDSuESYYP2tnCvQBsP8X4MpFCl0nOfPAo1
Fh6EhlWPiDTQAQyiKTSUqlDa05N3uWWrNPEvBGdoCBD9AfL2YpxIAG8dwC1aqcwA
MOo1J6Q9r5YPc2PBrhcK79SDoQZtgDwIhf25aIjyHRzvfu7VRJgwP9dX5fMbvwri
7ewSxSheHJRY2jV6s2+nz7G/m43rSWdyJTxUoAiHBfFi0TGoWgTOHr9sgEoziBhj
1gYYwHuIA6ksQy8jY8oH3QR9hdg4IBzYInRIp7LBxe2KsorDyREa2ajOUWiM/V8p
XMz/uy9oNG3jQnxs0mGZBPIalDp8vvbFTi074azS698FxyNBNlZft5GgxjHg22vD
WQJLho8c72WepLG6HegiVqwLkfdCmmkOk6TzYpHiyDrGNiJfUP9F4Ueu5hdJyWyp
f7TdlWn8l/rNjmlgmEX0qcMx6P3T4hcuXh7aqVfS/PhkboXrdZkwrS9ZFzMtLfx5
QOWspyUD2Ibe0v2DL8W4yPtBKe5p80UG/DiHsnuAAGhX+wSBxZj41dZaAM34vcVm
w6rxSI1TFZ56SW10J8nrgiVjFB2QBFGUTiOITR1JqaCHkOk5dWKrows0/L8pGmGk
UF9xaUK9njMF05uLsd9xP4jOCuwsOh9FANi5xdpJgXisD87kV7sHO1CPAFxXPabo
GqLp+IJFJpzTH6uA2D76ebsDw1mz18hlThTI1+obqbe6Os9nlvkQe0Ymq6e7octi
DKlyZ60ZLwWA4ZVqHp8CBlIMDb6hK0WupIFVocC+2BMJhBWOccLGM1nf74HP6UyM
QkWByQ6eXtXi1bZI7wCCiVu17oqp0ZDV7KNepvOtK8MVloFBqWztKlgSw6lgx67g
McQQJ1K9xOBatlgHG8TBLWFOl1c0eZz1WxqmFrj6ZJvLmhTATRwdNlpx/Fe2h0nA
R53Sk63VdC38sv88yzlUzuazQputp/Igg3v/6/BBOFSbjZyAXjTdcwhIuhCbOaRT
xe75mE0SwnYtmVOPL72PI27+yZlgrnIUoBDeNp8R7KfFzJHWK59Fl0ZFEZZQHsYW
Ed5wVmLRGMs7XocSiRYKehX1m8iXOGzsVgP73poG4QOgNsDJXw4XOHVXIJLLn1C+
JOwRGs0RQmrVqlQ0lEruVw/iavD3VZCN2oAgIplwWj1FcsgWFNZufggQzpsp/0yi
D5vCmAPZYvplI6jxeEam+/vjF0TAp4t7BaWECH03Uq+TngZWo3axMg42d7mA1kch
IRoKyqFalABBy++qDmrZjrBuU8hbFGu7d0UIFI+OkaVjCn2kpaTP6GHJTfUF7u/M
ys2AUgdNsDfNXelzqos6FA7F9K79jN20jL6C5xsqX3YFegt3J/v5bXASa+IvX/Tv
sCXJYQCHyRCR1NYn1e7zgL1JH2qX5fpImi1gMZZMoYyRQfxWQgVW4/AFlTQaHUeM
MeaN18P52bRd59CzUtgjVpot4ySrnY1aUXaRetpJlHcJW4GFSc9FfaMDIPCtr1w4
ut21qksmzrGGdNnScE72IuTjeEAbcG5Zt+oV+n7zhWMFmF1NkW34HJ36MfZJM1Jj
cnikkgLtPYNONXSjCFAJmLF/CipoNZwnnNqSpJOv50axtzuDP0flGiZ12BtkuQP0
12y6TmBRcJL7OOgUYEugolg7n4Xx2+tgNQc2EW8MTSZb5fNEgxBPer9cCWXIZJiF
G88CKba6GoZYK6/YARNBAaZjXfAXLks0lPi1Do0eJ94DIRD9fsRN73FvuuFGEJ7z
L2Keu523rCz7e/vOg0G2ABmOnvW4wkwWcsKr/8CAAtA5fznpIKK3m5oiwsg3WFGI
uD4QsCyFRDM3qZT7Y7Ccks/G0aCaKTIPLaMLY6on8Wbosamh3CjaO9HdeUB3TSlM
KtVGdt1CGDqsJOBFP8OPq9ecBClaFUmccyr4dHuypczAwWGH0pIaOuuSsVtcsN7T
1hiyfN3CcpKKGPVS2as0NYNIblL1bfhvrGKD1t+eMTfpSQJZ1dJJgb+e1DeEkFdb
7gPfCHMOGdR728tNopaj/Sx0YI5JyY6siNvcJpX071Tgos1OkjSLBVXXuPNblZSr
hdV2CrglBIQoSh0wnwiWJaenvC4qdNcXrx+9yx6UV1sVps4iGg0kny0+nvuKCdL1
Y/7mRzlQsMMGOILXHmQv/n9A5tlYIEY7LmpPgFlRljMHxoOB75m8S4FzrbQ/Fs3X
Uc28rmxwAUfB94Wu0CXJH0DPjk5N7DJYcJD2eajI3J5DWjGlZnB9nhl1DF5qpTTb
3Rds64k40HvefiueXiLWbxeHAVgHyqjomWI51BIOecYJmAjwfXG1k7QlDEs6xOr6
Cy3x11GFmEh6hHXZ27tsrGgZ6ggbHWATwRD7ICPyyLOUTEpjM4jg0jy3LRHdhG2u
cgregiXT2zh9JGhLkBLS6BJvdNsU2k9CNTDD06N+fR0w2yyRWSLmA+JTDdZxxcPu
xX/EDL97qsteQBxSvkW5rHGXvn60bDhhJ41wERyErJ5lj/DUTAiPC6a06B/Hy9La
4L0nPfPfvJTE/VyaQwYm6urasNBzlMTYPK/i0IEIQUbDUuPc7HY8BCuoAQM0aEVs
cZaZGPn42sb+/DLX4ywqZzjrRVtO5ClJEnRiANoSR3vSBXT+2iRahyX2MbwL285H
2Ob8VpCLKseMCXeGbszNXAsj8PcxT5oZEUtafyHp5c3zrCCmQN0yEFex/NEi5cjO
SDM6Pwu2abtfjWd0NvvXFFzqNefrHqT6F53JotjieqCkjWKD/N6G0FDtpCl1tln9
KxDYu0JHLtNMwZVHADII1WD5UxsgTgl3JYNEVwMXQ5pdJ83T3jQUbR8LdMpwR80O
bNbABEDMaq+/D3UHvwXozHuVLIHcUDJqQbiQpGPJ98RM4yS5b0Ya+FBK8jM8My4R
5zjBsQhLHwAac2882QkVHcjZ4omAuFz1qWl1SOa9NGj38wwHUcsBeNwjoqwP2zOp
sIInvq7QswAKjvSCtlr6pJZrHX1G4clcM1QGxe9ri9x/LHdXFiz07dHyh+1i2WOe
mTVwTBaZxXrQSK1srr6j5ihEMxZQ/6jk+1VYQX+DTsav/KJMCH0xvDOJBksPBMPl
cnvbfOCnVWKkLrweh3XKOVCg76v0/IWLyjFwV4MW225lXktmKfBHrwUDDaaQPWf0
H+fKJET4sP27oCjpp9HqW69ZiIdBKjxtunIDFFXVoql4yVSb8bbLMBxWPPcG+E18
1gzSh9O1OYSMGtjinVrM3jZsXvmN8pzWDoAnSfTxWnvz0kea4TBj3LqVAus47tbd
puZKMlA7Txp1E/HFRY9l9Xcs8+i1gy9bVHM1EEahTCL2BP8tFDo4QbfheQV8ZCKa
SEeoBZGHLq2D+ZO8wkrWvZu/Rmp+2nLU9/fh7NfHEGP1oMSD1ZAguTwd5+S7ysVS
1X5UtLnpOR6G7zyIVkV2BL9mINw+Lf+B4Ab6ES2NG5jeu6Fi/57Jrecs/EAcr88k
vwvYPl07sAF+W9w97Y5wWKVZifoMimxClw0fDde08Us3+kQfhU6E9/fRMb08FIEb
lojYeX3Q6JAVXit46s+spiUNQEUWqhNY0j1zcf3hILCxP1iwY23x1Zu1/+L3Gy6G
FfTy/SyjGG9VuHc0OU7nNbczoDYuGlZ903b6uKP4qpySuKeHUP0ex4bzoqbuaHd2
3VkVxXV84hpQQZmRrmR85M75NMCZE2jgkNSg/4c1Pni0oO0oKbkj0MiUhZfLLfZI
gsbX9p6ebwyewtU/y8vhIsangMODuTm9hv5hC8wsekIP5hY13TMeXkQ8cK0AEGay
wF0dCoUELeUB0gaHdak5rieGutDappO6O0Gr4zVNDxNZ8vjEvKIkkNzi4eFzUDit
ZRBe7xxspmCoy3W9WbaCaN0en7Na6nHw9eZ/S+gtWQB8LO6na88E8zY91440TA3R
iMUiab3k14wXGTLhlcpZ8YM78wQpRMK4gxbWf9MV2E91Qj/ui/+w39bT6+gu2mpR
FeYlUW9wF6KizOCBfE1NtRPn4+ekx3115QQtzb0nmwpva/u8RKHceD9IiWBgGhYE
WSqpKfR/dR9QrleUEJDyHLOEzTpcITSa5d3lWH/rz5TA/BMAY55rb7WY33LxepYC
xf8W0nNZnMRrNEgns+HBDbo0L++DZYa24LR4fITLKTlQpjqjOsnzMK1HOn2I4QBK
0suuFI6zIiRn/kRjgXjrgdzqfRfkC5IaVdA2O7OZpdtH+PY5wSmcFFH/bbsRYM2K
QE7I4Cm0WTf9b5oWBEbIpN6kGjqY/pvq+SDXB3qr+/2y0HBYinp0sld87Np5ve7g
zZnorfZ+RYf8a5dstKhhbXhtexvNKjJxvMSYDgvFS6f817EdvgC4y9mRzzq8DIp7
BTfqE4sQJgP4NcCTBaoaP79Yj2TQRNVuMnuHHim+uKIABGhrQZHoJZir0o+Kscf9
rdBeDPYu25xfjp7bCE+2oRCbOiwWB3i79dn/J1B1h/O9X2Egc3/UFjVh8YLVMGvz
2Ku31RuRVmNHNYlKA5hKYKZ4zthYEZR+kXVSseWYAXNkffPkagwvL0JtvjfTX5JB
twcCOG8F2U2FI0rahLjP+19FN0DbTbX+N6Ggf5cw/9uvK/4nQLRP43SOO4fJtzOQ
Gt2ISR7wnT7Y1Rkeo3jeWXQ2PaOBDO+hVOyWKo6kkckq++3oCQ3YCASMeQzlyZc4
2vKaakX9FR7E/2xQ7eqgvnOCO1X3twaTqVJuezcIUAZnTY5RgJ2wwGY+qVpFsCAB
9Y4SwRCGdU6vlxLJTQYSmbyVXLWyX9G7jGq6rAgXLQyQvCosZ3S67UQX/OMm65Ny
HXFIonLRKyYAPnXKxoundSwYCjpnSdVnXpkL0MIZDNTqiSjIMpR1FLH0BraWAGkP
T0KWQ2i2crEnVGisWeSsbxFbr0IlrsA1ngTjNNCESIp8N7JghO2mgDo8x+KF5wIa
5R+EphIYTXE6bbmKdPlD5IUwGDXyLdprr4I8iU8xi/LTwShxxQQaNokdMd0Aj+4I
2wVcG65/jVLCyIM7u6OJLLFWZ05vjwMF5aLVqJUys7PWvV8sj62ldQ8Gv/oRBDb4
tk90t1E4lzasDOTcWhMTYxx/Ip6dNwI2j+TsiP5/uPE2964lsEnN31WC/hQNY34B
Y5DL1PROYgpRrl3x3KT3n8KxSQhkK5E+zI0qu4Gkl0sckbOAbUj3D52RFRxhyZSm
COI7SdK/vl6iKkuXUZ4OZeg3a/F06jcVXXw8pvFoZZfpszhacTww7shnm87UNWC6
61MLLeOenucifMIPd9u13/ymkZ8CYmn8VTLsH5gfAg+NuRrVdcx6sqxPvXHThAip
/GgoOGWPlh2BBdOfFZX8PpX3Dl5OCVO6RU6bOjBZAOpM/S9GvGZMJ61JUTe9wAb7
ufwmFm/Mz/hs00/qOOlUW1GJ3OJ/GBFPRkoPCZyowFQ4u2CkBjeRlXsyikJQFFLg
ROfE4uNzUfRkDN8U03G8OK74EN4+OM508OZrCBE4n8QsSfl6pffnWezm6JVdtr3f
P2diOrN6umApS5PBsLJgOcXHK5mLtO60CiOzgjCfdlvtBT3p8IRWnuRwri5RvEjm
4pY71g5+GGtl/nLEfEEe6O48wwn2qhk5XvPwt0Ix+vd2yty7P20CxgGYnyci4Prq
q4qqyhcxyao3/L0UBYtQeXj7kIUt7+ORf/o5WSh4lGdrRv8+wB99JP7+vUEx+AOf
xH/UP9L/RmXc3jhSvxo7KMUXKpQjdQI/H2lmt09eCaTbH2DCeH4LRPSVlFYQajHl
BqOwz1tzr5C9feGEW1VWB1bWVAtvecI2BVUKiOiSBFc9O0oAmcZNdWcVWzw8xrD/
h7pwVH9OaOwQ1ev4ruS/E04bmL/O6T+fj6FlWYceRiQa5dZfwnCCCXd0YrZ1REUF
xQaWe1evwApbP54xDE00o6EPctFyQyAZDQAG4aFh5dwlHYigWft3m3jyJQWwhqsg
lu1ke0T7JJIgAj2VFl6JI3HEIpIFt4ZzfzMZIGdUMmU8Bk0vI1Xli2JtDW/Ml8u9
STfhoJIUVogvxm+llmn62m5lKE4b2LRqiJs20C/zYTXlWrPyqbJDKH25kTnODHuA
oW3JjJ3SR8FE4Cm0cyRbeQx8aalm5Nr5zxA4E3BLNRXXOcsjXk0WCvumhFlVzZt9
G79VD3Uy9LMC1085LHpOuI2OAgqDPTkCnCknX9Gc0dkVGY0EkO+kazHT8BWDVOId
2C0cD1OT/QWipiPTKiGm3+rw62xw3h2Af8eWaenmD3gz5A0bNTBALHRWOwjxMuk5
`protect end_protected
