��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����S�M�hkF��1~� Ά�``0Hɿ��b��i�<�1�SzFĐ�48��ch�iIQ���H����:4(c��_V����&��}�w9B
��T#�_qx35t���D��<��R*�E����nK�N���������19N3a7K�0~��!�@ըfG#�=V�[��&@0Xy8�U�N�
�y��I�S���j�kU�,���87��u�:]q�Ƒgh��8�i;�f��ܐWq�Re�R^Y�˒�
�1h��{�%z��1(Q�,1:k��S�pv�p�$�듮Z�����C;�y�A֚��Au��*��1�-�_��e�(� $��d8T4���z"�������0����W���j�Eզ�$f\��W�t�(;�g���u��A�j(���g.��=�kz�7݅cִ10m�OɅ��1YW��F�O�`�,�w#{�iR�{���X%>�w�?U4�re�C�E��C&�i��r0��vf�8�ԫ�ft�cY!h�����Ϸ����q�ׇ��/j�"(@��c������mI�kru��)��2��*��0�r4�������i:3a����-�������g=���\6A9l�6ιB������:p��Y�Y�[*i�29��w_�\�&�h+!�)�v<�}�!&��V� !/��y17�&�ţ�*�Ҕ} �2]�H�,�nV���˻u%x��[�n^j^���XԞ:��
v�9Q�����3.O?����Խ��@��5�RlCN=ۛR�J�%���oP���'�̐Ӓ�J�嫃C�EIg,�	кOY�y�f�����{I��xBE��e�[��a����-���;_4 �R�y�D7f3�ݛ���N�v��{,��ı�2°K�ui��:K���5rp�FJ�Z �ca�v����Ӟ�onHa_D�ޜ>��SD̈́E�8��>n�X��Y8|���"�UҚ�sq��x/?l��$z~�v���*�|�cq����D�%�N�[������Lt۴�����}�k�b9��5rG��IxT��?*Ԝ�|�κ�V �P��%�����x�H�l����7k�;���� ���t&��N�[Y��䀹�'�d�
D�}�<I
��S/����|��zĸhEI�H/�s�~��WŔ&_�.a�%��H�h1 ��czi�h�&6h�{�#�뻢D@g�CXXXeІQ}u ���؀�Ǻ]�� K�N�����B�jŝ`� ���Y�>x(�*�ڕ���'�Zql���kF���ƜK�w����
 }�]¢�M'��;�FXpV"j
��w�k|o�I�F���Ŵ	FMn���w��>wG�m�/>vK3�n��]�ˣqA�s�N���#_�V���6�v�d/���58�G
 1���;��u\��<D�h.�Z�pm$�f���Z�݈D��?�e�:�Y4�v��z�a�$��D�r�2��(b#8S�v`3�T� �Z'��g.����EQ�;J���AK�|�%Ǳk� A
��گ�?i'.$Ɋ��荅�yH�#;J����`\Y�m�}�Q�1c%16*�l,Wӿ�h��ڬ�W��m��j�A�Bm�$6C≘١�q3�����L+����%��Of�\b�ZµA�I����e�.p���?z����c���ჩ�{ތ�X�"��O�n��|Q"3�T�K�w�G�+%�XP_�>c��ت�S�������|[6������чߏ��^�?�c������OD?d�uZ�5 �nNټ���X���1�"ͩ����B�7�1�ч���6/O^��Û	�e�ld����h�UZ� �!��{���CW�Y~>�t���FT7P>Ur_z��èE8_��9����V�п�Ob:1ߠ��
B�K�Y���G\�� ����C�p��@�P
+�!�o�fr�u��r*-M��������5�qQ��5�˅aL����Z��oBU���I���
#�����Is�}�N�T�L�.-����,�J'M��~V;�n��@���ա�#���G�o�V��[�$(��X�Ͼ<wDY[��V1dk���I�z�I���ezBEܳ���QgDP_�Ԝ[�~���閰1��EhWy�js�*�RS��1�ȹOdY��L5�����<0��k�=i�<�K�����{��y"l�E��є����;"�nO�P8���W��!��qK�oz?����p�E�_v3����Ad�{̼d��E���ȵ m4�%�jR|O>���s�GLti
���r��w?�Bx��>7�����DXIUTҢлD+Ͽ��K��'�e����V�8�|�h��x
��'���V�;�Ŋ�s�0�I�4`��&t�����	&��\K�R틗��B*�{r�"�Q��p�$�������'�ܨo�Tޜ�FOrqN��z��Si�%.D�1��v`����q��H�t��O��00��������C*����d|�����O�]ԕev�J(���m�5}`ȣ���!� P#_��	��iW�e�
X�m�,^/�'o�9
Z�/G�[�w|Y{*vqC-��ˈ�XPUэ^fO��!7 �B�..%�i�#e��0���H�孯!F�������X{O>@A����u��Ӈ��ٹ����:@�eClS�ȏ�DM��$Q����J��&�v���N�`z��9��D���:{n=zO��؂G_cm$��]�D�<#�M�B���qgX��9�:��"� �c�t���|�i ���).S��2�e����&���РeJ�|�IY!�n0]��=���,]"����qnnd�a�=�b��!5�ʵ�`)��$y����H�����;xl5΂��������N�.��Џ5���#���V�(�ʨȭ�}�Z3;s���tC��s���ʹ�K���{�;����U���w�Y���1}~):"�]S�KJ�)N�������q){����r�ն�p*&vf�r8c;��qx�FgT�ߋhWy������{��9���[��n- e�=I�c�&.?�`ʛd�
�B\�������9��+ I0!���We��&r�_�6�Fg|�K��ڙ�����]�z]���c�<�?�)/S��"L��ٳ��!��$�! (2fK$ }�a���G͢��}E���L7�>���n����.瓼�:1��4�����s����Xa<q��PΉ�ӫx��"oB+����kL��ڸ�M:�Ξ(���4�6;��	Т.��t�P���7�=��� ��ش���^���ђ�c�@V�i�Wo� H���=X�{���%-·�)�/)c5/�