-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Td/wyYIEtg+uJW8tW/GMFiKfvTjBDsyYIK5WDyoLrRzlAierln2ZxQgeApNdKRnG
f1v3w2+zqwUoJD9XZV1L32mAp/5/sTAheh4PvKgxJUdBLUCh6aowAe6Rck/FHcuG
yB93B1nBSnFaH7KBF5VUSkhkRCEFfBZ6VtQXaUjaEBM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 27746)

`protect DATA_BLOCK
2aD/tD8g2xa3HiZBL6YjBXKylMgrpCohkc8zkn3S6BlC4DMqhf464Isjz+l6SkyD
L85+ygKqOjtHMHfqYtlJ0k7C6E3Edla3ekeS8yTiHk3w8AFWeqeZsf9z6urrZMIO
ezltYm6DhLx+W8eJ2T5JWa7H7vd/b8MiQmsExugReGMHcnhYG4RzjHQ+7KD+7o+o
pnN908TfVwEKWzEE6fmjS8JxUTwRfRsdjufDXP9uOK08dpQvBHNGf8eZV8utVH4D
8SgzHMsco1khhmeSVuxzdlTQmyUJSCLoGs0RFe5SGtrWaPY5aZQbJxTwdUKezwic
YpN01VLKVD57zfv8NkqJUc7JDK4Ti6cO+1opBi85njaU4pEWbJHDRL5rrZKaMm0K
TP3t05yPZkmZKP3dXzaVWCwwp9G9ONAiIl1fxQO09zTtsjcGAPkpxTPMkgk5mw+o
1a/Fv6JHI4FcjGiSjyPsCzFFummtPM8awYPMNOA2gFemgzktDmqTyD0Q4A/djOdo
SCoERk8e4C+AfQTe/q0lBnOMcBkBBk3ik8qwWop2yDPKoghbnGwY4wVOnucJo5c/
03QPGnrm5ZHtTM9FwN02lNp6MAfltmWUNvmiKvuCRVzAe8OvxwZXf4xAW0EyKfiF
w66ja+j5U46b1zSzMKJIX508aIVvnHOykBt/IdXbnpQJ28Pk67pnEYVjlFFuT3xA
LlNnoIIp/jgPa3M2NZ3wFYuNGdT2m28uGTlxm4zr8pJcvLwKlvpQKCi1Ns1qfrwM
k8hEbD8omi7f5CQyk3QXJTnDVWGU6wYfSorVApKK0s+KpQ2xRv0hFsrZ3DckB3Vt
oBBTdv0CrqgkouZ9CfUgB7dqPNES0ZGv9A5g6z3T7NZgS133cBgJ1+Vs4Ggkw559
tMQO4zILYat1wS/G1bHSOnhLbfy7TO+p+Ps1sWLQpgA6ukEPNq2j9fLIdoe8Rg29
QxXQ5QAOP/DxlK3jhdWMiQ6yr3IIrbtaxdNgQ1DHmyOy7pKDm8gDDqQNnqMAgB/Y
52/d59B059xnPJJWWu2KRetrUSxPDZdGnRQXI2pyn+JoqqAWuaUQ18NJLIM1+PDv
+DFVJee3bB48LeK2mqbVGgWQurpyl27j4FeVrUQrCU+dEkzlHC331b2+5iqJABeW
1dXmkGzNOGwfhSgvq0qjFnCmbWLqBcJNCG25ECJ/d/xdQjP8Dfz1ISWcg0pd1TOq
4FwJAJPo0dCoBrau1tPZkXinlD9b58jvj+N2m7GtWKBe4kJZHQNSQrGqH7XQ1vDe
4v8GcF6oiXOMC2fKZ78xprrTrJ3hMYC+f6MbhvGxMQ+jYxWavvNBruEwOOjYEF7d
pJUvgMvZz+tjlGrPYyIVFWLqRzLiYQJHTa3Z/Ptnl5NckuDNV7qvnfTp+E36y5ub
TkeoLs513Ipr+kl6ldd/zbFLXp7jZpajNTrwebbIm/XSSm0vTFAKyAZgqlT/vwqf
HCbyKLm07GhFmnMFxCWu5iWHWU6G978d4XJ/PnMdegHiOG0KHYbE4a8rEjhKz35p
8LK6Q32jvgiXtaAdZco9w1DsGahbrU6hKsQ/Kh/oYznCWRUv4W9IVUwKnix03hIo
1y6EEF50wACEswSw0qL4LwYd+TIsVAKqRdk7rl43HW/9crRDHLPNUczwGKJAy4Ee
amR9dk/mzN6It3kihLikE8m6zbB4Vh7dj090pb76J1AfjrgdPxoavosyawiCWXbv
+U4MAjNr0xZwoVkPy37Jt6hcXVs2odaHaTZS+qb0UtvQTkKi6AacEAkniU7Z/HMo
xQY/ETfO9pFyOnp3Mo1XDt8BdAMTtcix6xlLjvukZWYlGUEIo7Ltt0so44DV6cuY
cfgozkBkl1NUS7UxqOVNJEipE+HlEtGcc99ogCsqfiAXfBSd42tltjtQ0kgxDTiD
AGvL2aWeUtqgCqcsxQs3HB0qyDzNyujk7Rk8yWK6YMM6Z0Qm8XjMWo2lvreBemdp
c64CB+bnteGL9OD29ftmtbGkHakjymu6V32oPvItqv8nJGQLAia3l7L3ZG8aqCz+
Iu8+9oSeWLoXDRzFRyJNxwrtjJEV2KxRnDP6/RVBB5C/KuqZhNY2wOJ3jzLyGLYd
ON+5vLwwykKhyUv996eF4cP/rso36WNVRpkbw9DiQ3Xuu+qxDsu7mhkkU8XsmT9E
TLGPTf7CJ7zdNDErV/ux31ZcixRQU4kvNaxOdv3xMs4t3oFhUcHZOy9j3lgv2nGh
IgYVifwXA2+r09ThqpFuwh4c0lPBKPei3i3C3hjG9TTUguYz3qxhkPswAvGsuxMf
4LS4jJb4fcgLsMm94DwgWLMpvdaPpTO7r2+Sgd2Gn2t0K+n5jh36aE7twU9/yvg4
MEunNGEDwxvtfX0y90d1+wG5mkkBnCPqCBRd+ie+SP3mfpap27e9cyF0nnK6NXDw
JsjWSPiXa6VB1vcQPesFitSgUGdf3q+CAmaVhEP2epRwZ/b3ouxA8CkmOqaeiPo1
tqnpgCDx5ZLU4njeZA4tQO8Z/Gq99NsJ98Fy+SlgwLKHohK0e57/GEFpFR3sHSou
LOORRwg0oniiYT9Eo2DKERZs5nZ+6kdlFVJaIph+ieB43FYbx7broujLfAmaEizT
uDFeh1cPDFdqx3zlYA+vaotZIYAwxbrjs+ucnQRnw3rRaFcVl54aK6HKBs9np5DO
CYHvuX7CokRLuhgfVkJEz5RGWYZFsO08th1PC7mE5Z/SOVL9JhMpE4cZCciTKcek
wdlspcZxFRdnM57cR+oBZMK1pqur0bqlbL3QxWbRw92F/a7/Ce5DqwvvtkIOHptr
BuHqMeVhs2D8mbj4VLlrojWeZZ4o3PFc6HyDUZxKPPp7uzuZjcMCHzZpdaZGVX+/
pXLCSPeX9SQVi1op0/15bJiPfek6RSnS9MHsDPt+JoNL1aZXERtjQU0CmW1Oz/DK
gCVjuc7WL2gihbL7P4uxgt4dH6RewcT1Y1omUq/ME+0oOgg7V8dMcZ61tSYXN6EY
BUZbQRwgNr88kdRdcxmGzyLKe1AygFyo+DPMq76gc/DczC/h6JioTtCD1FRrIMWc
072Pw7h3/IMWqkQ8Gf8m5sGKfGE+GvOHjNlVfCPrHY2SdeKdn0cLysIX+3SXScsd
sTJS6tr1GMF5e8miO1S1bd7ZRI4fGd8rvK7adL3NdP+NsEWfLCh7YrsuVG6DP3vk
UZ9NX2bzyp+asV5tH1ORt/wl8lkgAiiA5nyTY6V8HuYg/wm6MtspHf9UloXq6tN+
xkDOLoUV21vRyE76LFasuzj+Ao8K9hI4sEHq4YA3+VkPd2l2L3i09zUjI2M8AL3l
WlKltnqTOpP8dFSKVlb6wC3LIl/evP1/VHd/MYEGOjcRX0JdgtLdNqRMnYBnx70C
NHt1Clyo2X23jS9DUGDsUj14zUjHsD/OCknc5RLHI/hu2R1gi+WyuFCdDz50zkkM
Ms1paDtNQtv55XeMsCxnSL50Dr916ACaaLe7D7N612WlZtT8gyI1IS7ry1sgRCaa
4Dh+3oIylA6dkGpZA6SIk7+lAfMgvTzzjXQA1Fy3tFgpJZTnFoJoFEk944wBrzF1
SU/BSHZuqFyuEq1Mj/NVdJ3D+JphxcjvfxxcSHi6q6Nm8Ss9tfLMdSeAfGkDcddy
BOmCEqB9Vf98ro8b6Ot0iTcPqNEy3qzIsGRO9as0zOhBzzbZuFozDT2sooPBavCw
A+E3ngO4mVLPOUbH4kW6VZVHgDu/zpFiaLcf+AdRjDitkEa3rjd1AsNbjLnIsbf4
8ypWEs6QWiP4q9CepVHGqnJ6yhbdKaMo96/HCBPWjDRhd9wED10Rnnjd5dLvJh9F
6iMEc3SgWLDfWSf2y+AH8o0Q3Kw9giwbOsxm3DN/FNrpNbe2bWLYcFum7h0DA8vG
U5uuj1HN+fIRRGXSg0uvqxrB3ut9MOseqol9J/CjdI9FqfisunT8t+kXWGBXT4KD
393vvB1O9MO76xsjj+X5YkoxBlSCqYYy7WDhJ8UmdfwSJwDj09CF6udHcpSyM5SE
ei6roRRmhjks+IFLivIal0EbxlUnw9QesSMV3pr1oGrCBolLhHH0kKY/visde25v
8yfcLEydlpffoun0RlWyBam6mRft/mEqbeS0UCu1JCXWrDUkwR8oM3vvD1VGyd2A
O2/K0mPhO7KtskoUJvFV/1pXvqBh4nmhKJQvKap9CfSXiAqv+wvwUaIfRcePnNSV
uEE/wjGBWcXoGOPBvUfI2v9tC8aNaMqKGBlYiUJNjpwoAp5aRZO3eqrZSE3zcjpV
KOOQerFBpGGLK1hupt7F/geNYsBOT72krY7bOZUAdZM8EkTaTUb9tY14T0wULjN7
FXDdgzlywqcbGYv31qWH0K8oSIBlpvlGBU0TyfBkxrVLS7Mcx0rK8ICr3MbAMXoA
Vwq8br/i+O8LA7UzIrysdFR/hGtxHmf4vbHyivxBh43QB8fc2XJaFsA+XxgkDw0R
CRPW8h7Pu0024byAZeCNHWftwGDIrjFtMXMHJJomJz3VhsfTqlDtsPB/aSPYXyOr
aARm3NgySbCMDwQ0isiE3O6YxEJQ3onamqt7BsVlz0EtejCScLa40lbaf/0tH+TD
HJVOmTg7toa9ZKL/v0Q0P0Nlwvw49/CmulGUTKl3fOhVqdNLHIXsYWplQFKd2UH1
yPLWVrviUAnlmpXAs3BMlmEhlPm8mLt86OcaJIXHnrwJu/4rRvko3H8xvZVp/PYC
u5sElznq0hI/Mrru3vtXonBE8pepm8UwwVjUnkYDFFlMt5m6xzaIXw36VqB88NkB
mRbRqmVOEfSpA20F9h0V3dwCeTLYP8QG1MZZrFKEewJpJhTasdpHzCeJIeOa7u8U
D0O9OqPmodDUa+hOzfiqM1qav7artbGzEKBYRG26u4ra8LscC+CtbRl7bcxgCfsV
2giZLClxxoXe5A4wYxdQSHlUHkQ7RxDnCTCc9loLTE5CvNY94WMbG4Hf9DvYd92y
m0ndLjxo2ZDptzkAAGdrNJNI1s2qo+p7dfoL9vg0DODcSHnHZM5aM/jw3ZlkAI1l
5CwV5fnX4GII2aCtsM0/CNH6nsOOSOtoL9JAOi4w83/2+RJ7HfKpuyTEWIfU6J/B
Z+rP7mBQRXjBMFMGWUMtB5Mws82w8nI4zlgXAjfCoSuUl8iKRq4s1Fs8EjYT+lVt
seoHQsQPIfIo1Skb9OY2t9mHhKzdtcXeMETfnSx5uhC1zykNmLutc7uz46SqhWUO
QQQt0M1sbZDq2IQKa8MbnNzBmXE34sEr4skEzS8Kd63GnscOpXED0itdt3KwJJRE
sx8T1kUkutj055LGORymNx/80vafRjfDPvwfZAgQCIHxO5QvWc9FeKCB3xJkuGfZ
Od+6ma+VnHUjCNFY414v86tYbHrfOaK8W6JduZ4RhmIhEKCQEkq87O699iNulc5H
AMKNlD0msVkQ/IQ2gdxWNi5doboF2SFxomUWRnHZEdA/BOOypjpHCY7Fdw8/6k+i
2u6i8AMt4RlPDhAvcy8d1GBXgHhkcSHcZSAUK/40DihvmbkS00MX3K8hB5A704FE
JMlLyDKnHBOKmR21L34F3+Km2xXyFdoybunUlVxU+F+RhTjOakW+UBNVK0wb+1Qx
yGG8c9wM28+ruPy0WK3WJFq87mTYY1BwPzWM7No8IJ6CZ8B17r8jy9PGPeOnZB+a
hXHsyhv7VCzC8tcUymqn9sd0Tcu6d4adpsOtBsLqXadXT063rfkJ/AjSaQDeOEHL
pt7XrF4fMkE4UYg7/vld0JMqSxHE76t9Pxl2A8bChKgLSf+SkyAwpB7pd0FdzKpJ
4wC9zg4CoJpNHrcooXlvvVVr527Dt7BV/FmVTMeEXGIOtEz/Zageoc2MTO2q0Qzf
wfHQkPm7sV4NY4MA4LYrzQ1/LJUSwanWZS+tlx0Y/YQ4aAaZlEphLGJSvHDqGNgV
obDMSsy3ZdSnLPEuyUQEZBSj751gXfd0iSaSANJkK+uTo3t3K/0kkNslh8VeIyUn
kzQMWJSWulwqu5RcE2uzHDMPXU1vKY6IPBHN3ezipZ9ZqnHDiD10G5VUHR2yxKzC
JLddeXNP7B9NpPKEd405JaXYm+HxHsIdsE0x4ub1He9WBujhTmGB6zDwB8kZqAeC
38VhW2lZsAKgDGoBM3MANfov0eihX9tCsd0QQh5ycEEUKt5oFdfAmnJ44YbkMzuG
yDLoeEV4Wp1Vevr3vOX8nnnifhbUUvGHPVGFrPyE4erAMkmOP4FaRxCRw7CJen9x
219xysKryucPY3VMxABHLeQya6qF3omCnIE0b450sJjDVsn7Qu+jJa6ijaO1gQQP
0NIf7TRWlxqR5vObJn7M0RihxKci1vWqY+HDRcmB+MvWaNOo9rop0Wg/vElNR5vd
Zq3917e1bd5ZlvKb6YvQ8iBX+l9AbDgq6/mfF/ZQa3sJq509jQhTHOjLgbJtwy8p
bcmb+u+7eImcFzylXnra4+Djgqc4xT08pkXxJBLFq2kStNSDXb0uJWrtf+AGUWx+
T2lBimBQDT8Moq6C5zBtNRz1yBYifVz3GLiz+VC/ExP47NBh1eYBsGNLJS4RodCF
rUk6gPRiIZmZAfWLZ5+PU7lRV3heuRA0lwAx6L1lVf1oZlSDEhEcEjZk4ydhrxsb
aSpGaeelHzMXQifNK9ARxtAsU3t07sNMNp1e7fBYD7LFTVE0MCjo70I+JxVIhO7q
DCN/U4Ml5mDWGSdyJYZc8rJ6uJ0+tYRZXywlI/9A4PTVf8Z1sv5S1LEJlwhs1TIO
uGAyRrE80U85RV3eWZ+SfMPOWF3EGpT/2qLIxygR+vtfTxDKcggjfS62l/yGDQzp
ZR+AkY0jWpGP9fH4YhGPuexZ/YycgAWjSJLjBfdVIQ/pHS2vmopmIiPZOibiymog
9GzwzI5DO5hQNj+n3pkjtp4s2USYda9UbciiYUQjVAGmt/T0q6BUjv+HLDFj62El
7ZiTID/xUjEqHgVljZi1hknFSDIRjybROGPlnyje/cwN80IwbEuUK5m1fC4SilHG
fZduyFUYHW1iKZw/rL35fBvYE2ddr301MNjY6L8fcqP0Uxwce9qR3z+dp2rXjbiG
xuk3Ct+SfVyMb8UZ3LYHj+SgVu1TP6+WD7aqn29zFajBX0PFOGrZC8ZDMblkJam7
Lvfy4lg4N/GdFCqFFLN9PAd88Nl2SlX1HgrJ4p5XdWThZWLYuyilFnNs3A6g5hHb
9BYnbK/r+9eVIXITRCdybtUJ/yi02HaLBh1qGsvIBfLAPDG4sfO2jfy84OKc1MBt
Fc0r0fvKAh6Ns3iXNDgeruLWYXHiDKxwYq9HgAVaKqP9IcRs1oZNQLuapFkf7ye5
SH5BvpR8MUp+66jzDJiW5xLEAtbqkycrLtDJPkDwXwHEqUFkbC8upF5qwp8airHG
kU5/aG5Nw6yEHHXOq36cPBswQHVZh8hBpl25e3FwEW8qy10V2j7ZdC9aekDSr2qk
uH27zs29fadfu1SOlkw1sK/SAwmEbyz+oM7r9B44XFE7FOgGbUh8CeNCXBwPavig
hnVaziQhelm837eed6zm84mvPWrKp1hnJUWBBqbnAwqecVxcwaOVC3xegSxkjbWb
y8nfPlf7sZ2e4SrHm2cXA7q5M/R/ePFz2WTH4jY6hEMwhEgQ8XmdHE0I04uTIUT0
pCrSjvpu3ggo/6a6kLSmsN24yCHJbd4vuog+NlFpADsKKx16hij4mMB4aw3SrTjv
ajmHndERiHbXyXhc144tWPLUJhjm3NxYs1RAWSjqXIIb2GZrqsXj8d9unbzq3jeR
La6CQtMKkGsCY7JXeM/VdgijynpQQUpiBMMpwFbz0lWwpdgXIhl5I6iWMqr/fggR
Wq5h1LJhmQpxUP/IWxjz/7CxEkbY1DbsFNeKtja4TXEDuCsa1UvOS9jACdnqF86C
jYy5IKNdmUnf3DLbyAB4lnuHUKGNWljFqTvDaLox+eBwiaS4mhysG+1Wc3N6cuhv
Q6F4+HvxrFf1by7dT4QnAHu02MOrfVBYsvt/eYpc3T8EWYoP//ZBDVHfvOAPcnIo
4jeWSGS1yquCniGIBpgTQStF5hEJijpj1LBwMeBkttaCaYKScJbt5KWrpwDjSciU
drl7Gk5fc1DNwS6OkkxiLOo6ts27ndt/gjzjjjZ8Efz16uBIxhaAluX2BtDwazwc
P/Rq84Izo8l14p0PLuJmOvx4Cy34zdMuSFDSMwAqx0Gx3pSWBfKHw8SypZ2wrrJl
nm3O+ACtnJyTkdUEX9Pb5Ia7gINUxTDcH6bfIgih4UdUGYeEq20UDAyh7/76N3s7
JoqfK46dgl17YCx3E1+LEoCY75M6XgoJDtUIIV00opH91GtM0MUfHfEcuRHCSDAz
1fXiMLZbxDz2LtLk32hfhY837NeQirog+XX4BkR3LfokHdwwq/RYAKYHg3O69c2p
iVLdh97/2ID6aNzJFe2Jldt+c24hbuMY8AXnSSyS+g9dL6tWzbgMxfC5nuK7kypt
edBpz/MynOVqMDFvD+A4iAOZpyko9EAmlZ/2YOsihNdK0KUygC0hKiNlltTVkzMW
BUMG0ajxy84VbBE+cheSoIviU9PRLl7N5gL/iEYF+/lew6Bs6MpOalHXJojxDhkO
ebBkYLYhG5fe5X3WdAl11+hSkJwq4tEFDlbLnNRnbl0i063jnHD/ogZT71V4MyIq
WQ/V6jhXW1IuxGyZ2EO47rEUDssjgEbLy9K+QemwNwJbmgRxAAeXNvnOIV1PKnQh
41iI0UjqeGCxUArUcKVACbmZGpCvcOkXJpgqba92wKswkKk98XgTe5YyQwqr94IY
RHaCncSW+Hml/SG7jj3aJJHVDQ+aY23FxyFDAdxYkHmkg2ccbcic2gWSjalZ2eqt
EaggRA1pUV9rmwSja5FKFUVrUBDrVXhNQmyib2TtmThNS4xcu55TMf0ho23e8Pf9
G09iBIDYMNOqAx93bFu9Osb9t8EzDwZ198p/5cqZ9g+PABs/9052rNSyhFWpD8Ng
oeg/FqHdYTHPyk3fu9sjZNDNTGoiiuhB+gLg4EdGp1lTkJH/7KVH7gcz/C+u/K8K
5RzYNK+VUG4VXufiCc3gJfmgpMpiSjzyDR76BT8pgdcle2LK0/h967akVX6WdRqJ
oAGuTX3I95EvYgohqsBLKHpNX5OQ9GVy9OkWXbdbjdrGOp9GlNdGx/dhxjoLayn0
IfQTF8Y4pRbQo7oE3fZhqnps7RlEJT+wGmSwkxku0bP7VN11/N0cqFE03tzqEjTW
x9QkQ2z8VArlrWzwv5krTGFZmticaYnshdJ5QGAdNTdAmVUmBITMiIFhkFcGGE7/
hynkI4FzcNqeFkM//orF8eyV64W5vqDJ4xRg9zCiRkBHEd/m2sOfLLaP5WP8fhdE
jiUKHkKaZzZIRsMX2Ha9BU3d2uWiX3KVUrtKSlk+QZ/+ULP9kK5X3rtT5e2lwBcP
9yMgx4wGDhhdihdQAQzy89hpcJx/iRc0xj7HV91je5FjttbpidydwjJ33DgFMJO8
Y8X6k/O/uqPCnERUWiTgE/vgxQQ2ryeW0NemhfUaTcUnHUV2XZPTHO+7zG7L0tQR
3/tpIQZuOlmgK2OV7D5ukJJvO8ZMmDCOY0T7K7DPOer0xe4JUu6ZEHtzX2i39X2I
495QvhkPTlsr4tFNTbKomPSiAsnZiuDKv47TMD2E+jxV7uDF/tVAou/5YwsXtKLq
XxlGJf8xEyvRpTWvHnPTweB3bUfTFDnPjJ/LCOoDD7dFynkXd6OIu6Evzp3DmHJ1
8ylTFkMVZbZXuiWM/sb2pFhJFbRWvj2WSCikSn35tP6JXylVF70NE1IjRI5CwpNC
LjIXevwbxR2AKd2KZEPw4S5bimydqvuTSV2wxSTjmnI7k+coTHnNgybWHaDXYBEI
+DIvZPVlA7bkkW5aFPxtoqPOuf6swnBP7UCDfDu6mWhdWtyUIvd/1ZNpTOQcNTug
+FBFzRv6luUhpB219PA2/NPzntapQt8Evdb1A+yOvLvuOWKAmJWi9TkymKPvJG9x
VpJT5BSLxm/VegZC2/wf6iaDbUjZHSZTlanRnUyunCngG8wz66XbIuv1RNJoFUgf
IPOc5TP0hRTHHjw8NkUC0lY5NGYq6QIZ0ne2yuejBZAlHCxhHnegPAFwPwinOsyw
SDgQeRBW0B/StHvrEFxBbq4gQKh6GFJPQ5HgsGqnnVAlb9rPr8UP6/MTmnvN9xbm
hKvt81sSIpF3Xkp04gCoMNXzpCZKFaM/f1+j7DJ6SQVC95LpHBfDccXpkmK8h2sz
9QrCg2S/qBERXdM1jVlTMLXa729iPLxfeSGjHDWrC5Ujb2YPWysUK/kZ1PMiBuKe
Ym6P8mf3QgiLm3ibSCcjAot71dC1TlfvQP6Q+fNDIUUk+1C1PVKYhrodWu5kykkM
U54nzuToQDpoHL5oMUpXOnqBGwLRW95+DLjkTCPQ7wWqbAvpkMgEtIGUxwYDmzjs
DCsTHYE2+2xdJH5USVdzQcZWxzHtLJxaIPC8WxvT3bBNi6X1nmppVQRA+Gsrs60h
ArEyDAJA47hwYN6TR4W7eDoVganjicXhA53KArlkSiZjzIiDqqTECdfeFbHAPrG/
J3D26h/cWIL+3bPyEg2vsnQQ8mybxcWeElOYteAYwgVJTiD7xGaWxxApNekzEoBc
VVEgoxfGvLv5hTnrsGWeqp7Q1A1v71+e98a7B2afZURWiQZogZW/oTEJiRa6AMTv
HxEy22RvRUyKLd/Hr4mHv+l3hb0kXo9iUL+PPX8FXV2UQiaSjDCCQMYEap+covnx
yIQEwJuceFukoQdlNjd7nNdc8J3RJIQerZT5CCdLqyHRxmhMFLo9XD5AGi+BCPGe
IbQ/m9NWSdL4+TgNnxinOFZPRWrUQjol1DNAbO0srx3P5dzPyn9TgdB9Mah7f2q9
3vaA/A/qVjNNytai8zyjTXJDi1NtI9LHC0pZlmw5L+dkDmOHFxTCqIkT09yAHbuE
sbvTf9941iz6IdiZbgWggp2o+Fn4MvM+hdvm6FSjDo4zFceOUJCBzweuTHgSLQqI
a7zMe/Bsb+bC8XHM7kyCMm18cd+8zjP84bL6ZK5unbg6vZC7uqnX+Ed7vMgpxTyR
VJhZ/LXgzkseotYiC+cO3ZmElPHi7PrPule/I4fANMvaSYNJ98HCPFJ1bIEI5z7i
yB2Oe+i45d+3jX8geyx+3vl0CPK4MLmGrgBU+EQ7D3m5qIp3g/24tuGKwuAid9xz
DPoHxVgQM78wqiw8mT7H4C0hafXTFp/8nAJBYJC68se5Ar59vMIXvs939EfMrsSD
O/UO2z/dLK3Xp5j/zTn9AdDdpnBdOWfByZm06sy2hxhfgAQpbtboMRYy2fRgLdoy
GM5r5fBBgV1wFwj68zrUVmNbpDspJDkpPyftoV2bYo5H99LXGpM7Ylu9SlMFfn6b
ZqiJEPEn00HQYGjGTIKqWPkOS4y5R6oW0QnmVrfjXURQd9j4kjPH9/WPb9R6InSc
QA2f5symoUe+pzdfpndjQqCZBxdNaKj89y0ogIojL4wMeWXhRiWlJw+VBcYMYlnr
B8Cej+b84YlNjTwhwKPG6L/qcH1oA8PjSVin6X9OkoM/tVRi1AefQhCb7dyMHcag
qhCcS9bW1SSKOG1I7EmPwVnP9F53ACJ3rthZy+aXVmX5TeUAKzTmAe/QU1O5olHE
Tlc0u2cF4ap5w8dlLek4wTWw0t272y6NdYOjyunJyJ2Lm9a/Yz+q8YkYAxSW6SQ+
8R2EB285AuPRGO89gIWg7BG3lcDcCFqZGu6ivRT2Fa2LXlobzScwnIbvEZ/BI2IP
ShPgUvggwxPV0adz06x4NCr5mQUCroCQgv2tNRLZV61P6pdyOkUQaurQxKgEjAQ5
Ro7n5xuFzB/rywwvQpv4iz7jL5hnDrXiPks/Gxpl93IPvYSsHtXJIPvdXY9u6Uip
QjY3KVTYef9CIWc8QvS6cpDzQRbbThLNVVK5+QeRDCLH9iAeRzEG+ujykFkorZFm
GvYzSqONGo+FPYjRJ89Dk/FhkbK+0OuDwWkdBBKe5lY3NzwwNvvUMi7WKlJArBCd
SrVz2x74PDeIklDDwgCOwV+l+3/KyxbK9SIHFDNaKaoWJORPX/QapzM7GzMY60+G
NvjiMi9bCvhIC+z+9oug6nYSs5PxvgzTLkTWgps+7TfZoFt5DQL681CD+fLsivxp
BZ9jQTtdrGgTzzVhuUjF+OGZar3/49e6VX6u9aCh4C0IPg7O3qVSgs0QOOgPYb6a
3DKK+u8TU+eDm3FmsbUY/WU5Pf7KZppmt5p9+sVevvWgNK5i1B5SHcS6HnTm+6Rr
YDwtBJAN4JipU//yNrqqwGqtlZOMpcyDnK4zTKKpMZG+DRFbJ61+uinj09cAZPEx
G1JyvAMTGyi7H4olJYwh6P9bv/YLycbC3do5nzDtTFsdxCnHpO1uAPZgVILXHiGA
+OhvBNQ//zM341TFF+xuzQ9+L+eY1D0uU+CauBcX3muqzoLpUtjUoxx6+m8F4eve
FeIjQiAvSK9Twyn8TneayPEARFcqO5CLfvyVxUcNjYsCbFnHjaeTO2Jk5C6iwXm5
YMGb9W233yBJqsqGUSVixyVxHK3h98fjCgDMg9Olc5pgNeo61V84I60LDO+at59E
GL3OqMs3OU+Gc8RSyYSpbkIbq12YsSlrXC+p0lzfZYrZYS3nUSIHtA2iFldKdZPi
HH6dMTEUhINs0gtfs8s+61P8amhdyUwRGOuqQHGZyILgaWIxmt5DyXRCExEKUg1p
vjwsumZfnDi65+LhBculJbNqgFKdoDAHilI02DXN4kDb0FQAVyRITQq0qDj7Kt4p
bGz/uR6SzFgBBm/ZHvfbDHUTOrg/5P2XTOv+uBzWEJVaGINwsvOqzJkDuRees1jg
zXTMVeEwfHwwpA7W4Hvzv0wo45dY/H7W6qBuxQYf4nTGYfRbf573NfXDANiNse8Z
mULnO0mIuMYX9QzO9p70z1qG0vpbegWJgvBfbnkuVwaCS4lGJOTLxKdIKkRjdxeP
SAtu1kPIdKO27wZ5Oxna7qWIW21R9Syb/3c/cpNharSg3mMtL8MYQKzuR1pAXpaP
R2Rd0TC2vBGWvfCRecmmx2mnNIo4DxVnkixpkw4hfZUnqQVwXHNU4Rf1du1BsBY2
+TVQeTFmu1UJVhfW6hccQGKLOTU8cAJ7Sr3vj265O6FyL0RcPqsgkHi2kgO0uMLB
/G6SqkUzGg+5iXnrgNoVClXegDu4gg7PYPJRM3ttoPxJA0zhtmGVIwcwPNOGck/N
twCc4izu/8tFQ6EvButNqKt8J2d0hzQZJcFRs7R20UK6gMHTGdJbRJAyGBaYfVcB
cy/VVGPsC825C14E/kvx1d5aCxBreLYYzgC1BuoSL2bJv0uhRhunQSz1hN7n6MCp
zzyObBymCyP68abrppH3oBXzRE99LPGlL/S4aEnbfKaPeHCE4GX766ajkjyZAmC0
DAHNgZsEBKMX60C6TMW/KLgFZneG3p08NezIJv1DgtaFxpJVv/N1M5KR/doKORlg
wpgA+sSIuqZXd+s1gONqbqReWHY+m19FLRwZa096OvDlTuOvFB8wTEOVPBuLVpze
fFC5HJmdeeGPPIMIhxk5ZDvnkcNb7O5NXumWUX9rxP28U5eiQU+ahC71wvLKNbqs
kXzTp+44Z8+qQglTBDgkDatoxtHsXK6ZxyiSEOPxryNs805g67Abk85QMmp6ux6E
GhDrN5oLFzkDhoS4BZDOBD8suKAwe1Grp4oPd4+k/aU3J7rhJrt/taOYghv3imX/
B8ApxFkkm+2eMSdTIOfsRWyoQ55LW/0dQnvdtw/ZZmqusETJx/txJWFKZ6BsQ1dc
jAd5dh6A8MCDn2yuhuoggJPk0DfvKRAWHGk2vze5Bt7BZ9XxPSXdnax9+7KehFxf
MO7h3H9O7+H1j0FtSGIp27Sw3DHN+57Dkk1SQXh+DLdWGIokIhX++iglAdqvuMg+
BxDnTCyitKyh3SI35ll+1Y0SriC/WSv8eTita3Kw3k2LpREmCDJfTMsEEbhaodgs
LcgKUWdqHesohH/RoUwlLL9CibJFQnDogM/mPfQfjcA4oGZ3Iy6ReRDUKqzXv2Jb
s67i3l4sqQSMtYMVlEHrY1lhS9vLTpPeq+OsclW9KJoBSeu2F6MK6AXqbf2Y5eii
VjHXXloLsgtLyTsFN6c5rjAj+pfem+DUvKZmP3cLD7xnqn84B7XDeym9o+7x/zG/
Lggt5hiXoU6Dvbpqad/yNTCeQubXAQdHJDcSAuYogweVDR1n7M5c8w8mtsLBlqHK
YkcK90N2O1PmzsMV+vRoG8A2byvDfiB0vP0K+v7f3j9a6y6F53xUbNPbMAJKF9A4
MzyMEcEMOw3j/Bqj6ZpG6NtAKXrW+oIiDg3ZcjKLIQh8BxtEOuKyUNyB1cs/Cfos
WHNz1Ggh64dG/1XjwE3XXsLpaXW4OuvvZInVQNEVsr65OxuHH5qeysY6hTbRVCF5
ugZArfvowHCCOcGa9zt3LRQY5AvmaVFJ3xD9D0WYLyFLMVDTgEKuj4y7GJw2D96S
iKRYy2u32eBLIoTld6Z0RfpQQi+4c8fp5hGhTFD2zIrXKQLukk8xBbiIZbaypii3
JmSMQZJqMKERvRPth6bqPSXUYwwucNM9Ja/846SGgHjijU30ERagbU4o0sFmDprN
RUmyFr1Zm1fVLl5I2RR0EnerMN7Krv6qCLM0KIdTYvkpRij7+wpERdPNeiYQ5C/9
2EStqqbIgZInito2wEj/wbSqwu78TiUwqCFBCaCA7PcFoKlZAjkgeeVX3Ow+D96u
OxWeuu7g1Dzz5qUxJh2GBvgIUaEBgvJOCAAVAXpIbE9K4h1RGoMXDkh7IJszGbXj
7ZaKd2vJSLtV6kEUm3FCavpq/HWzGQ7ZsdGzFRRmE10188+UHPPupBNFhotw5Quf
a4SzYT/akroUyjGTB0YzfivaG/n42yjz5hAw1rmTB/mnaiithovKgLO9zPvUzRgx
P9MTNxloLbWJBkdFO9XcRgUiyCEkImcA4X3fgn769uX7ZNuR+HJLp5hEzTuKWDcc
tqPu3tFyvKeyThTcJeuvfxUvHlPuk7zGe3WMC8XhZrK9G4z9az0BnayemnaAIzcV
RtgZLL0ztk1yu6PoHQrMxHV24U+UR89USiuexCzS5rhlBDU4o6jegTwTE2J33dOn
y4EFDCu/H2MaDLuPBEgMxWSNHuqpo4K8GmQ0Pb62UBPx7+ZgCfgvI6U1i2I3XBYS
S0c7Bkxr5G6VKFos9GzqJfNVGg85g3kfyxeYVC5Ob0pHvJEGduW+vvVmxiDXCtry
n5allBfkUjMffJdtECJCFj91N/0ssTpxTFHKVkUsB1xmUhOfyfnUJc8GZuxGVi64
hRs5THsdwkDJdLwfJ7Ooejkn+exzYW12K2SgUK9w/8Pkh+n03MuDlrXrJFBoqAFq
c16UU6FBkP1cjUQlfhS0eTtkXlHDU+dCwVXyHsWfaewqnqzLHSoTFUePp6/3zRT8
VPGxieuwnpJw7G5bm6SF88WyDzWKqeWkyJpw5PhPlcIMYnzy3iuCwlEfFhhUk94s
uF4azhth74h8Md5EBye8PD1Mt4pEOG+ub7vaoxb6PEM0+hM2fpMh74+zB5Hd2mAS
kltsysp2d5YlCvs4hr/NtBScNPAtPDV9hKPrJLrFFsLSO7EF56TSUbAW8nh6H2nE
ephSqwt0RR/RshbBh0QEcd3fKzo72guRzC/slWtfeShNZBrUvXqBoRgzALL0kzZZ
F8YvBSAZLC2CKKu4FQOPwNj3CJGq//N58lpGyVA/MdPrwpYBFbV11GnifjBu6M4T
gQCh9ywTItJfN8usuHTLZPwjdiub2UBaryZhI8T/ShCUOIDQZKCB+XbvE/GYA5Rd
dKemBf6/wRe+kU+BAzJ3z4dBJT+754TitYGf6oopOliQA5q+h6ien2PbHCHXbsbC
l+/lNFIgr3MBd5djHZmH1V6l6+HWC4Kziv+Jo0iIsyRguoyVLkEYvmg8lrvahB9u
CPY0LEgJPBUWzrJDFrqM/rzT1k1U4K+p7RoGWXiXO4OSuj8bYgvTE+9yLztW69T2
p1l8inm3/u2hG98NzH/FKaAPrQM1tuxEhgBqraswD5xud/ZjWC1hU3Xo9/fGvfbg
QsOIzGzdYwAfFY3kYq2LKjsZKSsVL6a98FpYlXKt6FtGAWO5t2oyftMBvynyNy8S
F5cr42G9w925Jg1Jy7jqyq5cSknFS+nZ9z97+feC5lvbAK5y3OYHzOi/GX233tlY
gn+LTodKREUwEMvGn8jEwGFPsda1AyQbv3JYuj4QMH2zfn3Ibw/+ShsD0Ahc1dzU
rIrcJqHFhNeeSX2S6p3YpHUOrmdYouZfeIfjKDhHmVS4LcUtp47PSGGYOnKIdiQJ
2krgNiG+0YuqtQXBteq9lWYHWpzZSlJaGXkIiJYmpFEdly57SZmcxzz7IOpbURVK
m+6KTfhCs6fES6FJ97Qpy/Ads5rlIRgPKkcQ9CzmC7HsEYTE0HohcFvRh43lq3RA
CpHqUshRGJikferoEcfwLDR1j2MZ73D9aql+/RUrc7j6G0e7NM6vJcTNAcv6uzwL
IxosoObCoIsym5nl6yXvXx6s92CI8E/ejnYiax1G4GVNOUo+vDQobJtE1yNiqT3T
ttbInS168UxBzBjmPg6Wqom/FpqLC+by7CyTPBZyrNCB1a3D9xAXEF3Qh4f3eiIM
U+fJ0s7CJvfMJy0y0FpCA1W9/jx2wGWHI6z79l5XnFC7ia6qbBogpXCveqLzT1S7
bR148idfxU7R0KMfxx73lSbr2XXCtb/Qq2z8ImB6IdgADWM2CxBpGRCwMruzZjz7
dRICtLcc4uhzrcZkFHlfbtfkYQK/pdubX+zNxjL1UBSCJFKncz7pQ9rbhekltITh
b+RsDKHAjzLJuOmDxUkmTXCmxuMBgtNjRqJ5wOzyBHe31Sd3HSkUYMOThtalMYN4
LVOKg3ZMHMoJR2tnYZCwXGTYXpAY2tNJwDQu2aEi0dcr+/DeMTLsj12ROMwcRIio
f2VNgfRKGx3paapwzslsThjmD4PhvDBX5TrGiGNP7Ma/+NLM//ws8m2sFhEUxysv
B4hNwQykhC3dtpE4N6+Uf0VJYnehTRJVij906IsCNXfFVITjtMn83eWEHY4AFJa3
gH6b1l9BTEpOdiwBuQ9prmeuKiLCYIqRvT9VU5UQdkzDBGe87zNs5GjEh4bEkv/B
xv/ywJsfAa5MqerJKplNFt8KqJQjwRV1xczKInhtIm4LW14PpO8UFktxuhW0FZiH
Wr2m+UqbKoXRHSjG53PbVCjmqOm7RyOdunX0/AiFXrGxbzMvImTLNKleMxPNZpd3
YQyVCZde8q7Ji6jyrSnpxnBnO9IHL26QKukNenHH3GScc10wC+0tXaZgzCAXhMgd
RfSAkv6T07ig9A1llTh+MPlsnytNeZJ4VLr/kXCQeEAmZfZ9ifKJvO0ik5dBg9DR
+BDsIfG9em3UmoWbiBxvktOVw4aa918L6sWXqA14rrzzxa0FJh6150M99yTsFFj1
gvaB9r/Wk9AT+mAGqXfYjOUHgsEpOWSTKvGutx5aOac8s40qnezorQsL7fo8lZfZ
mmzE16h4hvyCACBfgjaMTrCsTiBrPdkcsNWwMJh4aUkgvOPGXdS1kc8OqFt9F/R/
q0arN32EAC7gzGfl13yPRS5jrB9iEs4LC3N6uWQ3rZ6URwmtEM/LRAKSGzhIxzwY
Y3IhjyYC8Lrz8ZggCz3kYuZkCMZCzAYVrvL77CnkQg97SIMR81FYRTlgxDKlmzQk
RwgunnErLghdoIRT72ZUiK+HfDNUOAL0yThuj1ImnrVsYUD00pDg+rpsxyPJsMDG
CRG2VBeh32ihHf85s1aBqcJ0a8ms/6ojbRpeqFqngsJk+SLdSw9t2qgtAPLgQaAZ
IYC/8YLyv+y90wSSov4m5/sNNb48h0Z3qL8uzULqRfXPSvxzgOabMui3VqpW1wzG
GoBXpPAkqb7zri61mAQS1+KLziQ4j2P07iuKJ2iS1eZBFs20gORaXqW2rt5iwFN4
62nm7iVUmuoUqW9A6ymFH5ATQfm/vTuoGvND9xyDw68eVyDV6kFXGhNZcNWQOc1U
j0qcHwNst44cjBzFkqzOKCySZdz11i/Z/HYS7+duVxJpGLnt8ndr1TUEPyk1Lp2s
z2s44JDeUCVP+BwUMsp1/oz+LY2g9NWzojGJx9anR9kYTNmF6ECAmOTxf2/FSdtI
ouB1cO4ylQEEyTU4TN+I2WfneNjAS2tyeXUyyAtPkG6ZvfeMFifHOZdUMKJbhLJo
4JePdE2hzmbJSk0EgSpcC0iVBHyjfPhi9TVgHRKNsd9jY2umzDUlaOmBe49EnLbv
fo4mH1bo+DKHYZxYSp/xNT3t+vZOZwF9xLTw21ukLDqJzr0Zqs1AtAX4XhpzxMHP
bJ1pryvspMqYehOoZwiviiaT8PagmKsUFk7eCNCui9yCpYpde452uQP9GwwKVxnp
lsTcU9+qBmNv63xqmrJt/TGAv+6pfEYsQPHfuE5XclaWjYOFj5ke0dhjmbtO6xBE
fh/i9wmEIvoyTRI7WmkTG/pjQnrmMWITUjFPUd6ndrPINa7rN7w01F3udbgNsxWB
lsQMGso9LY8ASHjES9v/S6URgELHbzNblaT4SEgH1WtKv5TQABp4E8ymzQhjalUM
uoNTR5a///UCDYlZr9QN6dWglKsRlPrIZ4MLyHQSupbSWCVgdz5+lLS09xPrg88Q
iACC1ePImNZRggfs1XXQh4IWDCqeJHc5xzIu2hYxJAbZcXgipGYw6B+YvR3dWW2F
jGEMxrox9I2IHlKiMke8qReLtutsAjdMtb6VioWCWbNLpCzOPRmgMs4V688P0hJP
UXldfdSL13a1+hJsk5tDBGdS13Sxf8SVX6kJHt5eF09jIdvlgXlAe02K4Nhhb0I+
Zpr4ClA5CKHGHFkxhLl/369XWEC5f2G884sNy9aiVFXrJ8705IU3+20S0AWIue/8
CjqpcP5hhy3M6R7U1l56T2tg2z883+c82GvH93fOzYA2IWYLPWDIOYAp3nb3MPnq
W79iTaO3zt4YdnJMwrEnxknIXhn80OXBMu7Ulgd1Iq+ieNz4d4d/HaISUtjUdZ6t
bi4UzNZk+7zWwsZr7RYm39y6zND82qrydSDq3O21HSm71ZNc650GqfhMY1HQ0n3K
+MmZhCzKbuQvNGAT/6a7Uy4djLKkxPaW4HPTnVP8ysx/iXVpi9Q5pIdUQYvpmak7
RsGrblmAsg2MJzORGfsB0eKIaaQ12xzWZqrlYSkYv//9ovz/nPGnWdmSjMIlGTS3
Mwm5NwZ6HQm8A4ErKUZmonZxJB3K2VFRCQZ5ki6dotodYOkmIi5nHOQ+gdElorSx
x5znIwIk9E3ganmSN8OWA2yQitTFtTQD6AVQxNxf2fdrcmVDpKsexEQcjb0pTIeo
7/o+j1uq5v3TykY4MNuopj6dwSkku6wlfx5UrIrYFegrT+csKq59UScgxRj7jlxE
4ShA/4JgbfSNJXHLSO7KLZyzgXvO3jhEtdXKcEIilpCTWtATqAtD9EO6LXrt3gU8
oM6uSgDBKCabGtEF60uqz11vxolvF/GjhJDyw8q/9aBNbwaG2ZwQ+6fFZH620laI
HQvlE+lVoPEE6YBqP/mia3fitpu7cVlb9oa9NEdFOwsOfNV2xGBHTLQ3HINRSgv+
+7Mu34fAl46/k8dJrJB7pWKfP7STc+cQ8OD8TX8l9zQcke+upBCDBSEu7W3c8RRJ
iCZu2jCl3PVuUGDI2zSet6W6a7bFjEACbpRe68t1GLyHV35H2jtkAg4JBTkQn9Wa
nkZuzCKGI3bVqfSRp5GnIjvetG2iiy2mr7mRZvy2NRjcsYu+IHKfG4pGb/OntC6c
Avb3G5qvy1GsU7d5RGlfSw/Wb3ZsPhCgqbUjC47Iogp1WJSEqLMOqE0CuPl7NOYY
BRLN0twZoGrnLW7jHguayQmVjr+lmI0brKfitD59JbSMYOokbk7cHvyE9cSZUx7G
vct+xjjo/iJVK/lcXYA0jOWpfGGiKosu4yLtypDKtZMY8U2jExEdPvbB8DZn6Yyl
2ANpOQLneTw+NT88xipmsWTeDucJPpiTOEkw3CLHxN+jlqKQy8BBL1vgeUWqPc9t
jxtWn4hkNStPAzq/pbAszAE7g7OdukTaqLRrRc4lZ7wmwOrKlWku286WGD1zyPyn
C6ejAoiCj1U4Eb3WeAKp+JTYEVINDupb/lx/zBSWgY8szJHFsCiIRBqn7y1cEBuZ
ID8MgyOZokpQlIXDlKU8mtoOJEuj0WD2eGgWoce5j2A9S2XSQSwPLaVrGNw2fXLj
YCPP/NE5IRVZTdzlN5KnYkDcJ4GubT67NQ+17cxyv5tpttKZBeF2On0oYLirOKTt
Z5b42FUX2kVvFYsjo25KlWDIcJ6V9wQkJnIBsV94uDmBvw0UXnJ8MDOolbCKX2xG
LeczArvCb+OanUBo/y4Bk9Hu41fuyViOwtkQDzmEkbd2KILvPGPZpu4hQBOo1gl/
LWM9XPKY08A5PgpRPOkJS+z0h14emOMj6YbNrDlfB+DumFBNhbUTNypz2wxcMq9u
ZAZzZ9nCmuUhoKI83MraWo5c3TeVPOMj5RAX/A10aL53mog74R55ptDC7j6hQV11
wvgn74Awr+Qt/R7exTVAqr8NJIGmOtz4ewegXoWL0HdfpBr6V9TSCaiL1Mqbm5mG
6Be6oKdToqIOp5z6mXiKGXP/TqLLjsFbZQZbm/Gy8YONr6PjfiIiySZt2gTwDTFl
LB9HSravwmxE5Z76wf9kW8uEnDMYWB3ILrJkXjSsk8MzuddBd0hVm+mQJQTJa29Z
yssFkk7C0bGN0cfLBFnEHLtxriH0StVtYCcoaFZaG6Qzx3S0pfXkd+/SV6Pdkrjn
eZYrNldS5vzSeooXYcXeyson+yzK2drYtAF+r67h3IEU5ERYN8lsRW/bxb/8Pg8x
F3lWaVEGPcyCLi0s9xBcMIGViC7PpfpLlCpWl+awn/2s/gmdPF3EcEIMTdkdiCqj
lMVSQkC8PlBscEpRnL2uEAFEc5IZfFcbLkaAO0e2ghdFurgWzuxYe5NNS6yyIdos
1Ky5Z7AIHfCLvd+9/zHPauSAfxu1ld04Bv97vyPeqkyNmR40WSZvHdS6uoSYcAJ4
efKO3Ay7lsVuEpYzvsVhmgSi01rGximJg4xeMkgCmnL2Qnl7sjOHDRMD78rF8ZrM
og6h9BF2fkb8gbvjYf0IDyUHUUWF4nG+wYiripFyISCj8pOmd4oM1kowjN2vyx3h
Xy7IR8L7NItdCNelKr6+nrwCAwURogzLLKaADFjtD5D6nHiBkriNBKxsmnY7sU4e
5S7mMIQR3pvrjeQJIplTN/9rXb2UGA5pvWZXStgw9pFID3Mjh1qhiyVLk54iJ6Jm
aX+uSEpLjuWr1P9UfPLUM229urrEpAdununvlIEr/9EvJaITUIhpF5o9WWiA0kJZ
R5hmOKWW9IsKkZls6ofhrmYuBW38jpOwlPNt7HVyvbraa4pPM9XY1m990UTQzOCJ
E0nln7+jAShTj3EhLBALn9/XF7yqK22LdY1zLbaT/tNez0FUxii8qqgM4sYwlC+6
RNGhQbnBUr8DD7+I2JiRei2m997mwIzMZgVdFkxfeGnNXViIKFqXwfM6j+oyj4GQ
3FkXVUff2olDL/3SQv2jJ6PzstGK2hA7zKpPTq4CRYx/69VSRKTH2jDMpZxDWtXn
FExxatYsL6JJHGN1Ts7XZyDFVbpEVZHnP1iRHStIL/mbxZul8y6THD6PKRrhbykE
PfPMG0bzI9zz0GHg+4fvwZiqy9PeTHhF7UGNZoOC5HCMTDDc6HBKFERame2AVTsu
D7BsBdNtIGjJ0c5XugCmMiHdIX4nIk6AY0XqJ7f9j+vTabFOAVJ7/TPXbuiF+0rd
ckIZKf9T0/Hp8kYU4H9fjrJZ5Nbg7QUlroJOxEL4vwZzQ6kicIAY6kszVlAv0a0v
8p2hBQlXI4Ry3e0XpO52ZdfgAbcfQ/kpBiJKghs1y+JLGE/hrDeoIBPm8Ouq+bTK
wMqGNwNXLupeRpUDfZMd0EVBREt7dndMwutH7jr00wkS6QchgqbhZPgxbp/vQP+T
/NcWWWfgSFCi86RJz9mPSCCml0XgOjX+BAhU+bvLyoBVC5V2qtyALs1zPWE8jkbM
CdkAOCBZGikiR2tEqm5Svvab6OiptlNWk63x5TZ0DWsY6f8yWFX1Z3o+iWtzR2OY
WoCoTeUWnDUfhGmCXr05uE5e8BlC57zo9UP5eiCFWC17Zj8KmangN+/Mf2+8ldq1
RS5ECDuGzNjxmfCYTy2XY5Nmb05DXF43WAJLWdHKInNANPRxpjbCJsDXIu9afRGj
/LeTNq2p6VAyfzb22den3lM9EJNmwOy94v5Cf3TXxwRVWyuKlnQ5S9S4uYO/oGuJ
IXynaS7/i61AM9XUGQsHmQfvgm15ajykIu3hwFwS2sBTYR95Sb1QsVGfK9To5FXX
xQmiG4PPQJY7Eew7zyw4ZBgS9QF6kL7jci24PFmFJUdzi8aBCGBpaSOOFxp228Mw
aN0V2mupBGlb9tYSG2gqlNvh3Vn+4LUIe8bM5O0MBqCdIqy/vIdxKmjNFNgp9hSa
KU+3XKu4sAvTRcup61vFmjFfAhKD+rLg+lN8dBiVWlygNgPW5F1xl7zL/IygexWl
nZ7KtINAyTuSwPDMS7tH+AXC0Mv5AjxuWr4igM7s8DzP2kFItv8gsJSdqLPIpI2c
zfx0aHUdFFPMy4jnCi+TLX52IMneiHrVZjoKCSJFmQxW3kXZ47Y038Gcqt31hhiD
lk/rdTfiH2D5CnWXaNm8fNfsSWioAuHVMtu6Yyrj3I2Bwq+NfdajJy0A5Espf7Yb
QemxFW9k1dE82SaF2pO26guTt/mHwjXT6iS0YOnhNKM7kBrcd5Nv+9v2FWWRBROi
bZC+u2EmjnRVkSM24cuxxPqvtuUhBImUccmZHQ1i67pyx9QsmpGGPShu9vIQfzki
gPwr0UA2Te7YYP7Xg/jxKJi2kUQCsn7Gf1dJnbO6o68snZnrnwe1pIfOU6tfWD8e
j7iQlEUtKyFNoc6nSRw5Vz3U2gtSszaNulRqAbK5fhQkUI6tazk/4tpcgx78xkNL
8/EoMQhxHByVbzH68Ro8++YMrcqRwX2RpJt46qQzUGJSUncCB8SrBOwZjpqhbYa6
fEHG8sl9nFtnWdo6qZUAlhKYXy29TPMzBOc9rUADx7X/wQ9IcWqcNltuAj7a7vCg
tEdsNXJ028V7inWIK2ZIDomRmZQrfcRRmIAnUCwl/WpSWUvzpeDdnk8zKhs1IQkZ
xzdGvzzJ1yQ5ylxfYY+4IH1ecQko5ksiTD66+Kx07rs1mIkVzbFsFs9ppg61cyYS
Ll1KuXg0/9Dtuk33e182BbRQ9nzo5tvQvDizBEFEdL7q0PHkfFDecwTaVKyUig6u
4MHeXK5/0tCG/JSctRuN8xYZhLOOnWQXfIzU2zuAyACRUzf7aVALrSqt62/Qfmer
HG33YMtTxgz3SWaL5naWqxjoH/cr8JOo1j3hYaXJW1kEVenDiWz6dyUdoqL1wUDz
NSxyJ/RvKD58X60ySF1KvJLn0YkvQHyiCr1WezQMA28yost/JbPkh31dl5fyllNp
pwcGacuARTJDOVg3g75ju4CiDRsXZ227taJjzaSHqTWWR/7qunDX1f6y5Alq6moJ
H0SbEwR+vPdG87hVmZJhr13BSpLydKPBdemQDY2uiwHjWo9Jtoe/KtQ/IS3rjMAZ
5FP/b1q4DNsLmioI0w4Qg0blTYwonE/hFSEyG5L1OBhMLhKAhBsEbiYVhJCQNm74
Dv0jx47aCdbyKi1MUVNtxKNMpIxiO3iEo9S5Eq8D2Y924esZNRJ/X28fGRFH+szD
6OhT9uWejSwP2t4md7NrsPirUfovhS951aV41bn2I1H+j/9lzMMSM/vx6t5GaBiS
9HjbQCPoOsHDvG9g+S0U5FHQOLTHurjhqyKkFsvi0r5qhZnSVt4OTmD/MM62qGMX
ktgacNBGmBKu7UfUh8pz4whqWHRdF7/S4I3FDsxqwvIaYljMI1L6M9VKIrTxCJPT
Q8aM9XTtdVxkiXzwwY7moXun8Rb8Yis7njG/+CcR+QpShdmPG9ssGoSqEUdneKdr
J3RlJqb2Ox5d9OPPuOjLDEOE4HFesE1uhd249T4gJGqr6LqY4ME2ch1zwMosrKjD
TD4NrHVSKoY/b04YCGJDFj238vXOpkhajY3HndFGaXZij4M746thtkUQEY8pUH7e
2BJts+392qhvWV8+2APjJorvAdS8WYt03HJOhFQwSwQnIDx8WMfKp9E0AVG6mxuH
c1JnzGex0St/T9/60pA3IrAC7Xv2CwzddNPoA8spbIJz2KhBq2bNp6TgcuA+K7Ks
bFincVT2tt/EFZeoAevkEb4uyD+Nu4seUP/K50d8ABRYhjTydLre52MV54h8Yauf
ssSC2opPTAazkL7jc3KdWx87h1+OtZ07YJySexATYRNnv9mHHBWkRkAZ42V8d3J7
4YDUDe5DMW6OouTzeCcjblcrtfIJ7MQQE538ZzozJ8mD+M8Vgx9uroKNnOdXBp8k
VdKdqSllTQQ0/+altAGY42Yx4vB5Wa26YDDsiTCbUt0NbbYvWA+NG36XwkqZsEEC
FtOx6Il+UjehCRG1VNB7OCUsCxUqJx5o/POGgm39bBrd9e46mg0kg/FdyPvmqUp+
Y5CrasRcSnXvZoh9oJJ3y8ZijArQDiW9dOhGfgs8qVAfAJ44TUmb5YMt736ICi75
6zRAnWwtiX2Ui10S8GX5UvRy1J1gTiAJmU7CqWAn9xYNoQhBEItF9pLOFbwunaNY
MWLsPyGHuhcNzw/IjVKdZyqfU7jnktM150vm8U9o3ZHUU4885WhdIREIIXjmPrDR
KNTMUqG3+cR+8jV1NKG9IskAT27STPq2aCnyzq3g70oxfZzIbM7Q1337wrHKUZlz
51KYmbRwoxKLIsKWtF1s/qLK42m6+t63CVXMcTvjH4g+NAQ5cNN8bGtJMlSop2bv
HSbGlfBFBEio7RqkskbWhdDz5gNwUXnsLylzolxh8I+oFY62aMv6LaWlfjdsOed2
0j+7sexxPFnorPaSdJR4KKxvGkFQCFfTJC5GZ9VMGW+L4b4WKltYF0E0omDMrMy9
+yE7RSwCF7JnTT9crdbcpkTf4rmQgPJzEDw/i63DlpCoqmTsMc2QlO9CZQodcrl4
XW8cLz3TgyL6NuI4odAra73JsD8+v9vo3lANmuo1acgLsLHLC2mbB2ZEULNVUi9V
AIM9nmNp9cEplaghyQsxtfWZ3MWxHGMw1YFFIGb93XyiICWG55toTfnFR2Wo/bGQ
/wPoIqvRCqHFwUXm+KdM+Z3rP5kuAA9lW4wg/Rcb6VNAPejHqYVqP3NyS9C4lJm8
i6sC0csdr80eJ2UdAMK4AjhTiL4jO6yxHVbPa0peBjUzWxcFDpq/B3sPXzN82Zj5
KBLqWQepAmM+2tg04AYCcSJGst6WXpqtScTM+4WFhf4xjkZ0l7rj0v4B1vUQYwiv
X1ipbLLv+kEyeosEY0uvn+AhZ2DOcPWuUQ3owrGjuKgr5iZAGgLbjyL41avhXMjV
9y+g++tUp67TPiVVhzYF4rJkFWOFDwSbt6bfmmw5ypY+YYJT7exZxmr0Uzvpyzg3
zwmWpE3Ofk3YQ7ADwW3m8a/lOUr1Cbia9qclhL/U9bFJItUYdLPPSSEnsEWxEyN7
w3ww+9dJxprDjIHXupjlxUmr+KN98pB73prrsznuOAjfpVQ+w4F8dw0G85ErB1sB
GF4NbnXS7vlnDzpjucH6fCW/NAcb9NTATYCJRPx3E/h5qsOzeNUMoecJDSRhFxmC
h/NeaIYuDcfDOQj5jpZRgHDU2P3kiifNFEPxQtFetH3n+QLo+XLOuDF49elYb7HG
9JKI7S+fqUtm/eNgrDXfBPrajQ/bpd9pt/pnXL3evV3xgg7lGHSFPOQcTMvJ54wk
a9zecbXc8EHmqb9uoQPHm2+UHi6bkS62rlM/UFSZNzmV3yluohJx/xQRWhNRgSkx
ftfp70oyvTGr95aKOnN3KA2Xvjd2z/budLwWMutgoG0XkWVLI+/UKM9ZiBEQTAlG
b0+jIcxwQh4kRYtVCkelOL0yHrX4SQtwiRzeM7KMIqgAu0eoF+EJ9ewkEkDy6L4f
DZj/1ZaAIOoTr5B8QDXwrknbMBCFFs6ZGDRo7SNOl+b2ke2/h0e99TVucqwkRSND
+fR6M6Bh2aYudil2DdHsalTmlfghvwXf6FKtsHsC8hWiwCWlsBz1CMCDIyC3gW/Z
dhRLpDnZNOu3uS/LKdDrpTuI82wAfUdCWO2FPiM4XicoxW1S+0+zxA5idEd2zI3T
Xx5Tk14xYE7lW8w+bqGinO9SEKFBvWualMuO29HSfY2sMYV6RGHNnzerTOJiwXOI
NNiUSqjEImSzVKuNd8bKhuJdq+rH9Pms0Pk6Q9Ww6TIjDqtDBlCRNv9Uf1/2j+kp
9xdlZ9qKVYnpazh6X3fScUOtzIZygYvA5kY53K/krCaRyWOwonZd4c8cDVhSURl7
Im1MwIfLc+pTzLgz9gPbwu1UYOKlkZGp6Lk6/0QDXZRuYGD7jrjoVBkbR6KZckZK
YoHdNAO510mPfkbqobbN8Q/Rx8li/SZ+fhCoIMPx84/QD5evDnfz/p8Qo5203xU4
C8kKiyrnm9K2S+XIO1WqMVwNkhx7xZG5K2byK8sRAPd91NH+IBrAJ1+Vy+CIDzAf
Xk4nNv3KNevlC8SVS3v0wrisMj6yAS4eVgEf7GHIgw2BbW8W9PHIfMTAp7/8054b
/3bRibHk7gH+PTtIXkp7NDxs7Nt3hREcz6WGmhW+AmpC51eRkc0hiZUpRQNDnUEX
2EBA1CqiE0D/vNoYvygRhUS53qmbrhJEi/OSNsutz9Iu2NOqlrROKqhP4hV96A+i
J+RH5uNZMHLCvndULPLE6jt5xCu9ybYTxO6qE6Aum6JDbTetsEakx0Exh+DoIy3K
nypaIQikvc1LNUtCcEGGBli3Ew6FhON8K9NipoHwA+zXBAHJo/kfU+rOrOP/LYxH
vKW+n9s8veXDXwg7PqSeW5ILAGcpk5F2lcXlsE5VUoJ9+z+/bh0YpFPc5vk3Z6w1
MEl7zEh+ANZ9fHiPTFptjLVDf4hA0aC1J+qDCFtruvlm+ojGp6pfZ2R4LyRRVE4p
XHcuKQUwENYmyAmfR7zWy8nET83LG3vdhf+HarJPys2KZp05luChj3FIJTr8aZAE
9sswURlQ9dkKyZSeLfnygbZ9m21/WRZTYj/97oWoMZkek/4XSD+rpJ374oQkAEjo
PryWdKmozGrMglOyijkrK4T7nMXowoADkAHQt+EHZB+7pa+YyLNwgDPKx+zBQJGs
kYd1v4XCJLWJQ45x5boWnf20VifcyEqaZ8Py+jfqzvw5taSJUnjyWRXczWHAvPuz
hM116dNOBC7HupFKpnl+gjPkhGNJ21BFfKPdLrabFpidPMC37Cd29EdT6yR78qgP
J8iuXNQtR+JKLCYIAvaGSmkViUePssQ4r7PsGoPJKReYD5zbpucXB7jjEM9zTH9Z
UE+GsX62rviavIyBXkPVX85iESqmVlXhxDu8s1QW46j4whmVK/qL91sFMzjEim6T
ZC2+5cdMBEBgmLNtKmDtLwnhiOrjVles+BTBNPZso66ua6tvj79dL5l6E3kPTDeL
AkxU8aeEjJNyWgi/SXx4ZfC5mblCxmWUJLjAAvv4qznTGb4Hlb8PIPX65ymFbmUA
xwOB/mEPbIPtKGIGYowJ+xC8zicnwpv8zYYTxsrs9GL5E4dT5ASFTysqaQsKznoX
TqyZz2GSCC/Hwa2O5hh5KFFekR4jMI02LvcBQRDJ4eUS0Fgzm7Al5lF+mAYt+NDX
UYeXDykO4FpxMEjJno2gdKJjEGlZAVvyLrBgKOnGIk6/WO96BKYg+Z+mtO9B6/LG
4uGphFVix9s0fit2hBvaSvhDKOwLN7ZEMHRdlvI4TpXF/64kWJRQOrnwN5VNnjeo
Nxd2166gCFiwmlgbk/cb1yTs8oHC2aCiOHB/DBR8qdP3yQNBUojvoC6ml4hBFvkf
61CSgjMeyGzTKEn6ECec6wb+XH9Z4N+X0rc5/xcywwZp5Om+MrLXvIcwuCa94GXd
MlC1QtcVN4dMa2XKpbps0UDiTdBtGnj0uLAmyuTrrdD1xSdhThWwXFTFdROCizy5
P923qEM4ypLTTln3tfhGKu6IHIMdXkEexVMcobHGQYIGvyWEmNhD8BLRBGoNxWqV
7/BzKmff0tncpzZUna5Fh2S4Sk3uo5DTRfskZPcIicKLaKe5rrhsevWUsRnGpSK+
XQ/bK04i9Op7QIY1aVL4Eg9kVjIDhfBHgorpRmsW/+3+JIRVwoELJNZfap2vVU1A
e781bbLGhxNPUuAOmqSulRGhw/tnE4d/Ltgpuf4TnmQzQgOV9COlyElxMCtZXQif
hoKLkq0fHHJybASf2afvZXKLkAjSzINudgwDhTv1PzdwnKHsdmKUNeS1SrkmHvY4
Be2WTLFfzCqfQ4ExOuGr0vUbpe4b9V9L5rhhV+pPu6+uWF62hDk6ieEIZqrFmIU9
t8OExFCOM1YPs9i9BJkV0anvAamKiYzfFmMWvubS5C+EkwsQMFWASJHjNT+cVKQm
vSUeOuaYx3mof2Rg6K0KEQUQz8TEPsuom+pi6aWVyL0z+u9ETARJXWDZsssTne90
DfmDAS0Wdc0oEJkWDQt8moKHH83LLqhfyaZaJzy2p+8W7JHKyuCnY+E10y+SQV4f
jQncNu9Bm/ZRHZ2pi0jSuEiBfCkYrjeqG+oRolANAKbINsjy6uE5M6kTJbzoTL48
zE/DwxOxQl3sqFpH79wG1aJjbWCbcYmvdaI1MJMo4W1Q64VxDnAKw9GOX/Mh5MMt
umJicAJFFhHx0iRB5ghyBBS6td7AzA54JVfowignPd1Dg3McGL8OcyqiOcsVgj04
DWdywEMu7k/YIEAkm80ZhizCQoEvI3FhGlfqYtyQVoL7MHUBZNJJRk6BDEGpEHu+
EG0cP6lDFiszFNs6kgdYHqMF+qGOrU8rP+Ax7UH6/vPdCbstzP/pmyRlGNaugUwP
DoX2xvBdKBen12q0IItOVBs7AXVH3hRMrMf5kI9zMk14+WqsBYjgYflFp11oECHp
X0jDtiiwJh1qHGlYygISLrXN3HlFUUVpj0OkBHabOxoOsPkwGHEy36ykK3zN2MEZ
eovzhFHyaqZ8y6miAn45cdmD8Fy63aQmgDi0SEXGspGh2E6fpf0RrvsJ9aM0VxyI
N/DjYsKjAbkh6+ltao/kN8widksOR3Sb+NHUN78U4kGgCu7ptIol8/gKQa37cXnR
DjW6Tm4xWty7ywNIhEO08ALHhnuILdzSWy3nGtQcpi0lIiPVFZzU526MLLfFx8vy
u6M/KIp8cvfcKLnkTU70jCWM95p4m3FqSSi2w4JtVJL7JCYCZ3ib9lFA1qYZTnnG
7Z3IQAN1dhrt8TgTX45HWmzpXHNJueI7EhlkEm24HwJ0o6vi2Xz7pB8z88Gt+GK7
baKW1JyHrsx79+xnwcSbdIV/FD4EMg9J1bDBvcBIK50Ra6wJlaC2JkBU1c/VDRfH
Q7uj66Y5hwdZL0nxfgVWRCMXD+ke9+MRkHLkO7iJUaZ49lbJERSkbyrPnLkAj7NF
01cKzDtQHOgf3Tp55YZDgqTmruZqlGptBhPWoLIuqxzglZ2DAEILN38luipPd7Nd
kiRIp0oBsW4ooj0dAaoZaTVTIXEvnKh7U5YfwD0K/Op+T5VeppteHdEerG3xmM5j
NmtiPMf4kjdeA/tfaH4Im8ADWJVIPTqSi6NtihxKiDI3zUGg4wg2CHAbCBR4GGWj
+YKtq9BEtlhxHxkH7RM6ndRvfsRBRm/9++puNs68Byi5KRMIbtM1is0i4kNJ+ypl
DmDhkUbhv0dwSzHRHUd2ZMMAc9TiDl/yDvDI2n3UWulzTec1efRdDmLRFyuG1Wag
x6B5LNKFPUVAnrbZ/YrsCOb7JasYPrnoLXgjZTijwbHzozSabnrnjfYGGee1rbd2
sGCLcS+gAl0tv4niX+svCBNPW6+XNu4hCh5Yq2pytQhQNeL9PcSrYTcKt/nE8eZ2
hMIcxsV9sDVtWU1JrfSCFBPlhCIXXXk+jrUn+liAfWXExw1k/D7j7U8aTKpglfQ0
8oic4Mfsohq2qmBtU+Mga8wd9NCkUvgjkPISmuo76tJF8H/aRHDEUdqZvW0gpL0T
0D4rVz1zzr23xD0k59qmhCQGZAX2n5JueWgkYq6w9eoypgd+lSP4/4hBK0JS0G1K
fqDpc/flnIpPJOtdvBbueDcHGAV4YkD0r8FLw/o1a8CWo5pewjZHalUHU7vD2XVU
ZyrmkUcZ/4ryu3R9hV/crlhq1dZQ5OvySr2HlNVOHoxlY1hRIbCrM6T4VV0Oub1l
SpoEVYBbfKimCfZjnn2JLuOvcT3r7h2x9VYZc6/dezlnvEeXP7m5uzd9B21cQVPM
6Xm18MWY+mkGwNTAopzEKE/03z6GHUjXZvl9bll16uSrNPZcBCrUZsn8AhKFuVbI
GANZdZ1CYpYjQi2xT7ycdMVIHb2UciWCuQwfZb7JMKOttrW/1m8gtDNx8r3Ndrhl
65uXva3IYNSGXmGjP7t6oJLTlGYCYO7JuhYGnS13Sc6Pve0c3F9a1D2EmRm2hMt3
Np+jPwpmGGKgUyYd/DdtP3o5m04N0GjgaxoK2HuKg7kHtWujEw6nbn88aQymVh0d
vrhJ/8Lj/GNUELC3AD2+HUBngwncsRsGLRI6wiIMiQpGeeZkeU43Srb4YRIiwTxk
wnO8DChsElMBkeWLRvY8/3k43KfS9w+AezfuEstjOM8s5LeA1oS6X9kFzITodhVO
wcUmj7U3xW33PrSmXyLPWZnqWTLVVFkDuspmVf6D5Vznd2cnQfuELoijoLiaZeDo
kwLtotzf0nWyxRtptxX8M6qJR/X7RkjlJ252rC06cseMzBes9ZOJzRiYU71BWpcj
O2g3l2LXYfwc2H8dgSgn4p+IxAKSZL/QzF9cImsuasD9+raPAxyxMc7qRJPunlNW
6mQQq5sCf45418S7ppD6dcsaZydaVxT5fADPvvbkfSToJ/bvb2/LSqxp/zBaGCrv
RjYQwuFZZ2lDZwbQqNcGo5SUXTlTbEEmx07BrAA0OUpYdEIBw9dLuh1xtT8x/9Gx
M5ry+SXYSK7OnG7n/MmO0p5WsQU+FVzt19reumRApcvcsGJsqXPlQIMuRO6Yx8DM
wAVwkzxmUUVeDzZv8aRaoio58dAyZz5i50xGUiSaXFb3I0YmETBfKj+KIcVrHnYI
Vbep9kM+42Y1KYiccel4qfg2gszfkieRJTIQJjlBScueVQbLwyyBT6WC1O8jLPjz
AxwkSeyg5VCrqpu/Vsn3jpwWZA05/IbIh7IzOqhmkkxuzR62Cj7pSkQw08m5vJ+d
XbkGhsBBuM3iR+fntmLNmju3D5t6NTqpuASdFfOcFsllLpLqbVNI6ooyMkX3bicK
luT2BSISR+KjhFSoXofRHcY3mu7G+gJGpn+jSjNMlXzW1m6HP/l7Ia2w4F2PEW1e
YpMhDI4Qi40RIi102qVmMQHxHZh68m6WskaS062+WTG058gKq682zAa8NhxNSr45
z2ZSQQo2Wc/HmEVvPRxtfTzvWGyn1ujNrO7DPBVhDM1AsCRPaoFhEXqMbtw6KlE1
SunfdYi1oQfPv+kbSDkn+lhuFWynYkhXDzrTis33rvxeEUX9/Jv42j8rOSilTFQw
VvSdFDDe9y+sYLEwzllVIpg8rCqyCjLMyqUtAyH1cvOUo2PPGg6xq/lvBTrTq8jD
z4Bj1rrikXiRJwxYIjIUdJNv0RLN8SUzTC37NzPFrWtiGUXPM42UB1QRy1ygnyz1
v8Mmr9yN/3TN4w5y6HK4KOWSFzxJvXsxK9/7J+tWzKQbabrws67/NNmE82xKAZPm
TnqAczNu4l8f4YV8W3zOKYRzIg3r2Uq1QLYd6xpjjOkZpfOrBWK8g9c4iO3wC5oa
GZ89WGLy5mFMracg7iF8QDIOKfB0fsG1EO9ytaNo93eAQtiAg/b2+wPfBh558nuP
4AUyPD6EivL67lYPoYE8RbzhXZUr/fS5l7Si4NP8PHPNWDtuUDk4b1r8nKYRKJoQ
YcJf+nnuUhG7r5U0SF/auXQVZlAxXOLgpCG89HAHCyr1vbfQV0ki4wGljydmbRd7
a4NJ2KgO7pP9nzQQq54eTs3FWbCWEMQZ1HAc+ZGQ1uzWf+wXPmoFxy+JlVdYZ7CY
CEOd++IYMpTY687gXPoS/G08bEknUQQyduyZC8k8u6wDLYL9jesnHZ4JD/nr71GS
ZA/89NGMBPJf93rn6ioNXpar6YvvdCY9Ew2D1kVzSdHjHgmImidCAq4tsE1tjmag
ik29mzGJISbln4mR+uBUrAeHXacGZbH2DWPMfkNj7UyysEF1ZRRmJUDAVFoXh0NV
yoPh38i4QAjNYI40Isu+p0jjWZ4LiuFnE1Cdq1YAgFGhlf+WveiIuCPuVQ2sFkHt
iQqLCWfsnuA7rDti/ZiNyUKCnSc7kq7awLMiBHAN1TCv5Z1imDs5GiCrJcjP60hr
HJ0BBvLpKmXc2iItbnS2XmwAwwUq7bYypQkKvxgrZDHDLVT8DAo69C572e3bVylI
TyMQ+c1xeQu9KuLW6bUX4/dCY6QSeRAdxmRz8ZDCKVXVLaP3jzATPIgDWoByz4I1
H00oC0bDHPlinuqzvznipvJ0i8TRgfrfkpw9zCg92ntsLfd1ywsrcLs8v+U5ZtyA
ShA2QxW5GxJjIdgYnC5XRUkSWj3imTTMwR8n1a89kLa6vM+5mjG2GE8WZDpSmmTd
UaLnI7spLtDMSbk3TLEsbelIL9CUO8yqiEWvetpUnpkoxmJx6B5HZVX/WNFxDITs
cP0qhzxTVFBDUzpj+TrxmpFXzXke67t525wuIP3my0JMq1rEvW/1vXZs8GtChJ/m
57IMKuknKgN5dnE3JzYqjUfEt73v988CX1AoQ/Ffmndb1MQx6JYaCD6Zc0IhOnxq
DPfiWAhSujAkB6mA6WruOaVLdqoV6Qy+6PJi3w65TwTueAAP3g5ZjodWNnz1Rt1Q
a72L6hnDa9POkKQx/73yBbuF9RKVDQibYQHLhDwWEcw+UUcqas0UzwrBoegdjGcb
RRESZ6jNtdBC1rsnmpiECtmAaoHlAhjV1J13ZWEZHKBYkvM2fypu8h+KSGZ/faEX
dkkjFut6wil8fKIQLfXkfRtwzRTeqv6Cuke6ScJvC/Nfo6zyqI5y+UpdyZcQksJm
wQR5rmWX1PrqTfeimNUs06luz0yUoZBJcoHJDJCE8j+cvZF4UkMBsE6tWJr9w6mg
lKkfVfDxxXHWF1l3M55gc5eHngDOFuebcxcAOynrkLLnpSe/arEHfT50gR+fz6ao
yK+d19TOfdE3aNAQL58qLml0nsiAIhypUaGUDJpt1KIUsH5uNEhNYMYfDif0S3Js
10zM+lJ+wpI4YYoWkGm5IBqaNKpHYJwlZlcAEeYZEpnkBntXEJAsP0K2Kn0wN1aO
+N+HVpOzc6OvYIMQhN+HnF8P6wOT29NN2yb/uEi5E3ZVBg72f8gChcG/nRYkta3Y
sdTgsO52Cxl+hAicc2J4PTB53U7GQqkiRcTaI5J9LxTiITRPLLvrVUzeDm5EPysa
hGUasaqc+dj8/y+qyE9YZBAL69Yhoe9GByiAt5bymdStmof/AC+fQgRbZSq0QIu4
+V4g7B1juR+IAg0uZctAK3HNZ8Ld/v8Fz7OsSXOvYck2VRG67s15Pt58EaLqsne4
jVxOyPrGyQJasMpePwqnakb4H0cTH4Gr0/gIsWkqSlM+VRwYOyUemKnrcj/saS/L
Gh7Fgn3fRoB6Ig0D1q1F3tEzHNmsBpBjAcEuAsyFMKH3cwhNAaYG+xpXn7CZH5wo
omwg9PjnkG7oC/yWTkOGrq1mqaeyhf8DytTwneChlrhhrS6YbMNb2pond8TpsaAJ
1RqpvivT+tf1ErUJ+1kOIKDgKZ2zTrgWJgicgci/rmKYC1tSNfO08BvlLa63GhkZ
TkSc/tEST1J2UfvvoYvuOckH6h09BKLa3DgmsOaVFDxtpO2Ml/RMd059nlY+juos
LiXIVY7E69ydnxRUk8Ado0qa6dS3+kZJixtEg3spzZYlWTTxAilASNMWo0WxpX5x
Nbe2/6mbZ3tgmbcGxJXd38cYPGoccoFYGpmEoL+jDdMO3y4N311hhetTy0ea8bqi
f6824oGRcxTWo0GkahCr7XeJ5l3ae+zxYG26nsYOOv/6Nncryo7NXCyyb2V7UhLU
ZwPwZSEDghdbgJMtr16azfsd+vY2MnTt+vvL0zNgj1tj9HuZZfC2bP+MlMyTo1Xx
u3GGmpugrxdLBheQwhRJLIZb3XkuH3Ni6XGXLwQFCrv3Sfo63c5sMT6gYaNoh7/h
kgcbTVImF5m/VncUOPCadBiMDK5lhgiSWMjBQPlQT01DmBQNFyQp+zNImjD1bnZR
EGhmPa10mpkpRSxXPtMD+QxCEqPEkWynngaQDqXcCORf7xKksR1tv9+MenHjsLZw
Up/g/O6M71e8+mSWIwpRKoU7hvLpE4+gd8MgSIL6fK6slp4aTUWEdeVOOnIywpzv
tylt6SjWYGk0rTOOiCHsNWIoK35wKirUbFnm/Li86EfTpVVYuSfOTIJHzH5YjSpl
UeYIbRcUuMkj1hOurwKrYyjzi34/BK4WG+rrZBPV5Qm3dcx0lHEWnMiozYNU15dK
jUnA5JwBOBfG/nmrKEQifpDIMX1yLH9D7EjYe+7ldvndPbeV+/mUSWl+CwJuukkL
JrBTcOjZSZMA08m+ST8Di7h9uZTXOJwYh4w1y4K0ZoHst1dzYiEycC3n54UeE22Y
7rIiE3TsvN77oCdLuO4lMjCCDpfbMpwCFHAdYdSV/jTLTKiyToDUblOICyE8qqND
2K3qSt2BAhL1236kyP1+rJjq9Vf5iDZcm09xZ6+1yvpGjLBYWFbikDV1yN69BYPt
5GBOCB0uxNh78aaeCGrX8Bws9Hm720gyLbNcNNudplFke387rrNBHRTxnux5dpMp
ETGIA6kiJFCLlL7g592z00HtiwQQQi35mtDLL7lRTe9YtYuQVvU0M8BncKlELoLe
INZyqYOISL4Yo47dSEtKsy6xgol20yLVRSfvCc3RV5f4Ks9lBxWrUzncJjiatGFk
z1JX79mij3CptBX5AlzFX8xtzoLPiouKxJrW4vQCuqeQrKKETpn1kJ7tzkRdkFR4
/Au3thN3OVrmy1fEDM0a4/HajD8qWnLWHmXA3mKIv3CoNrDpPTgrYxjz/Wr6GmF5
3V4wCf2fynx1V7Ld83oZ34h5Lfqs2lwMz8nxglWOQEAr0G18zmSM0BOzgAyYaKs7
t03oCUB3YumIYW1cW9sQbrTePkKhn7Zsh2thh231I7IIARCh3kbFaq11R0BWGmCb
mRUALqt6Fypv79+04YfKECHJhUV9+qtc5nFHzzv3LWetJANvn0YnjO+hpz8JksIS
ZXNZwe2EI+doP64YKLrBGMga8GyxcFO7WqN1TJWaZ95xyqLO3/lk1xpoWtWzxPg1
Pd359rwLaIrF5AFnUGS1eHHQxqmrhqGLFYC5Nm8vLJZWCS5iCj5VnM6gP779TaR+
FrYGLKBiN04JWLLSs5ckntznGUdW0rRiw8IG0FX2nUqMERldTTxjZG37qV/ZCQNE
ok5szf9iznJ7DX6hgaonypolPxInvr6Zwrn3XLdJgWFbFXYPwdRaRQ9oR+zkHmfn
rulnJ/8O5dP9ke/l0CkZB1yTv6KKJmo76KGg+kJy43M4IvvIuWZm3NtiTo/fTITH
4O2rDxerXDrbTM4l+ChIZEDst3q0SxYhLZRV8d/rXFM/sg/gIwKkvmjEnrUTRJhN
I+eT2vtFB2vnzMna7ZydfyMnoBpD+k0fWLUCOGoyufKbtljLGPsURrP6mOVn3ZQB
9WW88W56k+fdeRLIaDcPaCavCv6YUkNFL3jelRov3YqcI9PhKxwc/r1WQuvZF+4f
nbqOgIgZ4Rm9LRYvZjOnSdmaH4x2pSQvznquLDFrxKOUWqSHpHS8oFFGrpWLHHar
a5GxTFch+a7NnCkatsWnwAvnvyDv+Ktw9rDvQCygVxgEy/BQAl2T0nT/5/ETvN3E
k9875EunGQIM1pWyib1mSpHk1dMG+ZZmc3usFsvEJ1vuFcBV4khzNT/GTvRqQ8De
XzkWUqJ6P949/MWcuKcWmSdpw5oHPGzYbA4PHg2jyjiFSOcPeWyhjL2Hrqf7+9JG
sBnZGxokF9XI/xaPgvFuBBmOX6lei/c7yF3q7rXo04OBlsufV/J31N3gIZtcs/IZ
wFtXObU+bOWqOue4Ow5bfYK+52x0gsiAMkUZ5IAEDzrJ6cdUvqzftSqjZzhch0rm
HylvnopOPYw87zWjsvM/yQxdawzidbrEgjwtRPmnys5h+GqUTtkGZjMTkSpalG+y
/G4JGdEP9kUPGLvQi2eXO2xLmBclCSxTJClktahdeMA8LeZSUEuMyUJ3x6q0sljv
yL+89y69yvV1B1MV5hXLXBBI+zymttZNUmhZfd2x7wEmLFQ+Cf6/YG5wAueW/PsC
NSF1bJsnwHbr4Fky1cC3wK8+xtV2r/MWvzlrqykqy3TTyp3m8upFujGXrjmw7YNE
A65K9G6PrdOiCFtY6rXFwXkX7BXQQfLI8mcohSPXK9ZYGECIkfYk0SFf69Kx7gw3
Bav9T9qUDtIDSgiQy8NhcX/QU37OXQsPVxlJv+3+LuZ4y9+GfMO+Tu/wH3FWLp+B
G+h+LrZuuYtEULwjOFnHPMnFIzA+JxWAPT4QqWTQxlY=
`protect END_PROTECTED