��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q���u��������=]�kN�YO�q}b��9:Mi�h浘	Ü�`�l��չ<G�|�����c�����\��E >�l�Bv���� b�-��3@=؎&��K�]�����06���p��q�}�xDd��n�Uv�.)fPR�1)2
|`��1���K����@\r�r��9�ju�s�jXb>�#?K��=GZ�ќ}�h}U��Ir�t���{�C�B	�Mlq��75���O&��S!�buu7ɆX���a�P=��)%"��g�L�#�EBˇ'�Ď;xd���+}�n8?�����5�x+B�6�U���v���g���&+ގ�R�}���(W��^��D�>����𷽻ۊï���&R��[�ƀZ6ORm~O��ǂ�z_��xЏ-�ǁ
�*��6��Q�'ep�"DxX��,��G��_gb�
ҿc�W����P�^)�()f�����f6��?�����~o��8��m��
r�m�~��qW
�_:uT�{B�ŏ��652�FuD)���j�^Y!o�dzvr��]�
�!tY��_{�9���8��b�?���q���O#0=���,}��8�g�R�b�[�ˎ�9v-�<oO)}
�}����7z��!Ǎ9Jbej�%��b�U�}�3+05�zT�M����U(1G�]�	��-x#`��A�k�x?�-����iD���μ!qF��H��Z.��P��d��o���M��l����~���d�T1L8�K��9q�/st��y�P3����|�$��?_�h�ۯBU�9߸'��3�����,�/T?��	��z��
L��4'Ir)�m����2�Yp�����iӦ�k���ڢ1�<�j�b�ɜd�~S��9��o2�l��B
�Q�.~�I}'�g,�,��Aa�����[bh1��&�J�w�k��:��[��'#�4��XTIV�`�}E3���O���wb�G22uq.��H��-%h]ʨ[�7��A�r�-�Dmr�p���o��A=��&�m���i����f���'��e%��2[�5>*�O>���s�`�z��{5)k�J��1��ݞ�W'���qV7~��uso�d�C/~	��2�oy�E�,jl�w���rrS��p����O;�gJ$�|�����$$�҉�\�,��8�H7Y��V�8:�	��<�Dz�b�����/2H\�� ��~��<���J�y 1�އ���u�Uns�|'����ջ�e�����.�/�������[�ٱ�c�Dd?����B�Q��|bW�#' �?�<_l�$��)��V�餋��,n˹����K��8�rY^/�r��I%���+?d[ʈ}*�}N��>���mU�up_�$0�k�&~�mxT+<�'�ԡu�^'����#�������j�a1[6�#�^���S�cpi�Z�e�q�ve�k@���&����� ��ެѠ�(-#�]�z�k�G�;̈�@�Z �p��E! p�� ��l�g�a��<"�������%T 7��-�>1��/o�Vm	>��s�+N2����؝64��%�D�5hTy��!|��d�~����C÷7#�	�ȫ��bM 8�A�rɲ)��0��M�4o�8��X��W�X�4���H՗�:�����)w�#�Ƃ���3ե!CEX��f�z��&�����x��8�5�ǳ&�Cy�a��'�[����G��.��i�%lEƶ\I���"���H����iK���}�:o(��LR�s(7�5C�ծ�C�(b�BopEL���~��F�(ŀl�o�W'-L{d���jl���%$�0(0\���	���L������Uǜ���]�����;<{���w7����Z�*W��2oh\�_Om����(���Ğ(h��r��v#����}Yۼ���yR�A�,��"ȁ����bY�;@�o� <��ޱA�$n��˓��Y�\��'I�s�$,f���J�>G�=�^Ҁz�P�G��� �Þue�����|�b�4�ʰ��[6�"�A3�*�RN��D�Ⱦ�sLC�ǹ4lx9%gU3�֒��1  V�?���؋0��n�+��*���i�Q -,�<`�kF���0�/7��������ӊ�LW±�?�`���ں�d��:�O���#�l���ަx�5:S>9_��,c�2�d�,k��?w�S��+���d[dQ͕��E.}b�F�.����p��k�U
�р^����쑖��R��{���9�l~�F�����=Ԓ����������&5~��k���e5i۱՝-3�n�W�C���ŉ�2GoV��L���!��������Y��P'�{g
����U�m=���U�o�.��g�.�CHk���Sb��S}�X�N:�N�MƉ�z^�p�2����۫ٶJ���;·�wU�V�6���P��do�u��E4��	�ӧyO�,��I���m���E�Y����y���M6ڐpz$�V�{�)�f3i �@U��7���#��r�ۣB�~����h؉{���t!VQ�~ݻ�8��v�?s�I��QT{�ܬ���C�d'���Ƿ��!��?^+�>�.I�.�1ũp=��t�Q���*ߑP:v��]E3���&ʃce���D����"��~�%����"��\�#��4aؼ�푑�����T�@{�}D�	�X@+�7�HC�f�cR&cG��rJLC�����&T0��-�b��=�K�����%�
��3z��Y�h�{%zK�a�5ul{(_
��EŞO���e`�y�-G�$b�#�ۏ3�2�Y�M�N�g+)�[��m�"������[*�%��s|����&!�66<m�\����G�:ky�	����VC~�h�Zi�X �G_G����n���2�5��v{r�v�>z���H�g�x:g�� |(��A�iO�����/�,l���Uթ�9�9��{��})~�{�0'6h��M� @P���������%E~m)���k����;1ů�@�g.�#$|L��ׁ�U���U��P��"�+�$�x�
�D��rA�T� Q�j*���.�vn�qFy��=��:�oP���#�ؐ�'sjɉ��>�ъ_|�3�C��,-��qq��g����;�wT���;�h ��^&�^.����j3"?R�P6�xT��x)�vU�|�T�j�rQ� 
��+QzhA�l�̢&:���\�s۠��f�Aj�����q3*�p�jŞy�sS�fG�8�[ڨ�Y�'��_alx�c.�#"'g'��Օ�a�{�j��S��q�?!��rn�Z�P���,C�^�tm&�{��x���|>�k�-���k�Qe,D��=�­� ���y��*���9?�,mLz��r�ŉ�F(�ssƚO����F���Ҥ�����M��G��������M�㭠%��E*!�~\�׳�ٛ���@��ܝ�О:�Y��f{�r>��W�C�p���
��7�Հ"Sqn*�C��Rd�Ao㣝��5ߴ���FO��$�?�����e|dkƷ��\:���եg��}ͼL�D&�^$�eV�U��/�<Q ����1��(���,)L`�1w�
��}���&ܔ�*ʻ���6W�LS�L�ӛhʭ"x�z �,���P�����U�	��ߨk��]=�� 6�̼g�bΥv�%Z������x��y<������>��������Xe*���k��G���7�������M��K�y�ω��z�.kn�_�qA<���l����8��4ɛ�h�%sx_H}d�3������U�Ș�g�`_ά���G}3`��ꪃ�ބ��(b�H����ԑ�玄���>�W!@r����k�`�I D,�b�!��05F&�@�it�� �;l�	�r���4�-+N��+W�����Q�Q�=�-%�d���>�tjߙZ5M���u'<>�C��ƾ��$�?K���oO�"Yqq������� �ũ�C���� <LD������a�EW�L�$M<��̋
T��Ē���/8ʤI�0��2�˶���P�ޢ��۷����*��+f��IE��U����2��ب5ˢ���1��8���`t�� |���[�ۮ���: �5�9�h:jI�ت�f��`��`%?�Zz��U�!�7������֦����7&�=�i��j"8w 3UlEDl���o}c��M�RW��c1�/�jtm���˄҈���1�٨�zm
�N����q�w���ؠ�y�s�Bˢ��^�\�J�F�ҸT�W!2M���7N�<�L����>PJ�q�������:�r�d�>��^$i����%�?B�W�H}X%��!�:u��I�wD�6��� JG�v0�������kN�b'�ﱵ�Oʔb�%���=��cY�~�R�l��@B�Z��%�2�]�M���a�gQt���)���`�b���uLtջ9��<'g��i��6zȹ3b��T�˩:x
�ގ�%����}�:D�&Μ�]�\�~SH�1c�p�y6G]%�3���r�oÇ�<�D���!rLV�������� C%�P��R�3��	L��=�=�Y2 V�S���b�n'q|��4���IWך���X�s+���uką��v�b�[K�c҄YE�R�d=,e����l7�bs��:�i[���WޟB��Gb=_�<[�`�  t�����Y���R�H�៳,o-H|�NxM�t4�}Us�	k�q�E��������1 %��)�������X9�)F�Q"�8�-�`l�����CK����Բ�O�<QdX(���20fd1 � �w']O�/��H�;��� ���Ys���c[~��tBiR�E[ �<x��\"�~`_L� ���4��kZj����k[6���KhJQ�#�\ޘx���G��tHs����@�z)��jzO����p���"e��mK
�Fńݜ�r�چ��wqə��:�[{g~6'Y�֐"�����һ�m�Hɟ4<���(
. Ղ��}�m�*�h9����^gwMvE!s+�G�]&c�JE?�B�c ������5E��0���Ti׫ircqb��;}��L2ʈ�\���Eye�L�p-�� D'wC�o���G�1u�䙭����n��߰6�Q�٘���.0�7Z����5(X�9��#�DZ9��]2�ةz:������H�j���t�:��ɧz��m�g.�4��M���9ٹ�����y+�E��b�0|�O�`�clP�b̄O�e��	"a�y?S��$�VdV�RM�יvsn�E(�C�'�+�b����R:���nas�ݑ���G�˨�Z"e���SƧa��@߿rHsO%UN�.��U~��0�=��̴098mr���h=��/��v�����-��WgC��5����ӽ��nfD˘c�#%;L�U\�� ������D��HҘ�	�X"����7����#?M���"�>��r	]圦�&	=�4�q��x�*[r���m�}XJ�=�<eNcA�9��mZ1{0Z�5V�M�+n͡ I�=�*팛_�S��`�ȴj��,3�/��8K�#�%n�s�WC�
�ҭ�Z�GԄ�l���(��7���N��u�����Y�k�~�1�3�Ϸx��ã+8eE�@�F�K��R?7*���K> p[�חط���٬F#|8*�E:� +�:�s�ܛ����W��O�2����#��+��L>�2+��)ȫ�
��AO/k[�,ʿ7
���[���j[(��}�9���~"󊁰�JB>�M��`��j�>�vߗ��'떍:Ԯ��JУ�ߣ�^�ظ��S��}�����}�C4�`n=���L9�������g��P3�>��Ě��䠑ڪ�LS�P�|Y���ﾗ�l���'X�Kt��m�9��%��I�q7��3K�cQ�����1Iy��+>^��t��fy�ڠ����Z�z��j��߿[z�޾�UG/CXZ�n�a���J��c#���+�
2�%�fgO?�Bo|78_����V�Ā;o��%�wȺ2��� wb3��0�l{��M�R���$ @zǗ8�0.-~O2��8?�� DT�3���Bs�����h��3R��sLu�t��-x�n�a�G��L�8�?���P��L@��v����r�w�Z�|��c5���a�K���UCw��;X�A��^���JAM/�����*��8f�YQ�
j>a�n�L����,v���m�r��ְ޾k'x��T��U�3X�J�Ŝ�Ɩ��ȯ^�w������l�&΄�F�����e.]���Z$p��%H)�U�PY�#���w���������9(̬ܫ�D[P�v�%ص���*Ey��\�T�������J��L�E���u�b����c{a-~pˑ���hK0&���l�k��d�3�`�qO��on�ʍ)�Xs��wRc$K��Ç��J?ʋV���߾G�~6:x^�����ж���H�p��C���jU�9W/ E?��%~��
#�����W�n�J��_�����\n�������l����U�*�eE�Ԛ���l�.�� .�����8��� ԧ����4���s��pE{I�����sy�T/]G�&�V���>�����׊3t�|؋N�ٮ�[��\H\�䚲���=�G���5i�/&�N�=wT޻c��@�!#M�i]��]BE5jR�=+Ek��	A$2��f|�=�{^<�~c�`�X��}�'-:�/�}��a�Z��E���{�����ˏ*kxc�#��%p W�4F�K�B[C���p$�}S��Q�5\��i�=;o�.�bfc8C�D
q.�����B���:���U�C�J��FgH �[j�RǺ�Ϋ�gs����z�8�}�D��Y$��
�D��o:>va�'��r��V��!E&٣j�"�O9�b_�إ�W?��B銁s�"�-Lx���̆5(FXc�_ �c܍E�?#��}}��i�)f�~}�F�eC,���.�:�Eqyt!�W��^`"&_:�N���*)0����s��.E���(�g��{MI>7������p&Hq|	��Ʒ�/d�&�v�b��hBe�����'J$q��tHm�}X�}H��n���"?�Vx�,a�4�e{�"��<ba��=���S�)AW^i�Ɖ�}U��HH<F��� BڌX�'��q��ŀ��
�]/�´�JEp��V1yK4o���y[?H��3�[���<iK��3�4MP-���Ŷ���~�R]@�
�2�S7}6*Z�g9>�\>M^�>H->z2Pxk'ܨ�Q�h<�"�,=`�����d�Kڷ�Ln� Է�E� �h���00��r���
z<C�vP�ee�����o��r�+�i��`�UjD�B��Xs�7~mq���-�siXij4�d�}�������T�Tov�#���h�|:&>+�~�B�ŧp��Z��� 4�TבZ����bX�|U|]d�� XP����eM�y�6ob�u�q�	�Y����ɘ�}��i�_�v3�8F�P׸���X+�I�%Ed��Om�;��U��I��
�:Tp�>8xMW�^�G3,���|ˌ�R|���Hߺ��F92f}��٧C�թ�}����V�R���M+�˚I�J�_���9	�<����C�η=}ȋ.GU��K���R�G�}� Q����2+_�CWIu��i��'��!X��Vڢ�����[=ʠF�9Jy���՝
95]$0"v5��q��E٭hdn� ڦaZ
Wj~0��@Ɖa+��3�C����[J�;�`���ڪ�Py��O6�)��	"Ҍ�x5�G�����
�h'ɡ���%�'?C4\"�R�S��K$<ٻ���cq$��y�Fٚ��z&{����I����T�Tz�ܵ=r`����3*7���ܱv'��M �Lя����m"EA�v��6� �W��O����Ôy @�q��*����R,�Xݗ��:\��	Gw��.�Ԥ����]"���N�eb��T��I��>v�%�̞��->8ߺ\�1�S8����5�À���	?e4�3]������u�
H��k�R�@���)��t���1ˡ�q<� s�;O|J��H{�F��r7y"�{3\���+�e�+Y�y��BﻟM�t��:[��#'&�1�c�f�/W���3�2n�06*6ëta�_�5�ڹ?(�:"���EK�`��  a�u�E���X�%�UG~�"�j"�:�j�ԥ�X?"�����W)���H -�|�3ٺDAWLm�*���?������9����c�~RT���#�᝹l5d���L	a� �����N�"g����-��QP"�Ӣ'�V�1����O�80$p�3�p'��MbՎ�$M���;�'C��B�=g�P7��)��H~��PK�����?�jL����\_��Ӟko�k���f���LAkt�O{\"�o�����y�+u���o��g�ec��I���4��@ힰZ���x�F�ی����F�Cd�Tl�0h'�D�Qe\�|j���5P�w�?Ne�٢�$j]��GTȅ�Y�<��u�PH�U�j%�hU���
����ZťFFGP-�M"×��p��d���:N<]cK��o�MF�4�[.�;�-K�6[��
�1�<�[P����r��1��������iA�\�fd��tEs�s�ʴ�`,�O�@f��n!F.b�KO����fblpM���G��\hy'Ȯy6�DM�)N�u��I}�ɂ�Ɗ�{�ZX�h��}�@�Nۥ�* ɐ���̾#�a�W'X�L�I�= ���W�;�q���䏘�Q
��AAjwm��^*�%���:�ӏ��ĨO��0~~Xc���e�<��%���':�j���Ο�y@>f::L��H�t�~���X���G��:�G?l�;N]�*@�z�w�}����o�Ǵ����!���l|�{w �X��g���@�{F�M�Q���c�`��oYK����~��H8V�6�Š˳GexB�V�4�\�*>ى�9��U��'*�'��[3�#<�p��FI��S`� �Zt��?0W�nzw��ؐd�-���f`��3��N;Ȭ5���l7�q��A�����Ӟb�2i�U3���͆΅��J�
�#X��r.u��� �K]E���GJ������`�탑�ݴ��*���֡��dJ\i��Ǝ8{�
����"����m�ȉ_vS` Eo�g1\�����F�LB������9`(Nu�fA畮$�ƕf��[0 6�����[���?������ �﫿�!h��u��z�
2�'�����s�2qJL�9Ӹ����#-;���4�B�#7���ݕ�?v�cUe��vG{"y���M�si��U�A01������2�g�7�	�;�:�I�|:��;ƿ����}�� ;U�Z����l.�7vG�5�>�����X�<�����f��q��i�; o_XM����|>����v?�˗ࣞV��9���-�6Ѩ�"k�����H�$*<�N��p8�U���_Q���(��M�����EЇ�@�%�������'h���̈6 !��&�Ԇ'��9�s3䘆����H��S"p	���h��H���G�*Qf�|� C��X:,�� �c��H-GupNs�9�������<�Q�h��^>d�Ӗ%�:*�B�Z.��[�I�R��萎P5m<��(m^i��g ��[o�-�(�ۆ系��F_�gnD����[��N:y ��֌��i�w�ڔ����J�U=|�nD�|�_$��G0�NK�k��sT��L�C�!yA&�h��bP�z�����Ĭ�\�Beٿl�^��X���b^�X�x�!�#��C�ҍ���䂞��X��3��5B@�s������&����q2���`K���fGE�sl��NJ�)��\KS��H�w|Y$���5��DלBf�Eh�EaS�,!�{�١F�D�Xb��AbS�%T2�P�<U��q��]��PQ�/�|���Xw��n��j�8T�Hg�T��d�3\�y4�ǥ���F�1�A�7������-9# z��C�Q��56e���1�� ��#�C�>4ow�0���M�'c�߇�>Tg�kE.�Ի�꣌��q;0>A�n������4o�ԋ���o�XڇR��҂��2��
*�oN# h�"��3�6�J*���� 7`7�?�=W�Iۥ����%G:W0EA6lҝϼ���q̕�G���8$���8���bSP6[��GH�)�4a[r�,�	�]_6��0��rՒx����9�)aL�5X-�d�zԕS�OЁ��#�`���������9����G:W��{�u<[���d���i��?��:�iI� �m[ �<^;=��ƨ��B��#�0ٹr-(�F�A�D�(i�퍉�6�5�2��,S�x���Q��KU[��sJĆ\FmB��Y�<�Tʎ��T�X�/�-;�?D-���#F������VIe1�F_�5)�p���@Dvr�K��sE0u癕����6ۆ[NH�Y+�� �L�@���)UWH�~����	Е���;��-��f�1S�[1}@V��d�B�U�\/z��G������5��W'4��G~8;gTI'��%@�֐Zǖ7⢞���c\��_�o��f��T�A�FS�_b@{=p�(�D��2�=Q����d���?�Ce]�w�Ќj�,g@�^�x�d<�k�5�/@%��<L*;F��m�e�:=jc��tu�t(�ך�P��<i�"�S�хž�s���Cm��'=(��7P?�["��Mp�q�g^��acr�հ5�d�fg�/�e���c�ѓk�L��K���߶~?[�վM��4=�T��ĉ�*�;��s�p��N:@��sy9��T}_�F�Ω2j�A��|iM��I9�g��m?G���(���L�f"�f����gB�3c�#�+?�}B5���C�2?�tE������Ng��t@3]N�'a�0���ߖ{�$�+��4u�:�P�)����-��<���_�u(�պ!�ŤT�&�HҬ��!�>�<	�A�^3a��ԓޯ?g�TF,��� � $h�R���?\���a��� P�k\�^=͕�ǰ��Ӳ`V��%"MI��b�<���8�*p�~㒴Z��o\W�>��]|��FR�{$�pG�P�(vq�?7EEOTЅm��3>�����Qkg�u�����J�<���NyXVD	\�\��oXi�wU���l��H����4��8;"�bAl�w]���uj]Os8��u�18�l垙�z�W��CO�&�P}��ǻ�8#���H��	oE|+r;m�oz2y����L�����-"�YZs���H�O١�n�9��v>��7���9�,�z�5s�q
�+��b�*�)���JU�FWXe������|�k7��ف.�2w�@s���rC^��������js����|*W��3v͑::;������m�a`X�%����RdINk�<���-E�;k?�/�Ou�+�+w��	��5�|2T�T���Sq����w�2�Vi��3�^r��VU|�6}�g=b�����ꏃ����eT<R��;"{��=<U��sʲ�k.�kzap���W�D�����*k�7���������5�sἱ��K�"E�:_�Y왿 A�kQ�nC3�0�|Hq3{�� B؅��r��ͬ�H,�K�]m�2�{ݠ�y�"��ǒ6�=��SS�$Q0�,d��p�[n^�Y�E�2��c�ӳ(�`7;J���<���y�I������ptV���>ѳPQ��� ,q�a1�!���z#dR'��1��Y�9uދ�� ��xd^�1�Ǖ̫��9���=YM�J{��]a�e�~LDX���?p4.p#����E�>4�=���o5����Y�}��8^��?���d S9�ܤ�{��uw����̨5� �WիFF#��	������͸Ś2���x?
?�7!3�܎%r��>��R6�rn����3������H}W-2N$��z����eG��J)�~&���W1�g��Z&��m��}x�w�,\yp�Go��$I�C����D�=HԚ���Ҽ$���$���QV���dt��5~���¼���A��lSF��Ik�`�?�v��C�Iڧ'r�&����7� x��f�h������tQ�'�-�n'sݰ0�W�=�c�C1<�a�Q��)ʄ�Mr�|���͛�(O���3�ù���7�4iG�7�2P}� �쑀���Zb�C*���Z�h�cu��:��Gț*�����<�#�b�Ă%g�j�	��c�RB��"��X�N��]١K @aG����V9���ӡ����?\fiC.`$������p2)��M�s�4[��,UZ�~X��M���<���/��}Q�I����h-:���Z�Ż�~����C�F��Yk��奚Q,Z��pf�aH-\��ܨ �ݺ o:gς]o�W���>�K5S��sn���DoN�C�������L���M1����s6mucğ�,#���;�slegR��3it�u��̵|�#�r��u�)�0�&���s�Uպ���s����P2ˠ8$��*�NJCɒ9�i$��_�S6��q��p�9K�6�{a7��4D[珱���|��g^���5㳁o�'H��$�f{pa����?l~��nôS*Bm�j��+�g���;�YN����8hx����/
�UϲúKϋ���,�n�M��kcc�})7��x+Q�-��b�mX��Jm}�Ưv�o7�Y�p�����hQ� �Gߵ�����i
�G�X���T_�z���l�ӦMW⥸�0���8`Tݢ�S�:�V6���9��\��F8^"ګ���:໌5�?U�:�ƌ- C��q�$���$��4j{?����-�hΪ�� ]'3�k�hP��T��~x��Gi�De�O`��7I��0\��[t{I��p�a���ϻ���Fdf���(���7V�b!�=t��=��K�Ĵ!����sU��3��|����)1�5'��9!�^����
���SslI-ڍ�؎ź��"��������۰��r�`�
=H�1�b���O��&I�:�j�7V�@{�Y:�a�4�H�W�X�����Um~�����S#�QfL���҃���Lc�6S�w�G�`��嫿0�8�ۢp��H����>t�`Io��R'�运��7���jW�Pa�Bb��G�8d;
3��o6��l�
h�o�\߸�H%�F��j2��YE��c��H���+�Ѷy�%�4Kg*k��T�5�28�B��ٶ��	ܛxvL#w�������Ѓ:h�"�����'�|�텫1b�^/�����g�Y����Vr͡�	�9�O��L��D�Bw��F�$f���N7�X/ŵ�7=y9r�#�����S�Aب�~V�pO��$%��F�}0�"�Q!Ñp�/��9W	R���0xN*�!�I�_��劬sy'��fW�Z�V;��G\�Ț�pR�	��&3�ϼk���)���s�\���@EvrdU�@���p~�v�-�'%�Z�@m<aW����SoA{<� �R<^J�OO���{�sׯV�F���z!��D�hS0����s�'��+�̻bLOL�E�N�4�<����%�1�? �#��B��Q�D����4������:�z?���0�Ŗ`����z���|�;!t\���?��D�:��̈́��L�.�&h��ZU,�K�]�S� X+zi&A�;b;��& G�y�������,�J�D�Vl�(�wg�V�|��;�%ԑ�C�g�jv�����F΂pH��w�ު!n���xA�8AZ�� �L��I@(ce �ՆN�^���d��|[�j�%�|	��̼�:ե���A�4�ah�D3!�͉^|�$'кw�W/-�G��_F�=�Z�ؘ7�|�d�.�v�f���T���$�� E����	�#��T�[ѓ�fCr�Y���6�Bp>o��Y�zr�F�1��z�"4geGeZ�{�О"<=�_�)��a�dD����e"�����O�u)^�;���TA��*��,���K>�WQ͑(���� ޓ4S��}���*Ҕ�����=�X�^��&z̑���	y�q�.O.Z�oɐ��+z�~�y��_�:a��AbX�^+�6M�H'�;��xHkc�{��$�� �hZ��J=ނ.]�U:���K��c���I�Z�ں��Pg�?m�Ȭ���w��@Sɛ��b�&1�8�Q�]\����������H�n�"�!��Gc�4�y���[Y���S�L�:*�%�M?���V�[~��a<�#�E�����U��Q�799Q�>�F�:�z����`���zQ��L���c�汙�����P������[��_ͩ�+U*ȉȱ�Rsr�
�(�I�}��[��y}B����UoM�]S��2׏�R��Lҙ��2����VO!j�IM ��od�a�La�lH���=�=�Y�+��ӍK���T�_1�wc6���7/�y
7���,��s ��\�El#��5��ihWJ3�@��H������k	KE���š�=܆ħ
{ޣs�^��a��Wh�w��Q���Z��j�J�6��@!�x�l@VS?XCN7�i$�a �Soh+�h��Yk�#9�P�vR���w9����(��7����f`:4���}�~�i>��9�o�ςy�ֆ�0W�a��Y"��V���!]��(V3}�,�c�=c�1��Nf�K
��ݲ]����.G�P�����ml��2#��ʭ�DM$)<SP��h�x�
cRآ<m׼\�|�M[2��զ��.���Y*//����&��B5R@B�d��~S�$=Wa�58��GP�	jm����9.y�K�p6jPτ~9㙛��#�Na{:�����9S*,(��`f��]�8ݣ�[����=2�$��b ��Q�ys�t�$��`��Ly����hk����T=D<��v�<&�D����?�b4
�|�� )Ya^ ��DṺ����r�@�6聾-�6��"=�?�V�8^'֞(��I�' �D��n+��6�n?����,[ݛ=�mC��7�R������ӨD�>���s؞����w����C6~�@ ���T�]�P�>)�����؆,0�'U��wZ��]�9E�X�6�/f�_sj��H�����&֪Ci���H�d�0[L#�Jfoi�a�Y�����Kh�\�0
2.'�o�	#���y�[����Q^tc��b�%è����y+jA\��˲�o��ҫV����c�';�i+��EEW�{nL��W(Lv�?���.��[��:�ag42I�k�<��k*Iv=�I�#��_�
�
Vu�>j=��a�F�T	^o��PnǱ�ʑ��C}Rf9#V��S
~Gq�D |�$/���@;	�{�-�����g�س8�y�m.�-�S���{�P*+r4r�`:��9�_�� �j�M������Va�S�:W�O�����d�g�`)���8������I�M���c��+H&�gTzB7�O��4�ɺ�	�ƌŀ�]��Hy��`�-�w�H�#��l�~�5�	ў��67�����%�H��=��,�M�9ՍE>kT����[9n/�q����Iϓ������V1��/�,�!�w%q3�\�E@]5nм8��'3[	� i�-H��rX��98qS��s������.={�?�o�w�п͋	u`7J�de�
4j[%�=s�6#��gP��$�!��^N��1���)�y��	�����&I� �}����-~�9���B��t�_�sO�?mh4R"�eVЎa2��J����#ϯP�_� ^��W��F�r�d�}�c�[t�D�܄1�>�(�Q���_s�VCH�P���W�\�k�]��<ڧcB�\/qb*k=�o�L�x11��c�)|h�`��8��>��"c����.ZR9�����rO�	Op��G��k���[�v��#����W@������輞y'S�,��|Me��P��5�h)a���jJ��TS����6�E(>6?�\%ʐ`s���`$ �z�/7Kaw?�4�pG���::�B�[���1���4��H����6*� *��b�~���ؚ�
�#�����pH����@�Cnҙ�e���b�~ �Dg8�my�{7�rD@*Ak��@ ��[ZZ"wo�j^X��טE�fkJ[E��Zg"��(�'�B�e���r��N|��lt���=� +�cP+i��������W��a�̱�����&�Bk���s�\4_�j�U�I�LI.����_�+��
�;�Q�Ӫ������|���6H4:PW���3K�����j���(�M$����U��z���&�SA��R����I|w[g�E��	��W��ߣRx1�����U`��`��,z��!�+!B|,���������>���p�����#���LEJ^���U������ءgF�%{Y�~T+�\џ��eh�a��,u֓5E����M�p�!���4R� +yʚ��i��2(� �$~��A��nfl�m��_�[�G�PtKk)v��(�Q꼩n����O'+�>����'?�����fǦ�p|�M�ӌ��z��e�A�Ҹ��O���Ը�:��w�yU�{��2��+�����6�r����V}��2gu���'�������T��E7��T8�^&��ѣ2��`�#�i�Pt�}��~��>�m6L�n�/s�Z[C ]'�H�1�*�7 ?�f�Ƽ��h\w�.%�~Kq��2��xZ�o���l���tֵC���>Z+�"��M=ڦ��
�u(L3�����.b�֭�<e���X�7e
mpY}�&Ho�2I�B�l4��K�Dr)4Wvz+�����VO�VM�kW�lt��"'��ua{/������$Q��6ӛ��*�+b/S���k#b-��n�tx�ήl�E�����J���ue6���|*����J�ѱ�F����!%Q��j��!�sp���"���L��/��_� ���=-_-��ş���߶���t�:��/�ϯ�ΈܱÎ���w��Z$��W|IdK0�L��M���{��������
�/�a�h��U$?p9��<øgDUh��n{mN-�؇n��^/,�O�3� L�����7�U2�R����/ �#�'#��L?-���U�&Y�8��ruQ��EU�h,w������"
�j���"g�׮�n1��'�00��IK�E%�J�lẋ�}��ڥ��,d�9��V�&}+9�����{�0������l�KݘsOJ�����|[�p�V�UK�N��#e$6Ӛg`*��"��`\ؘ~��jo�ZA��vI�SY.��L8���8�I^P��t ��C-2,��n(��;��de�s��MT����x5�1��l�H-v-M%`�x���P��)2[��ț	9�;F�T]JM��Z1{=:��%a��1��[�ks�'��O�*c�p�q�ʣ�FM�<q���i��s9Y�8��������4L��uu_����rYG����!"�l�)t,-k(��M��N�&�1��|�:|�dL$�Ρ"�x|0���<��b�Z�˜���G��EtP#y^,�Ze:l������G<qҠ��d����i�+����JRф������lyy�j=e{{��1TAkf���q�uUϫtr�s5����N �zRD�RQ�Q[%=��ޑ��k�،/+��
=p%B��ɡ��c�m�Sq����K�¯>"�x��jM��ɚ�w�Ť�Ʊ���<9�ϛ��~��&(� x�����G�>��Kذ,1�J�^S���2lR��%�Q����Z�/D)�⺊�BI�.���+)V��׳��e&$W+�8ES:�=(~����	��r+�5' ����ϩ:�s��C#�F�[���F�Bv��m� <Ca�Ge��HWV�"��-���SKbt2w��|�M�E���_(���@�q������yޘL�"
됢���,�.{3�v1g�\�~�dh�����GZB�V�*X9gz��=�&���T�%#�;���cM����[O�.��.�*s�v��z��+"�δ�_����*f�z�X�8�����\��1������j�(^e��A4}��ݷ�)�(%sCP���:�߻�C'&��bs`���U|����vyv!��y�e �~đ�F�ڭ���$��e���Uz ��"���	X�8�=��ڕ��7��*Yе�z�Mnd�\M�������?�?��Y�ψP�Ԟ(��%Į�ձ]e^�'�����H���+i�V��3�F�[���ȝ�u�U��>Ba��[�/(eW�}�w��_d�!HB���J���ߣު��I�U�t�0B�AsQs�P����V�B�J�4)/�%8����[o;O�q��k@#����I�۝�Qe|����d�ڧsR74����g�*��c36I�� 9� t]mBq3��_��Wuo6�Nq>����V�L%�_IY��aÂ�w)�)��b<=j?��=�~�{�����k�Q�� �;57��M���m3	��8�}�+�H�� +��w{h�~�u�.c���ψtћ�Y����}��W�\U�`��?�4����f����`_����L�lʁ$�%:(��VC�'�7��?�<��:~3����0�e@��k��!��1[�����
��E@��<�����`��K��@�w4���FҎw�����5��n�"�*�'�.�nY��)i�;��s}��F�3�AK+E�+�s�XF�d�I-�.z��9+Ab<O�x�ny���C`�%Χ����h�⛁<�S��n�}w����ġK��I��Ș#��|l��͸��h	�r��ȏ���s	�
��C��;���p�U�1�	��n�^a� t�A@֌B1��OJ\#��11�ק:c4J�O��@�/�eY�����	�"�$;�)���W&�̵R�Rش�Q캥E���D�.5�M���C�A$7��M��D!�/�"0�>F�Z�K<�����
9�E٧Y%F`E��wF�O�`A_����J}�,t�&���-�S@Z���̃�U%�����5��9c�,:�۳-[w���z�f4c[�B!�H���dnVb�I�:L�����]�i��#*��;���1p�޴Ѯ��|_��s��E�8�v��؁a�=vf�"k�tZM�����c���_���+�e;�Cxf2zx��G�tfvu�%qi��h�eZ+&&�!��ٮ(� ����
y]_��m̥��?jE�,X�'(���'�>[���N}l5�;&D��� [`z1�%�جs�c�쬶�CZ��GWg����cx�(�ő Ѡ9����n_ �"��x���F��8W�i�B%�Y7X�˧��~��D��.�O ,�l��/!n�J�� OVx�/�hBʜ�i�2��� 0�r`�d��<��[g(�R��J�T�`A��y�+����P13�,���#�F�����T�t�F/H�z#�X��6��N�f(L���ޫ����H�l4VZ��D��O�*`Z��Zt]��L�W"������z��4D>�B�n�Q��J��x��D�*�Z�D����ׇaVdj��Ö+�пN�G���z����bsI����/�*B��y�;� Y�����^��w�
��X��"J�/@k�I$ld�aK�$�/޵j6��A �=�v��.  �k}=_}QVN?�&i�d�l���CnQVM''��'%�ޢ�e�\��1�����2}�>�81:�>�����C����I\�HY�>������&p9�1	��0u�m%ل:`��N@%L�*1VK".��L�!t��h���]z�Ϳs�4���.o#�#=ҩ��P�yI0N.m�j���� �{};{%\+e���͠6f�>��4(W6�V6wF��a/_��'ҁ]�)�H���aN�rҶ��pى$���e)Y�y�o�/Jy
eC��;�&�:���{�� ���M �t�Y��&�"��E�/�^��9H���'�b]�3ׅ��t,eF��e_U�|BBsS��Z���RJ��^N����L27�UW�6�_�bXpƀ=�@+�ܚ�Jۦ[�1��ALD}'&�_�-��J�vH�ٜ��
�=�f��<ĥD���K��zM�q�e]f��͡�5%˅�m���#�4��kS�}���w=6���UZ�CC����B����OZ<U�)�#x������@�]A�z�>���ʇ���?�T.gsQ��������)�>iC�#������4�O��!�9<�vQ�+�x��������GƬ��S��/��y�t��-��^��oκ<�OQ��b������3n͞�a��&r�Ƥ"�[%^鸱��л��>~q5	:������)�,W����P����6��8��I��'��,�r�E�K�&g@��G;�Z�m96ȵA�3�����E�-�L,ܝ{|J4䵝�Î}���}~��]��Ϟ'��@��Ҝ$�܄��O6eTw�G	�&��W���VD��$G���_�^�L�����C�`�d0�f���J� �ډIئ�X���9�ZÈy�J�\�r��4�{���Ӕȑ����vT)�ӝ7����N����z��y����~��M��� s����I)d'�d6%nޱ�����%�&�|-��ŉ#/Y��x�߫��Κ��c��Ј:~3�4�Q)�9oq��Ձ=h=�^6���6�>��+Vru�7����	��������~�8�+}�9�!�Nn%5dB)�k� K�'���X{,^��⇀��̮%��W2L:ڃ`V�G�=��Ɓ2���rG�QƼ��p��k?�R�8�ļNcf�;T>�wu�V��Az�ml  E:=:��h�����\u��
J�˖�"2ຏ�*s���C�M�b-SD���W�ݏǐ�g6e��'/��IJk{~t�QG���S�[�Thᡖ �޺����b�vtZ��>�n�:̊�b3cɌ	�e���PC��¡xuC�[��/I'�&�ߏ�+�1��$������Q����⠲�°%�V���c��ty��2�B,D�%�q��.�
]w�N
��jLA�4Q��nמEƐ@��XMGM厷ޕF��k���$FS�sa�/CzJQ��v���8qf<G�_,�)��gfa�uFW�V��/xV�r�R��F_���x�i�^�Nj6d�~�c�GH�9x��0�2�q��vך�E<�ۤ/&!�騔&V���
�)q�]>��6�����a��Ѧ���nc��T�ϧwB�*X|��/at��J�T�n�����ʣ����;e�4�r��k���	�UɭYB8IJ��B��@ x�q��l���aRWʴIqsU�<R 䍇��N�]����n�g!�Cȉ8�8�������܉q7����ع�s�Fi�1���-'A�t�mO�*�xLj��+�����5������}�O�|�#����f�l��Pl�'�'�J��z��q|@��(�<�4���n�=B6wvnMS��_ 7�M�AnD�8��І��*зQ���>�V���eB8x�
>��}|ȃ}�v�2^c$�q�;� _���V%�(.� ��w#\�x�������(������N;Rٞ��o��M^���A0�h�<Wfb����B��<�;�ڪ,Y�gi��7	�D��ę�%��f~+KR���T�J��=�ȴpN���	|��֎�d&`�����M�����u��i� 
���c��QA���H%�3�����_�t�ӭ�H"���~���'T)�!n��1���L�_t�b�ա(��?|]�F��Vb��ѐ7h��R�� ��� R���p��nJs`�M�W4�q��S�蔨�o�U��@S�9d�����nB�=сr�e%���"(��`�p�]q2O�n�O�a��R���*x��9�ϐj�q�Vń���'X�I?$��F���^��}��c�']⫚�*�gz�y�Ùf`�2m�3`�*YK�X��&�(�������#|'=��n�u��&�����䗸��΁gQv��{�딀�*����>���o���'�	uE�^�Rp ��u�:�o@�p��d�v�9?&�2U��)wP�Ӥ��>L�Lf؄ʄn\�:B��)PnR�ˆN:W�BT}��N