`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mTXDlrbsfm6XwYxeaYSzzYNJiAd2CiSD2GfaVBL8XqTciSZ0kR4cc8uA83ouba4t
bK6fCrVuPExx2GYdCabmM6QSHwNeMtk6T+G5PoimtrNrbFVmiq8rF8RmSAx+5073
abFbZ8Y9PskanidA4CBfMYCdb7WHMMeiOvxiuxexQkI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10944)
zqTe/uptpDo4cXHDxfFi3g80HEVzAmHigqzRLjNEtWSPvRbA16KMTPYZV8xXQPx5
HXuoqRt5hxSNVHeQhad4vAGR7yHWdDa2aRpP2s7AMJF9HUHHzB5QNV+ZbHm95b1G
5KJEHFYoTmEQaMgsphnMfYtwOl794+BNZqEtAgpJjVlM+sGk8WSoWRCcfdDkOnLM
QMMo5WhHyTx4vwAhCitep5Fmf8qlxcWPqQ2LIo5ufMGRk5X0/tceZXgOQ2QOYqKA
Wr7bK5SaiTtZyFsIExM9vSC3e0M8ojhI3lhB0/9i/jmaTffMU6nhkdzNJvE7wem0
X8nIRRBY4f0q7S2Xedkj4Czw+cnQMK7Ij/2t+TLk+MrlHnVuIqHc3twdpbeIF8dB
iXxVpQK1PI3z4+/8oZnPzr7RsgDvw5zIKoA17KvF87kg/a+16pWlVEcf4jyWiPJw
6RjtV5zUjh/Jaw/tslXKjrNHX8BVLFNelVWFufOXb+uCV5PPYGGXiJVTMjvOp9+l
kO6aZnia8kzodl+hbc24ZyOjt+uRLoiz74QK2q9M3+FPBSbhQv0It2eFv0wyEWp3
KiAIkRq5cBocT3RvKg2koC9IOcXUYnnikRmrvN9R/minvFA0OXUhVjxK+8Z1CPG5
gYI0oR5a+6ZX+HhQ4fq3CrqNQgDQz4KSSF37Dc40pH3lS2lWHtXHy4OpJwR6okDY
LRKfuquNUlC4Tf32DjmDJGgoB8/kCacBU512Jz66lqwcOMOsiBLaZttRpqaVVmKh
KA9pheT6gY54V7kMSp+nLSumHGWTTilYhAdVfmacg14TfCBCu4IbZF7ZP1gdEV31
kraHWgGYNV3Gfz7HDmkfBayyB5vSmQSh9+XqLc7msObJ9SET/jPmnn258e6N7tQX
rMmD9VyMU3UmMa7i3tiChfQKyMAh8SQdCDwriIeFYVG+eIBQHWoMvzDrINk8rXBl
KWDzVrtJv/X2M/GuYz3TMqV6R6WE1BN7QNum1luP5CrTS0XAAUQgxscvzzubztyW
WGjCc+wL1Hb9mxZNUAA42WqGLd25diQirr/TBUYcQsGjiW1HsoeeQHLQ2FX0bGOk
1pM0P7e9ZANYepJ8+ef9zrJG/fq7+mGCKhoWfwEN9PkZNdviWnw1WaLCP25np+hT
bbmHOss0jsmM6Gpkc2W6xLPsqRrtoyG00E/fp2GZjXedxnM6PE/7MXGWi8qy7E9y
rItmg0T+zbDifrQzbMtSzRCFVt5iC7yq3McWm/X8znmjMU7ugyTTxnz5qBNE0S9h
Lc/tF0mBmWGRdzn/C6x9zuEbOr1d0DyCRqDuwwMJ5Dm/4WJ+T8X9yhhLXXSYqXXx
0Q6LKuVQwSNDd+QtEa+lZPri/1Hl0jAl+MOSbOhYHz39G9YNe4RNPw2IXYk8M5Sk
yrhyhx6o/3iJE6vRM/t/7TdQhC2f4BZck6Ljj26sR8VBKmL+5QMQfKKaQ22D0cDa
T2Sry4cNyhZ8gJYR/mbukybL6+Yjqjm2Kj4/RWXXyaZmEwu9k1VKOxGKIS8qC3sY
lah77TX1strnTJlpAJWp4lW7Bk7Ri1JB27WgALugf1wsOVjdN1aUJlZH5YICs/D6
9QdDIATjjRkNuimtn9s82yVjZ+xd/+X1YSMMkN0qo4xCdIx6Adk3mIj+HSgOgPOz
utVHm4om9T/JUP5IRoEJVVEEvhyv0gySUrBfmS0SXGVnrlZ5ABJcrmzsDETfbY4E
22uvwwaTOdqG5EgfrJN43rUL0Fddc87TbaJy3gSK7fGLDccad+ODS2HOqap+a3Rx
fS0SEi450WsetCyxjcMhlk7fq+MqMBapRKsv9cqyGdhdI7BrVw9qDclvV8wSoKgp
TBjUcwSN618t33vWEmROXqzDet4ZT/3h87TQ8MEkxEsnIypaEVS/YjKoB4mpk7xI
Rwba5PHI1gJUqdN2MhYI080xEDRZ+brNwGVMYppKiuUjGYURpQJv937ZreqDGNof
oNZjnWM5yDf7efIyYDuy6iNS6zJLT+YfRkP+ohTlkFACd6YbHGZjyIGvjtdBQ/aR
kTH7xBHadMGFRIR5l0y/F32fE5ewDKT7v78L/L+QY3KtV0EM+4+E5fR51ak62SlL
VM7tmeTOocme8jJ14To97U9LReiyg3yPDbfGMSvSNqJ3rkRbbM+Wih0rweocKzrK
8dsTvfq9QQ22NaXw7lkVIbLefUQdb3j7Li8L2pKe1NmhOQGMVBDzQM3G5SYQhKld
vIrpYvC0SmbdPlbUwqonjdg4KLuCO23kdVC5o7ofiS7BR8hKHaal0DqYC/gGxtFY
YoEM46dRRniL/hAE1TkMp7Aktd2nEco3NA89A9uri8Rhl0V4rOOyLYaTfeyt+3SG
qKp3OV2zNcPN9lMddsucRHboXpLwwaFkXgSujqMHN/wUwTGPRkA+maRjRWgJwPuJ
DIT0ESel5FZEVc91XclU/hg7KrgDf1FAZU26ML42hm93wpf5JzgRBgZoTcbVopf5
mCXm1/G1Mac42t9hhL5yRjRqyzMz0b9AYUxvOlyvaBtgm2Tps+prhz+a9FswZ9dp
ui9WKxW7xpFptzK0yd6Lbev7BwAxgwrZDLcxyh6W3qYmz6mEwEVHUM4L2cWuIiIb
ueOLYere67oChH7pRXARCJTuz9EdHtHPDxYHkVkBstk6JA9vAsMH4BKRPuIE0BSS
JLJSnz5tORjifFbtKpIFsapR+AbPTmo+tHYRJrTZkEYOKqS2ADgwmHpWkjKMjf0T
hlEmeOujsVOqJUkLaMJ/lBQZTdRcR3mfBOZT8oFnbZ4ovuwa4WU3wPKCdnH2YuhF
eJZrPaupdpbG2MCrhUvYe1mj1yTTYwbHnib8tcql03fORDOQtgkMKNZZsJcblW3y
gci0jVqW3bgJgfaRlbMWwGLSvFL+oqX+z46co3c8EHNmSCUrVsQ0WiSLOit3Kl4i
jzYSvhky/YK24x9ayMrNsuOYjXvfhrup+QW+2hxGubOIXB+ht3EF2ohp6m+VVYvA
lLfVHhQELYoCkaVMIVVVP1lGOLis6zH/UI+xSwLbnMDbCrggirBHkxX77c7ZHzQg
izmFYgeddURwp69AmvyVxCYuz+0Zjb/Fdabr6y/V4xFKSzaTK79H21IOuR5bz/YK
0pUDOZqVrns69SAkN1bYTCm/ATj4ci+fSUBGq+btaDKBip2fcJ46uy/oBjrPAeDb
/govnDRrqljZvHhnzaL2WfAbSrAT84/sexzRB21GXeXFG+m2oWJwhIl/HD4r199g
yJd5IZ2hdqVEf2RbUD/Ip3WhiSIf+KcfJkr2W+RwhLHroHYZww9O5kF4VASQVXVB
LtKxb3879FzkSCDMsAyXD5sL+sSnm+8AGW1LplSJp7aof1oSaPIj27uF05v0QrDN
BNJAXk/ICueT7fsfxvgxrLdihdiwdS7wyPWgd1RlocYy8Zqw1Qw8d3n0hbQVDboG
Z3aw6fRjIs41DsbYBZG4PaTbSPKEI4ZutnscSHEA69eLQ+rFhGpBRKbrYTKSnWnw
O+jvzsbTpaIS2Cv7ks3I+P8tB4GRgGsADOh1WsK9dhaEab9G63rsbx/3us+eKRpA
iDlalBFlTorkvXv8DbxyhC9yxyVpGJ+01WKOHdjH5qqvqp28z+1/jMvWuU+YIWjr
+Ae9jtz66YJQUJj4k67KxJqd2kw9RfoMKdS2wqg/DLQw5RvKW4EL8ZGLKfCm1Knf
awadgZdtLSiZNidAqMDu6CeiV1r0BHTz+hEV8JPp938vkTSd5/Xuf8u4r4Uw9z0z
0Qh9r202F2vlyDBhcIxhdqXg8dhqgEq26VHi70XApKLi8eUKJIz2CAACxaURbGgW
xoGuNIEyEqrrk76OWxoNbVouEJJB4DbEhtEm3tyvwqDM2Ndnxdzfydsf4R0r++KS
upqa/F2TRW/BiskiHm3yAwGpepNNJ1KWMvHLWE7Zoo+E6AjLAkqo6EzhbCkJOf4k
N+9TlcVgwZXIRqUyfwQmQ2WnYvcPWErts4icGEyIDtLWhx+tzdwtsdXOX+znANjh
gv4J0IanhRXNX1VvYZtr2iJQmMR20oQkCgmvpNdU25Xhewb7j14ZBjZLwodHm+Dr
Hjb+cinnGiMQzNRvRcR9kc6zTX00+N1ew8sEXktYJimMhrxOTOJt4JqAFrBz6BZ0
hnbx469hqjCCbnxx7k/1JVLUclzv3mJ3zb9yD5Hbi/mUniz1Scb7fK/UvuxkMBSW
rTqIvyqHMf2WxmTPS7hbW6pmY5Y7kCGff0P9MNspdzP8CI9uNo8do4eNju4c1ra2
AQC82V4tzMmbhrcYI7K6D6+tYumEnXSki4hkxN/j3mpDHhRNtzzbDlNCGEYwwqO3
2VcaAJioLIdnI7AfB2W9h+vnW0Guou1xaSnW1ph6kf9YvUTIylnFryOYtgWCytpi
Uk17B+TTLh4ZdNSLq57nJRbggKrWVOHwMiZcXGg7BTLrp8OfQrmUPZn8ynovgNjS
N81w6kV234lfnjZxopo8sAxJCZ/x8tZpayp3utCd7kOV+k/+cSlBPzfUdR/Ogpi7
PoORAeXRItF0IF8OQ6uuXXBHttyI4V2/OKAC4rHuQOY/Ev6mGtT22aql2uFmNLGW
wi79uIEpqmyOVr5NvRTgsGYM1uHt+8qklMKkGGRabfD7LT5pCE9/CW4e0MeOgp0t
d6j9ihfbaf64lDk0kny6CS34yH6315Ceq9IqkNATN/mOO1DIV/HFNMtKcBsBrNI9
PllFO9gKMldZ4XdiQgS3YGzpfY3nCUZSflcuvjJWVq7FVmkoK3kj0nQ9+14qQP8h
EpzF/RupKc1cjYmSWSi4v6b/iaYX0pZ/mqCBUsMCbdfMYeR/Pb1Y0ZYch9oJwm31
ovJpGbyQXAMW7mLLlmR2KnxXrenMs2J0UraVZpWjkaMafZbp0KCONwxtvbqfc6si
wEUI7EawbznPGHjnVEcUrv/JqrnozVYHrS6VGh+NBh/oYWOG5ltY+oUDPOUPFJ5u
Wz/8Be/Ybjq6N9kXwHjIqepbz9vjL/WZZuQyTKpPaL1Op6JcbGmPGQmfYTXaXyJ8
tvfX6oqPJ/FuY3QRSi0+ZtWGjZPxvtRbQpW4yFNfw19mr1F9bxomta49dEZxxORQ
uzswiGMlru7Gf2+YeU2ZjQycRwjZCdY8FX6LOggus04Ut/UregVs/mPWmjWhgbG6
/LEWcqqRZ06d8FJIh0GIEILklrq349hhgsT7ciWOptrFCpWOYMH9EelehvX2iYlm
Sez6xugX2TyYdj8BAiMiNE6PcWPJ3e09p4mhhtiRqpYtZl7CWTAX8tdhp2j3R2S+
ZgyChkdD7BMoMw9ADFH+sdv56m+YJu4xYwNUtx7QXzbvPJuu7N0u7eSilfFN5MXG
sbPXuT4rLGXMmlXWi2X+lGTMpCJTYgXantyC9h2QcY4+9YX87bI6gkkqszTQ0HSP
m57ozFJr9ODnRErnJdpafVSgkVuF9A5AdkjT08RpOs78MA7ru1rWfMe+heRvDGMg
lth1NnXSdqvxKxUQHbSSnBk1L37WPwqyjMt3tjp9hpPYxzc8aj5rKbT7PPbhcWm/
7DUIqETsn5XfnaoyJtDAIwNtG/FY5dEnTvONWldFSuujc3hDOWoKkbj/9BUYIEAL
WG7jYBQNcUurepmolzZCxhBxLbwWPXmddCPd6tjO28mfHTtwd0veyn3LnGAzyQ0u
h6yXlP33xI+QWVUpFujQ9EJCejpmJhEHnu33eoLwKSNzlYAKj01/3lsqDpP5pn4a
DkUGjnc8m0uPSB2iEc7UjJjCJbxnjcsiMKGauy3h7q7vttLeSiJ9W/yT7fGL4qtn
VbzI5OqyR2iRqBh3ijMJZEf+pdot1mwg17qNLMwLztsKQ/fLmd5R8sfd9H6kjkB+
Kpnu6ARf8pCohBL0VP21c83CnzY9AKZ3qWKWQrhgMFU9cYRCIdG/D14CGkk+LIxA
DlaJ+qmTKvkeOuMnBhJS1etMAcecmP3u7MnOioeAvd6j5ubaSaNflBvHBu6gQloP
lzd4EAmTeYoVrSun7gjihIUlGQiWjG6mSIO5ag8KoF8USIJuGNLbBZSw51z7mKnh
smuqKXa2yQDO16NZtsKHe5vkRWQPkezCZNMRXai/3WvRWLBECL7l8Vs89ArH7N8w
yJSmDrmTdmD8dQCk+W8ZFVTILWwXPinvK2OuA4m2d7zSx1uYDsuoqoR0kvJ0rk4p
KkDFSVutgcqxTJXwxfeRv6Gqp2xcnetU6c47xGeIrKRf8z+x3CTFcOF1t77IlDPf
SmP4Wj3BzBGHrTIa9EHMeOTbUkmE1tLC0DjIRXPStoVofZ5OTafACUuP9i+oOlyC
atYTTY1XO4QGiMTzDYRDZ5XOENT5mjPVpIov+QWi617B7EkXIkGf4vVc/vLaUN4l
1oyH4FLpFmSZXCw4vRL8fzQeGuXcGQZBrhdE5jFKD9TFfeUB0/75W9s0p6fvMedm
Xi4Utv2zO1I3rSv9RPERmwLnC3nMkK8xSliJnnh54QBNw4yO0DVVcC9KNPB6Kwle
q1AguwmLzabWjD2+eXhwcWL4X8yQATl2o2ktUUrQOvEVmgpcdWt0CT20VzBtsvWK
MXbxY3gp3XKUjADgfeDFBt7xxZwRxaXc8dv6mTWTSKJlh2hIlJ/9NrxmBto2jLN0
Sz7MDHi9MB5d5Iluhr8/9AEXCv9gyt0lrV5AaqmiIFPsZZ2KOafVDc88q1bKavQ6
6wnX1ae3/3oLzx3uUomU7Dpbe2XaoIs2ZsDR54I8RDr1uPB2SiqgZq1/5jVvhp6Y
f3+3+hp3WPGKGSUOrHLo4un2lTjrQUTP4rTfh6y22YbMXxe3Fa9QXNZtWrltVJfP
xcnjl51z4lk2Iew1z+7y79Yi6TB2rIvLTgF4oNAShkXkvT9Ui6i7xNY6453+0mPx
uvNu17EhwFAn7JmzKr9O2Z5AfbhUmxSjKdiSLaVTyiubub3xJoiPkWvjqa4cSBLL
009ObxMfaOQIYwSibB+/m3SobIH70fhiRnP6NCxI/TlavgFhO899q0zMOCH5vqkT
6yAdJrnHKto70cU2qBgWa6GWpEbu5Bs0pym19yW1mPnvITCdbqG+KZegCsg6r9+o
JjZvW2Wfd/Jd1ITx1+e3lDHqzIUEdplJPYev9Q8mMr6xZ8oMpCMFgov36KM+Ly7h
99vbAqMmE2+5jtubnGVDFVfwXX8zoMYbRnrZdbLtNw6w5l843ML7wqDTYHFcQPDA
neu1QgHJER9JFjwTMUmu0XoSSvN/q2Pp4I/MsU/GW5SmK/22JdSzSs4GKm1Ws0gD
ivyx6GGAQni+4IaP6kSfAAYF5wpMskHFbScfUF8bX9alxN3d1/fOcIxE3vnyf/gq
hwhJjVGGOWx0n1+0hcm4OjvwHUF6SfBlyQlrN2XO0OvV4e3mPzOfyaX6+hEizYmE
INED39faQz/YLXy6lf3v5OHhBiiZnsg4nbvwEc4zHtxi6KuFBcpFF5qzr+vHTXDm
IdjLZlBSrout8AYeXAIP5f0IATntaGNxvidnTILPrvv6yBeDk78DLqBzpyWT5Cpv
UxuHWPUIZk7tjcwXY7a63cm20WGzufqCZ0y8taD/B68WP0R3uKXXClnOx1DFuOxa
XeDrsCutpJ0+QeZTh/X4y+HSY4N+RZGoR5PE9LtE65gI1cZg+FxBRvusZBqB6L1x
yrS1g30DoIiT6zaMhQWaGidpcvPwXASG6Ia/t8P2srOPMtAe7uN7UxTV2jzZ6OhO
0kLn1bMJhZGc0LZ90zr5XF+axpmowCulE8/3zWM7yTtxSYPuDzEMqwkrEtOywEGE
6zS6U4mxlrPI3/HKcdqiO8/+x9NTrMHbcdalAwLpjiL9TBssgbpwm095apQJH4PI
1HsmQMc3LJgTyACjGORnO5u8PQSWU62/hICW9X/GPjEv9V6RWiVqf7BfhELtQljn
oBUS2OCaD/VJVt+bVEp+Jez8HUrPpkkCn5eSg/+7Zsr0g9ypf9dUzs/X7S9VctZo
WytSUqqdNK/JIIoFy5rbacUI3VX4csgz2ePzHJESWrYxh6oKyY6etfg45GTXJmz1
kh6X+TvsbBhVZ4ZID0JcTtz+KtRqcgVducyxvwHfWSDSBLytLzATAj4c2hszH2lB
UJg+HLGsWPBkNADHX59k/MMWkr0WVx1DHBvPVNpLv/vJ886OpHA60vQcXGgN5wBN
pFbAMf2BQLqlikKmD89fWEoboMVRa3r0rjV/5Qy9zUJlCOnWhZ7RxpbEFMdVW9sk
RjnpbG78/1IKcF3fTuJRbRakqg9lHPxJ0M+rHMAIRVyOVQuJeUm+GDv16fcylr97
sgRZEjHbC6BjLpf0I7iLiX4PCiDsrhojMN1i32wVbd7XZNh6K7UVjShje2HgEqui
xDOc2isdkRmnd5+O27Yok1p8PCCs3+CACiLUyK3XztycW6hrtX4NZmE76fbrQBtW
v46aw6p7oQHngxkNsZdWEu8hkE3gA2wi5R2cR132XPEps0oQF+BnR17wk08emdUP
gPrOVn1cJauz1hWwvdsgmW2wihR2rrwbekJTLQhsqnj4OslwttgqtxUHHuju4s8H
8HlOsinslv2ZyZO7tjFh/fg3GZXQvjdSAiWy7CFMivH9IxuYgCZO+1VpKyfMCf0c
4kfTuL+EXCGRCN+rbipv7iVwATj1CGzFcl2B3w4H90911j9wbzd/m4PgY9PMQG67
riK/zAQES8xoxEjiCaMgEP7Mr9BiyumIPILjEh3XjruvGLIJZn6Do7pGzK1I4/wq
GTWSVMv2FkHyuHRFszXJIh5f6XWz61iuutlGHCOG973dL3ByGFyIDGwdjlB7LFFa
Qh6BlEGB31+XIT36u8gzXKGiPwar15J4udGzodvi6zzOipX+vt+ldk5puUviK6Rp
ol7eMxAWaVkQj5ZUNcrkZVKyOuvsp1/7nglckvsKw/0JQQbL5cwBD7Le1Czmlyxk
oVixNOvex6kBTUrTWlsqP4u0BiASyQRUOIMmzAAowj7Hu1Om4K0PiDHX1ftMo5AE
egFzWbuNHCket2mjBthT7t/bnvirbzeiGvPqIf3pOSq6HlCtTNWu+P56HlyZI9H3
OojGIRhTtd6bMGL0n/7m1o/aU87F9bezQr9BRohmYvbsB6Og5T2RD3sPgd6iskE0
/t+o1ny+xivas9eWBTvc6RvV/Il8xk/LgjS0N9QpwsyyrzMqhP5N9SMY43mHM47/
+zpNyhqMWApn04wXP3X1xUgmX0Ve51NOH1CL/+z5RUJTXNRe61ZoxrYZo6nYPXHh
XTmthFpPlioklq5+LQf4nftyRRwlpTJllOBgpKuc3d56uTDwm6YCAC2VodJhQnp1
AcEnAM3uVHbFx56wcR5QXo8qvLpG7csqs8wi7uj7j2Ka33oVHbW1vF28VmAjMLs6
zya3GN54lcYhw5YgLGFOubKPYo6Lj92FDSd+QHumLZIjFNR1HEW1qz/CqL/LQgae
TxNLUGj2wArWla8Bf3nSdAicU+Cf0hHoEn/jKXZ3EpnYcJ4+DUWQwxqO1sGVIzgO
gA+Vz5HUeWRMV/stnhOdZ0uwVPkM0qqfTg1luyu3qsNV9Gep82fTdAc72MmHvbAG
B/tQeVQjLcWZwzxiLi1gpYtt4t7euBKJTsdZ21NE3KZBR9/W5jwlaakoN8D9k93Z
eyHMkN8DF77+HDiJRti5jEk1d/FUfZKDhrZbdxEFoxcRxWnuBI8T3KbWKfWHR5g6
YedTTcT33swtkvtML8gM6rzptyCniZQvGAbjGHBbD0V7UWNTnQtefm0r6+OTcjqA
Uc3hIo0G0VdLkyUNpTo8XpE43Z2f19n8sCzbsEbeS7PpTgvfc9S7ZCJQ40UfVz9s
iP1/0eFIliG81jQXhYdyZHkRcLXRJTBAkphZjoVbaQi27Oktt/2zRXSZxM4Qgj10
ieLXAmB2RDrbtzgCkDG+3cIf9l0rX+RAe18cLBminhuHChuDycugNTBFhgniTVvZ
UmK9WPBYW0A7lyxagu1x+w1eXU109hWILho8EJrKq8ozMUkEx1s1n2WlT+7pvbVv
csR+0SlgwKX5CgQ4e4VcTvlOgOktBj8KEr2gZdhj3GRjqKoYHAWu+SWSzzeWOe5t
UISrm8S309+K4ScGl44lzZLeamuvYDFBxm5EPeY+CXj97ZcTQDB0dlQlpUewjRRC
bcT5YA9qHe6hiEFNUJd28V2BP2EmdKSknSQDmxhpyObeLagIfSonJt6YBz+cwuyg
u8eyGl5ykU3EXxaAgzsCVaeakQF/8ZHcXNUlPirgnOEo1govW8xUZMZxbbafqlIT
ZVQrg1y9K+arVC9HnsvRYHUayagmNsQC/Nlo1REp6vENccAhE2NYkZWqWM6StSYG
6Sbt2w/Wu/L1Mjpin7aSgltKnuFzB2ctkYKrEArRvtOBe+8cG5VbVG8uJxcWzNGF
o44ar3JhWCEbdlm5flOVUpFDtTjttV1OURHw29mLog1vgZNmwRm31DHVHWZrXtun
9CWQTO5aBP0QVzx0qs9081UsxawVRfJqZcX/6+i9OoXgnrODWLBZUV1pq6KZ9WOg
mTSV+0Ky1sykhQ30FrWp6uuPbZh+khKXEJWtAYJzkZSYSEztwGSzVFzGPZDEZc0Q
B/USs67bEb5skW7QBny2yV5MGGW3EYTohR8y+lhDk8+Op6OdChDL9WWH71Ea8Rbx
/4ea5IbNfD1CcA+880XBfUWWru+xl6+UMcmXa/llf5vm1c093Z7IEyz02aYiLPFN
xvARdOSUUteFyXYyfY+unykKbITh6W+d6P1BYH7mkXYNYq8jNeA030eT+p5uZQ/x
OZdnFJSEkRI4QLuVY/iTWIjuJYzDyl7s2UTE4lVbjq3Qsc/r4UxTuUAS+VuCxFRR
A6xAzT89e7xj5m+WMetxO5vW5s15mEzkvsST+t5eYcN5ZalZNxfxxDeHJ/k/rSdu
qtOtU6Y3Am7pHAH3chIQQT2ceXI9YIqiwDjwaPAJ3YLSEwpzvqJIls+651ajc7X2
pAH3NJ7JmXWrCalbg2X8Ddmzc15peOwT5MO8r6niNF1TWKwLPp/xPfvWA9Wic2Q3
JNPgK1NU7ewm+ttlpMF+VVCtvdAk+ReqIuAaBfYBZ6KJ1sFXnUaZUCsBBb3xZCd1
NFpuwb0pwWh2y1a7JCkly8glpmcd3uOnqpIKeudqL9vZ8EewMOuhlq41ZeAc2lLI
xjdPduYgwVWf1iwK3Rn8WinMvmMQgUKpVzOVbDy6pVsunJDkcGiGZgLri0EhF/BO
lfl0ek9VnuipMO9F38coEVTsopb/gFGTDL84wCl0Kw36VjodgP6ORyPpfBmZem7H
ILW2PTV670ENRvdRLQgppJ9MMt3Xwku/PGXuOlyLI+iOF3DVNMjaQF2zu+EZNfll
iNCDTuSR37yZPq+h3V8rA7bKA5GpcMbX7EsNlkfqn6s1+L5wkGzfZ1yp9EpItNFA
HCRo5wLzAs6g7mOINsE7oqU+yZ/+vg0nLC6jeAKthxfAWJt5wsL62FrpD89xguyy
UxXxnAm6v8FKb12CT98Zk8FUA2dGVahpiX8e3mCIdXm8aPNJkHJofjXr6cHZCu8G
SuKLcbD0UZXmQbaxTubKiK4IWmOZB8UwMpuxEdOsFxo2relr0oxNwt6Cnsu5/T+W
EhtNqRSQCx+9DzjhLFMdTxyU54u9AFndjUn3rG2B09qu7WWhzOfjJaK79hwe2+b6
igzAyj8DgTKxZpMgdWc2OmKVViCPQnIr2LnHdZbgI59YQGzgoB1S5fOxCMcCw1Co
JxjdkSb2g6dU6xFRjxZY0BDOjf2Rq8MNOp+JsTGZTpTr5U1yorjT49jX+TaLtCmM
pfY+4x1XsKKaVZnt/wiuQhAuicR5v06vqkuuRJE3BxqFGmRZa1oDiMXECyOnZNmc
Ya63e+J3eaPJz4pf5nr+l8PEJLw1yN2NJbwSXqBKxBHilQIdPOFAyWFXp2BKhQoB
L4uyGhjLKXzn6Og8eqy41EbQL1hrGFVd3fc3mcCaCYQcPriqz+/vOQNJoPXEiquO
vfRlTEjmn51DiI1UH1lZoq7jKTCjedB1+gbZRNGxa7JgIdXVfN1iJsTZWfu0yrqd
jtEh12D96jWJaJriHqbYwty6XZjEES0EMBrc2I+7NuAzhhYQ6bU2zl8a7Y1IcKjA
pnGX1GMFr8WYrMfyVPDo/+9jbS5TI9eThAFF8SppjQanlf09WHVan2sobEhscJSO
Wl2djl8Mr6uPf54Z+G7YW02ZSxMa3GkvDd5U4KG1E3icUbxFwst8gg6s41wSTrK3
hozotNb3yo+/sIWEaHsFqQ2YLRDp10uQPCa0p5PoeMMSDKb9i4acy0fTZK+W5fwN
mTp1ixz4VnBBpHw+iaD0pGhfYxKBD+btQX8JdbAIdfw5bhZhv8usevtcJs3B936f
/V+KjBIylq+pGZ2+WUoPCjvvh/JlY42mTtBjlz2jtJPklzD1oyy2XrD+nPTCzhDs
oMpAzixqs3+b12zehw4dDZGBJLxqvV43tOSCGvvLBJqihPzEPL3ArpTZegMuI33e
3B2ix+M4s0ZELaGoi8/TT36iwnPNB4k12AzoBJB49v5Wpmo8t3CxVMu15GcbRsal
yxf+yDSz27NHwaAJOLkOjIfxSZvoZ8j0i4lP5Wt0hzKnSNEEuTD4mBlI6W6Y9Y1E
mgpF1CgiW6MCGwwRWJMMWMTF35Jp58KR0QA75BE4+ZaJumNUyo28gO8VH2z2wy8D
dCA0VFz9NCo39RNhHn1AL8J4EBQrdTQpv8Kdtc6YYqxZSWMo5bXIVfhKBNzMiFV4
N70iKAyhXwutKBubIOrswTXsHxO5Ywcf4vZf0tEv+JdVOBBNjEEztNmhKaKqmXza
8UyPXPlyJ3Hy1npsloBPr6sREUUfyBQycnadZTVa0h/pHG+7qxHhZleMtFpf+0kU
ZNjd/1mtSACBnfekRffU89vLtrmqdglBSm8lETyUf2mXbBxsfxb/Rspk3arUaUEU
bdEp1xxNiuYrxaO9PRNhOJhx3kANSZmfYFdqWR25ROY1Bp0854LVw5ju3HGFWtMt
JCPdH2guPSbPlzUyKKQBGz0S5YiWTA65Rqt/C5CY5KU7EdiBHjCnHy24PHr4wklx
lf/U47OBdowwrbVw1z6ZvJLJqNRv6NkWlEzyf9qrXyEPF34MP1gUxfpfudniapg+
YkFPV2JYdbDZPo2e3P1ZurxQvFiJvDqzu6sBSd6BgTv6GDQ/xOQfhmy58znQQ8Xe
I8UWO3XQKBIh1RAeo0zS359+IFnzPRX6F+5971MpN6IR6SUgcKLxghrAseH9fUE9
Fygqr++7kQ42cUVBd96tWuieYeJ/iQXjf16cFLISd1fDwE1rjQJTTVt4fNnwAS0Q
dbl5u5VLO5fl6gw6Uy9m7c0iSV1dYvOa2nmDz1R1pSJxHRY2pcMtqrjnUtS1sOb6
msDcxvoFeoYQUS8EQRYdcrgcPrgT8AWHmI4xf4m40tSASvuDLiENx0CruZXLZS32
alz6B9hJun4CQMJBUZggk74OSZIfQm9ZlHCLouHDYcsML9Nvm8umzE1G5Ypz0Onl
6rqQ9gtb4yPXg6Gzw97b5wIfFiZdvkBCWT8rkjWJRYunE2UMI2wVSiLDY5X4QtRU
Hr3yeSmC7sMoo6xy6la+YO/c0pLES6XfUYlZOV/q3uOtleFRD7AWAVQ2++7KLRfE
czE0MjJPOY2sfTWvP6gGcz2Fj2IT7xCdtd0gXz+q5UuLy8whpnDKWNTyfDAhpYsw
sYJ+TtHQL6VbI9/e3cZUc1L8yHHC8WwRfsa6jGd2HSJ7lu8j1MIE+iFf4JQRh7K5
LD3iRmfiqm2StzG5/uo+/qB7+W/VsD0Dt4twuFSUmeoG5syC2szNi/USR4UavxMM
atPGJVyjP6tSUeqibgqjGu8cfWUJp8/KSNVi6C7MBsxDXSwMQVCRPcaEkgMEStPR
qcOXguQi0fLvqYgMQB0Aa/dwijg/sRxPUvk6jJApRS3NPI328MD/yxxYo6vZSXdT
qSqtEbRDWc5JducW1Sa7eA20fo/KAqldNHqfEZYcxH83TAb6x4QrXJFJqBej4FWG
0b3aDB/Lq3fJC/hKHZh9PCAAK+wNodm22hu7DTt7Z/m9cObXVpHA9897U1vT4hk6
DmbiZQyvfls+IeiH888qnJrrcGzChU2PzwjkdqdJezNe35vxpISCrvS+4qjvpflg
WDmMzbGBJ1vy2qeUH8aOxQSDQDJuiwssnKOjLsVDSA9CTkzHxNcw9AdhdbkivR4J
cVg7QCFM7qAdHlp3HH8SBXC/kC8lEHI8yz44+pgRxoCfC0OgmBROshdVU6zv90Y6
ZYpALKnlzuYp6qqHo2b7KW1e+f6U7//3i8w2SuEDvq7194XAVcZRF5nUO4YY4F4o
wWcBoVMNhUgj3K6BY9q9zJpwURJB3EQKzhDwcWtp29e7DQUCwl36DI5YHvOetlPD
AG05yGSSB30sDYnXgdi1MExv6unkz9DtQ8UulbhJO6HpqJmwSeRVyvTaH1ZQrvf9
aVAjOyyXmKGkJmCks7Q4tkLGM1TnG8/0PkyrPmvA+SVzuYsZdHZgsswpWQbVS8W/
`pragma protect end_protected
