-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
M43ZbHM1E8LmbrOYvSUkztBsXY4veAyOYpyKtrxM2axRTQQ9CNUlWaf+OuQhnc2XVBieN9vcfDs7
2AiP7N1t0J925cUjeLBPKyC5zIN0l4M0h2rnHqrFtOIrF7Dth4A+RQ4jws+tbsmGpwpJV/xYATtn
cGx7QOz7gD0TLROH390r3BCDwugPFajuDWDlDV2f63xWMMA2Sw44dldKAgGNav5gfX1ti7zciaTq
JLaZ9TtHZmnkP2ugUjmen19DuaOYrrkL1J3aTxgpfNXpN/CLwCm+3C7/BHgwSP5pekzdzlgvMqPg
4IsE7jX7FmVS4B+aS8bCh9go+m4BZREowQfrgg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4192)
`protect data_block
+uBiEz1eBSg9UqcRhqcQPEkZs5vq33t+ZXeBSvJoF/3XLSWDucxu7W6M4BaTxS0PddXAdCiKWPOt
Trq09OVAaX0+5Rf7nCveRQ3I7e0RG6DwWO75jqt6W7/sRxKbaur9MYZN8NYvrGKH1fMr1CiuCuUe
qk8dmyMhN/bkj9kV+3kNxIpMRB8lfmzl7e3WNQh6kJnAoOQ2xX0XZQxXuSaTGgomqEcGWWtmZ5Br
9rA0CvYv3B6AAoFxE9bDtkb6pXjTTcFJJ97aCB8kjFvGRxiI0rdhgJp/162PXJejQdoGQPku2kvy
9q06Pa8EBauKfi3Klc2jXPMg2udrD+6nmWz89Cgnl74119+Zg2yCLCstONpPuY2jLd3nqvXo5XwV
tbwDx2P18PFhljhZ/nKwWl+bQMrWVfkAuD17KOc9UTiperGqReQL0EYtJxZ4LowZI/zpvYfebbQq
kDuMNC54wnxGNnl6i+nNt8865iJirelquKl3jg6P7Q7Vc39ZMxtQ6woledvZz77SDEA/e1Pxp1R6
fg3nUeOgXERQYUfyny53lFQYfSpXpZZLdxRBWNwBiwv291QTJLkFMlMpJDmzAO+0mxeytgqFTG/B
/tTa4trsShtWEHM5yYzbNUXeYW8RFgXezAm6Xu6E8fWzN9jDx7FixSCuAOJorQvRMpL26QarCeQS
RST+kb/LuLhLzQY/AtmhTQyeb/0iD6sDOYQTw0R0W9sIVlPH26VSxXyfZJidmAzNZAzwCnX/85cA
xEcJAOHnCjX1XWLfi3XiIS7lBriYotT/YW5X34+73zp8bp34MGzuzcZxRsieZ0pGkSgG5pege3Z5
AuHDzcuf/rVvb1tXJP+VEip5blrdr1PCzRYEbz2JlxiN5O/OTBNw6wQqcMvVKZPrcxCXZXBeyBe+
5/aFTSAZtZwfVzhno2e0XEvzF0eOlJguyw0hsaOf/XovgTWco9zN37sWG5xDIh1UQx687iO9uxGQ
kkvcKJVFq6yqUXzf633J3kwRiLhGWrAZAzz2d/5ELj1yV4O2pZ+l+pqyfoLV1aLvkI97j6wn58x0
eWz4gfI5Cklpr2lpDS9c9aQ37JAb1u95V9w1bv0UcJSAxVBBW151YUgA2jAzGmF0xiKJimzap4t9
xxZukxjDpTibH6pVRiBEc3cmo0G+XuB7P/DnYUodNe0S424wmkfrKl5VnF0yfwE6edKi04ZgCaNX
lgOu3dBFypeNfUA+kCldjHZlpNatzpXkSVPP8GkVJA/LUSfVyy2yNpfZjzT9XwZtSd9U/gwGLdEr
R9Y48TT5F4T0o3l8/Sh3BdcgLpcgSYt/xKNmrWaecAmDCWLe7BGFRgU9nnfm4vVECPdLIOoP5SHo
phYtbjoDzVT/JqPmoOkjfa8A02uL7jUdGHwlVcXAdfeXHOo5TorOo9tcEwGKbn9dxWBiOq5p8n7J
RYW4zDimDj+LvbniRwpDxAT7T/DgE1uGspS7rmNMEqfc8uJThGQpWMj6UIQDrBd71M132W40edJl
sHFNWhQQeMtVb2nUrdu98K0y5761nxf145ZI9j0CacV1IES1Jw0fgQYD/iAdFRtt/Vb9UwkQuhEL
L10A2374AeFycuCJ6oi71bZ+0xiuaM6OPK6wVfQ7Jztn2+HjMJcV8XcSSJhxJplmW/Ojypl+aUuY
1a5NXZZg9E/HBFGt2rY0PZj8l+HBlcmqc2FnrZg6kfPKPoBbNLcEgbMpWyk0quDv7F1v8jtRZoEx
CNKJvPNmZX9td6NFXL8K2KpTw/5mj8VeXg0H01diKX0EmJI7g4v3D0Po3GPuuIjn7s7zikBCP7uV
JInO22TG43IUeIYQ8hqEDCjzt2iLVPOf5wDaEoCQccUaEcp64+SzD0xqUqhRlfBdLYJyhPZRxBCu
W9xh3HCDgibH37RGZ1/pAZAE6g1doMQ3+B05BgC1fVwPtIKdJryt/GbvKBfS8KO4BIwuBf8ZCFY/
3ohQV1v5P5qdVfqrNt33iL7Swc19DdOp8OvPEjXRhPiXOqHArA3+4fBwYPGPnXMqWc2BGJfskFeA
veMKTmfToLK+LMlNsML5oWtKc/4itCZOOhCuSO2k1zSKUhKNmSkeVesBCudLfm6bWSFh7hOSLw8L
/AbISN7ym5Iw+3jKPUrLVkku/QnwKTQJy8qLphU9+swBcCZVsIoBsEO+egNpJzdKbr5Va2VFDAXy
/e8d3HqmMl1sLQpBh/PpR33IjPdjOwfMfnun3NDex/OHdltl608GAfAHVnWpuGLiv8MJCYULmSZQ
4fq+I0kk1Dx+1gHsm+1+73Fwcya08K5PSw1uD7OJFSA27gpMrLJ7zBI/Y2enFvAQjetd4Se8m6J/
pkt1bThGiZmj8v/+sFexuyJzy34Faz+hHygilFI5jikHtaGTGeN3u12Oi/ShDwQKdqHLJWe5zSVn
1u2pCfr9RdWnexAnjckWUGXunyebUju8WwRNqPZ6grct+38x0HE0xshBKlhZBgWWoGyMRU1Egncq
OBMxzHs5KALBS8WyXE9UIKcf46iPMkoDrQbRIFaICkD8/StrT61JR4Z2tS0DZ+KxMpB397Hk6yOT
+b9+ZZKlOr8Ud5Narbt5377F6Bv1+/08hX6dQiCNOChMbmJwmdD0C1VsLTs9aIeLQxbfe9xgAu3e
Uoh9VNwnedcPCadR3Qzf7mugN7T7/Iko8ZFy5B24j2IgVcUuvPz6FcETpG1hdEVU8uGfPeLgsRug
EVpokmweAZiFHhjZJoBTyCu4gwVsSSheCtBhQB4We0cPLhq6k7FvRxVJvUSwqv3/7og/d/8sIS/K
Cb17mIUNzAyg+akVO9xLJBiymYyqhgzkdffStQ2eaXt1/MeA3ZXNlT0wwgaJ3vBT6O67kK0N65fJ
bQ/DI/hcQvh73/8EuGwtI+Bhsbl6xn55nI6uxR2jOZFSOEdr5clnkoKO7BenNhlkDgZxv/oANg1d
3X2goSfrE/OkSuLGEqlXoU6sDiDl/csMRq3+fgHGy+jlbx2S8rY0krPvAzqjPgXPcJ2zYZBQja3S
ikVQ/OP/t7M4qyRHIM5sQafkA+mFMZKFS2UhXcghd/Qn2iL0HINrmsHgp+4RNyofIHHXeEZ9K3L9
qk3SRl7+E0TS/90vkQ/NJz/e9EJgb3SsbTPEksWBIMf7fsdiVgQaT5/nrsm0xixdTWWaQd9VRz6L
vukN/5qXADYa6HnhAPLulJ0SRHk8qLdkqlwL2ruR5/TYnNwck30pDWndFWCnLR8lj+e0IBdn4zcH
tYQoOkO4XEaxQP86ENavGlaU1EUGd1R+5iU+kWgwImEUbADyRO0OgmmTnZ6UcnBxAg0+ONY2dOxG
KFqNHMsNB2RHPkf49K5AJ1kf0Z9ZyfL6GG3nALMUKgibl0Ez2OsN459LMqlFbGKdoWE+Qj5BQfg5
v1SXkpcW7Q0v4AOYD1p0AxjQndLPIG7RuLqZZo8+rtKXV+SGc6OPp885ozs9c9WSqwj+rv7x1V8c
Oj51UDd8rl8Wr1o27er8WeIbsdXEO1CQrhluaaKU59lsyELhHfAbgYqYqyqtKXiPy/lTlklM7HJT
515CltXtzPDROLBmyoMs6bzXWjmppQvmMlznrkWDYC0eHABLCt3KrYqlX1lorfcGPSNB3NNuk48z
d6CTQe1Q7uvLLP6GeOHIKVJYNgBs8nVFsirsSXKiyn0DxJ52Gvu6yJ7tBNJlNzGmx8zSCYc6XeY1
9rNvc3FUuNNfYb0Ln7mUhrOFkH1+o3O/RFPOmYT/w/6v50CQBM06RfMJmR7aGt9ezkPj2+RWiLRs
vKvagKV1htAAoN5dR/QrMIdMW1xUQ/h0VOhQaWZasBy/kDltLn49Eq5B0owLG7txf0NMVxQuPHER
TSJlcKTg8Al4k+t5SZQG/s1c7ZUShIsTQ3+bZ62/fRb3Uq0zP+fISFiFVq+kR8QpQ9ihVfAajDMw
nxZrm4RWjXScRoyaMeFt5xS+5bpZeBkGpRzGYJMacNr1zK30dk6I37DnbadS03BY3NgKMd4DGL45
COCnuoXDjuuwvP6dhQdDOClnsU014IQUGgnuZ3ntP42z+1xnlUG7ICGpCxX/DkvZoJ/Qk4x+9Uxe
S23x8bowp7qkBzcx/qjFncla5PNbj4VAYFlmN+60YAtFRR4sG6ibZ0ZIUykWL6SrMtwwTDmqEPDB
jaj4CL3rYhY4NSst1/kgE7ov95S8glJuZDq+l+v8uFCay2OaDksGE9dp71Uc26Eyhp/lhEDEGylo
P2z7XmomywGMG4litr/VcuVPlS9o9ywuIWtr8q0D/LZFjDZ5OdHdHbXIqtzBjYLuSoA2z1tTKrlv
bsjjkuYVIFGOnN05iyhDddpycZJBXmZSBdH5m1UilX14z92RvY/8TTSDYmBcfNe1gR3EBeTr0X6g
UkXjr/HFUVYizFvTWOZdiBOmcaVabXlsVJtLT/Fk3wbV3y/JJWZ4mXsePPISfDVj5SKAwF7W4eTN
JNKe6wbPmKUmVLP+IZ0y5SNcIHVsH831IkvyCnyG0dKYtW7qaoPvg9gCp/H7R3zAd5iVSphWJFCV
XHbkUuzgydQKPMzSKHQ+k/Vg4qU8x1bBNoojnfBrabSEC0EuBT2HGukn56Inhu6Ie6KdQrx7kkqG
qxTf3RWitoei5ut+dM+g7hky02mwRGWbtPBv7NbUCmQXxE5DyqHCZRXdenAqyi+rf/Ogp3DY0gcw
Z5wNK5a/UKhaWyafFHGpoEI0c50my+5Zv/bSBCpAkS1754r0HwQO35x/jotDIhedCKq/Jl2g6nmc
8pGedd9/0k2yC12ZcetpqUOh2LW3hySR48gePRj4cz7MdwpIZ/HBi6yNx8oVNXhdzllPG28h0tqV
IgXQeBoETcGISJNri94LNOiAhH6NfADQOMbi61ujjOOoK9Y42eb2r12oNPxaukbrCMCk494IaiVP
vV3tq+1S3V4fVYDxoNiBhuN189QdorMlVFT5AhJm6PbpV/M3Nxz/Iuy3jgF9ws5agbN1vM7ze4cT
2xXM5pC59zaq4/L7NBTofRFSdZLT0Qtt2P3YyDu17oS0CYZ1QdggYsJdvnRK2on/ECNKCCs3mrYp
Svx+jRIrce1ePkghzye3+DsA2dPh9LYw3Xj30CbJKRaqdt2dcbXA4/kVaVJpymIudA8zNcyIRKfC
/oysbzryIemB9QjauCNHNsrlhFTwJkOmpll71fsXkBEoePssR9ZWSHiPzXoN4DkZLPRIFh2a823F
pQO0GzgDGUTPc+ViITV8uNz0XV36JvltoOpWtuhWHQ2DO0O8Puy5Fnfjgd2bjYWELQ0rcuZZEY4W
peV8FrUq+LPpfmdZYS7j07CHLWja5UXFbwJNFD48FFNjIZXRPVGNyVRIWTIJqVfmAJKRNB7FmQ41
0aHlbN0eXd+BtLJguPjCXkEU/GMlHdYiwImcH+gEgDmytXOhLABJrkIo4BobvbkbE61sU/LEU1+c
nbp7Eo52tTV35AWB1goGPLGo4upIeeK80+TsN8lGWqShAUfzs5dX1wzIj6pN/dcss2ahYKB4nPLD
/MvTZhD3o/eMcYyF6RY0YwGKjLmnhrh/Huq7DRHVRA==
`protect end_protected
