��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����S�M�hkF��1~� Ά�``0Hɿ��b��i�<�1�SzFĐ�48��ch�iIQ���H����:4(c��_V����&��}�w9B
��T#�_qx35t���D��<��R*�E����nK�N���������19N3a7K�0~��!�@ըfG#�=V�[��&@0Xy8�U�N�
�y��I�S���j�kU�,���87��u�:]q�Ƒgh��8�i;�f��ܐWq�Re�R^Y�˒�
�1h��{�%z��1(Q�,1:k��S�pv�p�$�듮Z�����C;�y�A֚��Au��*��1�-�_��e�(� $��d8T4���z"�������0����W���j�Eզ�$f\��W�t�(;�g���u��A�j(���g.��=�kz�7݅cִ10m�OɅ��1YW��F�O�`�,�w#{�iR�{���X%>�w�?U4�re�C�E��C&�i��r0��vf�8�ԫ�ft�cY!h�����Ϸ����q�ׇ��/j�"(@��c������mI�kru��)��2��*��0�r4�������i:3a����-�������g=���\6A9l�6ιB������:p��Y�Y�[*i�29��w_�\�&�h+!�)�v<�}�!&��V� !/��y17�&�ţ�*�Ҕ} �2]�H�,�nV���˻u%x��[�n^j^���XԞ:��
v�9Q�����3.O?����Խ��@��5�RlCN=ۛR�J�%���oP���'�̐Ӓ�J�嫃C�EIg,�	кOY�y�f�����{I��xBE��e�[��a����-���;_4 �R�y�D7f3�ݛ���N�v��{,��ı�2°K�ui��:K���5rp�FJ�Z �ca�v����Ӟ�onHa_D�ޜ>��SD̈́E�8��>n�X��Y8|���"�UҚ�sq��x/?l��$z~և��NU
�[�I�I,����#�w (���T���6 ���Z�ަ�s����	�K�W�̕e�s겨���	A�
@�<iP�H�G;8�^"Ĝ�I%�)�cã1�<�n�N�L����˟c��s/�y��y���m�U���Q�9 l[A$P&[:Dy��a״M�Ǝ+p/ �9\N�=�kM�B�}�K��y����/]c2�����`	$J��*�U��;꬀����z��}�b�ל��RH��%�q��#Tq���\)FOgR�=ϵ5P�7e����|�F��;[MSN#Θu��$uw W;g4�4p�h79�^�\�W¯�{5M�0���-���Ǳ>�<m���=�:�PR�/@�J��k�0��f��S �e~S9�y�������6Yr����؆[kr[�a����{З䐛}/�Q-��|�7��A����%ZPJVK��nET������!�lMB���1�IS+�Y1Q��@�aՠ����	 �X����sA����R����A�Pi�]��J5èļ7(̈x��V9�j
�:�׶�##���0�9�����4�j�^��_�es�"5��!4�����5��v���<�b<��F��MF�*`?[Ț��=*C���M��-w������
��h�lקO=Z	K���-���b!zz&2G�U֚a�k ������"��������L=B�g^$G�=[ 3��[0w����1�sk,9�9��Z����}�A�;\���+���dk����Q���]�_#UY���3%�c��	�k����M�#�!��|��{���p��*��6߄'W�:�1e��A��jO! 6�R8���hAܸH��������tт9羕�vi,N=��W~���4]�&�C!�ü��H�#9J����o�g�;e���&�V�`���\���u������0@��G��E2̓�X$�����e���7��x��9ߘŠ�;�<Ob-�m�Q;� q�}9��ٯᒢ�V�'Ie��T����&m��*� :;=��ڃ.�~Y�f��Inç�F�^y�$ils��w���iu�b]7��iֆ��z+:���֡�i��H��u�����e����}�"��(�?��QT�K��ɥ�0�#���|S�U���b�����\9p�U\6�j���Q	X��߾�/Ӗ�O�3���,�l3~A�Td��^|'�>Tt�����DNS���ϺML�)#�J�ԫ���pb70���j���VmumQ���r�oC���E�uy��҉6��� �$}3�W1ro!��Y�o��ۼ=r�{xxWn�M/�ɼ�o{X�� �/�S^�4/���_��̯̓���^� ��(��c�J��z<�$#���)���h�X�7$[7����"�"g�K�N�Q��n�I~*Ų��ҿ$��T/�~B���]�Q<)Ą`��+��\v^;�}�kl��.1��Nd˯��a�" `�cᴼ��!�f
%P;hR�}侈���D%0�])�1�Ϩ[��O4���w����Aڕ��j�_��Q�L�S�����ǭ�*��Śӭ��h-��sG�~�WO������\��������`�A���> �B ��0KЉ��_�IG��w55\���
`��$�����b�3t�H�����4���xϺ{5Nz�;�%��
l9&(�-�yuZ��u����A�n�&z���W�ȔH]1�w՚��z@���O,OG�i]}��擯���y}�B�J)��jV�T"�Su��d�5�v	Ww��Ǥ1x��{�m��+�8��@:1�7�B���&�̂2K�]��?�g��b�t��RsM���2��7�5%~ЩJ�?����bъ�!�C�C+Z4��/;����+�jz��VC��2��*7���*�3Q�彴��B*S,����Ԏ�����kދ�s_(�ww&t��v�8C�I�����V���6y"�G�4��� "���U��:G�'�!HF|d�\�z��u_�L5[�������泰����V֔�utM�!�����#�x��Mf�b�LҼ����{Q}�/ԯ���G6%�?b�Լ��� �=��( �#f������^ܺ�J-� F1�o���Xv�������<T���@����M�@��cL�D8��0բ/�)���M�E�v�ȝY_�oppb��x$�!IQ�`�6���Y�c3�.��D#\����z����U�8��o[��u�I��{��H6!!��J�e�c;���6�lb��d�M�t��W���:Bȋ�$\��Σ�糈:_:f����5��ø��J���̦\`��Ӓ��/]m?�(x�M���_����*��d��4O[��5˳�B���΀FA����D��D���¢���Lɢ�>�7�i�8��*̀��W��>Ԉ^�p��a>_���ޗ'*!o�����K�5rP{�ߩx�=z��ku�Kv\VL��ףLr�.�-�m������s�M	�/(�A�.�����-c��}�#$p�9�/(VDF�B�"��	��A���G|K����,�ϭ�Պ�ʮD��h����>����N`�![��i7���KL����<�(eҶ{�X�O�L�?� L��~�By�8�n�X���b���'�i�5�jE]��g�f/�=�L�v�U�TWLh\�IL�t~������
x=�`r�1��)�>.�[佃��4B"����U p^������>�e?�Ӏ�~3�OB��'��C��v���P~���n#�N�`%��������2 %o��Ͻ��Mw��c�-&�!Ŧl�� ����t\�|�L�N�/���WJ��"|�C?tJ�{E�UL6x��V��X���q�8���k�������.AP^U����~˺Z'�P�2Ժa�����#���P�C�����͘�R�V���X_�u��N����	��H���J�i� v�+_�pܑ��	Z�	�Y&��epMƷ���y��w@A���c!vvM(4�Kt��W>��Lj��r����\K����%zw��`���
��Օ;0���,����po��r�9�ikmt��Y�T���;),�H;QMJ����>����0s�x6L�{�����������_p{v#�uII��	���D����e	�ٲNSO6�R����^$�R��B3mJ�c�S��*	�My������Qx&FcR���'Ӷ@ &?-��C|��;ޖ	�.B�WK�x���W�6�꜌\z��'��!���ӥ��N��k���{Л}�� ����J��iV�{�l�jw9�������z�f��|~�)%�Q��YԚ"m}���̯i�Ly3>�	-rθUό��сg���G0�Do0~������ظg�_�	�@$���5`��*rء�q�}�S�^{���f����!f�SE�'���N���h�8+������[82��B��j̗-ᰄ�5��Y~D5Yѵ��G����Y��Mm��[ũ{�����;lU�{IF�W҉��8�ȟR+=���أ�����*�Gn�YP����6����-��k�iY�Rfd}�9���L��eG��-�	VP/���〚A��q݃� �@:�O��R튳25�C�A(@�7����<Q��+Xǻ�R���!{B�(�"�,��]3�f�������B1N������|�.ꆸ>�UWN�]��:r���h�I�
�2��f���[q	j?ꧥL���Eɮ��O�_�!������TK���>?��tD��/I�6���i4���=%�xK%o�\��9|x�g�P��Sm~�|`T +�{:�g����w����uϘG�L�z��qXX҅��C��7|���<ݶ�(\[��9�6�^*y�"��Z�D��-�3\�7��<��v-�7�w�b#X��c�.�%_�m��$RV]$VL�D���X�[���|
Swn�U����D�Cx����|QvRĥwy�=�֏�OM�[�걣����k �|�e{{�7�e�5x?þ#[��6��Z�����������?��%����`��0�g� v������I;��k��������a��k:c�a7n��$ f���V_�#(u�Syد�.'p����^���hϢ^�09�(YDY��B-�ż�8� �!.�=�'�%�����̐\T5 w��d$RtD��W�m�Gd��%��z)�P?��I6��.~M~��a�s��bz�Kb��ZN��������w��t�I<*D�+H}!q�m��F|B1�aN~0֋ZZ��S�2�[���L�[m���h���L�d�������w�ey��Īt�S�:�55"��%�~���P0�����U|\˱|e9ƨY{���_�Φ�
xo���9�'��yt�fpyU��
;��"1�G��72��,�M��/��JZ �O��VT�����l���,@)�s��z�Y^����*��9�A��V�a$+p��� �9��YH�\3��-���t@��ܼK�x�Y$����
�#JC!��I�Qt(l�2��Y����?�8������'�����܋b����FO�s�U��ܓ6,����@��wD�H���Fx���*��L�~�˕(؊������K��A�3�k+w�����58Aޤ��6�Xd����ԥ2�:�ۻo��=�P��/Bc��)�M�7���N�ӛj�L��WA�xܣ���SWj��6����c/&�Yo�6�vh~bȺ(�^6�{F:�_
���W�~�G�v��1�Da���X�H��"}���4!����1/�>�Y�p�ßV��w����к��
&"��տ�V�q+�0ka���J��@=�En�����yv���N?a��"�1��-�칲�%��͟��UWv{x��{3�:�y�ٛMs��F�|C��$Yd����X�?��@r�VA��t�ion�[5=�T��Κ�._���>(oR[��DW��Pz��:m��ǕY�C'�:��t��V�5���ɕ��C<�/�I���7�b�Bk���A 6�	`���E�i"B��3���ɟb�R�E�e����_�!8�
0>��	�.�2֬���tM0c�����){"^��<}�<��|�%���
��{�VS�ݩV�z�)��<6�+U�Tr�4E������2��˾��ڽ�P�O����S{���E���կ�b-8��!�I�m������{�����2���� 0�%8��s�y���T栛_�M���F���>�iX���t�WW�z�}ֳ�Iމ�&�m�nd�-�tE���(|8$MW?M��ޛ)6�@��Lu��ϫ��� �8�3��BP�������6�ٛ��P�>!��;��b�[e��8x*��b�i�4p��) +,�o1���3ޛ4���R-q�?��<��8f�CN�k"��>�;b�;f���!IT�&�G�r`������<����]L�Rw�9�Up��ɺ�(䱙ʩ4I9�$L1��Sy��\�G�t⸶1���hq�+AZK��G{ک�^k�$)�3S�rX/�"0��zJ(˃_3�/�È\ˀ�C���J�5�8閻�=�h" Āb}v���i��"��1l�f�;��;6E�w[� �Gc,mB)T9_po^���2�p����	�T,h����� Z��Zuk$��Ԗ��m���Z�[�(�*��>R�a5�t��5���A����"0�mLB��;�h �R7��Ǔ��{48�]喕mש��R{�4��0�7_��x0��H����ר��.��35,��"��$�ܿ;+	 �"0лLW��Z��p�,����FY���{�VT�T��
f,ءh��1��v��0�Q9D+M�\�*[��,�2v�8/�\p~��/&EKm0�'푫�v�o�������O�ݵ����+����9��]'^9����?�b�{r���h�}����b:L�b�Z��*j�VN@N2���(���s�Վ!9zH6��$y~����樫�T�b��y�#�}��ȻD�S\�fP�� ���	a�<����[����;9��}