-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aujbeVw+4F0PPf0nDSv4/C1IUZMCQSYtksMV9TnS5CnZpeVBUlzjbAQETIb7dv5PzK/kliJphPhU
yFI24q3z+VimAFeHU7gIQyHGE8RPIvl1b+0ndFu5vFCNR4SZDIKql5NzOlP1QZN9FQGm3aH7M/JE
8fydh5bMbl2mi576nyJeEonMLqsPbCDXiXpQm5ZS9dqReP1mrzGD+8U3B5KXLMUw/XYwRt/8MqDq
yd1aipB6dwXyWSHHRUgX3DObxcOP4sJN3c36VUB0Cag1GOvTEpyFYcUA5Sh3IcAFhvi6YMJOwaPV
u4qz+i2583Up4HZbeYt6LgC8OMh6bi9Gpepedg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4400)
`protect data_block
xlGPUQaPP9AnMgbYmLYk+6A9/GCJJs11inuVWCN6pQgU6Mk/rKSTKRkKlHrEP2PCpHErHktrOQGM
u+HrMMWeO1Wp4rw4cVBS/h3hiuX1JIKKFWNbQJCJcqL/AYH+D3zC1q0yDWROgevxnxuu24HTcBp1
jsvLvnzjVc2ByC4+/2Gne92OQBYM9Mnd4ZM/h5pTBXFP3A9HEXDb8nvWocN8sCS2aqcF7aH8mHYV
SqYfrkGGZPCxAv4EnRR5M66Lv4lceaCjTIl3XIOWp626wNjAgR1QkDE+4OTJ08sVLS+wIEveALBO
lzhxsICJODh3IaIehxPOMIlBOl2lPq4RYd+JF01Ju7uGlbbkeGPPCywHbFlUkmYzgVrCRC2ezxG6
5lQJm11+XXeBDOsAdePZzAr2tdRnCZc7WysvZvV84W1Ddy/Hxk0HAIyBLrz8Qm59OkV2+49jAb/c
6Vo2dyY/d1LNw3KolftBlSsivoij/xd9MZQxuxEri7dtZYpomWUYeXf1tPZPU/espI7Kw1f4vyG0
r8Pwy9rJmIFUzcU2iLjyovrl1emV4V5GRrZZrSxPZEZ2n6ouBM+jf+LHHSyp6YvnNSQg0bpBxar3
dJA8ddq/j3JtVt4TgFUJ1vEiEuHNkvS/c+43UKVWDFfOvQOr+Bw2RTHeGHOkGGDJOVnIAAeFeUqV
0IEgrv2sp21dpy8bwoUBsyXKBOI+L+D7VjA1NqDNpEz64n8JOjayLutVMbyGsQxHdAAVrVi8n4ux
i1WZuiEGAF2vfH0YOv4dR1SE2is34u8NVzBzmQJFq7xLSfW5uObtASzW/AGYTxXSTs6oNCVyEX5x
BUGcSWujx72varmOpl0tiuAVLubuOhNntFS5eMfcTRcZEKC0c1QV8F3Ba+u/HMDkUH2lVn9JuDLS
pk+ItA8QbQAh56cls3zMWUZS27yiau3c4IZtvb/eO9ReOtPtPx7wCg0Nn26nTtf5dtJBvWEmNQDb
mOwZDvIe25Ey/W8KQ8FjH9/6VGKyKc0G1YZDAY6pbthWaULhyzKW4JGGV7MedXX6KNwIMfb2X6mH
ubpY40ulP3zws4UDXVJj7fZKxasKT/ASQdr7xAT/CUb2fWgNjv+4mJRvRHsgpPnws9kpw06Fdb5M
Gj+ZQmurkTjfu6oCMlHaWGkXYqA3SF4O0waEOqLMOa8fCP1dC1B0ncR5HY2e0ZMQL2WcVOOVvVPB
e2d5vgTUjW/3DJY/PJ+3/L/BsqHv3KLpDSFt/ZvsVldcl4aMTfyCjfVdiBptP6MfDx/q7uYRFys3
lh3K0b7Zj808Wqk5uI99kC/JZbOBc4V8jgUKsmzyDhnRPPjqjSPS+BUZ+5RvP2pxViWM2awqQI70
rxIMknhWVLlpjVqhTfn7svgnd1osGnTUbKIhW4/UOUS08zGubnJg6TGeVO7dysl5dZnihr1fTDQu
fpUpl5a1tU8v5UJxjqWHPD4mK8PuL0TsoKLY2DL91fioAtp1M0jw6fiz6AXher/358xR7DStqFG6
IQQcxXUoC7NpJSoVohHy9qmcuN15M2rrCyVaC4ZWNPmwWotH5jDG7azK9b4bZoYRvy96TUsxtGr2
NSZFvFAthh7h4klT373z/3DX55yeNdWkOgZ7MkDNtwYSWpRTg7eTEBxhf7HLxqzlpitxb3NyVu14
rZnDQyMNbKvba/Yu+6zjs8w7Tr+XY75Rzjx3yrY4YoTxnrTFcZ0sujnxaeomv3Bz8OzdMU5CH/KD
OucVQa6yCoUWrEfc+dELqWwIQQzGYXkKkyfCcYjskD0yKD2KkAqc5qdpWP59r14qFXMBgVjoooRI
vlZJbjLX3xtg6YD2cu9BaZ0L5GIy95LFXSxWvvUsaQ61IR4fq+AwbZVb4YLyS5m0xUg8CSr9ZkzJ
yyPcIypdEk/k+POnHqwHyu2gHcYeQ4E0aWGXwAcPXVA98T+v98ndFA7B1z1DXjRv0KLnmmP1Ijdx
KmAmb5bCgnUCNL6VllSrBgmD4sh7uzLHo/KpmZ0HkD3fILQHSWzYINv720A7ALvxja7QheF6UeRU
cLJ83fD+RkrXaUbb4FKOXtkJmDq0pAW/NPnp4VGLKywfLw/Nf7C4yEyvkBR9UmuSk3P4OsDYDj61
Xi/DzDucrkdfZgwCR038DZ+d4+4YM+zKPc+8BG/RJvMVycr922WXtJveZnIunHcp4i1Ef5XI21g2
Fcqf4Dx8W36om2+RmESMTGAQYLtPNye6CVwlNcsRjMPBiHp/hioWeX/f/0DJyJU1Od57SWz/3izn
apgAjb+eIPcekWQZPSg72dB8MFgZZh5y9unRk+NHuRfHBiK9z/QR3qWBc6nRH/i2UXENrVz0To6f
rEyxyGLFNZ+ibOwiUxySYODDzhVH2w2zhpZE4XuNB+aX3FeRna6ihNVmBSqOmB4MGXSOFe9wFXyI
u3j/D8rr7Wo2uMU1TX7xwwULHY0BHRbTCQWJFcgBG51D2i5mvulkJ74NPmsOEG5GGSQL31MKbboP
w34c0KB1vA8wXmC7vV1fOvG1pArFeeuBO8rgkyJ8F1zdzc+t5MaQ0IV4UmrBtNnO3dIRZLgv/+Qf
qBCbV4a+K97CQKnq0/1gJ1SUS18e4jG7fJjyg86r46vAXF3FKLYlFlR0hDUshpehWCKZbwj+hBYK
1WcZdwJAW5UCZarOxAZPtUpF9fdhR4nZRsQlLCE82GgX6xD7HQzQ/8ff7RN2EYzcxq+89jSCtstc
9k1Fq0xCG4SxiChCcVtoBKQ+FTaLl8RGWEQ8B1WBqQLRaWYik7vLQBswI02jaLT2h6lmLw/8exSR
dRKQIBqxLdTPvi7zbJZ7WM2XsVdbEKa3L2BDGhd4EDTKxvzWmWhS7FwQWa3k0KZd7kJjhnJODsQd
x9s99gFLn/pzSwDtofBrq8U8D5RAcBZB3xlnjz7/WeogRlOULKrIlAjvuyCovI8G9zhEkYQ+BVc7
B8VhvNsZrhkk+47A3iZ91UbtHS36Ral1SMO3MYdPik3q5sZjTFh9r9OVm7EGgncmcwBA34U19T2/
Bc5Bq7uOT+Ia3Wr2SA/Anw46QVUyyKzXy6nOU6gVf9KSQMYyIu5iz+n+PiS4zfQHQJB1wPuEL2Qk
QOstwhqGMxHytqxvCihhjpMkLGw/oa7xlQsVOFO1CKlOMEL9cvEBeqSl/r0gI01h3KjgK3eyFeWr
g2J0jFr6MMU5lAKpqBMFAy8B3wlNXB9OG/VkeWP7Mv8B6RTrC3oJDiK6o7FrG9gMHq9dwPTlG0QH
nApji7BTB4Dbm/tw8xxGf8WTbq3jL7AP2a3aFdk9aL1SyFURqilI6BqvjINrXQbfNiErJJhW35wn
V3gCvNCHNzyNlTDNxpqjr0rZj8Z9tgMuBrLnHEY9KLg2ypHK8TOBEBt443j2/srMYOBIhqNMRlNc
mil6eTQP3vocBri2Oyx4SDEZD5N1Fm9Mc0MviptVqJKYHhhP8d9FIf8nYPJCz1762nhjcJVz3vOB
yLcNS7FyFc0ULM1p1BxSgQuwcatZLPXWK8hp7vVUwQ9qzKPTDYr6EMP97Jyb9BlvRY27YkQaxwiR
xwrPB5emgxZsAPIDrfvQg3fuA6kqnR1u86JK5BmGB1HMIk2QGxLZEGc3VDoBiUa3oQ36e7Kja/NH
4ccizV/ge4GJcKGbCMrvyLHk1aMgIf98KHqZhFEQICsd1o7u0ePT6MrbV8A2YPsUbw6gE99MOTNo
FcNVnv/upSLNY+pt+LyCLwiX0rMUwFL7kfnPH8r7rBfL8Hz37C4/N30/5vIYEcHOwxNEoNJSEPlM
B+a6tWlkDvoMUtWgz0H7YI9Dxwf3tZjX2CDklJ8KfLhozNYMQ1WBawwtUZpo9QZ2QNUuC/JE3/UO
G5vDsHBVVHk1bBbIHbu3+YveEOotJ9puLhVLJYJUuJ0/it3m9WDLKlmvKpC/P+z7TSYatevky4Pk
ArzhoMXY4KSmKgqZ8Ut8AtTozIegLbQvaDlT327eXRdN02RuYlvl37602EuN6xTvYbQzpNhjNHo+
JDbFzc9CLTe7SXwsRVsGAeVMchcthz8WLP1QioLD0FToudDPKjAqCN/Q1Hy0D8aDd7cvjuYIouZ6
7DLMGtQkVb0sxqX8EtuLLdJViNEvos9RGR3iGTwXNn8I0HbTfgadMelxbv6zNlehsTX5oJNCKvYN
nvyfrV7A44YW+3/9qr1cEy0x9wOHCcUJwTllLPfn1kz8rU2cui+4TnE2Au5/6jWAwLhdGmLvUXvg
9630DefU0RP8WRFoEIvLSYrXFt68m3R+4qhCs7j5qgZ9QYLEgyAf1DJ262/MJ+Lh4v3h7XHIzV+f
LNfyJQZSmxNaLNDryiGhmpXJbuv9rADqUFnHsItfwJNiTLQdQdHx+elpKz+l3gimP2gle02dgs/Q
+D2uF72ESkEUyUMpaATKrOuuXoVQ0s1L3YQT4P+tIe5mUQQdAj+4QARyVoxJJuAwnAOkytl7jyBN
juNzGepbad6WWCT5L0azrvM2v8/zVCvaucsRo3QSedGyp4pcrNWAw/DPn0FE0TJ34APxXfLtNoRn
WfZ3dGefGEfRX6c9A1v6uK9V/Xnxf+Ag/JV0r8r01g1lDONGyOWCmz+O10kHw51NBcYTds+Fpaqx
6DhV1i5Qu3FJeseP19DAzeHZbeaZv/Zo76TaLKIqwWtu5Xv4tWa/FT19YkaqR+/8Z2J+YGbcNat3
iKQcT3bWWb6o8QjIPClsR7wuT/owR9K3+ctmhXSI9I0sl4aCqLTynsJ1AqsMN8WbJN7faytoCvEw
oJTenY0tYHAKbKWDyK1liYGeNt3CA/9UOWuRbxY+rkkKgrZk+EKu7hpu0rJ5Iij3Xf6DGFOL5Xah
569vZTju8Ga5/ePCZ4eADzOCCXujAXZLpHBqdkkTK1l4xpBJ79Ayqyuu8m1dicH8Qte7Y7KuDzrd
VRTycIEVFXK3ItYE8UCWP/IkFWXqKNts3OFNEoI4y2jplDEmg4vG125WpScYPqAur+rwLwFGAfd2
AmXvvlX22zpKMcTstndLlNOtboQYV2VnMjsE708Xt9m93F5PK8v/Sm4U+U9rtmZ//qkLN8+bLftr
+ZhYgfg8r7OqSWEJ55/m+feyJJqxwUfjl6qRi8rHSOfjRhTz6arV9cvx0oT4eKXOYpBYrll0Fe//
aOdDhRk457GhC1mMyTpj0fRnZ4B9ezzfqRKodgTGXWqpPyeAIdrcTwt2lfZwJgfPp5UXGGjdVBKs
2LDeFOg1p2SXKcnygQVM2u58xkjBEIH7/pc8cA0g7RFy1Qqk5c+SQu9lsu3iEB7Rrj/NIf60h615
sDygrIw5YUck6IF9v8pjoVzSd9y9VmevGdXN4Qyj/21QUZBheRMPJUrs+0p7xFx6EDrCrOuKEs8e
CY/Ms7ak1+gT/g76/AN3akl4JvPF7ucyFHCKEwWma4NZOvyCU/v4s4yMmwj/XaY9oiAVKBB7n/Dl
pcMQU5P5z6hZrgGDfq8/UQ8oGlVXtRI9J/cSEhYabW64+b271ksAIg3T8pwKHKxbkipvEH2Pv9Zq
LONigJv4a484mlsv+AvEqufELUZAs8JGF4xVLDxYpI9pqx4BfpTm45snFMdZ9hDa0j0sDCdkk388
iBvKpajApxr+C/yxgp9RSVAh7+yJcIUwcGVyA/zLJpLRN5cALRoLmLY5Scn4lcmmO8DlKEkE1ono
ArSSWS0iQyfTRcoeeHEFrRXpEM94PQOx/7KnZNwtPX/JYEoYh9SqC7rXyA17WfdokrkFaC6X1Z6R
/Z++8xJWC1P+kRQKx0yDhExCAxamXa2Q0Z9ySSuRbeIgg0pj79TmOB3uSr2ZKitfhkhb+aRBJjta
wqhU9BBpudrr1cI=
`protect end_protected
