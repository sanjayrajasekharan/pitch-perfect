-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
yMZVM+Bif8P96CqvIBud5ebf7nKi+Wm6PrBYRN5/2fWkf3QHijLXvkFcLv07Ng5r
QRuj3N8i2rrK8e63iEToGzXC3ufukU3efvoAz66/jnAMPB9H48f6UImslIsPouZE
rE6akq8mIXDHMbzTOGmRs0v/Exo/CCJgMO+7984EKUA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24080)
`protect data_block
yMqj/HUr+9nqgebhT3Vy0bwI/SgfWJvPn4DDxfwtmr7/MMBnW9PXORTm/kL8U8Eo
MqIx3JbziVFOeSez+0IewzXwCQ84VUyqU9m4xT/YKexmYuFzAQJ2qT05enCejnLM
DoUG2JdULfAHrSuxp8FGBgr9JUFy4jVGGoC3iFY1LHGCKSHIgHMaPHJEpBlEaniJ
5vJGR9QKoYiCiiNpVvFYBXJdsR2WKZT3XAWoNhAkT0OfU+amfXsoyFL7dDkZqpJh
AEkkCzma3Z+NtJR9r73h0TB9cyDknAK8B8rKigHg/0fgE1YqCN1W9R632Xd9zPSM
/QL9tAXfVp8ILtjWnJQpDaL+CfZZ4DTMsto2AoOi/Wk+u4EKvp1S7t+XB6nWiXEt
Fy8RHXcn21Tv0dNV1NGghTcQRV6QVdK6SiOovBQJYAHI5uwmp+d+xZGX3ks4PMGt
xXGe+BzZB2NGNjJaLNhA2JAa9mB1sgcHBaQZ+e9I4JTaFfIHIria55VExbGtL/IO
vt1eob4mpYH6tbsesvf+EHVKlgSEb38VKS5+HLoSAVWJPUyRE0ZtAqoe4wImw0l9
3YSECVFcX+jsNi9dSYyteT1BWsll0h//v6mBCd2AF1YnqfAIENxyyi9RRzkg+gxl
Ol28o3lDwck1vILHqDDbFO9mzMuLKa7V9oShNWBgUU2exsLr1w4s4xcseQ8EMv4u
j9Qed/f2FY2qakU0lnufJKECPQ9EfPko8pyyjM5WdB7z0GEaBxVIk/ubl3khYvP6
Fe7rhY6JJpLyoJCCTr6wW8sCE68oXWbB65rM7SqptsoobcRfOjbE9vafIfGh/uk/
jVJGT7MA1t3VMlAsaWH5+MJsZjIBCYwtARafMhvUxacYy0Egzi8QV7rawkbIkmos
XD9MIna3DCtpWiPbMeeMviBesXHezzdtuuNwWuDMg4x9Frpexw2cIe8HN3kNiDUl
m+tteOSjlldVOYz0KweEpHQbXs3MEK/2jTDJ/5wSfOFI+EgzfUFUJ6VULW/7NbWC
OECp1VdoIYQ0BzA/Top+VeQydiSXoPwMyLFiyZfEuVLaFQuccaZh5Isi2xDmM/2e
jC+0JB0191vjqkBoqG7gVN+7FPNSJubCCuu1zVMwm545XLMDeUPRPQVjrF1Xtt75
JwAikjF+SRcwF6R5FhJ1msnalcA19cpyZ6szKcwj8HtQmBQZ7Cub0h6MNSrQY82K
pjCIrh4VHkRUGJDmD1tBBRFfs3f7n/8+r/cI2+ID/k/s+ql56d3OVcHLJ1MPfFVk
LvkRHSVzh28sGIudSSm61/crsWjZjmIQMacsI5dpMZAp4APDpBEmmXWWOm5h9wNX
ndIgCyVZVTmdtbc1zDjlDKyAjaMjOQJXbn7JtK/tgXXhtt4QbaRGF6UxrF4jl37j
CZodzO9FWghtvGafrf0G/jrAJgD0MmDVMH6E1zpXukYq7x+wQlv/zs+2XjxX4CHq
emaKQT9iZeI9TpcRhai9Ti/MJAAg97ypDNIgeqYoMauCKzucccZz7tGqsVf9NqX0
fNXkpQk7vP7meUU3R+eUCj+kgXtc5pc0b/vyhO9G7ohXULDOi4lLbPtD0ujB/CfY
hixkhAiXiSp0unHM6MqiCt+g7YAZk0XpRp0nzWsYlEUj4GaaLOHKFhT0z1UsyRcH
aLwRgxCNQvDVdqO5xxG3IBG+HQvie7bQ4SFm5yKCKldxWp0O9tK3p7qq2w2JxeDj
jAeA9+9eWaw2T7ncwPqan44M0JDHsaPiwzyx9NDMCS6jcjH07gOMO9Q5+dX9ZRvo
kAYWsCI0//dC1yESlLGJDjiD4e5V67dLnUAkhWsFOwEXv+knmg8Li/9twkSsc+1o
h6cgHid9XCKgSMdafV8l4ED+s90E2gCePjIEiw5EMOibNrZ1eD5+wrXkAjbKFrHi
CGGfNhFWlLmApceI/YAPWp58R72wccCoRiAh/RXp+or3KXq0vji1wQ3yxmL74TOx
ifqVHvl44uREK8y+NvJOfupJRLptyGEV5ugZg4GMrMKv82ohBcvkp14thLP8tXRF
p8+mGzkFzovdAzDSBWzRg2ux6L0yprdOwodnriNe4Du5hGzRyMwRGDYoxdKKZhc8
McnvVbfNs5MzVYe7WMMQHqOYh450Z5a+c7RijTsOIfXB+AWw7MoK9YOkVbgZaR8H
Iqd8fCL6MMxUhOhOE1cje6davz89w7OFlKHyY1pWsxaEfR2AKL+jJTQbDfCd2BX2
n6OywgCYgIYuBgFTfu9p4cHvLub2SAsdAxa9eF11l6NV8AgXCC/REmlQlq/KRe+L
1wNzZNadsQLEt3jdf+u8A/rLpeEOtdsh8qZHu6NGW8AGJ9wQn3+Jd+B7WsVHe9GY
qCVos4OTDMUbuRil3yAV/Hqan1WNqTxxAc8nDs5E6+oy2PgK4epp56/VaIh7fKCD
8/HODCEtD1H69a1waxnIXLf5d9gNEErrhYNHLg6T2bmjFEu+hopxyrYGwvu97CqH
PRbDOXJDEsSyw2zPd0zauxlXb0tDLUZ41qLdOY9TEay21wVjT3z+YxX0SAH2rm5w
XFqoQtKYBht0/xuxOxd+5FgDYpdtrubKp0RY+Uv4KzZxInf+CeKYIkoo4CSjN+Ft
JIBBu/3bhEnGrh+BkfYMHkmI54OPlR9qZxWgjlDooqY1s4gveT5h81TVkKNqvCHp
YakVe7pJu9t6pdbUpPIW20359D33a/ahJCuvkVJROgfdtNuvG1GOiSjhw5NWx/wr
Zuoh49q2+tRI0cUqDWTbU5+Tff5riUDl6rgdhwgnGuNGgUwktbzWHuXttDKFZVjt
fx7EMqEUIO7NldQ9/YPPjeSs69CtBkT+7wCk7jLc/NDiKfc3H2MIX4RLqpQB03+n
8p7ShFr4tEbbskIgNGquMZM8App+H6yRIYdeoRypQpPbTV0Y7TQhE//TiKwt5JLw
VBxUteoVWWR5thEe757NCtl3CSd3cWhs8xTQ8hYMdDZqAHubOunuttzfvKiK2e3D
wMuKfWSdRAVYtnovft/nIPrKdlTGF0XbVGDT8iTFa6YzElt1uu1P+ya966n/p09f
aW3oTYmmJ0ln5fEvZNZyRI32FOkpIn1/FAuyY+U2Kgzt7t+7ZplOxe9mnWKwRh7k
i6whBgtcn6tGKV0+JJ35NCNsaQFFtaOR6851J3yDM1/SewclqtTFA8BuCZ/LtXs9
RfsSE5nxVzkywYljD7BB5IQIWAySDeKFU/okPCjgr92s+zQCeiz3lQdIcPsWl1xd
MMMq74DOTR6wMuSwm0/OhHFkz8dL/kUVh4Ikm5CPUAA5BuKSCX/0eqbBU0TW6O0r
W1Lum0f2m4gcdHeoSYL2EnEqiRDNhRIXyPASxeAYtlgemrfWsTukpXRqLCP0Lk71
7CCSg4NGAlBGTSVDepJtg5mTJNBwOV6GBbs9EiPksHFADMjWehpgn/PxaeS/b1VF
K9FPUFLLD5+E0FrVzNxgsOCwKeLW9XTPl6hjEAdlJASqMorNObvfQdB0YhnPyZFJ
Uwif/fOEI+R/z/hdT2qhZy+TTh3uz6ziJQI+Dz3/nLbaSzL9ur8R55Rkoulm5l3o
qn+s2RI4GFFqtqyt3R3zQG7S5VlLbQcGsf1FzATCpEom4kyT+FFQlS8rkuO+cwIx
Gutuf3KXJonEUGClXWUjdNiNfYoOoEqopRjyZ3kbYJ0F3XGnpa0pIXsp59I8b5NE
CPr3kroHWmVOhRFqHXsy5c/Aa2JBUHUhsIElI4gVAO9r0BHvzvb6eAP7HNVb8r9s
aXg4any13APtJVHbvy3zfhhVN5eELssaPmJxppx7GlfVim9lzQlXUjzMtTvv1aDy
z7m9LZAH8H997D1fEzIMgyVYWi0/QXtsrmeRnqoqDdGkGcM9oeVykmHT2KColvmt
+mCmrssGIl+NigMMEwI8kG5xoRgwZp2yf6XxG4GagPrJlcMzfwX88mt0eMQBnpiV
CopBa+IOOJeAfDjXs2DKSWucRh4pwmzLQmnbtbuTqRZGqgBn5eu3/ClzcZpm7N+7
2GdckAevfcR5DCvXH5NMdvIueeouLuYut1GjciUTFex51LigOT3UGVtatZ6g06cz
5SisCdEfCeW/1v58WT7drODKF4G2Xn/F6WdHArahbqzkr0UVEYeOLRiOat1zBJZa
O87OZyHDTNvrD2cFkuPHHM8ce35Dvo0msOFSMWivUOEk5kKRYhW+75EPaRK0Yy7y
stGzNNus00AlHqGh7Q6XU3ks90tq51dvkM2UmipwjJdSP7IjQk7ZXEwtVFrx6mfx
zNqhG8zvyaxyuN+JyVSrfmf41EYZZDflRiv+MzE6WA3ki+6ughwL/sdWnwC9G9EP
CaECHVfEU/IOCUptHmSdXEGxBSLqUqyetJ3uaSHbWqdu8WCjwIKc2pYfJ7FvQCR3
2FLhDtDULzsTC4cszoNzMa76wh0YwSVrSGsSj+7O4VoqQtYg9UxYK+owp/E/sFb3
zkKgj5RpbaEPLYNwNGvnuRXgYYKfj2BWGad+p+46YCr7ZtgVlx7iL+KstHVJXjYk
F7YuUOHFw9q4NGQGfJyIyc5rP94tw2wZ8J4cJBz7mCXmH2FBNwV84hSSsoPhCuLY
FfC2fheFujZTgwimbQa1W0SiG/Pg2EcMaQ8sLWah4ohYBC0jbbjuflRUBUyNivnc
9d08WFY+IVxkbXxli8AWLXt5ord7cKqaocPDHy1TM2oO/UIrUNLV/HhnI8hysF31
k5j4Gm6ETtl0fTNUvGqrAHpoUqRSSiTXhzQVTFcXwukWZh69i+kqByXtZ30lWrsq
4n+iNDnwwWn31xZxOl+10H7gAeLWpLp2NtGa6fECw/37XdkOqoamLJNg6MirVY7y
Q2FGY7s7mGuMiTu53C8m+iBOgAUJz0KGN4oMY52tzL8G+lQi9e/h52jCKO/1t5c3
2L8c+GYEHda0JNeUFxif+IULlQCiF0VRDRgDGsg2plLQiqR8YJQNNmYnU9bxU02D
NIPHnSqL456t92u3pZofi9RTROazHUhtTtjeDCaGaCNQmstgsCy9N53h0GIqeq0J
vTNFcQkkWX1jvte6E2X9ZnVp1YQ9ox18vrc9Qdc3u1zyxM/5p84sV1f7Ot/CSY0P
mRRmZ2XgBhQjgd57wtFcy/gQKAtIP++woCXUCkqWA3qYsmVTzxQzrcXthHhN787r
zItlbqLCr4E7yt496JzgWl2gWc+mEV5cXeths0p0C3Fn6EX7BEGjd+pet066+pBe
qR8wY5WcynlTv1zeEdXDtcRurjsEbuHr3HrEzMTPB89ujKXhDUDpzHFWPiBJH337
VDQFj5u70f/FjIrQ/C03VlZQJS8IraoOOpe2kHfipZEyvZ8I754u43/99/RGW0bK
dO73pzREl8MDDHADWuEg0SatDuKvgpdVgD6ty0l507zw5LjEbL+inLuwdGHO3ErY
TMT6bSsRr3pNRvjd/afYH/dRP7oDwHkpAacpxppct5M9e5S0xeFMy2wnKM6R2Hqt
WJjREubzOt4/BVEvpJsVaUVnp7anOGXN8uCygZ8gejMTSTUiDZAZeuKMvKXO5/Qk
zVRtxHd10naKjVXi76E/9wSAzaI91JaJGmrXA+wTiLO0jbfxmzVYOyxjbmpUjM94
ZvnWnhiVM7Qko+d300A3jwZHqSs9v1+UZCOGh7nQKepjzbEUcdWc8pLHZp8fjzHA
Pr8kEhDEDBM/iUBn7NCxwlPVfLIgr+kWXQwz3ecA5YHFdC0P4u8S2NkMNYHZcLmZ
31DJyYHJ+vxY+RxFAI/JB62JAbt7cj86z4V8CaWj3q1QEr0Bt1+L9M5oP/d3GpJy
LSTmVpmL4b0gw/bkd5ypjZxINpC3KJm0UmBuMnt/xsSlSx/KDkcf63VAfiK0EgoO
6SRZxhnfaCp4thD3c9O9jgH1jaEufcMSdWNZANcVxUJLQDHxOIclXgK+MZBl+/x2
hX6Xd1xT4P2S7UUFds/2H2asOziSunxymmLYRhIOyFi6Z31U2LlMs8UaJSJMIkbT
iO+t+SJV3y2jGhQWlL9jhtbZIq1PnmfPSSP/Taoq4i6WDIspEFSlcJ2LMR8WtMAM
D5BRp4f+s5qAUBD+3a7whVhEm/YhW3hUgvUIxGRh92umvqj5SRf0RdmtbQ7R3mVU
BWsTtzNiUG319b9u96iz1pAskR6ItNckvjCKFdaQugZBRzbmXIy4j1Qp97OGUcNl
wMAkvBlCAmxFq1RHjoNsi+SNJHXRjxeoKc+T8mQ5/QomrrINOAXbqM727PaeyAW/
jjSHntV91bTf58DaGjhTIzuC1sJ+QJbyu2y/RiNt94BVCHN/alRxw6ZFM5yQk5eX
Y64SDIyv2oe9Lbv8vpfLzdJTL7Zlqw/Vse7Ck/k36nEbMzoc9hOdUYXLrXUf20TI
rmpEvTqQm9BAyx493qEifwXJ00/e7ojFkBi/tFolpS2xISoYlLFDjPGWdP0W45s7
xO3zs+Mq2nWdfnC9/MoqSh7sHFZTvpu9/BqOLXaX95itLeTL0xo2rAHGj6btVYB+
EDAemOLw3ehAbf1Zlnqsp6dQFqYra4BaRxVMUTeg+5Lf9X0wSpm61wpICqPwCk0K
Qie93wsnv+87ZqimWEMCzOZYMIG4r5JiNRR9AEB+9LWdxcHXN+zdejfftQDHz7iv
Sa468200ll/wmoWzNnon2Fa2yPlYEcY7NiqSXdIeQlRsiUVsu/NKWSd5yLxaa0JF
jaNcKHPGjUEMd+p86zOa+n/yS1Tf/cuW1j7KT7utsYNQXPMPjG1Y5XxoEuekyytB
vdfLSLa+Q7awrn55APporrItTn14krcXN1TbEqug7VhBxNvVgW0QfFnbJofhh0nl
1S6BEoaRdjAqcWXGk7bAMqa9CbsPlvIUXYHbRrmWIJ4cCaCQRQkBIDZ9Y9kWpT9Z
PTQa5Y8knhjYzITq8KZB6l0B0fl4Y2xnnPxvRJUwDRnOYq+6H0l3MPvPv+OpwYI5
mm8MwCS0FI10qmXooHCqXtPH+9XKV0mp6fc0sv6Pt4z4zri5BCI+liaelNDitsex
dUNonI134QKnrYRD79haAX1Kaaj93+TjrZcZRNxfAtKEol/ksuz5/3WiD1Vdzzhd
Xcy2gO7tZjQW1r0kKoRz+DtO2g87W0Qs0LMhmp9u6iaKyguoHOIxdTks4Rr1S7/P
1ZXolSu4SBZ82zbCeOCcUEv0pPOXQlzh+1pWVgznWvDL7kehrfgjRoRAjzQH8uvm
nvop7+Nleb3iExfTtOCDaA3SOwrf20xNVrWF/VSNBgWGhwcdPT/DxjGq7CCCJrs2
AOq+WgkD9+/cKZBfjBqmZPQPnBN0+RBIHB+jWC8f4TlLxZL+9PSJRhNsi6RV3WNb
8iWYniYkf55sX3wDz504hxQgfktVtVXEVFQm6ty28BNmtiAyADcfU7MlRzwxsLf6
YO9/gWCj0XnRetvj6ujONqoanG96Q6cRZjzUBHQT2C/5JwHbFzW8BULl29tJ1iOz
iNWgKpgt2rOyxOHVn1t2KD/dT3v3KJ/9wRZy9WxLejzJ57NEZto7bk94u5XdOCcE
FOaoUBYtiR8GICgL7lfEQ+aceic7HWdLqtmEMlECSw/4JSdCUWcLfgdS3fWnci2+
e3UTOenfFmndZUd8yRw/BhWYhDybW8I9u/xg9Kqtt+9UEtiOo+88Xtg4RDbebVmt
JYjDyFNlPKmYyB451rw77/C8e50Xm7AXJdSyUfEOg1UxO9Us9/dSy08dBsPFZ1uA
coBFQgXKUspk9Aj0UO4QwIIrwk0/YyasRO/232e/TLY5UkZH4zubMpeDinTAyWwT
ZVxSiKx1Ejaala+KOQ1aB7Ulu37A2Ks3syWlgdyuuBmQypOOd7Uxh+7XJ5o4q+3C
qbyKpV1SAb5UjnU1kIWyv5aZpXxwYMyhp6ieyZFx72/0+pIp5LDcIpftnj6zZbtj
cdSYE17+azF1qsV4sVWbJL2WgPMAL0Z3tzn/YhlbVEf6al0z0QZQgBC9OQngtAW3
OwGKOGk0fffBKUxJG7GhZBGy6VOUMWyrsziU3I6pym14+Rg+EGoi3Grn6NMJGu1d
xDirdq+zmDRnthL7fpgmh8K9KBZx/W6kF7cH8r8HeRLDTGKCH4RCUcoyHWvjzXcB
+U/guDT5S2jg2iHQQVisIuTBA3Lt+SWt1mVVysWWDXHKpnx5JopfVcW9wIdETkLv
Yv4jPI0qUup9KqItwtln50KbkaJiZge9dgpXBHQq1pihjmPfo9fQODN5NMoh+4zr
6yXz3A3vy3FzvFiVnPondJXdZhW8YtcGDiFm1gYHOEWXyIbbHqLGnhWgHZS6ljOP
DKqoXxO60X4elqPSerMDizwVSFteirr6Ho++4VDZp83Jbb4C0mbu+JvS3OfIhJFX
vEu1kO86mauyxXp48C4nNYgm6lzHTvwe3T53hoc8/uDwYVvsUbeBXqzcZsN6IycF
MZSKDY0aiWCjNF6Uo7Jv+Mzf/kcmCbsd5MzOArLYSegpCsB7RcURwQiM3nXF21wP
+t5+1/Fq2mHPujn5xZX2UNDiRvrEpXr1wa1ozonew0yMKee7PBOA0a7n0Ihys8t6
APbMe9WGldJs8V7IQk1mZzcVDVZjcuYngbvkcN10b8AxEDQe8aa/GJhqnA8YQ6PN
qQnOthVv8QKSO5Yiwoe2BK8catlcbseg8SsPOJ18w6kWdZNNTE47MSCV4C5GghKj
NlOpZebZbWOLyMKNXDPJubYjfdr5c4HPbnH6arKLrrV5Yc3Q13ZAKjag/S6+6V9D
OBTdlbRKbnXNAzzPNYSQNUfHLnSLgmp53IRWg2GHwZBgWXyvLKbD4qOCVr4IDLu2
Q6V+6flgXxdHQE9DRpz7Wr0uOidD5cGmkxDelW9T+6fUV7v2mE4ae6TmFGenzcUj
DpV7fNJ92mdxrx1rxjcsF/o5JMGubobRIbeOj/JekT6OFoZH51/jm2T1XedoCLZN
9IGup5wxAcq88LiWR3H3LCJ4un3DG0GP2pWkz1hpba5of9+9Mgd9gECY1nSxQYHs
/U0HGv7QO6yMbKyKSbYa3SdJFUKxPqGEQliGKr/UOrZdaKyMIH0DSi39hdXzNbBe
dJafXpAuZGd0rCqlonKj3JiDdNHOa+TCQ+iNXsJh1SDUY2FMHiHbAYuVSHd69lhU
3nf5uAtLqq+G9KaZy/KIlBvXIFEWzO1tJFPwPtW7ZFTK40RVmy9vgF5jkBmL1fWn
g/aW3ym73biwR4KJ3IXzIavQ0wlK9z6yeohVbjncn+ihnAXhF/sB4hLBSFmU3gZS
E3gkqPAbtKbP7rf0uReORuExGacqaW4v8nFnbwn1kAZ1QKjbwbAia+kPEl6ppi/U
CuYxUiUMpLTli4dQlpUfNoxm5xrP6DYtytO75VpT4p35uS0sv4ngNbpUTjhN8KuF
VUO4CArH78w4kUihBvDvTrTD2rOJvPV9fdIq7e/lyFvKExwYCUdKpx5mK/GmSphp
Tp03CMRiCIj3zM28lASYfVT8I/da/y00Htr0+lY4go/BQXg0yjPAyiyTUGSNC3J8
0AZwditjfmbypPwoXgS6M/SFRMWfJbghh9+VPB6zdM/ivaOSIxyvG+iK22GaoeOv
Ir0sJ9Z3nSQMM8/al8xgiHLu4rjRuZTMfZYCUduhgbCn74FNZcduWRP6R4FAaFyq
QgFqz594/1EdmQqAZBDq8rFEJJJWIU3FEPpqKDffnGnj9KZLUiRW3cB7HtwLBrFg
1DoL7yEmKzp88SZb88tB3qhDizbGT7VqDUiDiogBniCT4BKW4M11FOOQzzM1OjAZ
Al4tOIkxptP/y/H8D2hHEKD6jDg4e7LAxTtdGpLSj8qQKrktMTB/2RVF78YHVJwU
WtD+vsQp10z+l0ZdIvMljBILlacOinK/GaX7Uzemr6J8I4FTE+bdgZefXGB9XL6T
nKkiWlipt4UzxoW4DXvP6NLSmsfeKO0/Fbdd9G3CYq2Hq4vVyncJMxqWYBseE8F2
tPVtXd3R03WU4sTaT5vsl/JGKrVkJaSK9LrEGAvmUi6JQPiVh2r55pTmAlQPYxUX
kMbGSNoE8Xfr0D8/PZgYA3FNe7sQzg9sJtVuwdpdrw5vbAzW8gBK/KyUgYf4eA7D
bRBLcMMZ5fQLQpExjh6ZcMM/GeqOovglrQTDHBS0JOgYOF/8ave1p0Mxn06Dg8dA
l7Lbd/+mUuh59DBZIiHT7o0YmqB9k05yCUpc9zHma6siwAoBjYaxPnA0YuAAvNxv
wckVRY1NpYMTvZ5bWWBY1eKUjcxqbOOSXnWNOT4T6drseY8bi5qgJVKKXvpp1n23
CaYnxGA5Mni5b8TzqEJAb+4h7KQFvPuSULh3eZ+UTTEI5lqW8rdjmA9hNsOLUL8G
DWXmEFuz/qGUtkOMScnZrXzcoSbC42VnnYVXrkrkonZ87C1ZWXrhTMAWdtAWDJbG
2P5EqGXquIvzTedsdo6m712VhmkiaZzaixouy1KjqtdisYULQx7p/MtPL6kbXgAJ
rDLoAIgJmQIvw5Jslcuol6HbtmkXlvbsFausFNEufuIMSVwUOb/O6rJsR2jYwUGo
2XcQePtnlUlCXSWaXWg0NfaWNuzZYTSMRunkoqrAOknweFNH6ut0NHFL7pGvpMRz
c39Etb1LyhVFRgDodfbITR2qy3RZwV76J2jMDtWmp7t2A8tie+17CqnHaOOhTzNh
z9G5BHaJNTCDhvPumKHerNqAwlApd53UjFRPX3E8XSZuucKrWJujQCx45hTvbpJJ
mVQi+BAtfkkOtfwwgnJMfSvRvyQflv4Gtbaj13oGHi+h9l/7BXlQiqxrjER1rplV
nQjCLRDiEVUk9VussaVdzvqgKmIn6ijf39hkjT2z5LZ3rdUkjDr9p9UFCEW1FXCt
zFU9gMTtW0u/56McH7Gp+NjDtrEjLGvTEpfPFwVMtHUYxR2AUaQIIE/IvF3e7G07
e/hibRvoEi0XZaOFVzRXYhxMXUajnSntUOrl+7MpO1ZaHVW9RXl+Df3NFh7bRsgC
52G4P+f3ph1Aves42lEsrQ2A8/j2bjX8BCTc/s79pwWa+XgLwGSZjEA/hy6EWKNs
OPLduBlSlH6FvMFmreeUw5DURzBh5kYdWbM/3BNjcL72NcxmePMhEy65iqFxESXa
8V2yYQOS1LK7s9e7ncP1fBmC0T6SdmZGbWxUQjxB+UWHun1vgK4S1OPxLqOmR8Mi
UOfq1btRDXuvWqt9kkO0e8so8QgXQjP0lvkuaAUsa/bh+3o9mp0uYpua6G8JOorF
NEuOZAnkZJ1ULmMVnQBWjDeMdtSmVXaidFoRq3/3oAvBm2o+OAs97cjpgxfmiJlQ
RiG3bULB83XipoAh8C42V+Wp5kgJAti+2z6cA6Dy44rErKXREYKqcfIbLIsV0zQs
O3SqcTNJ5yOYH22YNcJ61vpZpAfpUDvCzLrhps1mZdPxSCqdhmE6IpyvV36wKGyz
j8XHJxMdgDqZkaUeaWzgORRYqSnOlZ7T9SaAGqk7JDUPvkXarENKYiNHFAvy7qLD
McNduZmOO5v4FBvdr7QJTlRUsHgyEGkrQvPQXH0IEt5nGt2IbOYT+yadmU8HIYs9
EUMh41OGjCClDKHCRSuWTrBTW/Gk3mcQGQX3whcpvQ/c4ZD8siqjHOTipAl12rMB
5KIegsRw0evK/DbVu1ZjQYElW0kLBj5kCwJGBEJ2UPO5teaLhZx36ATnzl7yyKTF
hBZSwcO8hFxf7f/yVAF/E3cxAsutowkZNTJ7YeV0m+Zlct86T8Y+fUm0DZWFzeFS
5kXA25hPuC+7oomWkIFSjh4ldmjNWg4H8p/fD7BsMF037BRal4JrOJMQVfkggMCa
K53DUuFnNizrOiLuFxk/nPA8lbYiInK+Ml6vnGjgx0i2wt5akJgNSh5JQVimbBdi
j7rxhb/bJEJfQDyGy00fgbcUVxIWZakvw+nJUtsFP1wtru2W94WUYMCF4umfDFmQ
cCdz8lGLIJI/ush/pTY73J7wrRoDfciNto3AVoJP2H3Ef4SorUS3AMjtnTOAnsO5
LEHt9JTgF5P2FSTnFXceEABA3HSYh+3IQjNZ5US/0X5PUX33HA/OlsjKns9+zNEK
E5HNjSoAUXVRiiH3lstF121oHAipJwXiYajKW3QEaV36f8HE13gGiU+OfXyNZTrL
l8zKdF7U6cOuJdZohXKq2X4UhXn0yzFIEv7yH9mqM/AhyonQsO78ToRzRhBqjhlk
10gRXhAJXQNPUogKeiKWNscKAEY5n1bz9etGYj6CQgWTvtk+TsJSN+BREqTBqz4e
zRJy3bL3qagSx8a09C9l2RLKt4vUyJ4zO5r3YnZqRFXKbdTY7dZ8m9dPVeY7Ast8
AI1di4ADlNI/l60MM5NEqbfdCUOY9BuiOwpCdRUoWXclZQALLMz0VDfDufArpeua
a59zNbOZ+nyV4fIW+5GncAZh2G5PaKx9Dt8GqTO7s7zE2F6cxxpwXXWa3f+Z05os
i1BO4kEnJ/m77OxO0fnpiiPGw69YMffL14FNIoxSe3ORivUrOxBE8l34qlmp+v4J
LdK9WkNb6ZSm+WmKA6LO6rcIF8IIh8+f1sz4xV/8YOp0zSIL/6Xpxfbwwtckgmwn
gs4/mUD66k1ajVrhPnMFB6USV6d1ZoFZk2ibV0HgM2gbroDIjNBYxWuz5ap+Th8g
Aw85YGGOzIR4qjaVz7Jr+gEbyPi9+6EXPruoywv/bP0kgI47cm0C43RB5IP0R4Nn
TjnKq/BWL4lNIfNG113k3MysSh2k6xGerp1p1jQKaSvjHzRGrmwnp5Ej2kuPyVgw
31WwmLu57REu8cYu3IAoKzgh5idZseSirr4PZ8vrc4QNE3oy5jla3gIZqbi10udQ
KI7vGzCt6OLK1GFm1cS11pK5G7XvOBNbNe9c8hj3ftykw9Bnwth5F27uhNzzi4r0
M6seJeSTDLFGJ5JRe4evcAWzO8cauUMYi3IveiwsoGFwFDTIx5nf2bZ9Pb3qRYjW
HP1JHBpmx07pZozoZqQkSqlkiYqyp6vW7Pw47Zjm0RVXhfaIxqR9crnVUOnZzbDO
hs2+1Y8xxeNZEvLo+y/+Z2Shweq10tWPw8yCHACbRmevK3Ve49VB3zgwwvZMiI4G
MOuUxQxNIj8Way8vgzUSKRr3inkSaWp/UfxgyFOwAGqSOhmWGI1krvmpReo8xKOq
ODAGWec+G9o/jYaHLulNBQ8EZxXeN+K8Xb8p4ZlF7HhoblNxEQxE4DRN2TCZOFz0
L1m6DomUxQaWLPFnCbB8XVWL3pEZOkn3rfkegyF/PkKYKA3DvLKVj7BDuhS/V0NF
33sYsuPrrvbMGhBfs7YsJ6TByL2ifHgv1/RZ8Pod4lAlownuWuxrJMYvOSpsKJgl
O4nwH3tBX55DLrBAZIIMCv0zNus+F4aG9ylBfQH/VjORU0VCyd8px8UVBcT8urT9
8lU1/Mhb77KiSGTw3Ryov7UdhiDR3e1kYR+EWpKBInUDuQ85YTM8dsPINE+PeZxB
zD2huIK6wF5SGUzcCG/x7qxjGwOHWYeE7S8ao8yD03ILLplJMYNyBpSRPz3SrEzO
cLYemTbrSkE0TYXsjtR1wp680d+u2RL8W3xPg7gy8yPAgi/Xme9UfvjIuScR63Wp
9Dn6gBZI23vuuXPEwQ7q7et2+q88WCG743ZVf2ZYGjAGxjyUNvdDDb8VfDUw2X/M
JBGSv2JBjU4Tv9KF+sCrtY0nNz5o26Gs9uCApIj2wUK3lLzTYGh8zNdh1voKH+FQ
jZHaCgy1cm89GwKGyQmxNHroL5EZgUFVQAZ/M7up+aZ1E5CGt6HxCGrZZWpmQvow
dHPObaIVi74RG93eydMU0KYpvqPXdIK9R5tx0YyKpw+zdTB3YjO1N7FKAf3pFNoZ
MhLSJvb9q+shgP2SXbrO4oKyFgfWrhP9LK5RTY9k6rgGbOK9Cm+R4hE9cJrTDuE5
ydu4gtd8rVh/KgjbwyDeQJl9GRAbwThTMil/ikcSMfzytC5xFtlHYUrX1wYmaMzt
Mi9byNIZ29ayZQqFutpP1kim1KxS6xDBPixDt1naTmUOIn1Nz+2vE4waVGV47hcT
dKT7IqGc6OYY67PbR6iAXAZELJU6bfGfHPrCQ3GEivfXyHAKTwFqTsUDqiwXx5ov
CO+7zqcyuTx1oRcMpnCaA8kzqyUGSidFrS4V07+6UOQXJUa7igdXHxdkRgB9KHOu
HpMoshE4RfR5aFR5ofvKTVaaX6DR/p3YRgYhk7UOmZazQoEIGWxP7Q/LhvuiehlK
jqC+BSn17p/KC501uEPnPGjdqzFwc2vq0jpO6BoCv6l/AzUhQIBJJV2P+9ZuafDV
ct9R7PbWuJoIp2JtjShR7+u/GYyZK2jvsp4PH4d2F0sbiJkOsB0d/c6Tm48rpAa6
FfNFphNyHdRe+QjpL8g37wnR2qoqo65xg7OVk1qCS4U5xoyI3OfoWX8abuJLmkx2
Z1fu+ESU9e8Br3A1M6gaceoe87WsopRQSqlxM48HYrM7+iuPasbnEThKugxkQN23
LOTpVZUSZcI44Q1C6hLh10A1fn2L8/2jCEg1bF8+C/GQcDTpsumNo+WLvJVXEg2i
sRogi8QTaDM3+Z92iMHVwCbjwZQgGMDDtLhzQxEgK5mxfCNcNy7jvslsmFUyRlEP
96trKI9r0O8Gucs7NF5eHxbAB9v2fGZvQ1HGOdkah//ijGE7EwCC5TtufdE10/Xc
cs9ag0D7/e3YKaaeoNAwgoX5hdcw+fnvnGb2VLByiF/vhKaC+FojwM6rBD3CNcQT
MHLDzWw6Knj+teoNt4nNRjVmlXswApLiPxx+JBbm0+aNcfOfX4b/nOxEh+5q8UZx
Exzbck3yhS4ooDmC6EJxF0LvP9hHxRWdzvTKD7VTPk1uHXeXNDS9yah/zq/oNrK4
hYvsXmBFzRUlkS0az0MIC7h+nPIkszYvzJdv3s4vhIK8vSaMrIL3k5ewkdg7iUDO
xljYLJjWtK/x/KkUoC3NtvvuslNbj/xT2giGF4mGUXP3ffq1BVoxJEr2je5oKIMN
vQ5yR9Kp+Jag2Defii3dxxoFs0UKseZ8ejp+14Nxs8FjubI05Hew3ggO0uDjH3DN
9L7LJrtBAsryXyr1NHsWiB1lIzIKEDHnz+X4vXzAKkx0k+OQpBc3dI5ckYUBumzM
3EzsZ4ec4Cb5uLaQL3xFdJvb5LSXcdMfNMqjC+omiQGvRGnf6A0Qv8yfA4l8P1IV
NqnwWUVBovqEya6vQdPwoDLx7QlDD7y5Dsjp6vyV/QKMtFWXdSfN1L+zdzM/lpOt
KOy92C3b9kzNWXvPSKMRsybdjYItHOvW2VQ1vQXh5FN70VwuM5R080oXDgofAOoi
zmpx7P9UZV2oEWOEsQ/lJ/JUygq3DGOO+KCrYgFjwBDyeI6ggLEe0N7NfH9XoogS
V9iPug2R5XMD8gkhzRPqHIItwYjbdeo8qB7OVc3ALSTu9Ak8q1oixam7+VH6RKCs
BFS5/De7tGwAPsIZvidWAymKOVcTka6yMmZOM9jzflPL0CT6Fbl5aHoooHRwqjvw
L42WhWe/cGGu7bOytJ3zrPVikBe2HaMMwX2B0de1uyMckUDmN+kT+7x47GUQsJY5
ZS2cdBEPNlSAsyeSG4qewvHjA3GR32RS2WmKualXzLun3j9PG74SkBmRh4IZZXtM
qa3a/YgWq2foyIZVtCwljaPIwqutXQ9hgLfdKKYCtI9Q6e0XDbBlB28zcep9KJgv
WhwlK/YGkjVAsq/RXf+4tbeTjehEAi3LzUs6ZY8ALdMFyXTV/H0oDhVm4mpidps5
LMAswjveOPlBdHcv3xdvm8QW62nlJXtqRWm2uhhXg0eHG3ete1AmR5BK0fdghvNc
4ErHDCMl7UsiMbiQ0QVwjaD1ytzLcbiStpm+g30SAMBTbSpGC0xVMCRrYhdQuW6T
+Vwpwv6CaSpgZGtd6Ka6TJ9NT7VAGgAyqUv4H8QUohnKz7tcX9DX7Hiu1e2jk7Sl
vJpP6gob8FsRgAcU4vDRVG3NsYjA2ysKFN2R7WRhrFbQOKWjkNiew+RDiUd8aZHI
wph4LEgujYRiugALJ6Mj5CXtuFVpFFV6NkYDsnFw9zlY6PO6Wam9DNZUMMVc3b7I
Rql+KtcEMoVBL5R5xV1SJgugukKdHqa/kYQ81wSVV/lnJhWQQUxYD9wBqyU5Dky4
qDsJ2RynrSW3xpKnzHPacM+os8wd5AtdbUNS51IAm8/FCQ0xLpMOZEDQd/CBkpv6
KKKZaQSRJYWEulqQhlPX9NixY2wzuCBNf6z9JpKoIpoHtwBPI2N5R3QQcHP6CPu4
iHV9TgZhA6stGjtzpHMsjhwlXsXyR7iLaM8LHmTcSWF/kdr8ByKCwyHTkgxkQ2ws
c115Vw5hX/sDjazPmaW1zqiInJOBirJNMcyWU1KPcOZApHN66BrANAK6dWd9GIFv
WJCPoRmngQIpEdcdg6cloARdk0+5lMkoW7Z6lvuH+r6W7GgKGWrd86XNhrNB1WOQ
yXJAJ0+Ao8Os8leA3SRt4KgrbZ+Si7emDC0qrtiBsCUI2+VDrcdsQrkzGhy+pMtC
otbONEycEP+6g8xaGxFxi9tWh11/gZc6aQfITQcPodEu/guOUednO+cNySaOL35E
dzRPP22AiJFq6EuBUBdU4DFgoifFoL182cBMqz5dC4ay565OxziePf86SRMEROcZ
RmG7m16h5BkFIHQv7ehM2Ga5xHtmWEZgtqqXuLS0tXctFzY6fqE4lFnIrgeXs1rd
HPbL2y6pCBZjbz00MmzRuj3b7Y5qFDR8Pe78XrCG3U+gLieBrywwFGFHOPmOVG4S
hg9263TwrJDPR8FRhuio0tmY9fv0AHFp+bkNNqfovWhJBjZ1tm8gxunlQYprqxt0
+EbGfYvL94DwYAj4xS0ms1K45VxrKr4aehHM11QwSR5FKnHL1IQ+AGPgFHZ4tnHs
dZgSbAuS6WkPOklD1GTyTAtiq9ZeSnhlXY3+jF9scsgINUGwlZhvJW8n/8wE0iqH
nXecxohpdUzXoXsh8/8C43hBM5Dz1YhvfyG4c3b2BMjVBTr0pfuHskQWhi21A7O0
UoV9oRztuiviX6knB/XopY2kHaWgtVPbLCpTimse8sULcf6X2StDdd6j7Wnwh7Hb
ukKs9cNAVw1g3mtvrYZ25qRn7PhYR2nbU2ZOzCrXeAPyPoydilk7owR9JZlZp89F
zuf7f2/hYCUIxWjDcFkn+qqEEhm3ec15fxdIf6iRyzGDRfsUqnS3QGdl6XsWJ0Wm
35qAmRWv8QjWEvTBUsFv25c8yNzH7Hr2aqwVyTRInRWdYAINzA0ULWM9TtB1J9AX
T0MnxxZFkLwD6V1i97P5a3bUWVNvThDRhzZWbhjmAugPtOuZccCpGRBEyuciWePD
u/ZRHybIAJq4TbF/RYiV4h+O9rMKL2MinNDYdGkU0G1y2BLerZ0P6wY5Tn1X2t2Q
zZcg43S4KL7ATep4B2bzcLOMl3xgFFBQBu1sXPm703xDVYzGnNnqGSHvzDfr0XT0
bmfo2PZN0l1Q6NvyFJBDIKByyMAXTVZRLUwP7BM5ao8aJe+V0GD85nmPMLPAeqHJ
HCZl5xe4GOizhN6OobSYjgABfrXW3oQYr+3v56lLZyLP+RrBDYtxSQCnGrK/xqI0
uRfkJiM5svtYiTkj/XhqUVRySBJ2tVwfXFFEWBblXcxr0ILb72oJEW4gRz8MAShM
Zh5a1o180gqAGVhxrMExZlLIpZtQzdI0pAMr9CEhwWmvnh4U5tl2+FEbgS9YpjEV
X2joUerBBaG1h7Xxfybq4axjsa1W/xKOZjbSboZC/jDyHjNYxjnsoCeabgB6mAZ+
jEI3YzPSbpXrT4zQbYQdTTf0g2HVYIxlGUqCsMceUcnHgrEbC9ssDD6tGOsVDkCD
JN19aCxrKq4uexXIDGjJfGkFJQvrAOFmy2n+GcNdzPB4a/aSDbCJR6mGZiT2XaFQ
q9rmbyBumfVKSG7eSuEQSW4PO7NsJ2jpSYkIcW7wHPyKCiJiRGxlNUvpAs8wOBzk
D8ApP1mLfdmvm7tNIfrWmEvx1K850x4008C1ED9ffk0nCFbJZmCrwCn11oYaFtgc
88qukOAtjw4k4lUkZxqHhz14xOwfZ5boZfALD0EHvs0xwGuazL2WLIXOrsYRslVO
y9N5ipAgKyenfsQkkICSX7fmxn9DZl6i8w6fzGbsB6wLMcjx94AMrVgtPEP7guyE
eMELAoFvPMwEjMrCCj9X9pIbWmdwSeKCQOEOSwiPS0o6mSPnFA1fd6hq5SUyzaQ1
z3XXFCxeKibC6qPU3WdhtrdL3KgMItr5SWRNpNX6EAKmGcsTXr+ylrA5ysBLKX5O
/5AtmM/ENowz1q1ow2Z+D0ovQaD9WYn6RRsUBPBGO1eDk/wYW7W9+RK9b3DvmGaP
KMqQVns3HYOZeIz10IW5bNeKBz4j5SkrlL+6lyDWlpQsHEezGv3yXlvPgfBkWTi2
naX83NLodbrsqAT4efTKh6Wg6JqP/uPL8/crv+QqWqdfke63C1rEVn1ydjYLD5N4
8YIL2AYQeqfwTE1UjIdXAJgUbStG7oVdC4jysQ3uyMHhJeLLjsz+BdZD9soiEUZW
UzM5QjFf8g7F3zLeaiPkR48pph/Pel7oAkdhMAlUwJOA/cIy43WWM4X5l0vi006A
2mjyX/BYEbuo0JQ6lhlDSavIVa6uh2jeFHs/X8XQOGXnVWJotf1QO/4KFkQ41KA3
m90Ycb7vQAyT3UWU7b6pk8lukGQ85tE8Dv3QzNJ9Zbwsf6vO/wnnPGy5JbT0bYpu
GDd7U2km6WWQRgBGMZchv4G0cH7qKhi5NxNpXp2K4STI/qz75XAViGwXWZ13NZDZ
ydgukXK2sBthCw0cYgv2lCDkfYNzcVJjzETvleoeOsKCGfpp2aWNoNd68xaemqEm
kHGjyzXwZ7o7jEn43RjY4gpM0b73oOVudX7K8bgIaX9n9BIXUX6tPZao6q70H0Wy
5xlAV8bXXTmihpYycHfS9anCLRgZarHjcvtgjuxkAxBPlwW+byEabLEp8Ul6TmcZ
+Aq1QQPVeDsfQocUyqGhcUsVxJPYnoNKwQFoAtSTOaeZw2ferPM+J0jPtliyfsOv
luK2ic3f1vfgHZVNnfBVNnhjyONQGlckNvgdUayFKIlIbb+MiXf09MfD9Ud6TvRU
6HQGr5Zyqz6eKlwp5XVoqCDrBOHfGh6o/n9wprGHN9T2aAotsqzw0DZ5csYd5/qc
z8/HDfY49WK90ugJrBhs9M0LH9WvCI3v1Yp4k2H6VntUkFfsvTrVZq5f84gyGOsS
UL787t8SWaq+yAZCEKqIZRNPvRAmP/2t7iajUNw2TZbYaY8FgpAF2mzRCGZI23Vt
7Su0Ceg4uw++unZr/Vbzwb2iOROatuETm7YTKsPW+lC3G/fRrFKDSTTfvW9ikJre
2tgRW8yAa8En+bgiKo1cPPKymg1uvAGFBacfEUx6+5eDV7vj3eQ0OoDaXggoiVHp
6qOjFRcDOgQITWem2ZPfctnJKyr7sgEDIipx7DqnZA+wzr/KL1byYD6oRJmaDKW2
xnGGrynMvxvE62qveayZqZ9n8PylBXp4CP7YC9ZA+C6QNouEDSTcH8p/6C+QviPM
jEav7vxwwkZHzZhTC+NgZjP0b+Ms34SiFkCjVBJtQMGqoQm5XvFIjTbICfZENFuh
aZXLLyYw9Rh5qU0SYOFAj/+lLtITRsnWkSCGStctDqnfAzsh4LlQXqzUb+IF7SwE
F2B4xIf3gWG/banDFy2J8ah+FY0rx9wirmFZCQ0rfpfuXGP+9mHnRH76psEdCrcz
Wo5KAj+qpCHgv9h+wv2InfXn4DKN4d8eBRJsvGvkGGf58k+IxqZe0LuuRjB46sDl
Ydv171V/w2Cg0J7AL2yZQGfPkrRbHYYv8RKktjXOQXRKQAPR7elIkw50xm5oRJ9A
/G2x9jt5OQg4s+75/JCO4Booh3hDr14s0zyQFvShTkjazQuYuKSnECWATZqJFXMO
204xWV4sWY3sG0xFkrI89fYTq8wNcqH6kaus47M7p0WTkSN+NgSLlm3+JR7wR3Wk
ge3oIc97xB5y5hP4S+wgt6qd/Y7DivKHSCTOTLG21A//f58l32R/zcjZj9U/3XaK
JApDNT0ONK7ijQ06zVfwDfOVzp+B7BR0D3Hg79Rp+1ykijxksAleQ+iT9U5u1bHn
Z3s8S56xIaTJOQeSC5AWpOKL/2NRxw4DqRU8JOnmzxy7ZcaGxhIui9mOPz956lhq
VEJCCZmmh75HgKrNWw2slepQzJJqwtO5ciR9k22jtoD4UqbAc5RkdS24EbzjNAAK
KUaf6z7OnW4k9Ti554pR5ihIqYt0zUbJLOrq8ra37oQy55gkKI4jGbeSK+PdT68y
XKa6f99Gw2OdfybyDTqs2GzLe/IFP+JBT0e0NcG7wTlG/F1v0IxugiHkSf/PCOU/
tQNuJAP5tdUKXyGJwxPaganOAK8r9ia/4GwPPzrEzXffrvogJhWGklpwNY0yDUx6
PwXltwvQU+T1ccLsB4KISJxAV7fZljrBGFB+7fPwPLRCvMipjCFP32+P7mn8KN0h
3FQeNCp0CO0eZTKDer8NGzZ6T07Pojt0y5648oqYmFXCC5YcLyxlH/tEWh23b8ee
K2iiXtVlPm4Q0agjXy6rOjaGASCNAExrbd+dF7PCoZi4nZ7CZiqFA28WZGZ0ydv8
+bsVbmtAUtcSx3u3eUol4RsUD0MHCQIoBLtw80CoOlt6pKxImEcfk4gUlH1S1Eo6
2GFYNnDFW9cmgI1lMXgnsoKwbCZ1/383jJdAcq3Mf8rC8NJZ4wWlqYc8PWYJWthN
QLyo2CNBXcS2rUBBrkID++Kzzp/QB10QBSmdP+OSIyHvVOyrbFdYs7s8zdGSSc+L
Mvj3giko/HzzJgHQ/NC48CUqEv2eUAMPpveM3oCYt7VX9wKdibZW9NHyOKB2Dd+f
+uzNMK/C/Gw7afLTzLBGRK5vmUDpIx+U5+GObSL7P7CK0auWjPYf1xc+PD5FzYkK
yX8iRGx9pYJEoBmC78Sy8oRz7JLYRVS7CDplIyhCm0wSnnr+1pKIqrYZ9/QQdKjN
PxIxM56fCldmb/CbxbmuSnZMkJkTHPgBrwAb2QGVuCv4NjAPWbxyRyy5i9ynFRyG
eSQ7RtqUWNAsetDY44PvG9EO8LiFvtSx99UjsBqFgpGUgOhb8FhyV4r+ZZXKtW3i
cepnG4YlZ5WSOB74YM5ncKVvaFk4gS3fp16+7hSJNKoZDtlv72QoEb7jvkHnHKJs
mLl+r3SD/7a6aR0Mv2Oykr0Qy8hJjfWtCEGadiNi2NS/jm2k5VSCryqug+esXJX8
2uif/I4dFVvIZ0v39l9MCWytdODL+8+2JQXxaQsQa68377FFUYi0CKzKoeq5IyEe
nUM8t5+QmeNOMZLKsb8pyFOapn9UBJsYgM5vYaqrMuMMOts2pHrjYNvLs16R3VmG
B4Q3Cs25yH3jo8wrVPKdNU4QpSFfUDYtqA30U2EVCFm9GbNIkxPQkkqKGkvmJEP8
2ohqesMeKdSe7h51zm1qJc6YSToTj1VJqBimlZeuHRhvvjIS9eJzXRZAFFZ0urWx
+7a34/fLHQumjkQFj9ZcIxcEFudkrXkAc9OFFWmozDA16esUqX41gvswCexE3K+M
Efsxt+ZUoj7OMU3kUwrGuwxOgj6V8IWJgndo6QqgzfPFCEeraDekmhGaLRZHiND6
QrLor2nnfeE2szBOqt5bSpfcTs72GfqJOH4Dj6rDVpzv7q9IdQBZGQd6K/kgd5TL
3IfMFE0P9csVn1E8dypu51kU18LFDS/215ZSsj4T7uZwcta2xqljobukWMK0ZX75
3bQMXHniSrc/X/KDqtVdJTdWFStLryTcKmHr1rGaVmx8+sv8+/ZntdQPAWRk/TAW
Lyp0tbcxDbk+ml732lEhuvUa71Tl3VFzSVd+xNMNLJ2Boz6kt2Tcvqrm+N+V1day
DAK6dQRlzmSGdzi0AX1EHfaG9+T6JT7IGt5IXUfNhRAZSxVRdPqWlliFt0YMlgZp
F2xzdVAd/H+U1Z3JILlxKq4BzV6psdCJRlvEItFNto8WIGo3UCjuK4nbl7T6CKCW
uKdVf2W4/IVpYK8mecV3b28PQ7ulieBJI/afVWFZxrGq8SGblt2/qY/VIA7z592C
Obq+1mY0Z6KBvtiFrB7ApCj56GR1VN/pfwrsMCH/s+t7D4d0TQ2/9dEJYD1OV4jq
4hs1sVZZiefoiLPlY/HHV0yUPZyb3B4sBGn5rr/vwrPOQfCX0eoeYHTj2pmF7F6i
7sFpe1ZNrhSlEqZVSQrZSbaZ6YgK3LnIF97x+Vzj+liLDNlVQUI2+p4B/Juy420k
Ph6n1w3yL9sYp1+f5HwDZY/sVZ9jxpZ3deHBxHA0pe+4D5ZLR21Cpy7AVLsakKAa
t1l32I/Mype1mFTEArZonrr4wrKtGgR8pw9hjTeFs/Jgd3NZesDAiMmM/CMiP32a
7W8puyVlrY7tr1AdUof8x9CIgSq13kOUGNj0cNiq+m8jzJTPIIIrK7uDEcgIWSup
+NqKXN3YHL+Awhz0Z79ZVhX1VZaFd9T/1b25plqYMAKNuTGPM8KzZf0zvk6h2+67
efKSREMDdYiqIVtVa0UQdlf15fFSOypb60S5mG4x98qK9E58rw80blpWV2US75Yg
BpgW2kqSsRkbK+zs45+0lZxZ19wqlgVxS7o9hxGuuOfsEiGEf74n/ZEwa/nTGzjI
AqTxs+gkALLv+Wfr0hnLkQ2cAogPkV5+FhHD6F53xOBikGWeOs48/Q0ew7HBRrl/
j/Qv7oVUIuI6HQI4KPmO6uPZfuC2Dc6w9N3l5ge7OhmmAYlDnZuu/N9kWxLH51z2
NQnlRcKXARmnt5902PUAxTMjDH/m+0Yi1JpEvKplXoZzh5/CQTToDepsf2tuJJIk
VSeGwWUBBQmPmmUbV/Pzh5wLhZ571Q3BdocwajP9xMDud9gvU9vvb9asqF2RZqct
G/Dupe3jnGDTQEGX4yjSPm0oXUDawI1K/hRGPEPwoIULsECPkSQ7di43vYadvZAP
7/9aFY2zUV/mWZ7nEzLhpysJlkM1T6NTg/H+eayz70T3MEw0mjA9HLohygDG6eMC
92gDMYIptr6UCqKyiDmsx2/YTHMSsfJlj1UQxX4aj/fJjVZbOhY0sUtjnF1cm6c/
k+a5K3ozx1Tx2voiXoV7wgQ7GTXl16IPZPhOizNTj6JdX5bTutiLlfR4Q1nM0cdt
Zv8CDfhZwmUtX3A4/C+fq6ejR0sxSJbLCfkLLBKpCRaxb05LfkD5FX4Nk5siv3F6
ghg8mhQKr+etUbDziLj2lXn012F3zHt0u82t3evT87GzKZbaoDSDLNFPCfIxkWOK
/10oXB9JxWNWSElvEU4RP/NBtvFWQwOoP8Y2r4poeWqUtXuI2MDJQGYFCbAJe7Mj
znuwLumS9lg4psbU2fpV4Zsp+730EvzpiWY31fd2vitvJuxtq6EHgWrgZF0qUiri
z1AAPR7IMerFniBKEFIQXtjnqoLwSPW6rXewxCeq5+oX68zESa1ShOZpIY3I1LM6
kVXV0SKb0W59nTcgPcvMtPGnpyEH/VDVmnFP56sXCRsftPwMpEZjYQBJVsS3dQAC
uqFBS1R0YE8hxHhisJ/i+/J3pSHG1dkGVjsykltKwww9Bebwj9Cm63wEHbD7Rz5U
qqDGoy2kcM2tEeZlKMj4Rnl2E6rCMG5e34AOFi17kFNbGaK8MbPLzX3QWVI5sxOK
1NOD2VhuABzCyzHgAAjb172+iHLu8x7yrNEW4Z7I6MGM8mzIscbDY0znU41E6FXM
4kRrpYAA2V4R4pVVmuBsbZpMwI9Z4Wj7HIBmRU/cuutI9pXugRZKxhuVlblsR4bw
3aCr1KIdMtmq3cEdvFw5RqstjJ2V0eaMEuzr+ayVoxx3T4/SKD4nLaLBnrdxoNPI
PC67SZt1sAwVX1SaEXWk4e8chZcdwMC5De8t7+Smh8i2ztqp9TV7BAt5O+L3U4Ed
1FG3vrdVIW+V9X1oGu7oa0zXU51jibD0bJl4UUIOGcahWpH8y/xmyw3H48vn7p7w
OLLsdFavtcaQYN+B91AbipIFphEfigsP87n9DJu+QBT+zaL6EiMQwA9u2mhUXjFl
/3rQw+1u9F06l252amvlZeOSg1muuMhEXCkypgWCR2hau53tTEvPXUFdrpyk2ijV
zabo89wOveeQdXIP0WoxFO8ADn3nZ9vst6XjQbrR+rbky0u44epyBnNty9k1YxVq
aVx5Wsb8JO1w4LbEwkfTLtljF4VFaCFifefVIO+5uMEIr28f0g7I/afL2aGQv/6n
cm9CMLvH+6LC/JJ9jTcE2rGLvJ5D1CrGqrYKIqmsjI6hmiLYrAi2dOfbfvHqd1+e
CYNcl23CunJAkpN+JQ2eX4AR3M5cm0U5KLdQyUJUecOAnoXVTiqh2ho51PIYYk3e
WH6DFegbgUks+w5CdW8YAotyRzPD8bP+BXUFaWaeRWtEqU7SZQdq2URMdi28niqs
IR5kVdre77cjEVD6bsxJapkvfdBYxzN2c98Eulvsp/XHXrRwlgYDWOaGJm66XFkY
xRB5XPUEOW8UWCJakKv8F6a/SIF8vAhzHf8Fbaev2tAm/AuSsVUfCzQAFrys5Ari
TU+r8Tn167gr3/O57qcan/LV3zzWjvGdo+15bgbdnIv0DEnFNiq+kAgI6hFslMCA
zz73DgzG3AUMfCo1Hz7CAvb4cANtu5kzsRa56VdE83o7hT21ayUKdnCKbeXMGKdS
XuIDtqJrxW+Jwg7NG0KJF7LwdyjEvsJsAegpSUY6gwV6ZPqnM20RPLc6HMoyDc2f
UHONwCoyrPVcOGr2sjomDpVHEgwhDjj93aYGVpfWSAexDCQ1ibzC1p4zO9X/9nc9
hkx11X0T7Z0u2vTKvKSWndoaXDToA8a/iN3U415bJVN/WKR09j5wAEOQfc9Sn1En
9rI2x8WeYI8DVsmcuBXHp15LvODDT+XonEIQPkc0jmOpRBAh/Ef49SiEaKlBoCSc
XOWbczifosSQM9N/k0dHQ9TUfj4LtT7vnVLN4ERFc53uBr6s3Lk5Iets2X8tvuL/
mBFW7LqL5faf80SHcwGPanBn/Pzz1FM8xvX2lBOLBDTxJ4C7IdXYHwoX/o3otlYU
iOb0uPJRQQ3Tj5rD+4C3DI5f6N7dHvUTgMHpVtNBmXPwMUTyRkvXfTeGLsMdPPJb
SYVg+70PGNIUrm0wKRiFxhp9Qid5oKSYaO0tmzW9AHsSHQL254pT34/dVGhN7hl2
H5PvjvOdIi2hgP6O1GkJnXlb4WBtaPwnKakf4AAf2EiQtDRfnQho0jjYvlGOpfB4
A3krv7x3u77ssdZtdhvtSg7Pkj/v8UyfZAFaUX0N6uLKXLoScS/awXa4TIJWJ3QU
p/Z27GXiyBdMXHBvqvCLaIKqG0zvDw8qtPi7s+zn5EUvSnrOmcfzhbyP3rl8rZ5v
bQvi+EQwlPMbXB0emqErRdUpBuIqFnfKBaOURVQPQDl0vZ9aeeBj8t4xElSMwLa/
DCmzaQql9a3DvMi3ZkSCb/fqG8R8QeT1y8xzAC4vFytKWWDhlvyvLnB6c+K3PdEo
YLfItStZ5whehxKs2QoozzpOCzbviQxnAR+Kji7uKjYMxcrKWSm57Zf7TpbsZhxQ
KuUpDzcexzdsV7XpaFuZ8bXi4ooShFTioP5Taph70qDdPlKVBlvMApG3/f1wjU6C
ng3ubB7L7YlE0ShZ+NQg73Evztuq2I0DBC4FdIVHYs+Jc82OxeMVp8iDMvY7UCGw
Xmk4EcoX2ANwgygCitz7D0WGxK1iunEVKeqx4c1ua2ATfuhTCtsyJcMUF2uGlCuP
/L8QufCtw+RfbA+Rg+kresKg5E5lQjP/fwgmDcNrbkShkWFVjubxPCwFvYXQziT6
atQqRKzqFnaeyljqVT86hls5gVRYqvfHkThpWlfqgHsmotlpogT0BgaPO3xPagig
hYTgE79ETYdCS1QdtVS3itckJ9cffN0lfu406QZG6PyvYsBvbUQx8h/9PPae3d7j
v09t3L/mooG4Q6GTuH1XOQ6h02GTJ7T9P8UaZFL8MAlwLegmxt9aLODs+SnexTF2
zFt09xbGWlx1CBrWPmYbI5jA4RgHY5w0513mKYgyh1bDPsIfHByVWW94Owp6a2Hp
86aGa5APrl9uavGnLw6s0YFboX5hXu8s+g6z+gdaVhNcsNXqB0f5oj/tJ+NmyR6g
ke18aFSOuv8aayoZZRiMCMrePeWPmym+WZE3XZoFqPlmcWZIUaOWXy0jOLlMTmRn
2WvPnDTJ0SDVeiHmmV4tcJiPkvAtvSypAxoEoKgIVd6J1ZRPrBhnpcnXLWCkyTyy
mwQ6vCbaeMpzX7ocBqBvU1YVgU/YDH5UrynoQWlZZNaLYu25guUtoKiiDlVfb9qv
vze/7vxMbfyEF5E7oVoAD/K0kzVID9jFJSYoMLq6HgplCUogLA4NX44jYdsuNryX
B7st+Pou73zrBJc1TTjRExb+q5WYP3OXXWx0xcaH4O75G7fQGp5/h0qZykeX9p5a
oVXjQdDH5qINZz6BWqRgU6/OaRe0WasCmSV5zFFIPa79pYC90M2nbL3FOfYRjcGN
3M+jOTmJvrCl1w3uhbXFE3cvFKGJPBiQSH7QdB8W+Xh4Wwtl/6P1LE0UKk1Yjnhs
Fz6gvo3fBj1UijzRSYRwFdds87L2g4qs59lTJIzM0sbN6lh3Z5saUJ2V04BL2/NB
nJ85uBphimn756JqT96JpKkDiI0HB0FM2fDMGLkWlTBLR0yHOulPLg7o/CdM2N+E
RGysGKE7Ucyr+9UipXfgxPtF8sO9Xs3KyxKGypYLhwtKFOBaDO6AgUTMNI+sCOPv
9duojv2KN9C7F0dZgxfk9bNKxn+czcYnDCrk1oC8WAKuiChXdSModMuj5Me8rtSl
oBm0u4CmGKpzYN7onaTAL0vBTMqa438G1XIwltD2gb/qZTzV+gGKAWq6NNBDOQtm
cwRJxnMfThMZwA7iRfE7h/EZiw9RIA9vtQhBGUXA1EBgAFLJYjHE+IMi7hvXqwTd
jtX5hd/jKpQlLP3RrWnkODFqeHxByRotlotGx4JT5nl2dkHopM+Ywph68x3nzTmW
bLh1jmpuVpGXpkmg8SPh1J8p/eSXD5/rIcEHNJU84Ajjw9RceLWPgXvDoClhbB0u
i/Xq9BvyNWyB5K6xVz1IurQ+IFvX90Q3UPJGTT1v7YRriMxj7UgIwxLjGwmH/xNA
4gRKr9aoMGzV0NQgEOsPhAX/245ZyjbiPXZjkuJxyS3SqTwPZ36JYpCbmTr+5R1f
Zd/IGcyyg3P8+1YqAP+PKs6unFdqYM8X4Pbvjjl7TfN6ttpqRhDKNYR1GjndHcwy
Hk84CJuzgYnhyAB/HYtsi693kANP/XZR9xHH1hLKlykgFjbiN6yaPfT7yXWMGj9h
JZH2dNoCmKEnKo11S6MuPHvjucGWtJikppp6fve+Echt1+ufWaTAiXWqOGzr3mdz
n9tHKmdCCFSNY9WkUgBvL14hHQkwvU76MhASfPBOv61O6FtyFgkRBbj93o6cgor0
ZwUL3Qt7NyLXm9uBO7HWema3jWjqIKXMnnphN0B4YTMIS26YNYZZ+0EsQTzBMV47
R56OolEZlI9osCMOpA2bnwLeY/VIGXm1bW4G6ZMN5pv1V062G4OHSFoo4MvQZVex
wpuNLduL5rbFI0mun6/JihkdyVhVI06ZDtHQ4DlqcOKb0Y7YLfgWWgoyavxqZFSx
nNMfl7wT/pMJi5FWYnTQF7nM3Qz2V5hS1YLTI2WOmbsGHpJXftFGR/0xPZek4KrM
E4iACfA2pQFIStlq5zULTsQBF1/Pp5DAF1GwGhxnU/0nOPKRa7LvyHDkXsuBmjeH
piYCakkunvBNhYeMlbCpuvHUq+nM9piC08TaKVdUtlBN+foQLGIBPQH93n2r+3Pt
8JST4X9B3csXBBEmiA2000dxRsnibnI8sn9boYLx31lm7wpru3Pxe95zoG9rd8e3
6svHi7hX65DEatwlI3LWqXG8Kcof49DCfFlGE3wqrNJMljTE5q/Oh+/mnbooe2Jm
WxYqtlqejDCy/j7gO2HzOhgMgRRcZZbX21vmaMpw7GVv0XFskc5eTc0zq2T+5/hD
MbwrNBxPSLNeXs1tV1myD3oFkvQCoyOa5l8r55copUAZvgkkTqa23vxCvFo2fZgp
keeqEzy4je4JqFcLALg468UXlHnpdVqwnC2uUvc7VjPDo9PR0GDVWSp1bdAtNd1H
nYYYWJ/dX233hs+oMkYZlez/dFzltes9w7jzFN2N33Z6ppd7pMHrfXBas9UoJ3nE
9UiIvqeUBtHpAmBcHDSOcwaN6lM3aAG1AMpPI4GAKpj7xXbGT0u0U9JYXKjW0cnk
iO5uWtXYPmSxvkkijLY6is6e0xzQNTzLXVvlqjc1swrF4wiwHhnVs8x25VQ9wWy+
GjrKOyIyu911mbcCtBikg4VInosJsEp8o+i6K0RjktpzpmAdHkaY0MWvef5TTYri
mE0Jkachlbk71TohrE79sS/F8QTkiZjBQJ+cy4raG0+0w0OCnAa3cEa1K23vCi80
gVfZfqkmQD4x5jGc1eTJy/AOS95scShLk9wV0UXbFXoWeWMoIuXuRQ0gxzeuqLwJ
FLS6goJr7Obi0rg4N54xvuMxmus8v92EDtqXrB/X3zF7uNxGQdEuvrxORLSDObnx
pzqgeQwe9boy4DHZz2UYFeNx13Nzd4A0TqRHICB02aMDNqMFVQLb8F+hZUx9ljTD
pwqoSp0tmPF1bsvu6mYDmOkxD4dVjhxHsr6b13+For4+YmU8A1/kxoT2MXPHAXxG
F+Oou17Ul2G6m3WW/d5PkDkkay3yUTYkmIwQ2irGf7ztUl81Li2jYQTZiPV5tgoK
HFSR1z3kmzFW3MZGdlfahqheaeiaslCRKEeM4/ktGvBkBDI8CgW5zjj+61XzDvi4
VWpOGgO3dT2xrv3RIZy3AUzXsA2sX7pxPvp2W7lip7YwMHosXPgsgIVxUoDRLSvt
1elIqEsi8NcyQW5giTjq+VdGYNvoGt2gRFGPaJvS8vmFySvIL99nNWirvZCE6leC
n/LXb+ZIEi1HR8ZfIosOyh5G029RtwGJAkrWl5oaPqdMvsaAUMWZMqrPuM/CqQi1
zOCuAxVswDYQoAe7UHN4gjbfpc8ypyPMhbZPbOS+1jZWEZDTu70PJ8QiiCJA8DpJ
wQCZbeMv8IvHJt4ZFQpGXApbHTSfb1diM3fUk22C0K0RUA/XE3TQVLx7G90bq52j
obiD5bFDm+RwcUALULyRf5lBsX88Y9rIKPMOiHlhfHo6W+G31blRbv53/WAdzx9v
DgGz6zLDQnYyqGnIT1BVX3Ap9mkEnqPo3MATJPSgft1QV1anLtXZFqi8CAj2ZEcO
S6Z2QTOxDAGVvErvn2rikTu7ctfFnhqKxnJmTFUgwvHKEXATcQSdAwUZUnmfDKot
rjyTXS21sAp7wLQUUNn5NqldQy7/VRHgPn8D2kF+kkfpJr61k/rihIv0lG60s2sa
cc1xktsLY77lfD3FpoOs9C8iwe7v4240l38GozhZ9G5rsfwVW2g/KNaEI2OjDy91
GzZ0sKV3JsErF3LCXZSb42Xgg3cGyC3up2cfUPlzk/hhEL8B2Z9ly2yznzoy4Wsf
9jjiYDv0weOxdXWD2iTF90QTtgHu9/DMNrSScfPk6sz7hwi43W7HIQz0TYxFS+go
2XUwYP06OJb4McHcUoRvkbDW9Jx7J+VtqB11vhUdLVZY6ghZTwpEMhbUHzfBP0L1
vJufsYWxcCJoF5dnRmcXooAd5uHrzJtCBENQI78kFpUB04Y6t0i0dXN0i/5tnqIW
nfS51vgnDRR9p8xKg5p1CwOJQv8YowcR0jVv8DsHMF+zgCel2zrQ2MbiHmE3sB7y
y+hV7ElG9RtUjqBysC1GbpkaQMqwFOUlQTykmMEtvqPk3vDd5yKZQSQrHCG/KTW5
g0TMvkUy3/G7P+m/JCxILz2UNC7KqDUXgu91hh5B5e7z+ZvLMWdI1nb/dxwEeTud
QTyU3iBiCybAPgBDiYT57BLBXWORBLcz7sMdK//+NRnbk14rF2PsOEXuJse2KfYp
t2VRIiEM86FYafpk9BLAxWMnkV6aYbwhuk3bgzgLV1f3KglUyPmYqozVzovzxqOJ
PAOlmKRQ1+LxOke7DFJNNU+1yTQwmb9J16Ein+BpEkP4Mm/FNeIefP1qLf8WC5by
K6YiQxbDGpczKbJ6/PoWzLatI+LaRWZy77Q+pWtLldJ6CGXXzmb0JS1ffI6k6VZI
genlRk6yzWNE8h49kCsxOB0LdxJwOVU84MRDUlbH4A0BQR6Xowny/RG+9l1ScIXl
aCEewWo5cjHvu7eLhYyLBNoC/2y7+bp4V08+G7RPfHfXrNlnYr5UovsxKtLiJOgu
hgXRo1ci5gxGOnNyaWg7zbfu6+Sg09zHnW7SHE/RSlUav9TIJRsRO499g9c0OfiR
6tKE62RI1GEeNPz0RncHy2ffzCKKToMtAqdERiCz9Zh42qrHvePunkWj/rIddpzC
6mTo7itSbOU7Fng68UEWhVloSZ2ovVW+PzUhL/B9WuE1+jF+bm9cj6Ml08EcaYd6
g15d0UhN4UVmVH1xASTl8OmKUvK7dFxuUuIvzn0lWV002sw08aI4GwyLrJ5FPv74
4yZjDROFdwG2o+VVIbF9PNFsyW9GCk8wYsAv6t8ESE8N+XbcurZutrWzaKtqEiFu
x/mF7HuLvYxtSl8yFn5DncqJ0FrlQtlRtyWKByjgiTRPdtpgJRopgW6S8MlhD9YX
CPBjjFkQIrbDCbKMeoQ41dxkA6hN97z1YMxC1u2G01MxNhJZw5Sy8BhJrG9h0Fxp
vmzzV3Y2V5zVB5XiPCrrw/uSvYcbe22sF5+12MyExLDQhO+7YbueAjoVpLQdvgtP
/J66igmYxebNgf9odoO5Map6yzV5+EDxuPVQb6mgYiiurOSNMIdtvu+AUGJoJv3+
sATZ/PwmAFOPK6maD7zWi+moFEWrm5fyAoDZeQP5mfFLEy4QiqfOTBlvWjXzef6j
VStDl+afYcsjs3Bh+hvsHGy0iTmx54pTd2yGemlKuMIBZMPG5Y3+euCgrV1xXFqs
JIBWjnL3bJQhbl04v09KuvhR3kgOhSNtgPAm3BSb2K1iAJIgkysbaC55BuHl+kCK
JivNFP+aLPaKKfifu5/vX1RcBnbvUP4ThnW6Ygbdb9m+hQvZQq8CsiHT+JGKaO9J
oXtvkEVR0uP55FFgOeYq1uJZYyY+rkJRuUkaatZy7y9Wdy06e9Zu0p+hbXv3oVeU
jPkO3tVICdWl/g7HRPR7jD16Ozj2NZCSuwt8QLoaCGdfYX1/Asl4C4tFHXiDkNy1
9nMADPIO9gXNn5zEyiFwdyLtg9HR1Kj5E+5Kr/7QEFA3CgcPI0Vkt7DbeNMy2zYZ
+yC+N+j8tQhoFizphLavdqzgexQnGL1PASB68ssOqbBPXiv8qYCALnllwlVhNFNG
avkueI6KaiJg+5Y+OiRdie0DGrayKyhzsvZW8W047ynzV3VDZXpPNnJ7RupV+tYr
zJ6FIeCxAjkaxtngDZQwVFpssb46p8rGG53xZjW3g80P6NN9frDJpL9HspWZQ/NS
VKIHoV6MqVRY67sgVbUH2oRPi1ODOHNbxSh8YK7umrTmGVeAJVyWsc7u2sofUph0
qF4YkH88+yVE8l0RFr2zuwc/OAgcFT0sZmYhcQf/OCWov1YU8WriDTwMunAsNcWR
RXczaGOz2ntOjIM22HpmhS/z7IiN2L7Fq8nxGaoSC/97Z4nkb26Zhm7RXVLdKi2C
TyHsGadTGY9djFSRDmFnNvTqCWtN7E445489CPiRIqkgixAxllQ59tP1M+Y/zQLE
x1YrQkCCVJ5O6viokckt92v3ooc7u1KnzBG9mHYBgsMzaTn4rvxU6w7uTfaNSMV8
SXORAfh7URPdlYHUCntNC1G241cSsWpVg4kzECE+OhM=
`protect end_protected
