-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
IS2NUDD2KxgepncDvEMWR0uzepHhUztJsybjm1YXMclpTLQBX3v0hkXlqWVQgRqk
iW2MZVVffPZtZ0DtDs9BeZbqOS5der5R11XNxaK5ewpK+IiFpYfkRNWb6kDsr6Ss
KxFrjDYQkFdRBcspDNJIh80W7xfqybsxnguSclrCLyI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10017)

`protect DATA_BLOCK
HSbpsC/wlI3fN99djvZya9rcOZpE2aS573oVi4YkT+DD2eAS5ehxZvk/iLJukP1c
D7wI4strh3UD1nFFRx5E3VVwDP07oK8dz7BPhemPwpuRDSFpGjKxklLoMZW3Y3Yw
vrgAuSL/TT/0GWco/DDI2GILRLdyawrt+X/4A8U13rj1idd3gE0hOcpfTzsfptI4
RjEoo65Fl09b0l+6gGSDReMTzmm7UOTIYsFJhgDIEJNCTWaZsuYmiZORlnVVjWuY
svWZooQpSPYA/RVhNh+8yolXyz7FgOqjMmuIa0LNUckECGX2Hoow+Lz4WMjQ7RCP
cxr6cciawFayiPi/SqiIoidtLh2golsp/UmQz1IKHnjUa6alKfPM8qXcxucnRqBa
A/5969brR7qR3H+dzUjbrgCkb4/cZmIk9Sh2pR1krJR6DbZ6vjJMxPEe0AdhG75V
nQ8wt42dXHjImAuhperpkjkHjQgvj1YdFIo0cNeulj8hZ+BD186+7lDPKYVa5JTw
7K0Grsj9fXW/GTlBvGinU+p4WFXHPt7eWbOMvI64NfARjOFG6EzliTlh+ygljBuT
KTgtt3IPpqGKCaQE5/ZdsZbx0s6K0CeLhNkV9wIeC6vzsWAiLYclZ/Ako7QZ+YvD
csMXgtZgc6IXZ1Zb0MrF5wbpOTXCLeAfjleV/SWg+YN9cUlyitY+wIcOgNQ8onNz
XyhWA2fokr9bRRbYK3t9JJ4fl5tmE1QSCd4APYJbY1tfOLVdm+Gr+/ssyIWdUh3R
GdQnpNAI3VRcyV1mLEwJRhEM1TvgCUXyHa4oaPxNpvazDGXbMDEG63omYjrUm7CN
U0gy7RMJcltwYo8848dN4zvvFLpkxjsSvng6D2ZMPLnBLyDkX1pxYekpVPHzOXhJ
9n5HDJE4FzOF3wT/vjtNtW36jzrErCiWLMU32BLumDIf2R0nsqFJQJtB1GcYC+5B
BKw8W0DgwJ0fjO4o5Rp9niDI6YN3E9ejLnazAYE+6AaGnoewVO0kZU3AeC9L0NjU
R27JRmjif+l/wUBq9Upu2Zp6fzvd7M44GmcpEf8uiIfbDBoyM5VkhLeSZh4j5rLo
olCyTp3VEQbnRNrcLowB85AAEbJMwqOBPobq/GdZNBr+FNby4H8TDR8JPz1eWbvO
gIGEv5VJON6NaqaO4fiv9qYIvXV9rcwl/z2dIpxBVx04i/eJQaMJFDI0V1iQ74LM
U1zOdQ04+wA+eXZ6Pm1vcbYxdhbG7SZ0vgebYpTc1RaIi9l3UIrCG8XTqFaOWNHE
I9i0RGXk+WJOLfY6GRYvpWRCpi+EVgNSK6Kh4MMpNn1Snx6YMIZDqj3GO0TZPKTG
qoYw6WMQNUR152z2Roit1xUJRBeEPYuZoUCwONzZsCC6WLiOXRYJYdXgDdVQScdH
3FyqUH6sC73qAuGGiukvRcOwRFYK0KKDPRnNLujb+wsSNmLwrexq/QB3SSBC93fp
tle5jIZ015Bw79Bx/ujaJF7Tw+YXWGowLWJV+ZsuYdK34y8t/O1w4xNdl0hMKG+7
OUskyYtKg5mfbBssB7rTi5+s5R9EqeCFwm/1NMrrqO1NWcWETHeNTUMNWCM3UFIi
KHlQH9Os0ikY94PqWgkCiIUiQE5Q0+dwL+RdHaB8cvXj+kG1i9ia4hstCzytI/UP
hE7tTU1RW9JCcUeSYLgqwwreTUqz6MAN6PgC68dmz183AIrak3cxHHzNFNYDUjtD
XAtiiQYW49ENo3XXtoDZw9KlOUbLweT+BiCnS9mFGAvh+wLZMSyB6aKlKmRdww0o
vi3U8sFrOidbZEUprVhjSv7b0bmEt0LvWhtsuDmzULTFe/02u4rjsZIHYsXWfoAi
eQ8o1yOao8UiL2YSPEbJG2LDATccJMJDhrTMiiW8KCIw/6VxBfHRuK4VR0R7PVtq
GECzzDnC8aDrUYv/tirX+adDPYriwgzyRKiLr0MxIYblxeyOHHiXQHUqg9r/9tPO
+bsM+gc1XDTeZFS8AaqdX8VFYi+3QdIr1iPpgUDHXJgcIuFt+R6wtKZ0L9Hdgdr1
4KEGAgOfal5RsWC9Xd0hwzrGct75uZekOFJKAxKtX3JAgQ1wXG1kxDfzw/3ky4zg
Il+sg0vfHynUiimKWdXs0GN/BlfPw4YiizivLySZU/dzx1XXqeSOnjVkl8Eqyvj5
ht3G/LfZ1JgLXNviC+piwEug6KZcI3VXhIexNErl9fx/B+5NbGYWQXUMvIMBVh2W
6+DenCTUBqE1HfTUyhClVZTvLURE2ZCVn0EHhAzaKzEg0Gzhi636wZqjNmZGD74Y
v0r6bL/WFmw3nXNlghphRDqtRWcEbUP/TzRKF6hhXvk15ux0qP9KgUTe/r45J3bc
FL3yH6u6YP28ckOSFxm/BsM/9yqQbYRoMnMuxrBAZ60+kto+h83XnDQ9iaifY6SX
T2dboXgcJgA/wdiODIQC2BnnvC6LV3oBjKo9j2BPM/6BeZlQuyMlc1imSrb4emsb
URXRm6rN60CZkJc59by35MGd9WvSjIvl17OwZY1+ECoJUeli5/pSk0kUSPAlDJ7r
jzJvu4g223zgwzP+qO3yQHS7k6VoNyU4dSdr+QK7s9eiByS2FTijnsiuN4uZbE9n
SPuZQeGjiNYzfW25WQOUr0EVL5Dh+7laLMi5g8gXzWwn7OwumR0zyNW8UClQ0+7u
qO9xjyAacYF9IgyXoZOJvRfvAaHVR7KH+BtDRGvxjFg7xVkYKUXddQjWAijr0Jpd
L+gaQVimzPqLeGa8QRET5c9j2F0RT06nlsU8t9yNUd92gupjJqlBRlQ6xuPygnOI
13yiE+fUegy0FcQlOFIF2Dia90s82Du6uODfJwYtr9Dg6ygDnM8g0tRT+YMWGeQa
ZFBIGxKUyLg1UoYfpLasSgoh4KwSL4CVp3alStaQasyPi2pcAce3CW/VcGS/kxwt
a1jS6/t8rf1lexLKMJOwXsyqvHdLAmCvYpmh2InyzwF25Q5oO9RmXdFHS9JWmTcb
RKiUX3Cai/NFy+yXUSI+AeBkAdgOXD8kZS2NWB6Y8cM8gl3Q713SPPO06Jznz1JX
auyfZeCkHzNvFj66L9vAIrU9JtTO0VD4iygXJwr2n2ocHfPgca+lLQQOvgIaWZEE
CJFW22oHpr7LGK2C/aHGLSJSRyBVY6GO8Apki2C3IhNMEK8PipuBFvd5vsarrjnz
NgD2r0OhIFYt2GgW53kIo/9LASENW3B74hrVMSiUao/l4rgBcgfBx3TJdmFCgTGl
aLYLqqRg/7uAZDHa9nWeB8L7U9t90Kg6mJiu3SGD2/izpY9o1Ev+zDx7Y2SXnC8p
xj7p/k1ov0eII38pwERb3b3AWo6K7dHU7OcX+1Ypgowir6f2INuT28x5yk3Dpelh
e8hAnBSHcPXlByUomJHhHo+u/jJEgGlo+CY3l+61HPjpXKexc4o8I2VtfT0IPcsX
opD0VmJRLB71F0GXDI0trX3KF/Nj5P+lnjVBvnHZJNntNRoCdROpWaMYltV2heAx
hNPkJXWrxXwm797j6vCBft9xc4NH7fSMtaOI1Rg+8RoUnBV1QhhEF7WH8GG1DjkG
J81g8sdBFXo+RHDJ4mdUeVhaf2vaYO8m+efyTZBzplIdhKuOlNq1ED72nEYpVhFI
v45+igdjMbiA3OSwz2WuKMjvVQkBT9DRQV1/hhPQWGW5srieikCSSzPdbrJNBfBH
yHvSJTtr6cbULtKTaBhXeDzTGDogaTIYf2UM++qcwdpi2x4llZO+6UPSGTPRJvDM
H36zxEGxmmH0yyzdD9vh7DF7ctROGXTFCl1d1c0bfCmsK6OP8pZFaTYs6mmOPA1t
jaXiwzo6/VoN/yw93lv22E/ZTG9BCxziBMvNyjBCibU7iQcdS2y+0APHtfpSCr/T
G86fTLwbTLriHItYA2zJdHeOYGbrMGK3w0n7AJlo2+r9qilrUvnhNYhUDvz/C+L3
T4FJXSsjUiAWxZAtRkuaODXXMoNI2TAexng9ENrw3Qis8crhPEMIPzvKf2hcb2Rp
IvMd0HPFi71IRk9d7beSvp76BFkMBOEFYBOpccyVBJyBHL4RwxpNaQmlhkKb0cOZ
AlyvzOFqlexBgmrtHrxjzfrf1Ud8NcA+jr/3TRE8mUJvCdbrufoQ4GIXQ2RPRDa6
dentzq71PHb9PkjdMSiI2wc8hjY7bxqKJ805NfZNLdBy4b78sTTysEv/7kAFudg1
1bM1D/dfnfRVg0sXCpgVCFxjSVFAVrxPTaxiG0Mv/oakia1h1JJOOHbbirkc+amL
OvUVP0H72SIB4Ihh6Kpm+QObXjuvJwO7i5Hm3TTZDmnfZCj9ECx1ekBbUDjRM1mk
Ra4Z+3vRDgoT6qiLksw7LySTPuKxm0VIkp/TD6IROIY0DZC0KEjkp5gp6ewL1FCD
UxAmv/++AS6gu60x5Cx+kVCt8Ev9Xad2wpXJbEfwCJShe3dWUQI8avaFXsJNwXXl
qvBb4PBQHvR6ZAOfyF+35nyeYCyki9QRmVKZdR4LEQyJUpz4wY6Ojuj4GOl5kXEY
qtxVLC1Kr3C7IKG7J+gGs63VnAtj6pSD8isa2ud7VS+rA0AnBLm6btncmneOo9b9
mr03mIIbqmEY+28h04xAp3cQSsfXQBgWI8MSVDhWKT7mvEV65+Lkf8Gj7gC/4+3d
lrwUoieWXnRmDrfAbAth5a1Og5Az05uG005rc6Rd9akE9tmz7udpFCoyZ7LB4JxI
TSio8Q1YwGZo2IlXUpVzOgcE4ZuWagUInKGClAg7RreoM/Dm93lAanNEOmozht62
7apZ5OS6urBamZOojG9P09L85yqWY/HNfSsfzDp7fxJzlWtawdUbpbMr5fMyB5pm
xdzWGJfxmBt/6c/5t8yDQnIFamd3bwa9niq4dmjBXghoXL7XaVk9NkXgeAumKHHV
uUxFjlP//wKnR9a/EBevsOhS1y8zESXlG1Og0O5bpPucw5iflnhqDRjY03+JeIlN
8t6hD8hmrxLfR6m8V2ap1OSpky6Ugsq+v4e3/hdwHpC2OsXFG5qjQbODwvDo6LQn
bdeNHgky7tgmeHl6CfAM9hYYcMxPlmdlw0CHMnd4uMiYLey4i+8QUMDtoiOAZOfl
DB/H/RHfzHXg+zxYvdkVHihT/GdrFURPFo2UB7Nsxi9uJv86rjglAUqinaGiEqwa
d+w5VmZNZUEtEVGA5FKs/nACrN0IVZTjnp6r1P28yDUYlrJ8AI3a4famQCgtyxw9
wHDxj65bg8U0qz/McgmUSM4kKwS+eiyr1H/H2JQimjk3/EHxYigoHQ/R4gCKljIg
vjL/J4QF//b4lFGnVALEKEIHqPTFk05R5/GUQD5HVfnRUqkSbtOQ3cbtgdvZsbLD
/kQnaF9UG2giDzYPcFnq8j6QChyFiSDYTDtZytCcSMXCD6FWCXMh/On7rZ9z3UR4
BcOAOqxWrDLGZiqSjdOZE5Fdpn4TGw1XP7HIomY3ITl/nQStKTQdR1PasbI3FSqi
tSP5QPbVwN0MPckcGK7SJKrXpmp7QHWKyU9RzxkjUWP1ePhrVfHX8jxf98Eq5ues
QSTlfymR//J2MeoiYlvR7fcvqUprq4ekPnoxhZ/3BawJGWwhotwcSzWgfGvyUAiR
9tLNCKO8iu2H0idekXFxfhOWW+aFD6ioodnbro4umAQ3feOsj0ANo4dNAF9V9QDE
wsPB8iNWwusOsfzqDm0pi1EH+Uf+CIIeCzpGnpKAtYxdMeNwEFBkc0gNbDYnvX2E
SK5eQpuVTDmbnDRxUo1g9nk1K2DqBlW99Wk3LO9qDE9uI4LbMgc7+2L+e0K4Xzw1
cAm6bLs/YzMyJGsRlL3NMOZn/UcRs9ElPPuwUe4PQ11+aoAHRGq4RdBK7GSXC6SZ
egS2cUZjsVpKvWChM3Z3GsxnO4LMUiGnz/hsiyPtGJ4xghsc6oxN/stHwf8N/J0a
TJ0z9repRj/OR7+zvHZ8hunwOc0p4E6yr+z/PuVYEge3bW6STkwbqYC9Rd8b3zNS
WcpgbxDBOX7FwhYlRnmmIbSNCpLczi9HBnqj77bcs8eUjUlNKYT0l3YTpkQtsAT5
ryATI6IUb2KaPgcTgjcp8u8yW+GWnVNotTxIaduyqCscJ1opYMyea4awqQSzWZPl
T+oeuHFojHO2fd2iYd+RCgnBsQPDW1l2IeDU7urqnuOylelihU37n+BVe7Esktfk
8pUp4/xZjNDT4Jx5w+V9FeVulSUfdpTBJRCZutXSJRAmh5WULcmRH+PyCD6zK0hp
dLfmS+gxojYwuq6mbxkpcm6zAdvL09tOB7Awi1oRjH48J5U5kzCK7n8hKRh9RTTL
9INyr6rtvSYoNamPZuSyUJiEkYtmoUbUUAMyym5A/q+VpkxQbvRyzXUBlkmTOWjM
7HAI1ZtQcK/BJqhRhyaFSmoXZLIy9XIKRczP2znyCeA59j/87xbbhbWif5GgfH03
KXLe9+uEz0XDQAYPrkvPBkpTex0TjRDq4+Kh8dHrF5yr6dhTRLDorgPB+7r3boup
lw67kcURqLnVbzhRpR4xa8p+GC3E/c55/GVt07cL6VasywZTqE1OAvXPmVmzyS39
9YlxlMlSDp9nCwiPmdZerw2zV84iBisNbK2lEkVTNvVWmI2VTQxDuktFdjk348mz
G0qTZ1PZfw7tnK1K0VqSQDiZeLDOK/F7xUhyMPWxUObMobwGiluBU2WF9Dto7WcO
durbO92rxOvH5Zll5ntIwAJfqxfBDsKP3t5rVlL5zeuXispnQVoJgOGehtANOZBV
dljYvt+7OL0u+D2RDobWgMPvHUGlmXoNixdc+zROGKiBTTlZcPezDVTTqkPULXkT
+m/by2cSOREfp0J+qu6jYmo1WuYfcZFNE2seRsCkWHwdP4dCPtcGN5UP1KcSGSeZ
Nif1VThXspgO4WG+lw7wOGxiOBt0xo6iRQ/d/cgw0CEcOE3GBF5iXt7dANtp5ZAn
9KVHPZ3IfsdmAEagXssbDYk26VkIF0k+19rmwdi4xTa8lYEi+SXvh4lcjl3xJj4c
Ksw1n7AdOkexSYTgL4mNIaW+qcKeuezJVFcWDUu4TBjmYBOD3S+M3NmEpALHgvj2
qwhM4s9wNKmDsGjfyi4r2kfvm7+bd37EJWdjtaQPWYB/Yru7VO7pBNyfQR/WTYnd
C2VsGBle49NKidLsc0rr6cW5Xe1FkXLKJxKyR7odYniGXEuRMoyw9Oh2HFHzwNC3
Er3hEwL0Lc1az29NXo3yMZLe2ux8GTenZDyOEaQLn0vnZRY/WB/sKxUnLX3iWi+H
N/QIrg5qJcjOQszKQxbY5NikdpO1nrmsc2ne+MdoQK3AMgj2OU2v65E4w66Fz+Sc
lUs83oZCSts7xgxGtjhzGoZuXt7CT+8NO9HLM6YS+7YgaZkPXZf0ZJJ/9jP3vX0B
MiVIKTy1xO6tqtDBm7tQdTxNiIKQQPW1F0Pf3bG8d3pJi0cjoeJZmYCqtDI+2NAb
fpce0pqhGeD5AdLlctszOC7lvjo9H/xrKrZ+zDR4aN8+aEyCxdTkCYTmPzIFJ9M/
w5KfaayyB9ZOYn/oZFLQYgjPaOr/Hr5em8Q+3rlgIG950iFpC/n9tPa7bIgx79uB
DcnBfhHkHdrronkVpQVV3FIfGwvpZwTrVRefHcSgTxTDBSkHIthYVMvTcoU8o8Ck
5iWGr9AuK+pdx7rpSybvTuN862Dk36VqwgfcG1rCCysyM+8C4KKWebkM/23WdSrU
zjzi+3wCK/qXV644LmJ5NA5648v2QMFrzOYtIoBzl30fYokFAyFqhndGM+h6s1iz
zcQkmbe+lVnh5S4ayHBSTD+GXe6QNiEHrexLCEw4l76WHly9QMdWu+jc/4jpqXpb
cbJ2kJt8+CFy3u/NHGQJ1g8Lj3FVSwF0lj9JPnz+XTibw0nTxYeyvfxo2VISjUF+
KazDUh7TgpP82Jin4CdMpjmb+JBEGms5daM2toE+xXY3TjnPW2aMsIZRyqWPKWEU
Mhg4OKNJpznjOcG8RJP4kPy1ovmb9jD9YAS8mg/lECYE1xxKmoXQDhW10M7vfug+
VgRFbk8Bx7twPFSx1groxZLvn5z9Xqz50+J3m8hEAxErcTvXu4AOUAF1fZFJIhRn
nLW5u64d9qZKfkMv/5cqoieu/V31DL627n6rLNXazcIauYus90+InTLEbvUd/eKa
r8uWSTYLmsSOSTJqQxRcS72QL+AfUvvJR+YnLHOYqosCC+Snp/ZDCVUhf9cHuvE1
VOxg4RVXr3hqbGXbtEsM6sBXo/yUTwr+WG+S9apND/LYssWeAsuNTbepnUN6/P+a
J0GTy+Cq8e3/woooH4CtxNeoNQJZpRVTn5Sg0Y19Mtm9n8XhsscJ6gP6Qf8sZ39F
uJ4BJbeJjhLjw7KZzE8LPsqENNbIMyR+iajqkP4AYlkn94FgpmEjvnBNUpeIZSig
8mDhh6zhZJmcYVxaNIbc+OHDondNdy5d894b44oVvxyE2lOH43uC0LHCAiOXvZQD
9W2683Empz11NKQ6ephbkP09pAc1qN/yAg3TxYlT258hMuHtsBFQWV0DVjFWMF2Y
Tp+0hRKucx17l6QEoIkzjhOUetdkNVA9AzoUMaeoiC/nR+QAHLT5NmZLI67AQqP7
c105ajYPCWCyCYEBfZOSun7t7bd7pAAriS2ct4xkFuMoU/Xh2S6G9zhZ67HnOErc
Q9Ah0DkztOVoC5OSuKQeypjltn2dCrkBuHqVk4b/dQyIpR1IaqnDpKe1/nDm/0Po
ycud6vJkbZeGZF2q1dMZ+ox9SKvO0PNKU7Kl23ytKBAfgjWPTzMUFNpm5KoIyol8
LCbwZ+CsD4enPnrPaTTCAdEzyDb9bQ0g5tKBX94wEW/gtlCAjuqEEyf/lDAYCiUY
DRvFC8NzVwWRngpfEINXGCog+azC7z5Tz8DCkWdvLEbRO+KTdoR9e+U9gZ73xBOK
OgBgUEDRBZ7MtCK5lqZKW/EXCoicxBLbusXecdWsl3CHFEOKjUuc6b5ea4bn/NAc
UTFpozH3Hld6xNo84m+M2k8ZFKLWKaBB7INrUTWQP5TE05dddRFtdZe1B/GT6Xw9
9GCJw3Hd/QDomXWYIuh51GT2jr5IRWBndm7OU/q5vAi7TA4VGmRE2ylrWelC66yQ
ERmLmL1YBmug6VsjZWQXvfYGLX8W2NZVoeF/fSX6aXxhTOO6mD84lQPjrJdgD+au
MJFuHY7R3y0RzxQZcVy0koqwit2IBHTEt6P6pFTxVN/3i68XZD/JLnpFikl10gXV
HSNpf5ndjURxHqVPlqxuclvxS/vB73K5+4WNLpEIgDrk3TZdw8Bi38CsmSjmjN3j
xxWNgDVfVceQuLXckrYGosLbZnmO/uBJi+5zCwxDqU/aQxQPSz8zDnAtLSeZ7Uda
gCQj6rab56pFInseFoGU4/ZS+09P6+pX1sEiNnwYEq/Tb0FOMkUg4aDi8KXuahIT
mb7wwLXoGsTyWC6rKx79ORgE6Eq9F4Vb3268XermNVcuhsD+JYALc3JHfZkTBr4/
OG9FnYznfwsu3LJymg1C3363GMsPAxwpNYSKAZSSLaP/fvBYpzYvlpxbY47PBpGQ
L5+Dx/gG3SHDWsRgVOk4MmAJrb1ZdYfiUFCaF7e6DwtGFPBV8Yy0vOb6MQtMZMuM
yWGp4DIGMlKc10ebCTIMXllVKF2bQuCIskAANKhCv9uWS3/Cc1YYi6D9yhV/7FCI
Bwtkp47XdeXHysW0WCyrrnFBEyLRr+7CZPD4C9xEvdwvJla9iDjM7hHiNovlQH5L
+BwouspGgDxmmBgp7ScNAIReCTlI0PP+McmhTBq7i8DWg8XEmXqVLcU45rSl7QaE
vaJ5rKwad6kIEF3Zb9dd3DjXIsxZUILKw1IMUYc6unVvd0ACYqdiF76gP+2fZiCU
fw6e5C1g/hG4l+xjgSbjpzWDhBjP+cRpzGGcscn3dryKitvswo6KEkFBbYXRPwBT
22/9T0kVVtHAtXWthRc6Gg1+flPiKQr4F8W3DOpk4d7Ah7ik/ylp5tgy6oO14SfB
aAImjKx9libGj6PMjO5EAriO7dljN5oKAHhjOK0MD30Vg6gNhrJ5c5w5bqaMdvPK
leCC9DziruEOzAV17jwBbVKrCk+uWHgq80rIQh6oPo59UexOk3eLuUWPLMTFy21M
vWWU9/emXDdi39gPNISvyDW6zg4N58/aBvS5wH4ebG2hTBeX6a6fC3Hv67RUROzT
t/AjQH4WzJUYO4jhv2lVIrcxg3TALU2co+GPSSLPGlD2A/H8085+4ahtBjrlx1ja
f60OoGi/4nOf29ThualSupUkv7LyfEkMBUQi6QM+MflpcUOvFpDuen/CNIAOXYO5
JzW1CAyAEhdKGvOb80mkA5AQ3op0ebU+JjYxwXRFG/9qQQnrZFF1bcWU1vFu8hBu
8oXdPH/gu+M1fockNjae6NFdQCbN3UFxP3Z0LA+1/OmuYBp1g+z1PM5/4SwI102N
egTBb/Wxz7gBpuIZ40PA2ibS0vVx3pobXTgNI65P1usW46HBY5jKI9iJiQsd1x9W
muCyKBOU3BO5suivVWsP7zRl1UyB24orv+ps/FcNrxDjN/tsufl96Cw90gp2Iocl
SbCrZ9OzKhhzaK3MAhBdOMULASt1R9Kc/mHrSshAXzB++2c2nbYt5ZoPcu+Y+v/c
QiGWP4K6F7yD5AFCvRTlO8l6yYZAP6u0MKV874FlU/vOjLBstnKeRjuEssw4E3cz
2HQCBlZ5WsdW6skd3C289FR9C3xK6zs2RTH/6S8zBwc567UjSQdIjz6FPlUFM/P8
ySCGyJw7btU4iO/JwCJv6zf23/gbYXP9wW8W+lVxqVKtmAoem4nfHZNXo2t1U8H1
Fz2l90GUz2FZ0Ktyk0iClIm9Jk6RpNTl6HRFierAqqUyXEN4BJPDClMK6ZKg3jby
KlEN6hcwpK6YhBPG2VQ8EYZLV2Dgxm9s+USC1B0GLWszIA+DM0rNKyVTJJXHlYc9
/UFHZE0g7SAk5QvbG24YHhasDHHug2bxEmZ5c/HnswLg/rCtFfEUR/r1pu+eXXVr
RjQ6HlHM8d8byFJzRnbExZw+ZmT82FOBvpFB5p60E0gSntGI9NMjHLJrMhNV+DdV
y31EnZNESB6v5WLxaLfntgTqcvtEprQLO9YkvPeTXUeEAC34b/nADP8FrRnfVo/i
aMoifJhJfk8VYIg3SPon0netflL/iVvKnthBeaHdi8FpHpTyYqq8MMRqUQaXUrfO
rej2HJz3FAYcu6mDmpy4LLT37QmnrqL+i5DAy9rTUqcbvGkjpNc+mISvas6JbQTv
zuw5ihOe86mHFe9pCdzIQamKdTi3KYgOYgkhtnUJQzt+PdqX9HaHDZ6Jqo9BS8cF
eECiZh+w1bwcuqjL8ShzGhlFH535yFkHc84CdEPgvnnLcMGBy3rJarkOI3y4Vt6o
0bS7bS6h8pIgIOhFFzUuaxzpTwR8yPXgr4Q49RLI3BQm+Ksomy7RouCGJRPQEPaF
ULv8QQ0NfKVuZbwPJQS1qqDS+z5Zr2KtCeYNDw/xCmv7AGd4ISsrjyXke9jzPH0D
sCpx39VZ9nBR6imcFt6Wi2qNqnaZaJpMZ2pavdI3fSnhGH9HSbXq0S3aTSYGTlzu
Ar5D9INzxhqvWeL4aPlExFP2yc4LR7EXgiY4ttHsYkPihDJX+l2KtaM72xO+FnA4
8QJTkA/NcDmG7PbxyPQxJ85xegpih62PAeoxoCot2t6ky2H4HFrFw5xEqD23hMgu
uF+jDttfUjf6g/c9HjMHxZ9a9/p9vKWgvoxfovQjGb+1LfneApct8gY6qMmRKl0n
gxRqNuCTztgQ259lh/5brOcFco1HlQpEwdwpS0eaO/jOgfAltZXi/Li2kRtmcoGq
pv4tcKlW/CwUY2Q1F0iZf6sfWr9oZoBVj6/Xk2Xo0tHhDjPp0IyIxEs/YLjfG6PX
j+tE4MYDBrTIMMtVppJUlImZ9n0QRQEZPs+4+toD7C0yB1OlJ/hnRjLaGdJ9gsEn
+9eP21G1E4r4aRSJ8hTFP05rTeYnKi6MJ7dnHKuRbI3H5JBMhoT9SgGD0VR1mOFz
hJGbnOvePf5hj62VZX/6LBkL8XY9JXphy/yBhUZi/zvFOo0aHMhKe6mzQ4kfda5D
J9A2Pk5lJ0Z+SCOHv5DslENZyvVIzSyy5fs7WR8uriElXl6E4YcHiCC3mRg8BMn5
wkwt5xrvA6FM6lBcZoOUEvexNRcAA+bJRSEP33W62Vw58JHF30kDA195bWVZ3BIt
sIZ4QfCrMzj0VArrBIWPAEg/KzDd+vj9c2lRnfB58Z26AABqdE3vlX7WMOH4xHoq
U4cQhPXMYOLegRXxs3pYt1WRYjv0U925YmmpYDW2MTVNzC61WO8A2sUbnr7W+0NF
cweFKStO5YvcORFv5MKTbACZ/CuDk4mKjRA3J5XGWDFCPoyWi2qzihwbHBLJjw5L
oYsQzsb2x+UszYCUPz+tgJtHjeaMoqZojazvze+9C9BM/Vyh0EQbqnfIFj5lnqpy
2GAeQNSYplgg8S7VAb3HwqiJljD6cHedkEwqFbx1ozeYe0Ugj9iAd94l4vzwTMNZ
UlvgcHSrfeCscayB89RQ+kYnLEYLXV86VSz+XIevK5DHP9VvnD48boln7MB77Sot
sSxA1XSU4+C/VN4EmldoEXGE+KabbDsXA9ma620ROc4gedBtVbtree+zRAdprGY4
hJwRNTK//ECJjafbUFj8GQ14oex34xAnvGdlOZa86UaQomEf4WUY73Mz/07KRnCL
9DgCdl/RKfST2QVpmZyaPzAYGcxSvtPwXl4NP9tVAkrrps1TE/NiXswAaZ1Kz7NX
/XIB46OMrj7aVtxts/Y/z566821cLqYgqMymHdrKACdVuX+2BNSkVprbE6PEk3rz
XnIZIdtszNxJNyCCTbQ59hfLkNY3orN0qZTNOL4BvG36NxthVmLUNlqwQ2etNy4b
29wgI3O6HngXULytqnekZyZrpPoubkr5K/5zc/04bJECaVNvUDVEyDQSk25Ni5uB
rHKNQnrfEdYeS7k+6B+ySILlHZr1+IksLtBRRKhRge1Z0hfbKSRShNB9cS8FjDfh
7DBxicF2k70kf/axRKi6ThuONGJ66fF2VJ0+mOR2WSUs4FMJfnwdzZB2G9k0ftj3
iXLEDCCIu4H6ggEet6JUG0dlkDk1UXr8PoRIXBiWlYI5NGwFE3lBqsOit1I5eQVv
QKOAb+EVtNMjeQOzzfAdpP+3JBEjuCIrVdtOEcduXInUXTxADRng6cEqkByz+3kh
MWCCfQjgtXAFgtnYNovk3Cs+p75R6BvqbUr+mmEgfjEM2VMnR5fz3xBFpTtgwAeh
uiSbokDghHjL8vrHSr4/gQ==
`protect END_PROTECTED