��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki���2p$�/�\�	+Z�j ��k��tV��N�ￔSX��75�#a����4n&�~;�Lh�@��R�R߰ZC�hÅj���$�n������j��kiSy�/O8���"�+֤���D��4�_#�k���zGR��u$��6�r-g�� ��i�Y*�*L�k+�����{u�A�g����(�y��c�E'���LczY��M�Xrw���$�ͳx��N�6;$�C���פv�}��A�A�:�#'C^���1ڌ��«LR������T��@�*FC�S[q��s^�����ѕ��8/9�@����za��}�{O��?�U˞���\1��ͣm��he�t9��ͤd��@;�SZ���]�Ky]�]���Q5�:}Y�F�UCm-U�x������D�ܪ�e5��CL^� ���ʅ�:�����i_�����롰U2�u�j�����u��(�0Ey�f;��� �����r��<����q��%��Q l�-{%�9�a5 cv{��c�n^���ɨp�5ERc��ӪE�d;���_l�K�cd�In�.?��s�C>P�b�O�=n�B������/)빁r�P$S.���5�se�̉����ʄ,�(c���9�v�qw�[�c��<�z�H�^�Ta�U\�!��dD'�d�ߴ����V��HvG)ib�o��:�i-s9z� VК"^�j}S�ؿ��.,uE�� CS�2�֌�/H(˅�ܫ?5t[H�MtqLs9Y�vE�#�ޣռ˚�	�Q̆�%}�����\�1m�:�$|���o���;�\"�A��[3G(
�_G�ma]��q��N+?k�M��yhi�[���ǖ*�m�����ˏ�R=��-y,]�J3��5�M����{��-�UT�F��'�D��:~��9�#~�s�H7RH5��Y�C�t�D3iv�L���Y_�����U�'�I�}�@��ɛ����A̨7v#9�_(zZ���9 �3��K�2�-n�6l���,@�N��r)U��H�yk�sò�9l���3�a���e��-��i8w�B����&��3���c�`�Z�ci`�
�<�����q�삑��?�8�Ml��y�Pv.�	������0����ܺ�W�_FZ�R�0ᣅ��_�.h�L��1zŀV�4�(���⇶�50nҦ�Q�~�J�3��Γ��A��y����!���W6Z���V��y5���\�Щ>ʁ=�_�>�fm]�3>���d����nk�fBW��5�8n� �d�
��<�}�*�AS��m��s
۟ �*c���Iٯ�����/�`��[	�Je]�ú5�7���n��5�)�n��$����P̧�rG5��*��e��M�yd�ର�9��8(R\	�OVGtQ,=��)�*(�L殘l@Y	d��)>*�j����nWx��:���=O����3��!ۀn�O�f({:�ҭQ�ŉR8F?��1M��c�<%D���*~%�������y�#t�{s����$��Z#N���cL�K�B��9QIC�	o�\�s�ԧ0�!|1?��~ _	&|�B��ͬ�H5>�#�d��G��tüu�?���5O-x.�t�:��dC�ƍ�>!'˪%�bo@*"�e�]�8ù�g�VD*�S�	��O��P���=��4���c�%J)��1+mlev���J�@����8OS�z�n���/��}�jc��l��ݖ9,��lss^���]@��&&��{9��hI��ʤ>b�,W,M��`���C�ys��w誘�d-��d%�Nœa�F��M[����^��/VNt��LW^�Mu�es��d�7�+�NKw'�S뢾�f3^V�8�p,��h�����t���R�wk�մ��uY3��P�ǺQH�>�|���f��n��`�**�0���A`G�h+�V�/{���CD���<A��(d�ɑk�a�O�3�>��14���GjL[��ء�:$���r݉K�Q°�s�Jz��~S�aW��֕�Z
7�S��v� `~ cX��U������W�i���@�bK�|��D����8�.��r���Ǟ7�s`����yb�0��E_�kO�ֽ�d�m��9#،VmW�F��߭}:)`�1!�<�����N�Ha�b��qB��Y���X�X�����>m�X��'�>�0�=z�vL>�Cg��ml3')*�2 wY��Np Z�+�$�*� �"��U��oSLBF�F��� ž4j�Ҹ:�ঋ2�h8��H��T�>��cď��9�����D��+�ꂊ�b�ϥ\�}����޸��X��h�=\��8���j�'��L���X���`|R-�B�/h`�8�ط����U�2��E:^�Ճ�:kI��2�<`�ȟ
�㉓Fi`�W?B�-�f�p�3�$�U�e����)����ߐ�z�L^6�n�l��9
^�P��[�� >�,mJ�o��������mѩE-�γ�e�����;�o���Iif����kqdk�0E,A`J��W��I���'�g6lT6U�e�JX��9L�x�{�g��{"Q]Ү������w��`ժ��M����4�a�os�ggL;NM�Vv �,l�Br�2��=��6�//�o Ϻ��l#���6�oU�a��/9�'=��)�g��{�)��}F�Y"��2Q�S����=+=���!�aFe�`�y�ЯF��%���P&zSxChh�x���AQ�����eVP�S,B��_�h6>X��5|�j�a�����Y�s��H��ݘ�Ae�xqg�(�EU���Nk�Nɐ��cNGb@�N����YR���-z#ͭ� gLԺ[2�{���J���#A����j;�OU˷�lԌ��@�P-� ��,Ex !�Q,a����Kp,�����*7㘊��/�K���~���f�T2!��@W����(3�N�|�@����g��J����q�IJ!�vwy4df���@��Pן�^�(Z��C�4�$�ӻS�X8���/V��V���u=�:���ɟ�ӛW�沭���0�ԜCG�|j���#�֬*��fBl��q#��֝T�
&��Sy�<D��]I�K��R4+$Z����v^��(��"�v78N��x��I������W��};%R��G��&Q���L_���A)3��W��F�gO2A.�0k����`�e2�f�Ƞ\�"1�����[K
{�Tk-A>��SIZ"i���%ɑ��WP��惎O?��}d,a���k�NA�ʔS����!��.l��
�봖k_�#Y�}.9�tg@X'��D��ts��7q�����'���nӺ��R9=:Hi1���vrt"�8��5�S��(؟e̫  �E�*��rĨ:�����&�s�I��[6%K7>�ƕ���T(Up�X��ق�W�fw��,�g�dT�[P<����Jg�^�/��96��- 2���9S.)��fU^I%ֻ����A�ǃC�)�����5� ��J��o�6�c��c�i�G��J���<YmfqQ.ДP��Vy�0'��� ��L�AP:�&}�ve�s��ͨ���� ���t�O�Cc�3�p���9��ú&��^t3$�唷�'�8������&Ј�:�f���:��cU�ϝ��;ᝧ1�bӠ	��g	�`Ga����҆���R�Wil%?1 ���Q��5S�����k��r�(�'{��p��#��P���x�Sr�`C��q��I��tu��4�1 -/��( Ur� 8���31#C���.g��Ӟ{�����9XH�b�+V0�J[�ʏʂD�
30M�o����T�>��4�7������M�t�JUP͋�n1��$4<��ڸ56��=�3����|��d�o#a��B6%G�[ļ� 4�>��V�ȃ�0 �r���Sz��1���RٝM���w�/ɍ~�!�O�ϰR����F�$��YCI&��ȴ�e+2e8r�D�V}y�d�ΞG[i��5��u��Ȍ+�B>���W �F�:�y\ٱP��	��yOIs��S���s�:��%=z�K�c
��ފ�J&��l}��؞�w!]x�[�&=k�:�̿|]:T��ȉg<j��k�wn2����RmقD��:4�WQȆ(��%�a�#��5"Nj\x�zw,����E��P{�u�I 4�%�unp}g��פyQ�����.��e4���Q`���ݩ�Àl��u�u	���L�Ĕ]�!u푣�v��X�fO薖�0�7���nr���Y�6Ta+�����r�}/�p�w���4̕UD��7b�XRy�⸹����v�{��;�'Lin�vEܲ� &���;^��LR����-YIϙ�F�~�� ��������ɦ2>A�d����}�0Eӳ���H�,��\�=��o��]���unVqr��?dˋ�(M?f�J��>Y��a$�B�4�+�;5l��"ݛryg�����n+����Tm�%'��Q�5���3��\�+�2�頎�8t�&i|�mv�U�*U�M��xL��m��O�0D�c�+Z�,+�o��J�Xd��]�/f�m�:ԁ�����;���}���@>k�$[��Ǐ�+��!�9=<91�)j� ��V���<#��d���%a�,:z�� � �2�� d�%\�TwppԀ�G)���U��A�3�,�"�CJ>���x4�!���r�TLN�ʿQ���AB��aA=+��i2\�^٤�LgD�is�vBF���x���'7��7=[��������\�ڙ;T����8�T�v�7����k��]7?��B�C��O^�-���Ă����P��e*��V��v7�4uu����0_S<0�M;s����eM��cS��\O��kZ>gSU�2Ev��.$6�W�Q���%5�����^K#ڨ�ڐ6���;Y��1=P[�����kk�lW�Ɯ ��:�_�9��$�J�Y��k�%e��]��LZZ�F�2aO��I�ɶ-/�A���_+�9J���/}w�n{�aG6S琉dts���ڣ��b8is��Nǝ!�K+0sN𱽊�R���_P�oFi�<� ��n`xg��p�y�&�c���x2���J駤�~�cS�V&���0�~4���)�q���^>*�ʑ��6WX<!�ĥ��b��U���࿗݃�=�P��X�4�ۆ�(G�_;�s�	������&I�6T�^a�U�in#��LIF��|%�5�����9v��慠�� �^���_묃6#�J�\�y����.uB����=A��9�k���Sq��o���Wi����$�� ȁ�/v:�����������O����<��+ꩂ�)?��9�Q����U��?��O���BBى}O#���������x[�̠
8�,*�����m�Bw����+��A���h�Z�V�5��ض^�zb�ae�(L�3k�]=be1��0��7�颇��]�qp�<,�<];�z���ȇ��J���s��~.�tzH��uX3=�'�����xna��$G�����y)��ۡ���-�$�X~���Dh����,��T�T!�ϗ�9���t~��iT�=nR<�Z�66��|�E-� ��Qِ,i�Do;/�}��ȾQQ�)��T�,WL83`A��͇0c�s�`ۍX6�]Z���G
�&������Ɠ��L4iyy�g6E�kY�^��`���8��7�,�qU�����*亵���B$Gܼ su�-�<k�; d�'܏����z�6��}�a(CjQUCA�CO�%sB�|"����7]�r��80h4q�'��>��8n��@h���T�In�ś]�ݠ-X��EX��3/�砭�����w{b�&���ޑ�O2[hR-�����>�u���i��b�ٺW�(ٯ!V*��=rI!�g�xE�u%�-�}���^����@"��2պK[��K�y��0s��IϑG�(�Lc�c������f��a��e�0���~ �;�ao=�|:�\�	�'���Ee��|c{(��o@�u:�U2a\����CW�ͮEsj��rnM�HK�0��t��G&5D[��A功�ɓ��bm,�0�.nlw��[�  �H�� �/O�ጧܬخ{�c�If�*/��m���h�i|L�o�q��2Ԡ�/�?�F��ږ@�$��N�\�Q���_W�Y	^�@,��J"<���Q�Hَ��d�?s�C���"e�(��i��@	�)a{��ﯵ�l��
!xl�=�GID$qZ�
�y޳�/����j�'���PϑG�5�x�e����0�6��loi�,o9�;�R*��)�kO�t�$V��Y�z�\�÷��l��cR�a���?��7��
��aJ:��p�ǚLԏ�\q�5m��U�:+�n���7�CUÄ����)k	���(yŚ����Qj��S
�B
����Rп��s�m}�dRHs%Y��Xb$�d��D>��:r��Æ������g�12`"�wcE��(�-��F�?�#����I����ꚍ?�ᦘ(�Y�Q���M`r2��J��[���0�Z��K�׺e��	?����)���me��?R�����JfsF\�4�ɬ��(94���N��4;��RfwV�Ax'oJ(p]x��|>N�RN����c�;�O1�}�gZW��7Lp�f�t7(�M�V�M��D�r��2C$:SM-K�},�L�Z�X+�`9>�H*����lW�
�%x8�$�a�Q�l�J@T�q��]˃�Ekz^	Șg������q����1���yW�]�dL�T+w���K�����B�l��q����.����N�!Ju �˕���r����ӷ�k�L?����GY��H�qS�Q4!J�g44� ���*ϳ���R��J�d�ɭj�,�r=T9�b(��sD�9�9J�e^��7��9�A��3>����}(����p? F{�up�,m�Ӓh��z�hv->wZ,���<��$�Y�߶���K*�|nQw0X�)d�CK�]�q#=�8Wa�%P��t	k?p�g��x�Iu���r+�a�)R-S�]Έ�Rmv��H�����FG�JBV�N��h��!�O���P��t�,l�����qҸ�b�`,��- �~����K����%��r�:��i}�znX�N�*)O�P�6��=C��� !rř��>�;ԯ�H���ıޥ�c�os�%��{��߉�ɍDG-����7�����k+I͢ ��'�H凨��d8Nrtaf��,�؃��#9�>0���T�S+q�g�b	��;jZ���cQ�k7�O�[e���_!�I��\���ڲ�81s9h<d�޿~O�����a";_L�����'�.�y��5p����@sU D���S�E�#�Kr��� u��ڽ���K]�B�x�<�D��=]�O���Y�~/�ni����/��b���-Ai~�V���=�Ë�T9�	��c�]����_��ܨe�N���lJ$����'����u���,�Ԍ�G��ǵ0��_� T&���&�h�rQ��ލÙި�=]��T	1���p^�~�YU(b�c�!��$þ��Xe�z�0j�eK_��uʾ�=��2'����1M[� ���4}\�H���O�:���_ؒ�`��=w�����#���N[�u�鞴qFf�J2l�����̄P[��/x�pP����/���X���J\M��Fi�M�'8ǿ��ek����`k��U��c�0��B����q�ػtE��E������L�$ї����p �.F!g� 9i��y�,�����@Wi=��*	�_��D2v+��q�lǮ����b8[l � ���
\%˿6�[���9K���~��?�-�{|�;�ԷU)�Ra�fXGAI�z�5�����Tq9j���������
f�[�^M� a����Ν �Z�!?��hܳ($��.FI�[0��~�� ѽ�q��:�p��;�P�X�X5zm�PŌ��9�&�����V�?�@Դ$�ϰ�$�os��R���E�2�7m��p�A"uI�
�.������	�����˞w?� �+�P��y ��ju�)j�yK���r���������ۉԷ	���o�za�E,������G,�ɛ�)B��w��rю$�.ˆ�]V@P#!D�}�/jܞ/����R�MY��AAK�c�*�.����μ!�=^vv˭d��cy¹����7��S_Ԓ�"�ؑ����:Q���
�:�
h nK�t��j
Ns*�ӫk�F�vڱ`��D��G�Ĺj�f�53a7�va��L�Ojf�6o�� W�FA�r/&Q��(��ʰ����ϸ����nUb*Aw�|P�������IgX��G�<_	�n�j6Q���b�<�V�2:�6��;P�.��uə�#���˯��z��PE�:n��G�v��3Z#�񝩹��v>��4 ��_˺��?�l�a"K�D�ۀx�K�v!�����0z;S"��J�tÄ8�V\6�m��V�ϖ�rߩ�����P/����`���n��GS�P��`�Q��fa�^�a�F�EN���|�ܬ�в�T�,i��w���X'^x�ɑ�U�I�L�����D��
e�Qv��6��e�tY�T���O��5�3����������zM�Ŝ����A&�]����X'�,�bY����Q;
P�#��;��ߎ�
�F��'5�����~�~6��2��9��ʋ0�6z>���FU�4f�S�(6,@�u���������1ϖѵn�M��О	����3��d2fn{b�?��̤LX��X]�4;!p]��ã]_�����z��b�`�~-h�j�B��XC}�+����ܧ7F5�9Mc�	�:E�mg��>~h����´<c��/��w<��rI-��oOAg}g���}�>���E�4&5����
d�Iϼb�"Wn������!�*�B�*��J���v-,�x`��9�3[,w�B��r�4��:Z.|Հ:?F=�J�uS�{��s�7�^g`�Io�ęY;�����d��;�JG�x���?�^� =����pY"�v$P��Ѕ��m�ܵb��D�i��;6�4P��&�m�]�8,�u�@�#����#�������Y��m�y�;CŹHžb�nP1z�4�y.dc��m±�����Ҡ��}����F�u��]�c��7��'g��7���占��٢��_<_�-օR(6ew��8B������p��!�c	��œ�R6X/8u�}��FEx#��!x�&��
H���W��=�od�u�BA�fH�`�>t�;-tE@��c���5;/͖ͤz�0�ǥ��J�9?��Y������l࣋��J$�Ӻk�ƫ�K�O`�JS#$�]��f�1��\aS����k�\H9K��{E���@�d��\��������&U�E����C��hvmʱ�����jf.�5��o��55����!���F�)ׂ}od����ж�I�4)�u��C��><eH����K��[iT�� �q�:63,^�l{�4UňO�4�c]A/(�r{KFc���A蒀㨽���}�#��]"�TԚ�$�uSv��D��_����aK��5*�xJ�uz�(�nD�EiY��,�a6��e�4I{�[�u8�	M��G�U��Qn�刭X�q#tjQt��
g��� ��#>GeA��2�ry,$�a�A�R�BA
���=���	�Ck����m�T	3��Á"�n�f�˫O<��x~�G�.��3[����nP��طN��%2=��QK����7K�ӥ�O�q�\�`��̾&�4��`�� ���������n�vfa��Ek��b�w��3s��$�-~CpYX�<aH�]S	Z]�R�{ۯ�zҿ������s`��99��a�uK����.(�<$E��>͚�$zN����A��$�L�^S��D�=-o�V����D!��@�Ƃ�U�S��PDb�%C�S��5H�s���+;h�2��I�y|t^g���EZ�)������g�v�n� 7q����e*���@**�K︔
�c�àĆ�B[m�; C���+{�X��5ٵ!��f�p�h��(0��93)��@<����>"}������C��Xn���]�Us´ء-��"�[b%=r+�5yZG1k�ڻƐn��.�Y:QC3����͂Om���`��I C�(�?��44|�ť�;�����M^�J���=��vL��Vo*,�dJ.;	�6�W� �)���fx9����W�90�� �iQ8Q&q%#�7nMo�jS~��J+xj �`t~��a��=UZB�?�v
��c�ތN6H��|��5�����cÌ~s�V�㞢���臋M@,>��$��;!!qL%����_6 �kg�S��x=��7B���<�-^�{BR7Y)�B��zI,���y�Y8!3;�o�|���j�!Y
�y�QI���\��=��,�:Y��#ڧ���z:�ƅy���C�<S��!��� M�8׎�X��	�%����\JT��2�s��}>�*���̏im-pge�<ř��lj�`�i���@˗�o3#��1�{!�wS��N�x�A�5D.�w���;�u��4�\|�	�̗*|	hUm��_(��pZP��x@Ta�Ďj�)'I���׺�i*|��}˘���ad�Z/����
m*3����R���e9�/�.b�6�UC�`!
��w�Dz��/����}K���]�����ł�3�aZE�$Xp?�"�znkyxt��N
�:B���'��X~����ѯ����qx5N��+ҽ2�(�����dT�V�G�~�,Ϊ�9���C!^�k3�*�f %R�>��_ە͏��:�¨�V���r����6O���(y#*,�'��|�ROH�:�#�<��)S�ں帛@SF��YF��������@Jj��-