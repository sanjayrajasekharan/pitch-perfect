-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rHCU7/oiuSgdtFGxAKXS2z01oJTagAlNi6YpnGWiDfmE6keZTUmTCPP55fLzUM/enRIQKr2pJOXZ
UDiJjiycOXfPpCWgOZSeHOIVlvGUioCcDRsHoW5RTmoVcurLnqju0zj3zugxOQCaPeuPfCXzE0G/
OAX3Vcjr1X2A6aOefqzu1kOHm4/QEkc5oK3mqavVmwBmv1cNYeLAg5t0fNPsVAdE3XSVjBTVFeu1
w+cv8vyPj9kbhmjtZeksrcU3dinXlbZWlFYEjN51oeTik3W4j/TKjMxOiej4jKiVP5XqYrzOzvrL
Mfu8WuBRoIu2Sa8oGv1avXDEWgu3sp+OoYPCgw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4176)
`protect data_block
HBm4uNfQsiiepi1UYcmRbW8Dmwbn/tvei9PmRNtR0UW2/EoUhdCpn91uHqEbSEVdNK9du0tolBDh
KuDAlTP7ZoGVVD6mXJ/NB7X/sFGy+/OihLBpKNwdQ58eIW/9MRlHKyH8uFIzDUmQORKXl1Zo8pj3
BQX74jASjJ6hxV27dyN4M8IDWRojWhWCxeXnDTaJoU2bpaHDLJhK2ATG/KeaM+fb9d+Qbx1Wf7yU
r99nTrYTO2en0iIK4oNT3dp1DEAjdHPZrAuloWjnwQGNpaEscMpcIL80bNUeApa/PstLNiYQw2iv
hySCNqPcjSfDjbBAF6z5AtpRt3Ksk1LSUiF2vnL2lHV3ebgNJnx8GNO+xxNNOJuFT4611NO4uOKK
one1YBTaxX08ytw6hDSsxVwSnRSCdNJ7DPQeNCSQvOeR4ole2mtZ4dYxL1uY30Aq0z/1SQrIpNmO
88j/3KLzqnfcFyeQsMnRSKLvwEL6SFfwUaYIeTwprFrFLbbhcrgJtKo065kwNR3E8qSmXqNXDMni
7XtWYb6/9dWvWh6s7imApbRhknPNYibdo3SZi93fCiFLMh0Dzb4rNdHzH0t+lEqQhZzZrFN1VF7g
0VZ5EELop0XOExtpnS/JBLfGFs37Z3pUikWYb1v6QJzmy25voQnvXhvdntKztJASy97YeXdcO0HW
zo6J2tDvmA+pfz3bG3fm84+KdRNfz1Pi+GRYfRH9CYuobDvpa1j066e97vsVp1gB1mXBcQV9zUhm
fxdgYL8QwlJLvkgzpZOBXNoNL2AjyndJks3eA7BKfqB5nTEp5aYIjbtszVsC13jYaxUbc/4IMHom
pnMDYFOdexaWdfdgu/72YblIIS8XrGppFhULiiSADcojPZA61gGLErSP2zmRSSe9mtKZt0a7PwtQ
mC2tr9preWQBPmbpf6N96d4oFv4vnxESskjUzrLXyqvuCXmd/+i8WZqm/EIZC5ugJ5/Bcx5624rh
n3m+TC53GgY2e2pOvBpGt+kKXVuhJjrZqKTm3sD7weCWM6liugm9mCRgxdTsHMCQc92p29IgLeBj
qUGFEWVDxeLplE6C6c7NXWa3omfDQTjJhADIDUeFdLydKi5cBdQqYqayWJgiIWzYfRhwuKgetFWn
qNohwuz4b/vN2umpjlOzgqeZF4SqudxY7MCrDtNl3hET9H0tRxTPamE/kWnhTtrPFnVBGJ3/CLm2
DlQ9HoZXr2jcXAZzgpV3T2T3n4RuwbZcXEPqhDwZQBnScIaN3en9Bmpp1lisTh1JPfGNmqv7hAZC
gyhQpK5EwotjO6ToqRS6xu8d+L5gOrE32bJjntkETaum6oiob39HITjEIW/6tnQSFSKPOwxjc3IA
tPJVNVikb8eC8vTbKQn6VzAU1cXGwPYzA4M3LfcVh85qcr/2p1e9N1waG7dVpKRPDK8lxcTtouxE
37QHSvTgy+qXUIemABARZXwwZCI9IhPqZqfCIk/m+uIxW/NYKzsHo5bf6zi4PdZGFg/7CYbWxC/T
U6mtdqU+1/cdma99JZVAdmtGrD8rfWj4OcGWVCaxU2YbHl0bf8VPk//fPYw2pw63SGQkkB1Mk7/W
hP3RtDlTrMI55rOWNFaLqujWOjL6abu4dt2Aam05aasINqU+iTH6/6TFul1MgKFu123am23kaMuA
2HFT5EvML3vq+CEej10K69uVo4JHhrVGMKoSw80mi2vE0IJ6xtfS2pqWlKJ+xMHhOsw6QDDoRAvP
BDeoCcnkEqxWDFosvyxYpmcNlfZPthZzzr0gnN8PK76SdZMFYzN4aC1W3P6Hu5hpm97h6qMILefH
4xZT5Q641QU8HR+3xxwX9qIH5rJy2qDjqAlQ9mGOq9nPXfpJ/dOr1eZGmGzJUoLAk/0c/anXbYl+
6dhpIGAHkdvXH9f+C9KUWa/mDT9QsAzVi4p7Z6Mppt9bLuAREE+DrfDhF+N9O2yf925KqZ+mL2s/
vv5+kNzceYGqCG2i5ryL9Fw6T2bVgGMSnHbXxTUfbWNFqXQRHrUzkuk65UBIa1fwyka64DYZgtMZ
POlPyygFFvE6MzUyfDYPp+59eeFxZpP6o197MB138wTQzi6rH1NMszYDFU4IRCwD/95e+gnJ8xLh
C70OoEXaANnOGj5gDjSej1RjVK89pUeJZFTfzg2zFzpQgUJTa2Tv1pQ9R35T6LJ3SyO3XFf8woi6
fVD6KTYUQXc6l4aNCPI62aYPgzKK0iODGy6LPvykIFlH7jNr4IgzV/WPUywwmZoKNlwXO5tzJ9BS
MVI0EFVGgREIW23G7HL1pfisrRpQ+peNBnPGPyPL8LVRBzDXx5PNEkU2Q2ZqkMk1U6NHwEYdj1F9
UuyWEyVBD+3vGnA/qR3RtDFJctZa0LqzjfiJaPAA1lwNL7erAid5SD43kwg3y0T2j7aN8o6uIwX8
3VjyJQ16ognhm8G5cuWHXkN+4WOjvHMwxLVSfMs/m2m+JHabbWVAGn8wlgRAAYQa/Um+aga7G36J
NHAlMiAsXMkKpoMsOgK2ysB8s2FLARC9ee2+4sO87PdA0VRzsQnmyAG8ZFxAe713QK3ShGBnc6Y6
ZtbQXsN1ZALtYMVT38T7mnZ5NoVbOp+Ut7ucMRQ7SZVU5Wh3W3dWimgFTDnMz1NhFgxSnjMrnn9x
c55cDUridUl21mITCr5VFBb53+Fjy/S9nLz3Na1yI8R1fkhpAE2IMwRKKB5Rdvp4m/V9fYYaZtdo
05N10xVmNtSqOsja1yRA4j6gt6zutkqWkxTzhvlxPx0skd1Ba2htRPt3F8FlRojtLxPHDo3AGRTw
5dGczC8J81EDXozKw8dqKo/lRghinyKlNuMhFuioXaPqB4YKaX8EPsZhQ97rCZSWlZCv1h9+QRbh
1Ey5rE9efwfhBoVGWwvgBlAOeemXczNHpKxY6sFF3ZMm+NDkTO9HZ6tTmERR9AJz/z7dWtBauMrb
GjlQK4B5Su3T7HGpufNq5tLzXNGD/DUn86FY49BxItLaoR1AEuY9nmFvz7ZcggM0DVzCzPeL4dMz
c0tbJ4aVsvOcH9HHQUimmFSZiKDBg8aU+V50PyjThaUU1nc8dRxfTJmex5s7d1fI7BEmjqzxOUv6
QduECxn6mIclghuhndfudGwa60wtEqbcqjb5wnoDNCZpKhPWTXaAM/4YASzsl1lu34LtsYZ1Ihoh
WvpPDopB3WTEhf5HdkDQJ+Nx64zfhS7PaOKIY5hmjfBXLhCg5l20CIn3E5Me+z2D0fOHCz60dJ4z
Qv7gs+SIaTKV+A1q/EeG5LImkJ/1NVpzjDJT5gQ61HSIRsjTmeFwf8FNgEgQzpnb5IMNU0msAG12
68wu7aJSPD50arC3OFIfAzuNmbr4m04vCO95cij3a3G0Q7t+wLTxB5WRjocCNfLw6+9hG80XuERs
fVW40YwgvE5BK/GWw0nqYzScr+EYVJNgSqDXK5SeIQsMmP8jV0nulseiXn8lBmk4WWDM9uAGV9Fk
MhJUD3zVD3NxM9aGtZrsNAbMJY83kvkBoJ9YfmYS5GsATe7I4Dm2pKSZ16Rrfr9RghIj6EY4FgiI
qabdDwCWCc0vcXxC886e7CE2i6cqkp4y9R3GoUXR16GOApciN4ayS8p6NnzESrILEWXc5DEKA1fl
4wi8DvAsO1iC3ggm7ui7qcQ5oKlUjSM9/6AhmYvnbOZoc+w6Zkb0XUZXOxuZ2luYKSE1pYq6miWr
omt0N5Y2U+nmCoRp3CButdDV7yn9bRVy4ZN10113FXj5n4+lNXfx9SfHT9LH1MKULs7ACcoh6kpf
QBlEg8lvrcKO/2WFHc7kliFCyNEerr4D+jKZ4i3BFVMBYIBE3S11LMxmDBGrI7zVhzna7T7nMIbs
FDnWZ+AulTTf5hSLoCndSGDN4H9mNm4HF01gYZ6//hA7K/9pz9yM+nq4ea5VrmABtPx8/iQrxe5E
/lxj584xoHfzdcTtzuXBccXzZlhsofFYldUScPGnlv2PG6CgQnwGJ5VtXP4h4ItKAry1zBONpZPt
89F8xiwVfJanIXD/yW9DV1jHtC68sdD6KRew8Qj24KQ12UDVvMhnAAO86NT6w9lt4x3EdzquPeMD
0Kjkzq+IEiGc+E5zb0dJTaQMrboP4vpJnXrwjf1JidYkm2TEHZi0MpT2tsoFaUVCBuMrxCig7MWr
jo3eHjqwjsBtldi/eEODt+zelBFO74ozRCAj8fGJjlqT/BLrA6uR6zNy28N5wnw7xr7wfapXj3+k
oJeMRMWfpkKZJ2+nUUcW3hFjfM2ykSGN2S5zoWG8huKyd1FUpyIV2KRZNuRGE95TFLTG/AcdC+ec
gmJ7mE2m/LHquingNJSPTBbPFGAzMLX4UqGiLSr6kaBi15OSOpXdqRU24HqV2l3Ad867Y+TUj84g
Wwv344h70oA3kVhxqnyDsnPmYEzOIahLa/HOx7CW8AyD0gHi/9L3KwFUvPjsGS2MVKQ8moCkYsKp
9XABDGiUOEdA7WeKOX5ycJmChvh3uqln/HBTENV1o2laYJ2lpq159tEZUn1VCP/ZisftlU47BSTa
KAnMHEL8bVqNotTcsEqvtuvrWySa4Y3zqfM/p7uQG/PYxbYFf6CWvwBEWPwTrCScz+YH5jVYTKQG
NDlytYmqFeCIIUg0soyUfIwnCMUwQHVZdqPH3cZzh54G+ZCS7fnmm7OBkEwcUXnG3JZFmQeb4mMx
xsESVRVupao5izU7rcL6UZ327z9zQ+NDK3TsZp4JvMumZ7Z9ku+ehDAwgNzrVGQFlIE52Q7i2fw4
7ZVg0UpemxlMknqrPGEE0wTSBhdBLgeOmDCEt4mUHGrOqIpoX8mdMTqw3Fn0jkBwbyWkBFfzJRyS
n9w6rAwB6R4ViHwX2YwnuEhf2jcAl9etWzhPzmC2Wup5ZMpsUALdVgHJ2DDh5qwo6Sm0SdGUlM0V
JwSc7apBi851LSIF5HBFLhZ5Fc6p4bbxl91czyOi/f6WAGKCNWmIQdFPX3QbVik15KNjwWshtpNd
tbUqwExsXTmimjh57Uz4w8D5U62QHQViK8Wc4J92B+e7Wzlp5TxIp4XE30FQxWV5wddnfll1jh7i
0mboxUh/JU6PngGkYfmdd+A+JtALCaB1MkSLYRtXRPgnuFfLJBvzlHHO8a7A98hbMRSWtydQ+ft6
a6tQ/U5YIu6r1TgM6zjVLxqiVmQT0Me2+H9HHTboDGrO79eclcA/wpBNf6TcG7MMSZDfB4+yvjXD
YmxEzswgqtQCYF/dyhsSo/Az4Lw7zvmJTbnbZic1OExqkH65C+p+swIFLEF61F/u1JfTv7A+UN9i
yI6XyCGyjTZd60n9akc2rkxVT7SDtS4tr+KI+19QyTEde63iYQ5c0AChOHjJYEcQrEidOCfw8/aI
DeezfMAiQX0XlxAZTV2J/xBCJZIat+ako3AsCFAcJAPlmEe4jSY809GJE6HhKpxN5+8F1NZrVLt/
PZDyu0k1Tf8GkMlyzKUUlhFou8TSMYmTTSi7Uv+6nK5KwZIfOVwM4KQBchJVPcnEPyHYADqI8Yoj
pXAHQHBx+4FB+D8Tv3/N
`protect end_protected
