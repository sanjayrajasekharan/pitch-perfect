-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
KMJ1Ii9FWxvd/cZtzkyA+iAMY7bnLH0bDZSkKpWztst11zEmvAwGHplYsOwy9HJX
dxSHv20hZ+Ds677s9ZVDgYFPWo4TG8W7KsjxyKowzF5orPm8KwskXcLqfOEVLbVZ
nWKqzDfU1z6SmUfwdbNb+lYtWK2+UzE/NJZKgi32dLQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4162)

`protect DATA_BLOCK
lJFFcwbObxZKmavjzuAvnD/70hOwgBM79GDC9UV1Yu4IoM0VCzkV25MFfW3IjePW
YFljEZrutDT/T5ScMXqIQ1yGj0leFqBh2lxdCRLgXcTVqPy7HWw+dvrb34bXUdPj
ym7O5EifndM/bJHGeAbeBiXR6YK81r9gynXyTRcvmSiHdvHqHTfl/afnDHcZLlia
kZ1CbCm62rZx3IivqOgUv6JnkakgyuLWz3fjAKCnu94W6my41NfwI2YgiBY7ALZX
T79/oCD7W9kCFIGddTLgFDo/G42ZyU5OLI0uL7Qo1q7IT33EOyJoUm1dlEa6F57E
ZZTna42JMvuOs+/aN0kCumDHp+njKe9EETIaw4PsHZAxMQ42fTB7hk2qeiWHo96m
196eZaXtUM0MiJ6OVe4vzEBrBkbfVFIVQAoWxdnyz6okkv4SkPyIOtaAx9/8oq1C
r6InMCg9ovIuoBLhZgbelyhfogkb5dP8GCsXlGy7cf253SVnXJDsnGPksu/S8lNa
CT9nsdQhnpYTyObPMWP6gjuivH6DeDYKHiTOBSIqlDCGF8BnwYDHVHDkVB7WLvRh
3UwyBinqyCpMHC7KeYDv3V92smLHO78N4/7cxur0SEBVzvDfpXWzQkplw1t9E5Ng
2ZPizXB+/SnLeN7yvhNNqpsdCr1KEIA9MqgKG446ID/MIU7mJut7bidD+pIrOtKw
6C/0WIcChyI1vAdyn4/i6oNSHb6paKDTb+lySavaXcjxdYojv8vbKqgnAlh1jDtE
P1PtV3ZorTU6co/cym+CYC7wIDg/bjatEdKxhAqx17utjrkJy7yoWPtJpG0kWyox
hN0Y/bhcdTP3DSUhYX4LNUMXPrO0rK/9WHqW503lBPhcCrYxuzsfgx6p7r0+C1vS
GlhwsRbvDZ3qs993ch7KU9b/dFsKMHGkwj+r9u/06vZc4o35uLE47O1tB4dZMrmO
eF2B1yfNu6LY9UCxCBX3Ly/Sp++Si1GJryX7i5M+WO5JqoaWcA7cO3f4pHJaUAF+
qF6Yj94U6dmfXny0p0URs2Bq/V9O6fWBBvswrtVlVZ8dWzTLkqc5s/swh4HhwvE6
93glFxJWnZT68bE2QA/zSmygtjQnRTUi16IOAvHAjI3QfhC+7gNGd4w9whnQP5G+
1FJXKako9SkzEPrUjeBJOqsDh4pBkIFYAt63i70EZE4jAjIhVen+mQj429NL/rLC
BPq7GY21d655P7S2FiNaohU2pnYAfM6E4IhJxbtrixwbUBRCLutStdYaB8R+Zbjk
xi3olB22esrQ+71YM1JRdP0mMnXy4xRxGPVF6ID34+3/Sp9Z/2CDeU+vBBaAK5QK
XH8wPBIFgoNiU+I3qFYEoglrkQ8E8x9iNZ1+gdEvYwLCjsWEDYaxg8rXcMih5hp/
zKX66xXASzs/6yBYrCZp7oE7IvjSQPNq5p0ymNxy4KNCD9L/87TFtzhf3L0vIStT
/TZ1QL+jWEO9YrjZ6IbH3L2cqTaadbSNyN5VwOaRhbmA96bJia3pQYBtGzM6DkNC
ifkFo1jB8GpEFuQVQSoaoyEctCbCt26WJeayxgpoEFwR7l47cdLOSUK+kBg95L7j
EPtdNqBZOIZZmrVCri0QduJQLMIWs0DCzLL0WJk84IgTRUoz3jFGBfGb9Q4hDco/
HDTVRvGV3MZ/OmAtAdq5MdC6iR+xPU9s+/XkqwXcooWFF4JOM5EMnqDPdj56/3ze
OYkJlaqjqnAWCrH6yRUj07Th1Qe6Od53dr3CZGxHOMFbw1fQs5R2QFSomnPDt6Jk
dtuvjkFYIpsqu9eePXmhbgq8sKb1beBGk7cftg9FWJ9oKOlaTyGOkragStwTjHuI
jFYfRa+AGGogQELub+fK+iWJxs+7x3ieTAgOKQbdo+3erjGgmEZkKc6eAPCCOqpc
asIJAvElRaKfeMrTCYiV0EdaKqtTXl8oN9WeY38FdcTMC5eaoaK56WHmqQUFG87H
nulhZpq88xt3q10mlbK3G2SHod022RIHCO3rDSWHTYxBdZQWZlvytVzTSOJFQfla
qfpiw3NtVQAMQGbLsghTwA+sFlKTy/wKwMdSxq71ZaJmxcnWkEkbx8rD5cILMAkH
eUkrh+Ifb+yDT13XiTDahnna8PLLVT8p1qkfWKTLpwwJaQDy+w82nvTV3w2fTQbx
mXnwMs9S1TenhMDaiFmbxdBrLLeblyyQgI4XGEn1U/+6+E34FFuKwz/Ntz+EALHt
sNAYOABZZPRCqwG20oVVLAJ8/kJe7tc/P9C3XdqhO2cM4EVTiPAtCntwYtge1ccl
YDFAUkF2MNFfgL4oGMndEmtvDo+Q2KWHEfBteUorAHsDC+dZlzkBIpyjJp7OP0ct
5lCtyvJxa2RDDkpJjkaGXZAzFuxB+tcbniv1qkFvs2JEQa1LQTrC9FhqI09uAfxO
Ep9wiwf2TGFobELnmAvoHWA0rSezn94ZdlN/D3PmhyEB6cK05ZShk/Tv9K9eXV+R
rgCflzkgf9FNWJlLAlTZBcFBiaYavpM5/jUU1infqn7Sa5tUok1k8E6/MfVH63KP
is/spKQE2SObK/+zA7vSkmLzpBgnydWP73Ogl4aLXYiKbYTPXRXiE+DfYm5esL+i
tyxukgzpW3RGGZb/JZkMr52/sY6708Z+F7zkPHEudqg/uUi4rpcsGaAcaemhUoDj
sZmdKeNt/iiE0LKBAih+bRuzls/EvzzHL8K1ZAupLFjZUka3/R8m8VQfcFXI1ChG
bhJ58zVBJFdz+OsiUG6A/Qm23+u0av7+QCaD3KEtpwXGT8QBTRkvAjsSRWsQoNjp
D4nAgviU5gxLCWGvtFfw3/wILCWF1c6IE14qjPD2F/cXYBHr+7aWKaYMB8JOIlBs
bRu+56zXdmnCJFxt+lyrJ+Xbypa97nNBIO1f5NwnNCXvCq3lCSBvl1IfTzXTvNo4
k5o68hiHHnwL/jVTBPKYTEXduGGm4UOJyTj03+Tvx87sfcb+ekBrOPRrqFVQR8kH
cRxlG7EAKg24idEShtMeoIyRLYyb9aCvAUzgLOX/dPPgKOWmNvyD+xoLnE/8Bme/
sLeV6eHZQmC6nLdB2+rLfgDm/L2C9qPm7QUgRbr+IHHmCCa36nCQ0bcmsyQ4Mckv
pm2L80dDdQv5V/SYrnds/DOVWngjk/H320EuH3BnoCBfK4K2NA4UtetsDPhoryEG
W9t/JVYcsmnlAb/DGiinHp/e9/ooGBHtLM0eHLgufo8RAI27nSqpTzgmhidZmaX0
2OnAwUssQySk2wSWZq1YWtcaagh6epTeL8BqXtZWG1ULUuFBZD++rhYoL3IW+2GC
o3HX0mF+QOutGgvt79PVqWuv2+8f97nijTxbka4v14EPX73IhPnUMGdyNXt2CiS3
80Zg1otKJJW0VjSNjGNIkT4hyDQ2hySupD1CFyJjkKfufQBn/ELXLbyRW6PkSlOl
ye51dIB9KTfbG7YRF5x80X4p013NhvvXFOKSYAiiK+BZu5cF32eBZWnU7p186t/d
ja4UZQZbwGgljDnDPGgWqAHJ71y1+3kkK4FOEWyTU/aEAxwepN59sQMPL9d7hE6L
58SKQCFqTvOyPpLwUaDaG/elCepNS2c2LaIdiEx7QMvnBdTeDWcZDbT8+hJ/nvbo
aeJgjjHJmr+s/J8+BktyCQg3RLCk8QKvGGgT+SFEAqrHh4X7YfuNDalD5vf4qyrb
66OGfzDx43JjjRaRHulmEk/v6kWeyp9wO7BXV+P75Bg9aTUEugxjb//ukbi0+N8x
0W0ibpAFLfK2knTKLGBJSFe5DlL6yQ6I8f76Zmf6ZlJe37f6OHIv38Kh290j/kbb
vwUQ2wVPOtSpVNRMm961cknUQksYee3uti6yJJpKZaZuj72b4L/SwMVst2wsBG2L
5YP1tBUc4oMClN9itqeaqvr/MZY++2wuv2l9IAgCXd/U0gctRKSdfBiCKDwP1tAn
EY4onMFkZm0x1Dpmzh94xi/iwXkAk2kCRMOLHlF77bj+i+d7TdQdCR3gONUpNuR6
0vGip4HSpiVWxikfWpNSMZd7boVW7SHs14ouRubEKZMhZyoxFKFr+aUvQq1jk3FW
kWSjJ8xKyNvHiTGCPcoDbqSycpU2GzanPfPE+0pdrbVVH+lfXCg6GbTzFzPn8bCR
HUPhPSmDjte7DRvxf95I2K3fcLVlULocg/7lOtTmpr88Z33ue4Ny3u2fscP///xo
61ldSHLgmLXf/96hdnvQpdJoNn1MaufEYPkyIZkvuEUk5gPRJRg4gI4T/Kisx5NP
aAIkOxp+zCo7jwF9GMT0XHzMGNHV1z6TzF0w+I9isnL2NBBCRfrkWF2ocBtUwli4
dg2ffSDiFsDgjjA+wzLwT9zdSxnQdFkVgtPaoTDVugeduvBcIInGSu8v8s4a/Ga5
tTY60X5n4PR54mfQtCBCFK1RRHnO3s7gSKrMzHUjc0SvQvV68sD2oL3MJeVkXkDu
Uwa/IWUVcEifvnqv2S60XwblrjXlHIQ0AcX2CquLyQCmecg53rFq5qcuNh6F9BA3
LNuIvhYkMau2t9RP5gBw9pviKpdS3nKfbQj6ckkXQKikB/mPT5+xs6WAijvjPiYv
IT+DQxdr5Xv4f523aDweOfNiW+d+KIoWwNp85Q2e2fhRacOpjSlEVBnyWtDSVquM
EaqDRG/JTxOvplHkYkviLBLOBJA8UaEVrsA9mcFKz5HiUNjX87USP7gZ1uUyn5my
WZxuH4WxcONt7CjeBzvYZlQbBH8t5ulR/g3RKLSwfNdtPS07uZZEJGci2OvyUqni
SGNyB8ecVMYYCINxmwGwn7FWDocrZj0NdXvmUfOXFS88QMBMyik2g2wxrqAL65cN
VrE9aO9DU823IywlLzVmWReUvLx2Pntq6QnTrIKSnEExVFFYZDhNe6UeqixN2Xes
3s3y+MPdyRMlcsguJE0q4GMY1bn69xGZpDviHGY7zpZ0PFJxdtPUZ/nieVJv++He
7Y1zSFF9M2nIMWKJNJQJ/lAQMp4hThCxiBag7bDGKp3TcdkVpWTnDUKcis95gtkQ
ZAbqfDwIJn2qFdGPz97C63Mp1QhJiGhOodAWxWrIOkehKYDQSqrcOalE++Bcigxk
kNgWRn7yb8EyyP8EoAUs981hTqr2F9v7tmqBriJlkNG8s5ELneBmVo/t5bTuo+so
obntxWX4443CafpuIgWc81USF6/LUBC3RxXcPqOXBbSBHYH9XXudfRe/S4B6pGDR
pusKdUESwuvGaPcUEjtBdYFwg7F9ePDH3Gv/+zyn7+I0v0ZXm7jzpEC/a2qdnkAt
3G9ynRME6WRg8/EInOV5qwLCKmVSPvMA5/5UFUgxjoVgIo9dy38UFPgyRZLVSn9w
3El01bxVcnpBI3i6nqTS0x8MiQxGUeZeTF/kSRNEY2JvGobP+IrMoQy7rE4xmO4G
Zt4nEFNo4nqOyl4I/HZOcy+2NbDp45ia8TVMIUkd3k602kVPYVM66HQjfqaRHwNF
d+u4eFbNwP49rYqFYFk2AiXnlMEVkUs0myQeLrBh1qVZ3SK25QgHI/BeBcbeyugG
9zjESGoXVtpP5Z0dMrTm+A==
`protect END_PROTECTED