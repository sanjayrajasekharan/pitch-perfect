-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
kDSKBI2/2XO5mzvKVBzuyeZBKw2aSeCcFNEqIQLcrKs3I41I0GG4watUqoIF6LcZ
Qp11L7shy+5Lze5+JPqD1yTUzvicQ+QWUW9tWDiK6X6r6tqmH7LUp8NIe2U8IMbp
4QkRYwJsewd+2kU59vLSIDQhtUOkSl1XKSZbFtHR9WL4Ib/1Z1VmTQ==
--pragma protect end_key_block
--pragma protect digest_block
MzwNwZk5ROAp3xKi6agkP9p9S2k=
--pragma protect end_digest_block
--pragma protect data_block
7R5BSd17GEJAYgWqW/+tuWCo3HlSxgTmCvH8+lbbeEL2PMZ6/6vdGKArQZa8MB43
HpWX8m0C4NKh7mt2Keedja5TsNx/N9BdFmfMYPm5nf7zWZrbXxSD/3lqW8/eKO+D
KfwANewzrshQeAdRZoxH/4RtHNpMPIpQbJ4GDvpdPjwkAV65WEFdvwKL7HuadRXU
KIEULmkSdadmRxNmlU2y96/lihtyUboXSk3BFcOHJWp8i12SXA0ZGPYDxCiN8KqC
ZLgsgxthI1px9+b1QRI9Jebrs2NeDloLoF9d9iog2hokGVajLjzWNPEWi5xmcgD/
Jw6VP+l3TqD+fFwQnC8cX/C/L4iUSDbEZxK/+gHiEt0Tgm81bfKnZEjzK3nmZCLL
eecCx6RFD3lYAn/Utr11Mi9q1wJF1xukt6P7GYmjhSi7gcQT8uYUaG7OUkuZOior
xauI7EMsWjPPR67koFTTmb+oww0iuoeS0u8bwoN55/RTHRV59zUp/d3oLsq1gU23
dJ1RUC+3niSeaHRjoflS+uoHpyIXXRbCg9uz3MmRJ04K7702JbExfq/JNLcIYdRe
0MZwMM/yIj3nN3rrWIiOYmIt13i9odTCnLPtPzG4oiPWs50yYdf61LnaTxp4NMjO
Zj2oiaAoFHM/+tpAklDONcmgoLvOO1nLhH0SWw4ia8NPGgTMVcJxnucZOi5Y9twS
OaP0Tsig62FKds4RbHs6sqEBq2Eahy5Ymzaz66c1SFFGoXnz9EIUhwJWh4+TzcB3
GUuvawU/qzx59pWrk99SEDC37/FRr5F0ebLRcOs8vBGE050nCUkIsCr9/lBfXuZJ
wk/FIBANRipwJDUm/Dkj++6x7l/qP0tjZvORUl3WBTOyHw1WsPCV8uJLB6Uhm++v
N2P75n7AdWmEPShodMGkC4GmL0Kzu+zvXhphnkMwNkJWhTZBzfYQ0LwY5cW0Rcxq
SukSYlYI43x5nAcdZOyXWhnt+07icXZPwRdNDjP0Wj61qDL9PVPqwoUidGkqM65M
eCd5k/JDbz5qHhJE+ttWlAawWNcIUFPbF+HkMy1b/uB18sxO395kK0gSfh+TtxpN
YrZRkM9i+9MHfaYM5d/rmHH5SFr0IA596qtbQ6NgEKN6WZhWHIUWCURlbKIQ2KmP
TxluBkvm4CFUV0VbksppUBm0aepWJHqJpbUWJlGastq94hLDwHWjUU1Di+WQSO0D
ffqK3p1ylcyNmwUSS7wvudj51kgufk9+Y4ULfHWzqApzIpN/2gQU/gGFzqgELnCq
f0xTQxPcnrSnu4eXGdADzsS/h6MDdTtowqKQDZfuzOBsRJ+XKtvYLw8ANZFMCjVe
doOxS7lMLXVgYHPbxTAJsBuFPH66RjtREBywHEXbWdsD6+j00gvO2EeTdgox/B7p
+keqlO2ABCtVUhQP0WHThhy+55J1++WYLirX0RQ+dF5iGoSh8QeFojSNkpSk1rLN
LPLbA4/LwVlM16ZwioVTcf4HVrg80DifHkKlE1w3g5ZmWQusI5s4OwMLb+j5YXRP
80dUHLc9ROny1KUxDMKrUU+j2th5vBHvqxu8L3YaK4Nen1kp384Qx6x9CvwVg6Rh
rbf6HnK4o3e9LbSdRRuvmzRTf4tfdfh7SvvnQqHgQkgEISPE7iS6eJx5cTFcguJH
C6ISrnDBtcrPn+uyulGMpFTYeUqhneUEaXNMCf8LdP9J/FNhmXkZAYLefAN2TqNt
pmcGBPDqzICGc0mueftvg0+NnJCpgfxEbfT4DG+ZFK9VxrTstzME832muvyk0voc
P8j3rkV8uKkMWzqiz9jSVR663X1yG7zyl7FWNoC9Lnzxnqc+KpI60A48NHBeea7O
zm5RI86nrep07z3UyRDA9vcHhkAhrTRGS9VO3LLiKjgHYyndBe5nyzdtRqetOf3D
wcco9EckU9jmygyBQf6TXFjKHcbUf1xl9ofYfRERDi7pXOHyqbmGK1MGWrQ9quYN
E5pg3tnZwC1+1atIJlFXyiKpUDX5u4XivwI9KW9s7vGWp30u/ZlBA5iewfRgb+kF
YrrCnjKYhjzXOoN6qMc6MjUNPvsRi+2MyzMf7sUisDzdWnJI0Wxh6zk75ycqAz0u
zcw24/toJPJL3U5w54bZ1IaW9dfbEajhc5UMhjuxO+b4PGOt0Jifs9Pq2glSlple
S3JwsZg1gxk6yNg7kb3fwlzI+HThZdIxxqt3OsVfDqPXTES0sce9WgxqjfqJytkf
w7dBiy3KcyUZr6QYOMSwaRy0dNMYKbJLH4UtiZAGxVNCDiQsna9SJo1zj1Lmmt1g
UcYGAhSslXBkf4z5FdZa/QHzCyTKedV5t6C3AbEJafHED8ejkk1k0Vm0OcIODW0k
yMrIhuqLHWiuZs0jb08GtTv72Tw54uHNn/Z7N+l/puiydw6j5EChub9gbiMMNHLF
7ZC+Il332xSHyYt2KGlQYzQoBkwlGeWD/lhao6Jcn2GQEOPHeRCGg8DuH1Xwh6Fw
27Srf6MLAxCD3/daH8gHoUPppMAZ1/VFtE2KmkeryCqfrTfxucuqz/hap2GbS6CS
EttznNIwfKQuTB3tUnwqgBkty3K+pjSWCBWDSnvNKi/k8wgNmpZqpWPjusXuXN2C
K8NJAc3q082mcJ5H5RtxNb+Udio+eMNw4UQm1QLmtedpG7EL/7jobAwlLX7npZnd
RAs7N9s2prfvyUAhUytaDe0wr5sgmZHDBCUfq7GIRE3rXQ0i6qSQs6BwhR+b5SP/
c2u5aEfgkHuTC42XdM4XtvrMpag7j3stosvoFlm67xeUMJ/iXCfTPvQ96PDgtC/5
QE/su0svYPMj6Y7mdEG4DT03kghKzxLZACrZe9z6V43b8MsLwj05KkY4TJJ842Q4
mb2F62aSTH+jZorF9L/gH/CEjyZyxh8BSD2lHfnfaVIpu4BHYEEkNmxHl/cPqY3j
HOjYB0c7An8Nc46/lzlFNkjPsS/9wLDZZ9bDqodL6sDASO3Sv8TeAKqW8jsadeYN
SrnnFc7KAyG0L62TXiaGyQE8oHLoebfDX8HafnqOLV3bNKA+//nMlX12JCUrhnm8
8QBT/DCKUPSKwTlcFhTVFMnyLxQo/cfrMX4Mtqx26xnvO6bpeBuO1TdiyiUcs2Ug
W57HLPomgW1nTU3G8B8iM2ikvs51ecRC4kljkyoxIVRYzcIy3ci9r7+M/s3PNf+x
zTDJTQ6tMZZtaoLQRu/WuovMyEzcNZFRrOS1pYqxT49auxqGf3O6G0iCezTB9mbj
VYSoia7NYXHh7Atbpw33qne70dfUd9zxPcfsmA6rwRPNiyWnO+sjiXl1TzRBqm/w
/pS6Rr/f49D3YQJQD8SSNgnAswR9YYhs5I7QY8KT1/p2OKaflpRz216cn+DiRX65
/p4T1hTh8J61m4DyVp4dhTcf5l72u82dudQ08Ke8Xj+8L8NoXltyKwm0vDgHAGGA
QfS7k56WxlYnegKgCA72o+etInWfkfCodZ2sLAImxeXr5eJYM5u3epdkTx64lVKw
Q9zx4swtmjrG3+5mboBDHqM1MN6Qm3tk0PwUwZSSo5TQnb83gTBGt9A63jqliqOc
7H6DpVtxKa1HQ4xyCik+3vGaL0727HtNNKwJDXmFZI+EFcgaY/elAXMH7EBrgjwr
751RFxXlKou86t6idZbGL9VmLXyDL6C7AgT6ojMvO2b+Ub3QDpSGuUC6XCXNvSd5
44lzYDzt9IL9NpxctMPEweEZC+uXxtZiDMSVvZC/Kj1gAKmPKdodMnFqEg8raPSu
ZT27dedLLhXabwW2pISQzkfnZrn2zEdALwZweEG/3ih+l/BiQmaLLmH3docL/Ef/
aXWDya5awV3N/bx47wkMoHQzt62+qj9FgjeJBTNFPuSqpEO9X0Q71m9wFYN5LXCt
5fg89X6xAOFGX74aGdZ+6YIKADK9ovBCS4WWrSIuNZY4u9rF3LljgUwpXqREtYV5
aCPilq0qLj1yaLvUe9mEA3Z4lFcpWfYpKF1wb0ZnsoundnX7TZbtd/NZuadqnsmX
OY96aU+dInftAoiM+Os85dekXEGTp8T/lqoICJeDpHbK54wNpIOwHcboXJBS2n7z
f3tB0ARgTRGS/vwGosEUgjWKnm37dRxXUP5e3YslKI6G2Y8mpFqNuHwsHf6W00Yp
sDf83XBxXMnGFXNupnnZ8AaTZZBtrRG3Rn/snS8VKZvl8sUFcluBiA4PaN0yCZwj
uUt2/zuZLplGbmtRnRS0SHMwfpMWNyhkauHbGAmHaJQc5i0F5LMFp9rzGj/1FH6g
TjVV2df3GUG5+JQvhb7DcE+AID7acH+CZc1vKaSUFLWKZa/TLxqK39F8z58ZFzmI
pfakW/6hke6EVDv1rgwFH5lKXhKHOnlZOM2OCli1FV7nJykySuynxynO2Kuf5TGH
I7hH/TvfZoFJ+L8wW1fg83e5IQ+eGmmVNQlAf1wZgNUDvxHl8stJyKquwo7FR+vm
nownnl0XnlAGq7PsnF3k33+qZWd3IgzaTeTKQNSLe9+iHIgvemKiw9C6nDY2qsQ6
jHu3b83xREuZOTyValV/CHaIfnK6awQS8Gh0UaL4rLndWTp9LIaf7+yFiQTreW4C
rLjSZ56kS59+mwPArdMrzennvvSV1Q9R5J51tG/dA4YGc/jKeK4ALEiR1D1VFyjT
i3dGrLqGobuTlPA5TkcgjsZYfzLJ9INLNeulaljg1h3zshns02zbLTuSL+gjma2b
3idXoCvXYbVh2NDP5XHL0cur0Qg/hCsQdEooxNN2Obzvazle7Xp0yHbB6o8Z4UFI
gnv0RnjBXXMxeMR9YnMcmcFCPS8jfD2kee2g8kzD7Ly/SemBc4qjtTAvi2FX3tdi
Ael9Vn9i6v6I9a1chs/95izNrOTnJrdAo00Jt7trZXePYa4tzV6b1dxakEiyv7wB
SEw+4YBu+ADaHq+ArTGZHPh8WMD1UZL1KbsG2WMnXQ+azosMDOFi+e+qO+2jc78I
FQYnfMP64XXavszARYjSfulJ95M/UvovO+KFsLCJf6qvXIzNSlxru1EhbnNVpwbO
/lRh1knC6QP6jIcpqLLSNAd1QB41tB+CyXC7IZsHKtcsd1DhP+FkKIrrZ8VF5Tmd
n2pfCOVAhLcc/rleCmsPZUaGf41SGQ850hEZ9vRAmHfTugXjcLoeAHrOD4uOys9O
e0EbSVf/H5SCcGVuOmDwgPP2ND7Uxr4s+aE793A05Xww2dR0Oi2vLKwsQ6GGS7NG
VLAGj27YW4P6Yo40VgL2sgzH9Pgla27VqtmHSBEpfY4wLnED+ch802xtuuDix/xH
cSabksmNkzx9NMfUiah06ONoETecTTWqzS9V6ZSYzhhmlWJofj/OY8aBVMNB+WqH
v+TklOERHJMg9tFUkinUtHZ5jqr6+VVzrnAGIpDHIKQUUbWLGieLYOXmGY1laEvu
fsOnftjW366n4PuI2maGayBmrmWIm8SFzV/GR0CqYz84VB5sMwZqARSl8Bee9xsY
f852ity0ptdD7W3em9oKtD6DFRx8PicmPVs3aRfBuMkZt2X17+lZGhPeJU2d7Hi8
EIR2LXEI3sZEpQrLdr5OkPyQyIl45Wdg5alo8lVrCqy6jmQtty0ZCLFitR1X4PEw
iWa5EusNJndRuLY978P9hQixNxwy2PSlnmsaqdJmJqpy5YFGhX5q6Vt/j3uFsIeD
wDlb1KBGWKX4hPqzRiWq7S0XjRVdXjbiMxahicoZRl0z1bOJQqaypNUmVHMVC+QD
d+h3BpNUP48BLoWj49U+jH8T1NIu/OAdrDgMbZDEygNDNoPGeXtKmaL/mWaXoRI3
cM+NUyOLm8Jjfgx6hHLoGBKooHlkMtl59hGunhYZdzrC/vuDiVoILH9u/2tTSH31
wpnoj8igudN4IgCunWT+Goqdux71Whz8Af6xi9EtmK6suTcjJRVEJU6SNixKoEdf
JAAynaQgGQaoIieiaTLg0MT7GHundlS17/G7d3Bs/OzSWKuSSHQi18SfWlMjauj6
QwaamdPK9PcaUU1BcR2OrBFVLTMItfeVnt1UI4ZViaABqjq3E+t8CYK5P9zDl6gx
dXIBJpVAh5Tv1Y+niFH3O+vY1ko3rKzRQB3utRB2uCtib1I2Suq87focL9Tkq6Xk
zXjeJwIJE6wFpJxtO59DOEsbMXE8WFoq8be0i8arjxsowGmI4pOMiT8JzInLXaMI
mtQnqH5ymGWRzQNj6pNMd2R/fhhBQoSUF9vsJW3PKojeU0cJMGhtzn7CttlwihWC
dfYpLcR/oOqs2sOXYC6SonZ/CN5meCDEWhQqEvzfvoNstciEjc2vGsu03Q0pLLap
0vT/uAnuJ1874ftDLPyQFX+a0huPPtdOOHza92BIRIDHscsa1NMdqryMn9JyY3vU
F9PdpFxbEDJYiIUR5/gVOQbtxGMhL0qsKLCSHgyr3B7szdVSEOUPKxIzoH8o9wZj
pQmZe5M0H/hZLrA8y6BV+hg+BLNOz9DR9AprHxUBax5kF/OC4KziDmeXr2b/hvOT
q6vp9poecDKigzRQe11fLcaT9w9VuekwuU7VkTc+59NojEGoaEbvvAaSkb6HbwRD
IveB24xcQHz08IQpCmMVtP52nVLwaw4zb6vOWeVUlFTqS5sLXd6xzizBpfe3LqX6
O5JwxSbeXNBmRMbBU6kU68avFsvcHwmA64GALV+PVKqThPAiv/P7C9V25X80Uw0H
AZB0gjneiUFPTyBfFgE3dldfbCxZvEwKgHaZ1wseNmqWs9dJpkNs5E7dPZi63g8F
k80FF378RaV9vl2cusu7mT7qhPodDS0HZmbNIUO4cZ2UUIE3A6VxLu8bL5nmVNb6
bTlCk8UpIwTSs2u5cR1Qg1PtLvz431Ahh4uTLu2GCbEsfSnzCaeOB2pAMSBX2kDy
DJuNKYHnqkXui9HiKiedUQi7+uItdwXyRdDqwNl6ffbMc3TvXHisaMLdob1CNEWS
GJVTvAuhdE9qE8R9xDOYRQk03X4CSscRvs8ae+XmNrQoX1IrZaU+Q/yXqA89KUP1
S32Iv+xnNi0VS3w/6NrLwMxdpHqy/aoIz3dNHf1oyZe/mo//8QwOu9qv50YzkPM3
q1ECAToo4mzMXlQ4LnQKRMgeVtVOCj309AlZUNMS9UVmOVx3bd4/5IOBws5QIFP2
aQdGIc3lp3Eb5hCDdpO9Zr5t0IQ3Xl8cZJYfG3RCkqSEZev3D+QhI+Hyl5/ki4Xx
2eok+FhVIzh+RXcUCIObUmgVRcN72wH4FuNkzhUYhkCSIWTRGCmXCSCsk7jB6hTL
JJAs7a5H3CanVV7iymECdY8yOn6WAkKX9rf8I+5AoTS7HQlO3M0JL6mOcH3v2g6G
PPiil1YXKHdDXzi8V7l6b43iJwKfQ270sm7T1Ytmvo7rGcZ5Jw7ZoqkExn92wc20
C+krD/7qQE6jl6tsvu+p0xSOXVv+SZX4Um/ZF0WyA02jPgAdj54uJFRnCuHZgzLT
urtlVhJ0zhdg3nUh3FlidfDOQfH+/rFQC1JVH5vx6dLCcDyEKtpfS2Naan4FvOWJ
i3Gpf+jM1LfW6JSZzmb9zynXoWxxcXd+sjCNfLjAwLvUSp5gYbsJWCMPborrUS/R
LT/roMntdi99n6HgS3qim5wt0d7jPsjzpI6IIpfDqS78Jw1semV3ZR/iDDnHOf94
WoTOuS3t0xvHXhnI2yBseh1eV6LbTcP4jNokuhE5OxbJd2L434OqQLChwqeXqTtj
nCSTakgr1XVwYokjQrWqXZjA/t46oyIajFAttKW88ZvhWd2ieMEjgSgV8+3sj5M7
VFo9S8Z610ryG0cb1m7qIp3ppYlY/k3NCA5voFExcnV5a+ZbJ1Pe+Z60qU/Dan1K
1lOpljOZLgdD3kSvoiC3941QwzQMEMBBm6QebW2RfqvFsVVEwzdiXDMhZsAushgV
cmU9q1F2waD/OBJRzACgdX7D1BnN2k8aUps3a/Y42K0gAew5Y8qdfB59ecmb6qW0
ODUEOUzMpkflkx2CY9kZzajOP+B9a8JcuZgxqkdJrOJDsQJs4E4j4kfyLbogT2Yu
1G5x9zaE+rhggVYzu6iXJeSG7dxIVUw7e6I6mUXZocqcQOrFLZRTYutyZgFnVbTP
oZFKddi9MmJezKIVrreOWDIW+vR5LQwAIBGoyZkh3b52obx3Y0PcKHK5Hx47FUv+
KdttpAFKK/YEY8H9pZW7V26X+qqgH35Hgfa1mKLIbsi1e6UHnrA+D8I/8NJk5wFx
C+J/vUcMvcK5FxhSwOM1YfUxtH4qB4hNmeYyu/zDb7XXNhBmpQmofHHQnHljTPzy
xaABhqQ5hWuWYezlp7iHbSrPUb+Hm1dja/Y2UDGasB5a8q+WhYF7CNPUbWdoKF6w
GCXpwS3GARebqrzwfscx7XsH6IAUTgo0PNhfI23QWN9zlKUSEQUofXCXBG907AYp
iL5nx+5HYSTZWWAjPBNFuy9ilENuX/vUZoM9NcdDIXgQZ9huZEPmvIn2Oi7Jj/qF
6xYwGcg+7e4JInRGj/BsNQOI41f3S0Tjnvs3YlCICe4A0o8tSC0vbUou4cYLPURj
BA2bVRRuvYw2UoPoYHOQGzJae40oTz7u4LQZ+6sHZDNvXw4QHtb3bDLaNVMJe7Cq
95qVcCAFEH9Qv2r4C1AATwcrcDKvClTtw17+wK0yE/15dZnMgAE0190BXgHEUJ+p
3CtCxvvnXI7rWnq1tQ6+ZaAo+KyC8FF7SsP+5kkTQXiOoXLGTWmB/4VevUKMSB2I
xg6MbNgWUTnUB/4KwUhK9GX1csnBk61bWs5Zgo1bBsE+b5aINOx7bESVT3EJMlLc
4vdWnbEUNTMYZ8bkniA2cMS1ca3MPX7hUgRXgvkerZuRzHc1oHlybpcCk5WM1ZC/
bY6jvvwRPvdJ9akTOAZYMudawKpFQCx+iMi/MQfOYuQP5V018jOHY4aSpZP/2teX
r2wtpNAa1rXOquAkGrQehxQMdAgEDG4IDrRABaR4xI7TU/tQUFUWUVbUKSteZ/e3
QaSiHGVE1h/tEQY9cXg/sQwcHM53t93ohWmaNIUQ2xThoV6xwIDQGzjVGN2D63cC
t4lyMRO8/p5g8kDXrOYvM3B4dDAQ7UCJEcnhj69Un2iZPnqf5z38UOz0QXEVryS1
s6gF918QLlI4Anq761bm1M2vpMho6+jTOoQKgAioO0Sb0gs1iELQkRAK3wNu4Cf+
5HmFXQ7oKgNjDGIT2B2N2ynMcHmwJPSJ1Qk+xqPqXN+sSK6tQsv8IblW51rvqmOF
Gr53hZ4uUbG1fEBK+scpSfk1+S2k1QxAImiwq6kBFb0OfIeyqpy74JOnXuzKv5Ha
xO+vbeUT0wXjAGGRM8Ihcx+YbWOugDvuz+S4E2ehd6GVmJ2JQYRuFvW1jza0J2Cm
u26I3ElrfQmFMP8224Rc/O8sz6JbXDsOS1aA9IXNRphxcDdVzdXGPFxIYuocXdnS
bNNuk4Z9QBBiCJojVRcqvlLffjpFkvbhZzcOZSqy4xcNpNAbpg6Ywg+xenyQyE9s
5ri/k6YKMzCP6udaZhuvdpFIh50tSTkuayRVg4xIq5doZCmWwPHjtnyDdBKUVvfv
Aaqdo3ClfbvBYMbyq0UMGVzR4uihRPHOgrwEWU1kvxpzy/nPboF2cAyXSBXf8RXg
kkbOT4R2aTR0QOMSZ0O3NukSRXz+cKYW6/5I+04Ne6lAZErlrEnLHR1+gr2eH+OX
srINS4iv6rXojLvnDG6LXRgZtmbCe91Wuu1wp8xNUED5drDJ1ZPoibOEwd/qjGll
xdXc5abFw+l+gqBTou9hz5oTQ6yXmcfykMtGCKFDBGHAe+MkzbdkvO3+FYj1eWvp
29VEbsQ/3avpPI1+a9fFN2UGy2uRTfWNHiQ+veiux0gcLpV6p0MDC1w9ovyWhN68
MIwgUKOrg3ao7x39WWmHoHsYqF0yPorkyphrT8tjLTJWc1BZ9fIkUUaZK6wQ4wsP
0qRni7c3c8+5InbolZaxlghpKqcVMAZYYEBpEu77WkWtfuJHgQq9vTgY9hycCKV0
UmWHjPaenq8VeZpG0imJXlnIt9eYL371O0s8DC2dKRbOx/RW8VlSFcF2bVoJvo14
kb+q6qfpbxm2ieUGUn5RGfsA81pfwb21EGfhiD7UHMaXfgEsig+AZ0TOQ7IQf/la
OqthqnYkLKCnMcMZUozPSaCcEr/c+Cf6XbM3gPtPbTdL6B/me5DRo08s2T5RZwTN
lzXWP9A4gCFKbKok7f/6/+wLpbGYwcIJlGCRoKGu1dANdqtmMoRG/Zp2/X+wa67d
MbW2S5Z2zzfi5YCrw/WPS9CZGhj/YEfMzOexGSj1o/OtuZcvFZ3bsOhzcDyJ6T0x
L7nCsaTcN4wmfDRY9flmjuDp6rzL3E62ILrNrSwLIDPsisx+j56E87rCYsLpk/cL
8AZ4pK/ibQR92TwyIFzNkqOXMtVDqXGc4jGNbrFhuytlWp/n2QCoAozu3t+cXD+r
n0W5oeoglultTe5OvEqGK9OX9CZkrUrCBxduVZdna6p735ySRsgRG0Gko0yQhHw6
iOQ+77b8tJ4M0+CtGlPmBYrWaorOvY5C3pNU4DrbiVt4MBXiHMU+BcbeUntDvub0
OcD5e5qKoOZ/aDEVswfc0HUZs5gE3Pztq7gDksuiQLy64k+zrogNCCuL0/UcTPeU
Y0qnUBfNOuID70teEPhqurNJDm9DMm75hRHzZ+x2uUGRAUR+jhmn7fV8HnsGrl39
V6AXrVWuLw8IdWC3+KEtQ/UJQgdBgCpL7Wr5ZMLnWbCbzs7yO0Axj8ltShcXfUcr
eLuEKdb0DMsyqbcgpnogPKtw/tsG03J1eXHRTjnfxtzNRrgKgVWfrnOM3OiYmXtW
e70KnXfWKuBv5LcpK+7MwgXdI2FaEtvDmKCcFKVUuRb6/57eb93XjkBcrgA/rNvu
SN9g8yWryvBBT3RWx/ay5RWfjxedC4p/4Q095qPTgilVsBhvCydYYzZbpazhJY7W
V166xixCxcJ+zlcBNS1C7JbX5twQD1RzApK4E12R4PwlR5R9Mr+TqcVMOm7c51u0
dsGPKCsivvqYINuB2cEkjrV9Rsh+GpyPtbAJQW5YOFoyi+6dYgvYVs0LZpWumex4
NmnFxA/Y1fk6WA0lMdeW9NQazuPKxPK0Uagjqcy6yeWCv2dtMV1ZGYED7nyUy3eV
MJX8Qna1QZYT+HhUdZ5sRcrrToSqtkJwCq55IeoHLSm42aqG1Y5c2eY+kKVZwSyc
U0wFSRf1s3oKRBrmX0O7GZWoOIYRIfmv9KPtuxFqszpie0Xi17Rcoe9CkL9Qcwcg
oCxwa7rU79Vxd9BdinPmgf7kLEvoWpO4YwZNwxMcVOdlAARTeldci4+VOpuR4Tbe
C/r7d6Nq6+7ZwygUt+WkL+Rio2ID6auJ7IvR3viJ+Ch9khYkNpl2Jd4n8mvOHRSR
VZNld1FqPT3np/Kpu900bbRZc46W7Fr1F/w9IWwGDIKyXG22MX7ZqaKqk7X1Xcra
tDTTmXhn1hhNJeY4y3VPRJ23yESmz/X3Macn/kuNKjiSOnonYNNUGaUxnbAjh/E6
osCKuHGvA6hovGXE3l9IXTV2IlhV+zMtEmpsHkaiqbvmNLF+l42SFfGIIhRijdE+
3X4eOY11G5hRIWOcS7eM6VnfIeCXhfV7Xpz1zaxE7wOpSirnoz0FbMHwoC+5j8aN
Cumt+N9UquBd35TvK8pNZ9uolgzSbZVx9W9xgmq35rG2Qwm6eecCmOeOA7X5VZ4C
b94EyrGG2E2FGc+uKFeQ94L2ecVE4KlQ2FF00Jwcvge+DqfhAoEUlwHivPaU8xHy
NfCVpq6YYksZ0lGpTroIPoygfADhpgxY6Ht0CM2geOu2aMmaw7gO4BQxBNdPgYlz
dsoS7wHimyaPvSDnm3AvGuCQtXr9bvUN2avG4/+wvv+V3y5dY3M3U5x7KcQdiNZD
dRoPiN1doSmpKWyRAEkz0ymCaQUQnK76rA4TVGkEi5YhqOtDKh4NJwTSfBEH89SY
SJYrEMTDFfvwu+LtVmXORNu/3byRVDGeIP84wrijd7mHV2mRwAkmpOnGOxef1JmY
WAAf3uylHICuJUL5UimpK29bAiUQEIr/BRsHoJm7XnVgLbDJiRNm4DK+I78Pf3nU
anUw6ufcg+RsqKWlhtj9RYBbvqFqa8mNTFozj4LiCUquE43fIYR1PQB8HECIEgBn
4RdV/fQXH6+gAzrNXqRyCzhGnYfeKN+ed1OUmorFfgzTrI6kNZe2ejhhSq1fITI5
Ak1bdnqF7c2+Gj05wMu5yCs9py41MkKQXlwesyBOvSelIn8jluQinZv8/Xmjiepd
n9BMbWbSPYpzYcwbeV/OWIQmCO8cNZdDenkurxGt6WUBo4wG/3SOrWgmcJ6mNyh/
17loFmTS+bocxIv8v9w7brmltZAPGyws6IaLUnUiyzrpQK8vRlDr8kGRlxmVE2w2
pHPB7Do9yadlZBC3ow8PowAIXOA7O/1mHsp421czUjxCgfwJuc4ovgt2AYbDK6LW
SKDDZAo5FQUCgLGOQ7eLoAArocbV5S8U/NIt0yHa+XhOEGaLr/8V8EtzrjzmraJt
u42prsloPBSJQnHS9O5upgYdPVv89TtHTPBxgTp3lSxpv7y5bT/mzqnX+/fUcy6D
lEyRNOG5x9F95mhW18sC3tsGWt6j+PAL9jj1sHFJVYe8h1hw1V3frodSgKKNok21
Xe2dVlJyO6UmbKOQa7lltMoPWR1c6i6SnFEwQxp6yEjUXXXoelgY+WHGX2CzBHAV
lXgdFheie2oOboUKrAcuZEZqT9W2Plaz0E29WI+674QJcxY7PeE9PyR1R/uHCUhW
WN0HmizoPfLOBmlgA1xkQ1S0nGCX5/5TCNuW3HSiHlQ=
--pragma protect end_data_block
--pragma protect digest_block
QBmX/TaSeRWXt+gTuuWsG/THCfI=
--pragma protect end_digest_block
--pragma protect end_protected
