��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@��D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE����.]�����[�J	��o��)�	�V,�Ñ���+��3�Q��D�ʍJ^�"�q��F)���������Ү�'7�6�K<:�;��j�WKӉ���&�x�h��^J�4��j|mQ�p�A@����:�w����~�9�T�d_Z{؄� ��>h��g/gm>g����	q��Fu�D��,ͱ���h�R�����3ɣ�n�q߰U`MP}�ֶ�%� ���$�*l����%F����� R�J�a��t�ҢvF`A�Px �Ò�­���C�U���"�L�~�>�u��>����}��{A���������-�^�ize�}$e���	�}[BA��6Y8�8�c=�S��;q^zh"�O^E�̾��O��.B`;z>��.99Cy��
�/Û�mDALگ5�����3��hT��2`A[�����,����ʜIğO��N��@����A���!���]��8]�/M'@��P]t���~�g��5����kH��ӛ4��g�4���>�2l���VTpg*�hl����� �/��B˖�)oB���"��������!�	f�x��~Eq�!�p�B���%��<�退�5�t@��$���1�������݂N�Dq�84�<j��G����To�B~B@�A��6�,iA�a�qRÞ�
E$�,&������3���b��r�Ԣ��!Ѧ�,'�Y<���ʗ�e���葟���X�6t���1��Lɔk���4��a��Ll���Ȁ�[�__I*���8�lS�Sn�D��4�'+M�d�A�����⫑s�c:���f�l����"O˟�O���zt'Xܿ�&��Z����Xh�F������ݬ���Ɵ���r�/x�/��.F�Fi�&q�v&I�5n�-Nc�i�b�T}b$u}{`�N"����+QQ�vD�?ٓ�iOi&�EY0�F2��`@T�s{f
����&4R�O����:g�^W	��7�����28j#�Od>��,���B%>v�j�/�~��f�2����Յɣ�_��S�H��*kF[���6/h!��Q�Fe�D"�X�|ȯzl�Ϗ�ɍ��dw�������;��*�f63rsT�6�~R�+ԍ#8:����$�Ȇ�΅��K�N�=�"��_�@Բ�ݧ���E�*2�������V�g�"*��ȭ�E��!酲��s���`�-ܯu5�����9\r#|륏:.�DS�2�|�WK&�팄p�a�d>�ҋ�3�e�=�<4�3�h/�F�c9%>J�ӡĀG��%���('���u.�)*�I�\pt���+a>Ѻ)�3sA�8G=���Sg����eגՙI��۲u��(sS:R��c��F�@�ܥ�M���������_���Ҫ�Og쥌�2�gp�<:��VS��^�?7:����6h[`��vJ ����8��i�%D��QT�S��D��N�{⎳�� %��>b0z��pw!�{�E%%���Mt#�c5P&�=."������i���d��b5�E��_���ǐ}���+�[�mDU�
�E���9��E�DQ���e��N����u����4P���4
�O�� ��\sʈ�s�����FՂIy�<���	3ٵ,ʸ2ȱf�,�	�Å���&i�en"y1蹉�~���㣣���ȶ��j'�!q�K�RI�źn�~���D+�������3�	��m�MЧ�o���h���W�
����CV����VA!���9�n����`Ws��x}8H'�b8�"���Ȧ%b�&�*�����	)1� �Xz�c!%�r�����e���O��9>�w����-xH�V�d:ߪ�ȉO]�����bi�B2�F8���*j�A�i_ȳ���C�h|����Jt\u�`M�z[1ϯ��q�*���2��Z�w�ҟI��:�\� ��RhNX4�E�_��߶�a%�;�Sv���N@4�V$�1��)����.��KG(lO�o-�����BX���Of���ig~6���ήIo;7��a�E� CI��i͎Β�Nx�Oz��=5�s�hf >eB�?��0 �,���.x�\���òĜ��C�gK��x�!'���T����T��.����.�'���[5�?�F�OV����K��p��T��xS��>����|E\b��J��;����M��I���S J��4���ezD�.z�M�q��`Q��E�쪆c�$FM~Ͱ�ɐP�O��NuP-\ë�5�����}"����k����
�e�8��IV=����jb&�i�O�A�9Ny�@�+e�OX�i�)��C�еs|�?�����=�B����uj�ۄ�<��#��`��"0�
R�b�k^�$�䉄��� �8��0]�ܢ��K�Ү�uf�
C_��L��9�	�4�e�����m���;������v�M�dH�������� &����C��(���*����z�����yWC�5���Y��Gy�=J0"���8�R�C��{�f��(=d����"�������_��k.��"�ATH`6�<�EU0�Us�g����T�Ԕ-�"u�/���qu�[���S$��s��K@����.��ڊ1�K'ϨRVͼ� ✛M�/ˆ��o���|�T��É��$�P��<rH�.�v��<cKt}����0��9"�<�^v�X��R���&�'�{�Q�~�w\�#�_�).���,L����q:��D�.����v]%�ܺiX��N�i3Yl*/��/��f�`�פ��u��o��Q���Rqr��em���zVǏ{	L8�� ���[��$ch���V�
{�*�+�Ӹ��#
��sp"cX�8���b�`���VE�Y�0[�6�)��@`,����zD����Z�EBw�>��=�;�l�>{4J�_�8��>}৥�o�6�� �}��%s��o�4�0f8[��0�߈�Ra9��=,�1~��n�[��B�n�گL��~>_�	hi<b�;��g%�W�s�H'�v-�G.�F�qK��ў9��<!��Q��2a���s�9�S�n�#�G~����[�*��=g�iؑ���s��u`���29�]��[��M�(+Z�0�}�.�R
ޤ�?�e{z��U�2����}3��O�9L�T{���yo�N�GgI���
p'���H�`ҧ9�PSx�8(^G9�9ůhN��󯏥�A�b�س��) x��a��At[wt4����tu��Dz���u���eyg�E�z�k�Ռ���&�
4��$��� L��?*F����i�'��ZJ�����{8�I�4�Q�4O!�	D���E����)Uf�Ac+B�#�m�B0�B���kf�1�sK?�չz׸XRyW]5��^�m��b��%{��`�H�3��H-��(����'�p�i.���)��l�9ݗx|Pv�v�\�@����kу�߅r.L�8�	���*�Ŧ�%է�.Mfz������xl	��E�j���F�j�Y�^^��HD���[�g���R�)�BQ,Wɒ�-aiXm��`T>�s�~^�Ofd^��{&��.8
��y_�� ���tZ ��x����A�st����F���g��l�˺��5�ɘ��&2W���?�m��S���ڥ�M�<�?���0��RNR�UTv���#2�������#�ћlr�D��,�@�d0� �+(DO���0��Y=��Ŏ���wn3d�>��!�眈��.���E�{w��ǛS�7��㟋�'-�=�mz<qǤĚt�p|ƌ�AS������A�I!��#�v���z�&�V#j��ݝ
)���	���H�T'�g�A�������R./_R�oԹ��T_���!eҡ�ҲX����aܲ��P+h��!�u���>��>��P�G�wi�y"-NY R���+icL&i�� ����®+��Z�n�����j?J��$uB���'?�b�̩����D��I^�ß5���.���aՍ��Z�s&l�*jѩ�Rg�����Aq4������H��Pj����ʳx�|�n�l�B���]��/�d,�_�0F�dk'�c���vA�!�4G���5�T?Ƈc^Eӻ��mR��h�� fK��˄�\*���ѳ��uKD!����˅ڪ4%R�n����W��- /���=w��3�{��M;�U��78u��]��J��ȁ�i�V���nj.tf��>���|39<�r���s�_������
fyP@V��W�O-yxX�}S-�#.9ʰbv�z���3^��Er#og��R�[�[�ϸAb���+��!	���8^+?\�ʂ�v3�5�\�S
v4��o�"o�%o�C�	H%
zC��?;:,rh5��bv7�"�Y�P]���|�56��6U��h��s���!aqTb��L�ۉ���R�������	����c���@�\4�ld��|��bA�H�.m�n[w+�-~�e+����	}��B��2D`>�����W����avU���̚g�=�9�vOEN�9*��0
@M�Iܻ��\^����(�O��.W՚�4��ϦZc�Ɓ�C��ܗ���+�3��Kӂ�r�q���F3���q����f3�~
����vx	�K���!�WwG@�,�I�j�]����YPP�0X�R>�8�5X&�#���5��v��㈕Xi��*�o���BH�VJN�(��zt�L�l?��V��
���|]r�<Epj��;�����e,Y���%�s83�@��{5L��G�̖��(����UA6�v�������CȎ+i��Y+����
�o��m:�VK�ߌ�51��ɍb;��찞v���f�5d�����Z���W8�lw��b���M� Q. ����7Ͻ�*��j��<S�- �?��n�H��l��"a֘ߘ��Ǜ�|�Zq����w8f��Dj%��K
�{#�%x�O�Լ2�^b@�k����}>�Q�*2�x��6���)&Wg��Y�5��]��cR�f�$�1+��ͩi�ض�c��n�y9�_��d�O����m/"���Y��w�A���F�9.稓��&U�<�͠��\HW�L/�K���s`.�Y�Gث4��Q_��9�̊�o�I3�����3^�e����d�c��*���y!�m�8�ܼ}3�,�jgb�'<����5])��RXB�<h�6�y\��~4�8>�1�/���.�3G��bS����2���]�����8��M����}Z��H��ڇۼ��X�<�Ӥ��n�O!y&: ��c���	8��v���;��j��/��6�l�a���������L��g�8F_cV��u�f<�����E��Xٺ����Iϝ?� ��Tg��(�!��ivm�w.�����z(�����K�W��g"�UM�V�{ʫ�Yp�+ h4�8�f��z�%�Aa���+^�~��pF�bݭi�����T���GB]��'�����}�!o���pT�Qv���^����["��=�b�,)��$�"U����p>T)�L2��/�����ƇX5�T��J��7��|$��2~�����F[���u�wПq3�Πl~��"�*D����}7f��S�	�趯�t���p�b���I�J�d����$��(bQ\1�p5R�V89��u�r�I�⥹�ɗF�-�$�b�"��(˸�	'�5-���8�(��){����o����M�0i�(�{��l�p��}��o�P��qz���iF�P���wM��n�B}����C@{_'"fr�4[��[�ǜ���u���-�4z{�%Q�+Z�a�Q����A�M�֑i�6vi�R���mT��&�)��"^�.ZM����yP`�oW�,#X!(���#���� 0\�fY�����pa�"�F�1L�t���!�6��}��mOdխq�m��=��H�#`*�$dN"��H��̤2��)��v�
c��[���5�_@|�r�Q4 =q�G��x>l�������퀭e��_����n��'#�a�$���P�J?�P���L��(�.=������:�b���.r[�o�s*4��Y����ns'���3�@�K�.��D�;ַ=-��W�"35C_+�
�ٺ}�RŎ'@�S{|�2c�c�l;ST~�k�(���4}\1��8i�W�1�������>����OC�G3���>Y0�u���y��E3o��.AD���"F�x�ƪ��mU� �r�x��빩���w���jR»r��}b��ª�31�7�n�F_�B}DW��e*u��$J[aJ�k��ѵ�<����i&D|�A1��y���Y���_0��V��
G� M�l��'�ҵO��\��Y�b�&��N9S�v7�9��&=��K	��*��eNwa�%���
T��
�9AqI]�-&I���`u������=�����.ɧg����)._NT~�a/��hG�Y`#�)t/�橚MW���r�4�nS��^g��Ws�b�-��)s]f�sx�ng��Eʘ����<�=*&A:61Y�"�����@违Z	9��kDG!d��0��e����}�x�ء����P=�-���&�`Z�A۪
��[��릱$a���¨�+� �i�܋)�Ew�"Ae���J��B�;�|�a�+��+��h絳�'*��<��̶��iv�$al�G���HW����^Jb�V���0���x^N-�N����F:��P� bR:^1�O\��q�`\q����F����x��QӼdI�?B�%��:���� #�3 ~�f���J�GKLݒ��<�4�^�j������jk�E�/T�H��L�f~����j���ט5�!�b����:}b�Y4F�el��v��=$�y}���6׏ӫ_g��+1Ӕ�8�@�1y������1{����!�6R�q��`/���i�4s�v����l~��۞_�<�q��Z��Jœu�3B��P�m6-����rK?"V��:���f�x1	�yb���9��:��#��7=k�f�ϫ+���qI��RѨ�<w��N�xJ�46��ҳU�I�=2-i3�ys������ˁ(��\=�}�����l0��b���bz���>8�t�Lc�>��L�ǆ����+*��_���S5�j�~�W�*댃f?��x�,_������&?�eD�]k���qfW+��R�+���e��2^OyYi���h�;�_���HD=#��O��C�/ǎz/?�~\Q��5���I���w+;X�L�LG���iG4^l���Z��V���y�����o��c-Xt��zLF�-�R�-��:ӊfJ��XLF��'�3�����{�e�Qqu}��:�iw���5u\`�y��|�Y�\W��N�w�mF���*�z�(eUk�'�@v��++�%�ݧ>a��@��Lh=��'nlP��?L�q��,���u�V�a�̉6�C�y�{�������Ea6��;�a�N`5O��M3���� X�iD����A�NX���G�S���@s��R�Η7�{�`~���W p��O�A2�\�������ft@ȬK�8X�����أ��y8�D�ي;��w::sr0�WU�'rH�Q��������̆|��c��J�����&�9cs�]����ISw��`�-'�~�kMY��m��{NQ3���lI�2H��r����8�1�ؤ�^�M[D��y��ǰ��bU/��
���ߍ\�F�Hy������ʏE�,��{�/;~�:��O���*�i�����k�##�hR2��@����m�#h�Yk�+y*5��?��+1��<L�>�_�7_�{ @�84Q !����am���9C���0
ն'��w82֯�a��/��2萤@rˢ��??UuϦ�S?��,��2��Q`�=�x�ȱ�h2��=�z��䉡@���@�"	�J���:��mHB}�s�d��F�L��f���4�XŬw�2�{*�s��>��O�hz�\�%�N��+���E�	�03+9 �	(Om��K_�դO�h�R��H���f0�aq��h�ΧM5ڮ��k��J$iN��J���|\���=Xo�������I���Mi��{���S�YΦ�q������ʗ�|�ҷ�Gg��TB�:��3ٯ�"��RS;%x��uU��ݳŐX��(8���9��C�zpl^�2�/�E�C��^�+s�:����i���ws� ���'����&9"�������td���Mt��YI�[ip��w<X��4�3��B(�5y��%�ٯ�X)�o���P;����z���EAN=�tu� m�X"$'�O��N���+'"-c[��4D�nq����K0m��-�G�����h7.���-﷎�>W}���X�������e�y���K�����]��6����S��<��X�k?�����i!�W��e�r��B��Cmb`���B�Df|�J�`�c�vv%?�-FpgD8 ���ba��W[���/�W�ǯ_��e}��le�jD{BN���X:�|n��w�[W��2N�����k��ހ�;Oy�h���7�@iÜòY��d�U��
]^%����8�=�AF�ؾ��zg���f�O�Bd�>�
��3�G:��P�w���ز@�YN֮����|���{� ,ax-h-��h�Aދ�l�h�f��h��pQ�G�kg�N��0V���[G��6�qs���sVU0P��:��Qa��p	|x�a!inK:}���E�/�-�jEo�m0���a谐�}����B�9�k��B�-T��w3
��maZfYsq���x5QU�����ч�#��~�i�|�N�Z��SJy�3���Vg�XA�G���{]U�����,���4:�D��a��dE��0S����Yg�W޹��Ӓ���d�A;��0�t.~*�Զ���c�qu\!uf������is��+H����x��V�h���,��������� QLP!pQ�cw�H2qr-��
�ė�8��Y<�/��h|��Jw��A:߇'�<dzW3&��Iݯ�j�s��t���TТ9�"RmMy!;=���[�X��*�̵ᐎS��3�#(��d!n{��B�s�I�d���Z�#D���/��Wf�P� ��ٛI;ЂE��bhB�n�CB����q�ۤ=�@Fh M�q��T��'�;pg
I��m���b
|z�aBm%^���A0�+��o�L�z7�(At��i�N0Q^���`^�q�z���:���#z|:�����+�O��z1�֢�}�⤏�3��!��V#��Җey�>���0�B��G�:�,����y�
���#ƌ;���z3�Q���3^"�8�)���FlJ�1&�q_���Dg/��^��5W1�m�GGoO�e�gl�=a`Lx:���.�\H��oV�^�P����q/����8<����z6W�p��#jZ#��=�ʁ�Y�����0f�e�A>�΄�!��) �2
�������l�������U�u���Az�m������xbB��k��,��
n�K�*�S1�z"�蔻����9�ߪ%���!-���\F�+b�7���+7��yM"Uc���`�`��y@�*��7��࣑<jˋ�5���A~����"��K���W�t���LB��� �%�	\]4���Au<�o��L[e�2L�_8�DT����K� v�����{g���������7nՆ�K��#�/Q_;	�h�Y��%ʂ�'�i�k䐤��z-�V�)D����E-�(p���d��V� +�:����R2�sP���
f�B���HVt��{���b.g��lɉ�>�R�2�g[ ��{cė]
�"$��훜SڍY2dpnU8\��t��-n�p8zI�k��>>'�:�9_D�4��#���1[�E�#a�5�=��=�d,���
�u