-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
hZjuxckKbhvu1N/KV/ubVH0U0M0faaddOdo/vUoYZMTZ18BI3VFYRh4U6gWEId6O
i0NcujiNMH8hYJXDGEho3CW0UeNZWugB0JotNemPMX1+Swa4M2kCAKEkHjeuFLGw
goHnAWlye6SI4nvEG45enduiF7cSewlZUfH3wg5P7BDb9cWsZqfYxA==
--pragma protect end_key_block
--pragma protect digest_block
dK+PpNc6sAu5gZwb6OMkyQ/2TO0=
--pragma protect end_digest_block
--pragma protect data_block
LShofJ4xR3kj7BpOE3eswR3I0UJ5JffuWhvujSw98j3izexsHZDl3kL7fdgiYyF5
OKD+OG1E/KD51Owr3Tk1kVfXxYCnQmh12piV4rvqnwpdV7YIFTtgoNhtvGgfOopy
m7keGtj+P3rcARUtu2nqEBRzgRv0hc1vN4kdXe0VG/NEu0CydxrxmA4iAgkdFeXE
S4Khd3oezibteU2fDFoIMmDfrmMJ6MmuJpU+U1egDIq6uLGCoPq2hQ49ymbX1f3a
2eEkPjAom2ANbFujJ9v6ijc3k/ub3O4q1gEffrXN6adK3Sg5FQRWIsEGf9gcg8LX
6vxMw1tvkRuzqzXPTZKNyqM704mYe2Cmnk+xkF3Fkap4Ejpv0eo3hmQpLsYnDV5q
YkbYBze4QGJbEg1+I+Wf8jD9xoRQvaquka5pB+CfpFQEACNy/dJZVLAFfzQubyni
wD5TTlWQXxclwsapANk10bN1+E2c9vVwSkr20N1jb6O3oQ3OMen5/ucyiBW8gJAv
naf4yJquYKzKidVZ+F1cMO/QM5/Wkdss12jLBNwxvElQab9S8Ythz4reAg5JdMIL
SixePpCofpzpWHsV4MD4lRz7QJq8LeVC2C525tGCjs08abz4Rk5GXYfaNgrga+ge
Bl1BSsZkq5OIiW7Mg6uNci9fH53PwCghm412D8p+VLpgszWSZEq5pHJYUnoluLoj
4toWmPKf8WXS/Z+N6ZLCf4k2+GY0Z659L2nVdamN6YAboNbmFJV2y8NnMzmzp1BP
RvV2OA8HQCxkYJncM9JWiGpLhKiU0frK3RZT1nm3SyniRMx07YwyYFVgyCjqTG/0
/LdFx4vVdUXiFLD/2LQDX+N6pNJ5bzOoCEJlMYIyOMqdGSbO16NoksFfHUMhmIu0
LpmXAtvAzlzS/1L5uIQRNrVdKfG1VxBbYG+Y6bojbc8oSAZ03ri6G4iDJSdBq6Vq
Svx5mJfVNdAjJJnGaFxIrsrqkAx0+uZB/sQhhvrM5ppleNir2GH+FOIjmkqTc/tD
/Z7vMyskTeoX3mZP4cY4JzTM4q3m5qwnFpE2k8S+t0WA+nKAwkorC5QUhbOEIt+2
VFj9AcoIcC1udpan5YrXlaLa4Q0UzWR9fZM/38M8QUENo3GRNSlIC9RPmbBLAolF
rWOuCqs2o2ZkKJoOkrwppoctJwTCdS6k3dNM+v3m4P531bwL2stHrhZKcILe2/AL
Fe6Db3y9TDt9F/T+ldfw0PHOsIEgCJOSbLmqgVWGbnjPsYVk/aqoHkPxdCTNsyBl
bWNcq3H0PffbHR6NNWSeM5ACpDvtJ2r5WadiZuXWZFEGp3uz06pe+nbTRk116TTG
FV60pohovhI4/BRZ3nyaYRUq09DEaf7Qr7UNCjDyVInNxnd+ILHcsj+2Nphd6/20
UQHR0ykZeBvpEE5uPM60d/YA97Fq6Kvi6M6xXJ54DHe+axtNw0kJL01s51730Dsk
vI5uXBVBr0UQjOALE2CZutUviI/UtBAfl0nnc4vpZ2NfNMw/wzQHcpaZ5bY7Myin
RGNJPzW8qYtnbMKT5MXGgHmpwy6wWsBxUDplT/48qOjnGWQ2t3y1fxaePktZ6F4H
soCeRavdyv8oQtHE1laidV9ZuQhv2ItFDCsgN5qdp1PAWfTz9L1iHXeG2lpyl/Hh
ZINxszju/Qk6zkQgJ4IJsC/GkbvKeliox2ZMlgy9+Bcm1JkUy7XHlbmX8sTFJEbi
xIbcg6rskP2sRYg8bzRoDXZJdjZap4UAEvWANevNZInUtIzWzcdpQbhuqjrwkxg0
hlIGhbhFBmQcCry4tk/b3Wa/kgavMWzAp4ycdwqW/FYrAl/cjkMdWO2xuKD34aOO
6WwfiGc4HhOOqAM54sV1CmLon5KkV7VHWez7lEAZRlLntyX/YsOiZsbUlRUP6Z/f
8/m+TeUpOaWYRmyHonyXxjFr7g3tFToXlqi5tf9HDdOEs4CvE/wJ3Zrx8X/Vy3NP
rOcyjqwFK/SP666hUkGR3vU4t/xq4zK6gjZlvM8xXdq0ZlEe1wKfP9E2Xlm0aVJT
h/n/cT3eRwh2ldi/Xy7WsRRZf3ZuxH2N8O4TQ+2X76PQ+h8RxNYk3M6R/N5FMvrg
oX1ERw1kCrMCY3zL/5UX9k3tHqcOmyu/OOew6/EHoik3d70dDnxeH+XT5VeHh11s
SkuSKsDZiU8hZkdse9QsopO/AnOtAL/lQ+jh7cIfj9sr4eBxbnhe0hTGAmbHvXML
kiT6jB+0bklkwFWrbk0qJu8ZbxbnHH/QUbBlxdtOJhZuLKnLnrBhcHfA8ZdvXVPN
gCiTg+r9QtJHx2zpEGdGFJszGuMds/zXS7fizMcxgAYcDOze6h92mj6dZA4GU1PY
zDnq7hZTbgoVz/Z1Wy1d0YYhNndfJUKjqIQ7YKhw6nvS6EMucLS6qPRGwCHT0E1q
mGqUJLlc4/YBngBcJIkCPxb203WSdz0qbeTmIbjHp3T3/P0OaPp66AXambFVaxhz
1gnW/IGE9q25Fe2Du0m3Owo+3RtkH6Hwwci7qHcRA+qxR7w6Xnah1qmt/9BOAhQh
Ojq4S/H+M+Qe7t3AoHH8QnBEtkQnRrWmrhugukWgLIFsYan5oHqo/U/kjtDvGkDs
fNegM7pTCHhfLwbKq4zDkQ5+s5R811cuMhpfQ6yLu31bs11T7Jm4u1kXzHNB0t3V
chv94ray7eS5peg3mMo9/l/1NIpwBjZ8rGUia51F3K4OjOQ4+S1oo+uM00OHWHmy
13tMK5McGk5JtzKqP8zrM07wsx+wyuCv/s/+5SpZxlOHTzYp6j8div0idsxc0zUm
+s2TzX5XFs/eg2EGpHzngASzwrgAUkPVteaAIn8upgXaqpNV/vBFizpTIHbZvY6A
iIN4h1Mt/V2GJdxSTcylSyZxaJV7JyxaX993SHM6u7yvdgvg1GtuKM/vBvCZBYu/
LJ0IQpjavnyfaexvJS436srSV/JnItXVP6PVRN0y1A+euTP9LLzWTIfluodEv7OZ
c1fQwlW2fME1/CX5DE3Jxk0BFlZryDomsNeVBks5Jm/tdBOIpvGy3n5CxVs29bhC
RciYgy64C0/yIBrJoSgmPTtaTAs/1R8lkKg71BpjxikYIbXWLXkRViMROFHw8pDh
0zsL+OF89lyOa9jhyyRlUS7crQ2KHqXJZ8jZfF12CmqpqMTEQvNnx77BsD1zueUI
unypnWIbWPll+3BbV8B3fPp6UQ8WGEV7J586iNFCtvK1zxUVyWd6CbxxdScs4yBg
GJfycEaRLu/c+pbo7gQS7PRvN3a8qgLKcSH2xp169qGPrWOxXWLMLFAuep+tm54B
WUJvEVj57vfT9tWleP1A4tDCU8Qai/uK3xnVZRE5t+WOVP/toUbjuIg/tKUZ++qa
Alup5aoudPaWoE3BqS1dCvmuoquBcEu5e5mWfiPj+RO8y7iNe3ccqJQQJGwM0Ter
Pu0//YDwTSZyYqurfsztf54tPsu5OmGFxPQTcGGymTT8VUZoEP9XApkbwi8Zh8HG
jZHpKNnW/QIC1XeXiMQyzkwcXRjh7J62JIZi81xGeras4ND7Mw7IExQbiXLdNwhI
SxeqcNvbmvyzHl8vNFLxDxeTlmdIxjXod7LwLOXFtGicPUKtzXPsKnHozUKsGq8U
rqiHEpa6LUmvMNlwJonK8L9HRLCo495tlbahU+HUgXxb4+SRyyvnAjy6AsKrN1iN
6X/1IZ3oVutdtKRH4V9MrTjWAVbWFX3BRnE0X/slqqSRah4/utYwOX+NZJY8lZnf
zjXwMT2z29litgIEyurHpkupy71Jy081mLbmlkwCKpZRuNWULb6Df1Yo5KlHCOVZ
PV3nA0YSHm8PG6ZHFHR276X5tpL2ZyZ9lvqFsyNNGlBhgAL5BgZRlDWS/qegCtqX
VfMZGSVRJdyffNdEE8nsnJHw0UHVKsfWkITerm+NewaJaEzZpOzu990HDNXaZ9L0
MPFnZ4ul7JhXBapIPQMVVisjGGt51SBx788aHnceoJ/xmyUI9i/QoLVUEpSc15Ru
bxfhGlhs3QWrsDrvrOWtbXab/dEXYjIW/4UBh8c09+gtMZnZSdcc1Vj+P4HAAg4x
lZPouSw2K/wAqXs83Mi5HD0kRvr5VsCof3QGW1H6iybT4x0b/daNhs8D8UChrZiK
xYEA+i0639dz4aXg6Ryp90lvw2HN7CU/GwJ19fzKHWeIkfwz+0vgl00k89UFHmou
3/Ffgk+24FdEom1flzy5wp8O0jfwQu2tFT9HHkwTnTK2gbaD5KkznLPuhwkfWCHZ
W210wJac6irgW1269ZK8Vp0hioBo7ghcpN68WmIjyiN8xHCBOWVU0IHoGX4ouZ7y
PEmk6/2qJyD7rxSz9ZdP2CSJORpYnHjHjXPl7DA5pNQ+qeXh6a3/mS5KuBoEeVKz
6AV/LW6Ct51WZjRJOTmx09wj/+xv7xYUEkI4G+Xp9YNoIjb88mVkzivJao/z5fZa
v3KdRY6E50lDdD95MPwHYBzSaRRPbyXYkKT0NLtemXFQzCp2kiCUtt036B4SaFjQ
pWbW/p1abYqxuXqE1Jtk494H+h5A8FSYIrfhZJ9Juz8DFCdLeLFZFBT8gnxQ6TC3
PgjTWtAlDrB3/ukoslBPmgpQmJ4iqVkem0Tual7MMpB4uHHheSVMfAumMsxSnD0T
AHLzp0IRM9MZlqW25OuN9nPxEZ3dBPB4Zr1lZ3yDWu3L7cF9awoZSwiXiQLDEC9f
HAAmC3+ivS3Y+vg5C0OVNgiSGkJXYI5J607zOSWHxNzf86JihDQYegENgOjflwag
pAFyojT7CEGp0WeS7fr1Qreb8T7/Kao+a9ziBM0RQYPsfZy+9GsXsYvToEG/ydNE
YIVCNxzJJ5NqLtDmca+5iJmI4BmrZxvkNoCqNxSNBwUnadrPg8rQE0Khd09R3Duy
MTUUb5R+GeJS+W0ab49w3jd798NjSvaIYqvd8TvcuB8s3U0WthV8kpOKAQ+GOg77
FBPJIEx+FCK+19qUrY0bngzHV4dl95L+KMTCQHcWPLrZuj7Mc6DTWBuetEnM1mfS
ok/pTdeiQe2VPiypNo3ikuJxMu7md8ecaVx0YRzZXvuuCiVuiDk1zShhlf8SHhXO
TTI8U0VwoWWIiY0uRuNvlyS1eBugTtI4oHCP7TowX2GGLSoX1QRTZJLKg9FRfij2
dyGaERVigu4mxebH/58XHgqYSi1qMxbNGLUTZ6QNFWYJ227f3dBdtxME5oxltizu
pdgnNE3twpVkxXR3YJU+B9Qgd3C+AfcV2GM4yZom8Cy82B1YMybRudIHn5A7a+ck
ZS/M4TKDkjerMl8LTTrqBVIlwvbnLPw/gkiSde7rUrVmbvftaxWOyshV03GZsUr4
lQ0kv3bYDz4AmQJ6dsRh3nxKSWnfcCBRF3kU3Ztrwt2S+X/coIU8wbBwkScM7EWA
cu8c+7CzMFJIkxg/MQ6vrb2mCN66sodMht2pVL0imvLZxhV/lxJk1E6vmJTn34Ol
HMbXeHqvrLUcGh5dpIazizMJwQRDbXgb56v+LyhY+H/q7mvBmkwhubjFgBInuqvx
CBRTdlCwRhg0ibBtIFxZOx7XY0CPm8pZbYJBs5MURGLNZoGpIe/RyxzjtMHAOY/K
QVFcjAoUQxrNDbOd5PSfRPL096fF8qHb5274klIYqZFF/d+xIP457MizYnnEYg+M
PXE2yWxWjDMaJA6bavYANUWumUDBI7N3qZhMxqzxCsTf/3/Ofh7tRTzKhV7i3TaH
zeb9aKAqDu+uDL6AlWuJqzBgpStvT6yK/oPRvWjPlTuoqijDlsIwFn2AzvkvIHdS
xrKxoTZs/jANcBhPv76eI+il+U8V29Y2lhqyuN9giYMcd7V+M4UjARANCOd1yMLe
lEPtq4UXAQRunshRwljR21kjiq+orxjCuAH3rMjP6j4yaQ8hSq5cuh+lqXkMeCsu
FLZML+2lcTmjhFhJm+4hM2VjaWo+WGPICIm99u6KDKpUsvNyHWXxsxrM1YSOrLK/
IR1qk6XuV2SVEZ2O4y+91Ig5rKNbS4c83+kQ0/1v3TznAdgv25zWaOExRqCWA4/S
yfi6Y8Zxmjgrq7y0HvsM/yH2l3x3aKKhbhALTSGrfoXoQHIFlzEt47mTJLRjyXAa
b5krvYeASc/5dSCrAkmv5BVl4cKAc0Wtj2RUKtfITvDrGpQ9NheMt+2wfi512Ct0
Lx2m3B3F6BmHF2o+XhpMdGLs5YV60lVhYaBCUPTxkQxpevxPk8C3alqEqWVAN1M5
y3hNZG5mRTn8crGOtllloKr4Ami0PYKoSrJXmQ01B0QSkHyBchsmheGq+6LCyrrb
a7SB0t6svWgeuccHzerkedgjc6s6hIHW66PL1iKbIQ/AIa3nTGkT+PskyUr46s4X
eMmYYVn66i1jlm6R0LbPh2HlFZslSoeLEowyUmfrRT5ax+90j3f5rQwI7t+fmhjA
pB0x6N5fd0g366f8CYM+xuAV0v/dQ2n9x7nCx0WMzmJ/t9lCYt3ce7nulUch8pTA
l+jmaf0Ct0KrI3HB+GOEUPNCqdWqDX0Kd/ATiNxH1E6tEPL2SIx5khldLYiJ3xZ0
nKWCosCmzksKeyp/nmVIJXuW4kSNEcuTPnRDhrXaeidatfmInK6EwxISHwQdh4O+
7T+QmiAJXWgaKVHRAR1ADlApTZvoURpM0riBq6/R+ZlvLLpjoHDtMD4idFOVnu7G
V53NyUH7yIa3Swj6gjhTNFTdEAxvUsB6N/M9oEOZZpyATl3/PHzZm5dIgJmPVU+q
JMNX2MkoxFlNWANfyrtOa1nErLYiagLEsjgfFcOEaKamV+dCQoBwFfooW+VnHccW
MLM3Bp4qffwJR4dbhIKYSx2hH7Jos3XtY1+3EdcXSFV0+RE+79dQtlAI/1MRqgiW
jnP/WpIvY4uCDw18+6Ttfhe0yxG0Qj1ON57A0m9olHSw1wFoOfWap+aykKaCy70z
IDw8U6udC+1T7FVKjn8wRDylvn9SY3pvBHMjGBtxsPyZBqBlM2N5w/nkGjZmo3T2
rS4anCZYoVfMDzRqYDwIyNDGQleJehhoBhcwXiqlC3e6zPpm2l7dXS1dQNnOVpJV
Fl1FdyecM+nf8p0fA+7b0Jvx/N1sT1/fxTIPHfTfibNAQyBI3i4Otb5FS3ASfxpv
RfmSSDqYYgpa23Igfcp8xrXoukw2I5D16TwjqgJWRqe6UEqa2vUvYULwB3F9E+H/
ZwDCpa4z1K2gJYDk42aI/jSgoIa3rdcNlOnkOTWiGugkvOZ6vQZWGS7spg8VXIVi
JMECONkj0o/BwYd/Osi09OK+clBMLGEezsYkXaTypQSEKMxJDH3oN95DrJ5eGr+m
e7VR0azkpx8yw6rGuBms2jYkNUA4B5LEXy/Fm6ufNQl4oyNYNK8+vIFFvpcw488r
qczDo8Qhy6fQB/3NVbwi8tI6dFwojcz8ARHrc8qiM8sworNcFU0foNCa13D+PZN6
AgGGZZCLZHYL50uUCdvVA/6BYPG7jczv2exdg5vDsjH8Qd/i2jXWtNoypdsvgYeF
c8VHBrAcTBJKwk7j4/6g7A9gC06EFEj6Bvlmf+iXOYlH7j56r/nCR9SLPt4YxOH+
UI5EZZHblwfyCJZYXajzzBdJjT9ub3rCAZTQjgidnoVgFHsJaFjvCPthOwu/DTVE
KRyCaG9mFCQAwR02EmwaJDDuJRv2JDb6FQZVV+APLp6PcwVNO8yphye6GhgY04Gq
CHoB0CVJOgH2ZaDW2kcTSg089EfhhpUMiaNIpmWlGNqEAbNbW5Qo6I3b0eJ7jlY3
9yPURMWxhlbLVzhqvNh45q85eUBb2WA82MTpbBHdgyApy7ZV3HgkQcfq7h4tolVJ
fx4I0jersa1LqKj8c4uk98GbqOUT6tkPG/r3VlqzqeW9T2/XFHRa5mbZTPT+Quit
0ggphHNtiAQA3ABcCSmZu+JCMWcoxJv3k/tdAdilFkxxHUiXBwQuyQmLfRO7x9mO
phl4LJhiHMfwLykG7tN9F/nyYL+5Hi7k9ssj7HFIqzoj8cX18NrSPGLuV/Pn3i7v
+4kmbXVJgST62O6HGluWFRCjwYpBGtjof/Z5uiBDc3XMi4hu8w1srO+foFaTs/NK
R9taeLUoECDHkRHZdFMFuTUMlmUKkyOl12eZF1ZByUbqVsYD/Zo1y0F4bS3fasXT
UUaAkGEmYzvvlJPNpqpYc79q8dVGLoJe+7g53VOTU7djfKKeW9NjYilYttAoL7FB
e/xki1FmUVAC00+pO9MhYXBqhdqbuE+bFAY+5rE0m4bCDZ9qzKAat0Ugzprk7Sqm
B+r0NJeV+5D4EI4k+hQB+2twZIzjcBtYUdxBvOXutzDS1mNnae6fy16I25m2sYa+
RMCZFprPlv29sVPdymSsrdQjv1snmE1LqoNlX58pv1nnQdeVNTjb/3NlEWKUZ+Ku
BcoW3vRQkU7QGIlH7aYvrulhF8VQFXzHuqEzLVeydtEG8dxOcZQ7RDRTrunkvRLD
vZVIU2GdUaBE2AZ93JRUQlgkNjm1TPXKY/ExMzRUbu34Gm2X9e6EUpXoIR13gNhd
nQlhCeil4kZ5tC1UG+t3rwOg2URpzp8IvyDPV/tKOJTBrYd/7TvW7lUoDGycJGdt
mdMnEg/KvHy/JFHRZTqGdtyqcXOOLy7XCKo7ofMXnLWHrQuFcR8MiHARw7z0ihBm
ton81SxtnqA798bfA2xtZx+l8h4ZDzl5AmFumkqaiQM07qL4U+Q9k0+Mbhl+k4Aq
45zToooRr6Gwla4Wv9/Ib5+tffh67oMSZwTzTCM+eGU5qtqad6Hsg9ZERl4FzNiv
RuIxMAeLhBjp5hWFvZLIVGTOax/l3UUFDHQWpySvl+Nh5b0kDwEQe0C896spPoVb
lqVMfqAGAw4v4Jr7KUdchsurKbVhB4UF77OwIlUGyaCnBZ4mdGxtOhHBB+vWGu4h
NnQYXX/3SqyFO4o6WkRwesVpWRgS9ya5Tui52CefVMnwkpbJ671WEgBwLbpHGCmC
lyYf2kQCcWXjMXDRoPxxxPYL6GW+jJGQDjRKFkCddch5+dLB+4y8+1nZ5AIqM7Ab
stbfA6sFY+HzNMlTE0MOdI3Tt7l37/tfxv6fYSCQh+nqAUfT+/SehTdp6ptxCVUk
NT4S5IPEC6J2BSUwPABhdQ5j+X4j9PQKZjcredGBbjYYU4/krhUATBUqTYmTzb4e
bc1mjT+89vuJF/ev4z/11vsAj/bc0PLujue40W3uP20KndqMy0ekSZx50gzzYyBe
/rrp0oLFCZZsgregnEowdENoEJFVpgDlXtEdbljLnJy6RQYZOeRU013twAkan7ui
0RlkOq3FWEAWkYJB9D3FY1AR9RV6qiGajOezgF7yUJ488vtUSkVaPiR6FCBKz3ta
pveozp8jQ06Omgyj8KmIbaO/7EGRW1pkpDeKbeb/s1hTTbGcGAFsCT9JpBRN5GEL
CmBgse5nZ3ReVJlUOg3+LfUzF5YsnjL4PGMy8Oq6JaiwASHtvSjEDwKEs1NSDOG/
hBGMKwnD0JvJVU5ZZr2eLBY0C39Pqe0SvpZN69JbzPk2BBvcMJW+cpwjr7qDrdQw
AbdJQfj3w5UFc8Pt+yoqX3xF/d6K/B4l9EDpy10eOX5U2RUDLNudjreWTuP5XdeA
IXLegFrJFCGTiftbSvLLE0LSXD7UCThHjOhwcqzw0l+5Z0JnP6Q0oIC8bR67cIBm
UVbqBjPB49MMM75S+ZgNP+1wjJR12/nQVqpuJjAwBHTSciTIvnMKyhE4gGX4x14Y
dM+95M2ILqkq4iDeLnRK+Shia+trZuWHir4eBBuAZuePdKNKZznqlSB/5uTy7mbD
v4tqWV5o1iEZl/r8KYFZeb4j3OSYXJQm3U7qEVhYHFrJPsA39MKhsuQnp81+wiL6
lQ2XgpRx/yUr2COQC5U0P8BqQOJ6GZYbU2/JeztW1svgL6GTVB691BN6H4wo9gJD
RrCxMsyUdsivfeeOWckD78c2wi0IrNwQ1pxNN3jsSdIHIhg0R5CgUakeVEYHClej
Y0qJ6UnNAfHzqaNlbEv5pgIvshWjirQRNpKv7gpmdlScovbqSuXPjLXRh6QWhd8b
5Cnql273RANH3Rl5NOeXv18m4zWc2HWU4MP4iI+BeVfNUj2HyuvUCJyAnY2KmrTK
/TM+vZxOKK6GhV9GC+NdhChEobTMtJLJUF86O8EjmNegSUxS2Y7yoHV6ts7QNEDW
9JCJYwgnoTDP5XUl8LBzKljxXzmR3N552K5vLlp0HAnDjEZR93LY/tSQHV6LTX90
pc1qk9aJvi0pIayzLge+x/4g9qexfVI5ehJ5rr11Rhbrgi0JLqAsPGWUY6BwtkI9
JNqy3WOfCHYnDjRj61xBFfu0gleLTWmKivpyYhF6qC1CcQINoA62HA/qmglYKwVd
lEXakireaGd3YPSuLkhuHIFfF1azouECVbKVRxcow4EpjBHG19xyhO5MwSrnbmnk
/CoPsQ/kfoMGo4gHfHZjvrXhj6NILjIqR/xtR3cRZF4HFf3GFQDSsdvkS1bq3u9G
hwi1qv+jWKkfOvs2iPr7VmGICS2lAYHVRsXab5NT5hjo1aBjX8jHAde+/iVkmN1c
4ZP/+d/6zca7tFZEDi3Y2jYVX3wN/69IlxKjRf5lOS4CIUmqGAYLC3Ys+kSDBgWp
e28q/Lu8ljXtW5hvoW4Dg2ulsOJ1CSvzwAqBXgVdig/aPH+cfjSJ9sn9de9l6l+V
nN0aQDvgwGWaKKnNqP5wga9XtCj0jr142kYdxdQJLimKBnVBKekans3rEQ5yUYx9
JOGkAsm6RQScyz46AdTqV/P8SCxkugUE+1R5NzVIP5Al0fSIXv/xj2fEK9WqtSJ5
wj8Cdf5j+qHCmYNFYTGvWB9+HS7sfi19kMyYYvaBhxWwTDR02i/yTZV9KWdd4Plm
+y7yVpKpT1kugGJRg4GpPmnRDU43aDyvlvAL4ZlU/9WLjItO31UvR4IkcTwK33FX
biT9SI64JwuHzUuVjEdpeq12ovJes1hUQt0e1MPfmdJ/IQxQG/slJze7PBYTvbM1
xnkKdgGrsT78MQh/mZ29J4qS0eljActrJLt01luZ+vx0tg0YNe7wc00NuOudt1pl
DF1adzLWPn4XRYlMpt/XlI6/Q2m6gBOHkmjzGK80eucpvrI/GrH8bbtGwqVLVxdk
vfZPoAn8Zp9AIP1xETNAbI0XntnhzlOvGECVZtPt17LpF68cj9dW2tX3YfIvGkaB
OaT8QYFUVPXv2CDDexbGTtav7NcjIltCsXqD26kZwyFz6WefiXjnKYh7e08ukWeF
dLzPWGAD194iB/kpqvWQ2lyOzuT1CdX3fsBvpgr1HhuohUHcKb0omcKU5PqV+bml
OeHovXemMez8837+InG9/S+ptJlp283xh4s+zi4iguOCkJcwC8jruG9ke1nCrgmj
mQOExLEGr4xWFx4nA4yV3C4IocwJApBMtIX3cBLcLRN8KEJcrkaFEfMgG2vYkXl/
htqDFjRmDxflqPFh2t7PDBt8lK2YO6IIbNzOe7SMBYTSNG+XJ8fSYJ0E9q8Y1Lib
pP/65WQK9md5WqKQcACictHnYvm1JpldjLKFZLh+tRx+fOSUuhF74VSoPAFJ7mKw
otZlHLC+CO89X1+0LL1P04M1kRiKPEjkQch4BOZokRVQdLTKlsB5QoGh1HnLle2K
EWYgz7KgepE8PJuOA/3pg9E3FNPUkb0pR/DgwymF6F7/QBuhWPXyoeJTkbh8ogKV
zk2aKD42rzO2oJf0sh4EVqYo/YRXoISFjOktnT8zk7bjESUecuR8HRiYCtsvLRfJ
w2UaeuAb67JhSojPFkWB6d8rOYbhRICAnsOfVW7SlE8G8CsPafj6fD7vCaBofKAH
fHEFfGFEgAFIg2GZNlowB3ZCjMlwBlj5BTJTtwOcfOn+KZlFwQEQlZJz1ftTnnPX
zOu+hRcbc5Y5s3DwcD9Ul+xEi0Hb5p3UVDb5QHgPWX6mqiTV7pVCVbDGhURlGkt5
S+0fLNMpU7KQTHJnYIHh6Jlanur7uNsHHDNiLw70/71xbpOM8BVzJB3EMZLiT+ar
bsYvoXptWpCviZZ18T8/yXlZwj5TMXfdPSKihqsqvix3X0ZAIFzNNlPYINSCSCGl
DD9FSCVto77+GMM5jRhL76AyFcnZv2WV8Q1uyzrbtYaCfiF9VyifDlvrOvWP9IYS
rbZOHmqO08FyyFTTXHJSWIqqYXL/NlgBUBIEcdNB58+Y4RWEdqQ7gt8oexbj13Le
o8ezrTwUVyfcOWx70cL+5fKhoX0KerrtMsPS7qKj02w2tLdC88h/ij1IhbRMAyi4
8RhUpVTVsDhdW2wkfMe2I7khLv4He4qvIp8om2RW88WwPPNfzoQYr5ORXOzmLPuQ
GD0nJE2EeiWZMzJwkmJOVtgc2imsBoBd2IMro8SX9Rpflf0iObiC3HMJ32noJDdD
7OBxh11dP6kn/AlMNE7SS6+qz/PfXjRRUpk5D13RUIx/7v3Qg6W82jPADN/nAKhC
M9GpztEARbhPTH6gd/RelaTuFU+NBUsidFt4vSAaNFQ/aemFTFPI49eS1YKezdF4
N/xEi8r2uVFohLZpeT4N5N3x13CFgB351yJ6QZuo8Knu3Q+r3k6ITOaDZ+ofCKsT
FfjTDGXNj32eN4nHblOaT/fsAduIYarcf9/wuFMRewIkH33Jk62SpbplKPBXikSW
OoEpNjb/dpUnDV0HdEWHb66jfp9KJb3Vq9VFnYYw4aLpg8GFKdYpoqQ6boY6bnSP
d3gSfhLIM8ag35Yjpm4DON55IzcWSxLQ391H21z+ExKwL2s/HLGxbR1S/QYJkGCd
UE1bZkiuQooosjgsPT1pCRh5YUXBpZb21hh0RBw1yWFq/arYvmb7NLGIW4pqTQVU
rtsRmkagpOjEQjIUPWBxg6jgev158E0cJyR6bElJwA1aN2OecYWLoGtbdnqDcBr/
aJGGTv77C28WUKEaf4lF5vCGga7XL1tW8J6Y42dldDO2OKQzpFpIsB8O6kH+45S+
FnUJ3F3AFe6sBUmtO0ZTf/VzJPxqpo4r9qNA4mdg81A+ICEveb23AbHwanQejq5m
haEEYrNMob8Q7cP9/y34Bufs6DlkKsnDzAa45HHuBwIevzPP6jnE8dVdXYJ3FLXS
lw8AkTkIkYHQf1eSqy7nxbDT1dnQXSuxTZ49m/skPphHcrtA1hN/DFU4/AKkQHAU
HObzOH6CiLT470rJWT8XB8/p+eL6WGLR1wNf2CTZnc3pkEM1cW+v4f8uxTXbvvID
L4/uTPSxYHq2FjcEoV43IzCxQJPHaxeRUj8ARUW008WXIVv5vKN4mE8WCO3lZYZL
zAYRmPQljONRyL1gud5youxcn4VyU/XGn6kunK+22E+bnHSH7DJXImvJp7cpbBxk
P7j4zb0Ab5rJE4P7x/Hm3bbwoEL10ycKegC4EB0qtCs4/5sJ2mI+3OPxd7Kk4OSM
ZIzmhAIjgBB2/pvfaYvdz2RJfLXoQHkr5TwVzUQ0RRUdvp+32mJcUe9TQyvV1XdO
IdI4djPSlwuk4pus1l2jTjl3cvIq1jIGNs1VFdoPgTJzuA7qzg8wHhmDdzCU+B2I
2dgavegWbSzNalkQ2z2CzJE8FgvQjqC2ti+jplCV70eNulaoyylXx3VIacLeOB/i
/mkjRE28rzoEe8Hf8IGuthLSsImwVNYSanlJXP37JnQD/UAuaAH3hj3Qr8ETQHlb
mZdRllR1vM/NXSs6lJ/2v0eaQe9uwToKKcSTDqZGBM6/GLv3MqCtMJlOOehBiJFu
ICqnwyBJ8QPHWOcMPK/3S1PmUXSQjQ2q5tTZBbx2N4lstDLUpa6SuC12050WnXXP
beTar3DV1z0Ige1lp4IXqST46Lxjx5/BU/vAK0+2GKDQBYu8IE2ddEsswIWHPMKJ
zcSMSQrNaROxP31EMX4ku5S911cNM4Nl0qb3fUooMLcv/YSzBK8tS9zZtIqp4/6R
Huod9CBEBPzcWi6KzHxj/wx/TQsxhOTtiubkzg7NPizSlM4sH8ax7grdwaGIJgx2
lpgvib4f2HSWlsYcNne6uqe4IOtD2YjZFY5cyLI+73PaFYQIzW9uNQd3JTTfU/OZ
tzCnCgmXtWuEcyweB4J+sVcad2wjimhqYADAKmVJ/LmnUNH6pY5P+I5n0lvKgPd/
BC6Gs/mbPcqWnQiqU6lcJGOzGs0kNbqvaHXc7tSmzucaLXJjuEWBo3nD9DLmFL+x
Dw9GSVR8650waLxWr0ktqQXS7tcv9kWMcVp7OBrRwcMZQARlxg3zVOJThniLbLNc
O3iLOQs7wYN4sqdy5BhUQO7qE8tEkPVspwJlH3a+MWACaDSe8JVQyusU4NeOWVkF
K4SUe7ESTRjnEKfwAQ0hU0g0mtsT1POP/h2u0zM1rdNurymg45fMJ0pPlZhc/Hhr
hWpKuj9JQ0ry5hG1264SfCJ+0EWLx1APf1c5wm9uQ2sUFU6uqPhJtTbylEazWS8+
KkGu0iGdLSmDS3rL7i5dTfT4RZ2BRjv0SRUctjer8axRbtpmIYL4+UxDTb9bTma+
e2hp4rqNZtVUavTKP6CCtOdc5/GNEeqFRXMRKPDzkDWI73G6yxtyNwoGgYw22fks
DQeIGpMEPtkrVtgf8ZYnTKGTJ7MoUJAeykatfhTo8fxpkd0n15nV3NNKM5XmkdhB
AAs9fucwCqTxCz3FNMIPkg917vh+p3OKNEspmZN/MzhKuA/Fm07g6MaZNXXJZbSL
7D/QpjIwxP9+nFfGFuqwvyRWUwcInGSY2uEyT8xiZvwPHcXPyPRIsTo2DVrPl8FW
iyReNTu7MoeEgq3DeSi8Vl4WPx3tqUlqsqjK667zX//fNVln48k0V9vuAQTEdH/z
E1dcDRqqgsQdi1NaTBncCiDdWCAvo1FSAd6M947tYuUolWzRnNUFletYDqGsDful
Op0DCEg/ZMMQYfFVDTzRrKSJfCjlTI/Zl78oRrQO/sh8JCArTnv2D4D9w/7iG9/M
uf9TG2OoCe4cWG093cWGwqI2Zo5rs62ysPPkE2Z38ssVYGC80UR2RM5iIoxDVlVJ
sTok9FPd6B9zvoXHGxf0kIlQNKnOeY0prhbBlc4jNm3d7j6gEvivH3CYa5bWezR/
vPD63nNnh517EZALgboS9j69UhcOAjBoIs/BCEd6psNfHGirjINcWpAxCWahTa3z
oMM6T499hkYbi4VW2XJuErMMcozrxXfNVqZOgx/Lxee9fowvCAbGj7GlglUWJkYL
pBRpGNgQw4iRSC5rdViswelStglJQ5/M31NPjSDWtF5GoR0C2sjqFWG+ykAnZq/i
l8CZnmHU0aVlnQkHBmJeyXxot5j7r/ZBa/iCKTbQJElAS9l/QZlvpGYg5BV2jtFP
SWJq6zOD3d1TbNnNKSQbzpbY0OniGJjH+rLgyrO7xJ8IT+kytC+Sd+SCihOZQgSA
zj5acCkBgtgjVJ8eWUwHj9F9pHvicpDFUpsfjUdFQfiyA7pOaEzM2k1Y4A99HThF
8GqwFagu6g77j8J0auvmBxt1ELVsSjp4QLvKIuWiUxnyE4ZdDcEwNjn5c3f/gWbu
VlnBpkCQiwlKYfmYWrGxoFr0GjSt5Nl2ahzo2dMgSytd8wRgK1+C72Ejkp4FfWae
6iFmsqfWi22mX2r2rIuDRB1P6dhWQblo09PRCi+r5m1y2EeP5GdxDz+N7zeJ5cxb
Y/LXi0A/5k2cOoKghALsAo5hJcHrXUcZcW5D1EIishkYinEVbz8WvJJxTjjycVoM
ShKES31qEYvxVqVb+hEOyIMpICop6FjXgmMM6952Gs+9QBYpjWLVk/yeFKsNuzul
/cyKfXBzvpsdXH8mT1SuvjZY7RseFQhKWJEq5UNqy2ta+CBr7lbPM/FYilBpsfjw
JkDhLphCTuwWdwpCZ+G+GwtRwutzGosKX/GDBpTpYhz6id8xWDCi6IYWPydFr7+W
zKkx92nKF5wAbjaWIDxzIL55MKmNEs/5tQV1LphxVGNhVal1Y2uhKAi4QcuMUYwM
32IU25aFzEYevVL08VBaqpcJc0dTfFG9GmX3WySsqQXYPpldjsHMorSgYluX1n0c
DI8splgVy6UzcOJUTGwHzT3ZRxvO6re6pvl7vCsr4JOgqB0MldcP9nMlJ0ClGrhZ
IlfhHtlEFC5/U5YLSepyuEJSCvH6iTuEEF8wuqmmUFylUYfFesO4XO2dJ1YlUEDN
lX3dIgmhX1CqgYPOZs75esSe83sFHBdm6VGIyFRr1KjtCj4detkGTCHClc1+DNoa
YGd8iONU0smfkLVMdBoBLWVbLcNY5f3CV9DBscY84rAIWYFhIdFCtBBSkm5RFtrj
x1luvAfGvelhFj1INY91jJW5+F5TAnPhW83BxoRuJ/Mme5iua4wmMkZ7jYdv76Jj
+l9RkYdzPLYT6V+dqdQhUJWn/2M/2hdPV18bgZRnuOWD9s+jtBNwlpw2Htg+wrCF
XG7f20yGAZxzbthgoPPP2n2GEtvc4CfcgvgwMTsxu2V2SWwxcb9Liqpnx2lde+/R
hGfCLzOgg/llL7+0YLSPaTaiRwx9+lAm2AfMLRQgcHGGqjWB9AtbWmPPeoqJqGGr
gyjkzjAf8eaVTW/EQRgjGrdwYkGNXechSLLqWRUH2juFIcUEXf1A5E3nS5dPb7oN
07kG90wBVL8ohuFKl+9avt6neo7ln+fozX69oF9jgecuhOE4yxuzQOX6KNQ5E+dk
dOYL+FYbosl3aW87470S0hBrDsXZUHPvijq9VB3li7WfNUgm34g16Dj0ND5q3fHQ
81dVZv5tRevxKE89zWfu3GBNVFoH4GolqS5cqzWj7nKubJUFFutv0EtrKEUCdVaR
Imw7cDTN+AFqCuFsTMbe2CpQg/N9JpR+LbsmpJFTfyLOkT7eCOrFf+icuPV9Aovh
UnUhvADjcDGVxIogtRTb4JH0lfUTVane3csD9g4FE9r3TU5kOoVdpVuIR3MYM4L3
HJItHStoq5759nGjOs3/MkQejmACSssYtWtm0If8BTnWZ2O9r+qQuikE0jvu3Xzn
hts5PuwUPl0TKdCdV/9AiBZOm5oJAppnLRN3WP70FoNBn51+Jws/Np1FyQTw9BpT
Vn2sAidCQfr6kJRDbJDsuNcJHZADX1c/a3t3B9C/Ahz6TxPpOx5BvNlezAgPbj+1
NRc4Zb10X28ppSKS5Ucpbuw1+p36iMpHgx78Uoler0Spu3kXN8ahKnQDBD9V8E/t
2R3DKKA527hL62JS5o/4GuAf/zMSqeVJDozr/U8jfrPB8RlXH/aB59Py5oT/zbb8
q1sSeKcY12K5Z7tS42Bp5JRZN1GEr7eJ8H60p44rF1bYPQ5ah1/Ad5xyOjE5x+zZ
4Wb0Bd2X7mdVZqr6TGO0kDt8uLUx92OwB5sYCyFx//B0zLYaUz1EBC63thCSVhl7
yxq8pHyL7pwYfR9nCSd7kzj0p8qUWyzRidgb+kBMA2iFsNGQP+c8EcBJ0DTuDEeL
gIkr2wdT6MWD0JLstkQEruvY3qOTIJInyh8NViePH/m/5brOyu7VWTn2rdNlvoia
muANfwkek59akokLS6hVL46SSdSCwSG1eh6Zh46EFiAAguvVNstLqWBFDwmBVMHC
gFI96QjoMFmOJmefy3YTj0HmB1m6p94C6p9Ud9OicQORT8FICW4DvNQitpN+bhXQ
bcacIgqsrfK/fBzUuyY0TbSbJOFCD1scQndk3CcOMXoE06u/dtLaCzKDjPJPqE+Q
J6gZN0y/s1c/+88L7XYF13hv81z4d9trqsi1ORghlAdYET9qGyF+vzplaRLzWhHm
NEP88V3u7vuzmwOGVFK5Toyut7rNxaKOnQpeCfVSxldmhNFeMZB2gIh6Us91dRVg
Dn5KWHHxp6B51EsSiHGBwSRukYd2AwMTyj5aa3jdzp4oDMENLMlWkO/Pxypi6mkO
UgoyqywMJuttvcUqyW5Qk8EGizqjbNc9jKPedndpqw0wN1TDMCC5EGbbBPBMfHQI
QnrjhcgEHxfLqPBKh0e1ElxtH9VEBY9TOhdOmxRTfglF0ZmS7lQA4kuYZu9R7GcG
Ko1yElUqYjOSVbs9/XhfV2oB4C05cOn30GYj8G/skH6bkuUZQeZR6TZ5I4Votv7I
4mwj75JZs1g54ct4UnrLpFXeW4YF1wTI3RwQSXnUGMc/wBDhrsHQ0bXUS+/y7+sZ
9k3yhiFBK/KiTDir+iBL7SWWPBD7QJfzvJTZf1YlOfUtC7FyN8SFmC4hQN7C2Stp
yh8RaRlWzGvBq1fP/UNDS/fphvFu0vu2bCGa/b+5Omvh4brBqgirAfsQQ5z3qIFE
rDptY3++WARh7gZ/3irMhX+JIchRXIoXtsyM/1BnK/AbyR0HgUbx3Hg9xX+/eHKu
sW08FMgHz89G3kaYmnezIcsvrA0iHLG0qEDO8ySBRIY4Vl5q8lj3jvGb7xHTZgB9
5UxrRT182DQUQq7xvDo9Izu+tn9FZgH0bP5fAJMv5g2OFfcyfIfelurXbv2lcZz1
tgBQtpXzXAG2XjIH0bPQdd6I/Q71ZB7dmfFJY4vzXBiiDTF9UV12luxEMBxlqvwk
2B2+BpwfHeO2J9oIHgo7NqMj+6vJaoGSEJauC0HJB7S5rt/BUk1tyLcUQPAVdpPU
TNmvhalSWZfkC9JaCw5cGu2S/+LD5954Ut8mj1rVQ0SvC6u1AOtlTi1lQWqpYsFx
FhD3MvyMrpQEfmmuDBMEy7puqo++YoDJbWc/6dEuGSJsJuuhZ4nNzzX0Ot9/7+L7
r+GH4qHcBpX5ojzzK2+0x9wfQ287IEZzxgC10SEBx3eiMe78h3q1i8ZYQjURqjz1
OlzlGboSsQsnzGVFePxt6RKlanSBxfnw2J1KeZ5kGjKPJcuQCa3tmYAReqzXjja3
dEOXzalbYJzIcVA7vChBvLu7LPlj4RCCqCm+cIAPWocIE7xE4LeQd9YUrJlMyLSS
26EqBIYg+nkhm2R1CfSiQ/YPndctIScK5IhdV7hxqEdUtFASEL3uG1yUclGw7pDy
3yLS0+LDYSuMfZ5s7JXwrUnVMBQPANdRAa9p9jZEjwmUcTb6djqqtCSoLDZLi3ZX
TmsnOO9ANB8rnd+h7sZof1GZiZ9MLD4wcAHvvWtr3878ezD3SdR77eKfH6MuKla6
rcRy3sto+2PAyrIEFK9usmCtMGqRmq4MwCKjXQirKU51fXSb+3SQy5c7jLDttU4H
OclYAEl1CjkM1snDmheke/jWJdMbaY+67jl/Eb1NoZS0yL1ecuv3cJKbu4WeHGEv
O2t/PUy7NBgZ4tFd2Q0nTZEJ5wlHaCnf2gqiaPxWmwv6KNnE3PMumjfjC3hgNaxA
sfz3FCVlwzWvzY2euyhDYv6dFYwdXj6KY/LdJg1CwCOxSc58RFWP6z7kxnIEzMnT
xZ9r1R6n54+e2i6xywd92q8AhDSg+NV2BGTwt2D7siQy9VWe6Xk618IDSZKqhwp2
/ePPxB26FxcJAJuF2fBNHURtSffOwg9kcUQ6l8oc0GKkvn3hNyqKuHgg6HX7RbdI
Zl+l1SI5vcpwXHkPxkZl68iOjiINM2U8IL0RW5LX4Eyi2+C6HoZNWlsPcvAmF1yq
FDsg1vIPAFLXl7Fa0XBsLeysaf0HLoyZClAre2GNmvMNY9TjKMaCvNkeEfqtCrx0
P8+ax5TubxCukC4d/ZTkJmQkUibds/FkX4udoAa091W7qx47HvDPts90FUJ+lTjq
jzG1zF4WDUTviVXzvL1aA6k0SpLRspiiY9M/dHsJa7acJK64WVOVdgnFH6hnWDT7
QSOBPBVsGVA8HhowTwBIaTak2xnJCZOz+FP5AzkuQdTXDQO7zYixEidpPeGamK0q
B/rGED5dNcB2UcUyt81Cm2dsThJ1EFCZofBce7C+2e3iQtaNxfxoh+gsRpm+aSag
vyWsAVzStSrrJTSH2pkSIssP6Qc/KfzX7M9HwiBPcbX3UA1wTVgZQDqgopaWZ4qv
3GKjIES4yfDzS6T9/zdlGY7OJpqsOyVqM2yXMrbDExxIohR4bobcvN/ktt3aY5kK
GhHLW4HMpuZn0VGrTQOuzqFJeYrTxPBcbj9KbBMrrbTEKyQ47+hmr9NIS2zvlnhX
Y21Qwvp7MCW1PrD03nFrYg9N2rJ7HxrWxOeE+IaIp7esVWwVy0UUW/eyI5wg0kda
asE6PBUcfJseGGFOBFnFxwXO9L+ue6eW6bR29jWYQ8vdGLOzT9aDlb8QeWpixfMf
CO0ybOft8qNfWQXq/MAvNEDb200RKj9CXz73iaUM9zRwTu43MOjAscSnBtRxYeOj
trv+7m9kKAVV5QWeOApTbYp++3M+fmgjjN3btA8kP1Ce6JumdcqnaEutRP8WFKJ9
xv+2t9Y4pFo+pCVgjMk2bpt9l6pCWYpsrOzD/RppRFmmkZedGw2rqStUPJZuWYvx
lfefYMVcIaSaTMDfR4tgItoohAWZ4JztPlHLQcXtawCXUCFKtAh/qO+UhNVVqzOH
i0aXR0opmduKEPZsouxo1692moH1Zqzvl+uIGsVGiIrwbvZqGVjyHEVtvwTKE/Bk
zJ+id+8mK05GMPINciSsLe7Xudybl7TB6pdlGU6Asa1G6mhNHx0kkrNhlAQqLPah
OpDN0P04mYu51fAegumBE9V9vT9Uvo6oTvKYIaUzXPCY1k7dSVV04jK064WwlrzQ
yEp5LGYL7lvDRR9xpn0pEgmZUnopcE9+gZH18snoTO2blCn1CgQ/jXpLT17zM4S1
y4ip62G/NmPhw8LQ6z1HL1dG8IacEjJdG/1oZ8GcY2NrIRJhjE5PB8jvjPsx+r0D
IahAqlMuG4R3eAxh6QqWLcb3GiMXl6KquuwklXZfc1kjNjAGWi3qRzaf8/ttIzd1
u6TQLoZ3jsdSN5exAd5zcTkBpathm+Sl41NP7m1dgLR40fGJaLNRZa3VHx3Z52j6
REEwM8HVxj4me4w+Dbh7sSOzMB4BKdmNqddP/aNqMXiKMmBxPY2VApK9IWg6Wl2n
tcX5Edi2weQ3QKjmLla3kqusaP9LDI+q4A/qyWzhqDGNG99ICcdnqWKC9H4DnVsF
h/B+yroFVZlfcwvWeOlK5AalvMJsc8zRzXghRXXKeGvb/RpEYNPvtznaJZ8uz5fe
prmTrEPbseZvE4w7zm0eoPFLjp7g/caX9eQ2p1HF0DKf8o4ljCJLlRZyE9FyybBZ
gcJTJ6nToFioucOuTkt0fBA7TtuzYBlRcXHbFYicp7FxEFD/X4gS7izyJWP6h0Ma
L7q4PD8GSG4PMrHItvoy4YLK7OHGT2x6OsGgECIWv3VFV6InOu/S/N9kGnab3mSj
6ltNpuSLTv8pecpWY9pIOcG7Q5otyt6xkyVZPpO/UlZMZwUTxgueDTUv6Zpq1xlG
QJmEGKUeYTYpz/FRyxqreGEPtaMAe2y/JIb9rkZcSEFmtwAGjoCD2Jyyw22bl1OR
dfTJwLMyR5p9NPj9tPFORz6CVqxHqqNwqxvtL6msIfDumfD0Okr2ZijfGQDwG27Z
76OXtwlr0cdgPkGgnd2HAst5msbbgRM5KFrtsv/i0a+uNrdr4v0xTwwdDUNOAtny
y4N1rsttwM0dk01UKCLHBQQNEV/KmsfbQBIh/O84LpbaZQJlY2J30Hergg7Ss1U5
dLa4up+XF5JGJ4rw/u1gnOsbLetF/McXCJ5t2rxgu9iRnWoKVNCbb6v2c89s+4X1
xre/SPwg86fm8o2c9ZWrfk58XLA93QLskZLxwahr6YsRVJUiCceiMdRR47S6odNL
WGYzTfeV+56d7XyTioLRo1dDHGr26oHc8kK7UzS/keJSFUxb9Lb3sx8Fkrt/1PuW
+ngKlwbuuiN6PZBnk8pwFyK2hi5uxmo9DlGF2X5uMYij1MIR+a+PsVuVAzYZ4fgB
VBoA8yI0YuDvWUF/myITVzKaBP3ZBPO/qvb8uyffy4deeKkEfNXjFlVRJpNW4Xj1
ZRi/JuDR/i7Fe9vu8kS5310ZQDWAeZzjSCTB0xJwr4Ylw7UZeKP1E7xw51ZE+3Fe
ikU/AbQUhvAlqUT7PzNe+Ouri3CHUFt0YSBZnG42aso1+EdcI8eAZSjg7/8IqWY1
jl69o5jV6PsUO61f8YxODqm+BEHYUMzGJJ7zyuFhmEhHplf+qR0pYyDZOZx3YOxv
RtOjmwUvTmCcTMqMTiVTU0muYKoR3GAt4FC+5f2dMmOCPl3Tycit4RMiSQVoClr/
mUN+fBnzxesbdYW+ewO3lFkDPlqbjLqZR/nHZ60hhynFs8XGyELDvE1qR+MVe13L
XDEbkKqP6ikdlqz+IKlDPIPxwOWXzMhEvnLbfh5VQMwmWDdCH8/p2fHW1A//cZaO
B+zQbVcj/8PFU1BILqaUp+UnfterybpWiShWPIABk5PpJOVTH6pTTyNNtEM8/T4y
cFumX7sPJb9PJMU5UZ3eAIzIjqkC3B8F92dvAQP9Wx8HkQWBluo5ZOPAaY4L7B4c
ZeDBaUx2bqPyz8gPoixOwduZ+tQJkHJdtD2SUh/Ol7hN7BNMPtMkdZY+/q8H65Cd
rB7CbzW2y+UbtI3maAMY5y8i+ToBsjR6Fe6RUHuCfrxSf8/57ZMXVWPul1PYOZah
f9rIO47cW+vFaW9SPmjxi4fzRoesSiwkxpzo+I76/mVWrdSJEKwlGSTzO8LlDADj
CP2zevnGSXe5sDOxxdPNQmAnDDLHmbQs0Kz148M2VXKPa4pEMeS0jHVly6Ocfeu8
uUIXpjKLUwbr3IhTmEoLnBj6JrImhEdELdKi6ihpKA8dX8MSJJjaGvDQt6/FTQck
NEPerZARNMjb14w+aKlWX2VEqRzn6bpa9U3QQ3k9WsCu2vFCNlrq2GGZAI3AqvP3
6YzLNFi7El5M+isFo83gWOgx5CKaHEO5wq3KcmcjSUtVrynVoMwrPreqvAuFOVyQ
hU5R9egaTf+VXxDAc51tKZh6lsHPvXd9rFRFQU77Quv1754InuTjgwGmtGgdLupb
mqDGjW4pS8MXNvSOMN9M9WKHXdharbR7tNlqiwzDI/bdPzMhUU3jKffKwKPVsmFa
Pp9Ox1B0IAbaHFf/CdZo6ZpICcdWh5/TBlfA/+Ka3EUFfT5zTD87XcK+7RX2zp0O
W4S7wpCExvs9yPi4RFAKBcpaqLmYwiSbEFKNC7qH3vYz3XUaMHI9VX4Sze/VFwXz
/aj3b/UBauTYHcrI+NKzkcZZQxkhTD4GW+AAbqemOs+Vc92wF5+5ZRgQHT1PtPjc
RqRjwEpCvlm+unwM72PyeSN63RJQ5+ZQVhwvrgZeKMKS8qQiWmpXbUL2BEs8jw6n
CbRMf2wkCuYMcxD4u+Xv3Ub6pec/lpMmdfaSmCQ5TJvOFgCdCwI/sLeQcVZxjozo
7xz7l/RxG/Pbay8irr8B5aEATcDjvpRpp/sQujRH73m+M4NUIVZgTxvXhX2GHtsU
bqZQtxG2I3oOWgaJvWC5ipOynxfGwmd21YSesVo4rvLuezMbTaZTRWbxYpOD4JBo
Ol8ynPadXBN2RHywLLyXUD2lRZp+e7udPruBKHXU0yGSw4kOQz147O5/8qdWWycD
HgWLEU3e6IvOLxOBELFK1LZGDPHw6SzsKaA5B7DFnKtbqwuj7gIxXZNq9ptPfjTV
xRTXGQjB/WZx0og+r2cbuYn5YSKTZSMPGSuOhhZ2a9VRdsNIDBTyJHUVRtxJpFd+
EttOtKY8pJP0xefkD/CMT57m3v4rdCT5kB8V9gKNZzO+a7bemeniTF8RWptXTusR
Xj73GRmqNm/hOSb0LOJLR0Lgb/5r4ee7b5BJGDC9wyEmGFm8K66Pfkru76DqPJ3y
fBX+16VtuwWTITIP5rvSFH0M95GBlQcGreHgo5NVhad39F6oiQyncU16EOor2/Tu
abKMzqPshqGSKkfbwhIfyhr++VTVQu6YzPjssZHG65n5NvoX3RWdiVNY4TvVHrg8
VibZiT40YHAwkl2+p2Dnb9gjjzUP6DaOCzXlc8WsgTXu7otELbbQQqRgL++dfW4Y
petxKqSB6Fsi2BwJukmcr8fTOMGK5yD6CI3T/yUi5z1xuWYBD06jsawJ3kC5cFQm
i1rmIAO813lymIINAkAwb1Dt8CPjqUm0MMilovqWoGSfITg0Zfjf4ohLgewX2M1d
Nv1JROWbrswwPrCZNSs8QcRDwNxAs7wgK14plkOlw7VkDjYYrLHb88z+mCZQQOiH
13FfyvYtY9RUpYIENnxLZdZEFJ9VpmaVO5Dn677/fi7RagOIwOlFJVtCY3aJ54op
H//SG7KFvGvN2xc1NXdHhIggwwzXGO19LjMiPjIwt43Fi0V4/+SDRhVX/DHP/wtE
uK5G8EUIDO1n2XeGyA3T4kDSr2I3ZOh1T+Mkm1hM6anGQ4TiH0GqRDIJnp9WnDdb
tYtqtRlvfRI3muJEkDFQPOF1es3tQHJAXHuDsoIaol78u2AERseA3DLxdxag1xWq
fyy30UTkBRqgITRElJO4Qf+HXZhcZjkP+Gjhrj3xNB4ehvv7WQVigV1/YIwZQI47
mlY+ik/gGTJQ7VZ+j7oizB/D9VxApKcsY9eRwM7kmlGH8vpGro2Du8BGWbyqMAOA
7Ts3ekbGISQTy2pAszN180vXX+R7UBpq4QE13e70Uy5V40XX0NXKbZSKak6Rs85D
mSfZNH80Bs9AVUQiLqpIZUm8nssRyN56B3jwYRnG4SShZeab69mweYpvupj+afww
KGJsgnXTa+RmnqSZhHTDKBgaieBvSBGQOhjTn2K6OoMIE3cOYCSYpgCHPfCUTuoG
PbIg9dnK9jSz36mhLOpiKP9BTgM8gjgtDifhAMSQ8vAiwGzfnKHSkcOdVzaOv/CN
AUeD66b9TsrzvKL45wddLNu3yA7NckYV312s8pV97mv3MyFrILbqYm/ELH9zoRWO
tzK1i4Rnzm1FZSy/R0CknRdxrX2RVrHlmiRT1bXh8QNcHZNSGS0CsmRsJ0XcTplx
Kx2mkb6EjM514yTP2xzdq6z4RDaP1pJNfwzxpp2CN/M+bidI/FU2WRw8/FspF6Tl
/H10K7Wia6w35py9udam4N0FGSdAghbtwraSm7C1Is5KziJ/V0bNZhX729PKcbNL
nNy7VsbRe4+vw8DsffwW9gfNophiCd2SMNb7ymiPXlKh9fHyJhUhg/yID9X7RoMt
jHfXLNb8tW4mGbAcQNxC/PZi069G/Fjbu22ZcNQBCIG7amDDlcfyQ4BMjk4XopIP
63AY/17pDaDvnMdNcRQz5lowXDLApZjZHkOqLCnSQPAnyB8ItX5mloT+DYyyj72g
k7RWM3t83nnA/TW+jeSOuakbLXpz7eCaOVATiO/NzhCql141YSQA5AEy6e5NBPcv
hMdcy/V4NX3v+55dB9tH6Bs4wQUoehRUhHSY4rtEnEQmqAPo6Z6M2lQFqoMTv8FY
VoCtihRHlW+zAHgeJssXAd7q/zWRVAeXdxAPbusKi03BWI7UXdV7LlhVrfWPU6sV
dqGT6tqDDK0hyk1jvpud4zcktyUPJs61pHOcJQRXjjjW+nCy1onQwD2Oi5ZtQ6SX
e5UMuZNM1WnaJzKjS7x060LtQ2Xhsa7vK85rsrcInBgun2YJSKrEv/tuWU7sRTV5
hgZC29NJWt+mRxvewxYv/3b8AVcfYXZAe8SERhDMzRRIPf11c5by59ekhhv9CTv0
rqgyT4hc+F0rFxD18ejeJkouTiB7hOg/DmBXPYVwDgGXYQ7FbkzuUW8qQhwi1cJ+
Msn/vKBriHcTw4QKHc+I7733Jl0/pjZxHDJdjeb4Qgt9EtjdN05pTQ+E/d4JIgSZ
HhB85PI4MmebMTGzoVDYRSTlR/D9RwtJOOMb/qb573DX+8XkUYKsOAjLft5lypbV
xO1veGcu0yA9EC2rdXHSKMMkCAQLZDddtk9A+XQeDyxByMjCdcdWgTYbcJzf2Qag
0Br0DW25qZRONeJTLloyJlU+ZXYOCP6UNuwoDGAFYHh+yhDhbYLfkcJVkuhAXhue
6GZTpuQf6HYvctBBpOY1WPWIjvfO0Kxdgf7DEXaUuRgChp2gHRLDhESYXT1exQXW
mAKwt3nDYaYADtcUpDhtcERm/WQA+oUCFXVm4PIAYXTRc8AASVWGoSlTYbopWBR5
oy5iEKeEA7qy+Suiwl5ZTDccuf2e+o9OwiWAuF/Shf/rUaSw/MBAC8L4E9OpcW3u
p6b7F3HvEPTyvwhXjTQO3pIufumxGs96oVap8s0pA0K7v4hi2GtJUiPXjFu/BawY
Zlh8WVVxDWLPeGdjVEhnBaYyl60/C1hXGwHYv2C+4fCbgPaOTpRH1sGls8/9lbzR
ecvKekH24s1xNQ4voKitfEDEI2iLeG5L4ViYmpcbU3jsENlXVGUvmWm/VaYJTvEA
/VIl71J5bS4Poq7GopZjVL3pyZ4OIsZKaIulTPQxM56ZGajSwUbtlLk8FfEDMgKx
ZtZONV4iL8LezT5HkLBRsufS9Rr6fHECtSlm21WevNm8v64jcSmDC9RpRGUUl7NV
mYf4b8+cpUOTqWhZohfTUhOUNf56IG3h4d37pGBAns2kfcLSmOOX3DJemUKURoXZ
6Dwd3Z4Dm80Y6EgRnPBClBFa4o2NliWkdec4KvZKa2DqhN5wGoPnP5WsJf8ZGzdC
d6aEzj3R+vD5zVj6N2ePQ5Mdiq3iwkh9+t2a+AlBmcKeQUkQcT3kL6NTR6beHX4q
kfnPkPZOE05NblbP6stkzIG9LCx4x2i0TtgSZyxu1+PGEycHsVB5t6lo47JXLtt6
XaCM5mxZvV+zI80hhEQOCUEEfbyN+k/Ph1wuZhxpTBEGvfola4rBJcMryu0kUQzb
w8Gtlyqt8poXX2hmHMWJDnqNBuxWSg9vtrYRHOheFLXym9kG5QaIHUgMCN/MAGVb
3qsDDZdrTZaxxSXtO00uO7AejqtidSl24dQWOspkeWiBhgozaOQN+JYsKPA8Hbji
OoQXUbzSaikBh4xGnkM0V2VKXvSwpprgsZQijKDap7l8pSIENOfUf9LvLsA/oNj5
ZrjHq+wV+Hj6XJTfAQMtZqJ+F+YxilfPHGhaTKPHXII+p5QIk0/b48Xy7lBkLHX1
qYYTuLVeADkDy3/H5dOtouHly3oj9Z/Dv17MOqEMNwSoTucjuUfzd2HCBreaAbER
Up1OdNZIKI8hoqtach7YaHNdN6EGE83ZuZm2VVUZvBMd6TZkyW/RQtNOQdNNuYka
sHUMeL3JnqlGMuQ1XigO+GXUubB6xjBZlviqnmOuPlmJq+lOBvq+Daj/LmpABDzg
mXD8eBu1cA8Oly54ckazcCfu49G7tqXMwUckBMpfGaCIqdBu6TewlOaE0tb7cap6
qPCcgpNJdujnnvKjzrh/5EYUi/4ezmYu23AgItrvKt3DuAP7M2N2KxH6c6AnY+0Q
eQPVceyEJWxVlbNxw2U/JJczbONnirO8CrXgSyFCVKykSDaxx3ZA2rlXu0bqdbql
AIAt5DG0IVA7mVd9+ViOXdNkx4ayMK04yi7TRtnDHu4kbhI+Ea6nWK4BnaXcK3f5
xsohkPYcF95hqiuLlzpPgKS3KXIvKsl0dhZzaNQFCErJwbu+tU1dOzbMIwOsjfCP
2aSMmkng7ExG/KEi9UQz+KzxrZ2Un8bex4LhUu+yD42KKHMNfr6fQlz6xYA6kYme
FAZG1rqrS4wjFMmsrkgX1ZIGUcUTfGjMSmSVgVRq6XMYZyx9stkhZKjhoT/Nio96
q0lio55rp9F4KREVa7GxWBrAjP1l6a6sL01R3EZolqXiIltW7Tv0CwAJucUydanE
xFpsfSJPJzbcWXSD4EVg6hFZAUmLQYPW+y/qM1zc1uGZXRV/viG7Fsh564lB9l/b
TjrmMGJZ9/m19J20Bp+6ehzpWw0z9bScHUsg+AL8azBuBaZZ6HHNtRO+hnzmhegH
dtqiIkY8Fu9csyy0hrPmwDb5RJGtqsZ5NghpnZdF4GoBSTJB6S6Nj0dgu3D1HZdr
FFh8a+futv6OAw4DZTQ3okACJOClR5KMGZM9th+w6AGybvxqCY3ODmr1TC8kpQ9Y
JlXDXIs/0m36DjM4H5dIxt7du7XqBHiszrTGbJfqFgMtXHr5O91sD7/Hz49/8/QR
9Vlb9GZq3DklCYEdQ+H9Z0Lw8Jhp1HV9QvQp1P05LVLQiTUvVtDgN8qMzeN0uloA
QWzYPFTKoxFh3/K2FeEj0cYg44fvxrx6kXoerv6keiKF2lcd0DlsKqIV17NwswDY
ncgZKd9hqTaLVnL16MLgAX0KO8yGkX8HlHT5BTteOkf6QhuvEanmPRyeSrqRD0Hg
uutrSl5kBFxhukfJ3rp+khTwJy5oOYqCWQNWFAxHgSKULK0VuEPOpOUuHzYwQDfd
0RsTHNPaQ4TH9N7ivNGmMxf6fZzLlTYrZ8uLrj+oP+bGH0YvZd8ztR23UWfozqV8
TnGuO4wj9OpwwitCL5WppUK+h97OWD+Br8p/ZRsifzNxI81RMVsHHPwY0nGHepWD
KD30K5jlYPrEXZjtaU0zHWBQ8ACuvmXIULv1SDn+8NrQJDXvtBpnLxZE3WyR81Md
ek7PvEhKJ1pMKTWXAcW+grD/J9ZX2EMqFQJThA6BK7s9G65U3IWm2Dv/yuVLq1p7
iqm0t5zwXPuZEjxpviKrwSNNVD9d/Gw2777Uv45eoXjBXHQ45G3j5ANUSZlyG++r
HPY4FecI9KaLu7Rh7H0SId0ESCnFK29dWSmnl7WqW7WN0Qfl+Tz/aUxK8sPCLKa5
DTapKxSkZJaoQegy2nbKv7ypA+vf1jrc+l0K3nTVjhKThZ3n9QU8FSt0cOaIBn0K
7yPbZLs5UQDMTfjpHGOMm4GHP9JmQHoGxRyiXEBFGt3G5QGkmSVbNwZCMMzrffI4
4SnBcRpFbBalEYh4+V7T7fNOA0WitSIKwPNbSRSdsVn7bw5o5pj+BHBpyYl+zljm
KnfRXSuCry0lpHJ4R/ZOF8ZnKs+842bwCqfoqy+3V+I1zhxDV55kk2mXzEJeW1ut
mDMvTAWO2xZyiXFrXWHWoTUadXnkTPBVSdN9dWKMN0P6Mqocbjuj01t9QfXpdTgg
X+r92bzzKR0htA+a4/4muZJ5rzNciqfp3lYQltN7j8Nw9jXqLFfVlbxxoc/Jh2AF
zfijIPNiskP6Ge1BEB1A8Ve9KYq0i14plIFl5+MyNr6ixJqaqejhVLOgWANRjISt
vf3lYwlMvgB6rsa9AHtaWs8l14LzI7tITLeluIcGH+P30iuc1UXAtkPLjIdSJe2M
5+4hjmqgczE2iLW8FpJ4zVcwNgX434k+auxo5mxuaFE92DHFYvR5KQ+JHnZNj5RL
MwM7qjQSI0JB/xGe8b7xLWnB5a8xgjizIjD5ZDCEbQMSU18TfNeSh6Z5aRmCtf+8
atm+nbACmKbJxU+uSPiNwJLVcCXmrD1bxrgxcTvwfOvXmkSst706sYRu4HS2DATN
lV89Vz1Po0u6/gSy8KvTxt0RFQfYp47V34eaA1NQlEOOMQZ0d+AA30CbnxzokRYi
z9JBzph2iGyBWov8o8vy5Nmx6RVLxnrCsN/my7V8VDIVMCn+bJnDds+DkmMQ3Fmj
IRvYUCPkAas92oXBenoSo/fpEn1PBw3SED+h6r1eCrnxHARRpq8Xsx+xlsuLb4Gj
VnzI8fxO6eq1yjpoDJNGMrT9qjYA2s6rjmCLbXMa/AKyc//3erqJCv8LuXt+qoGW
4M0pfNqHVFLoCccBpZGSPz0p9uzYqsx6AFQnr81H9icKC/NKoz1OVRol8A5CEvmC
aahSSCZyzRIor5FQ1epyaemzZG5FUvaVThX6BBJtnLItT+I1/5FkW7O8/dK/nIUj
THMBDTE4YJ7GHnMREtyiXAueYo7G7g9WssBT/2xszFFhu1lDqdQUBxMQ7/YTIw6x
f9HfQQsOdtBjuur79OEamgBmNwIE6DlfNkFv2OA3wdGuZfwrmhyIIjc7LUo6l2P2
FK/Bufstq/584/GXFQPP5bY2ZtZNMhqoz/9uWWdrxVXvol0klzJLdBimeVDIYW5D
b1mPJt1VBrG5xBqifrR14FWa8ukYlebxVpURfdQa3HzARJFdry+yph2N/SsHZs7J
Ey0Hv4IjM1XxMxwjFIzks9rCtWnEm+Z1T9LC0DpnukrZxz9V6ltTQArMAAayV2iG
TVh6qCZwT6T+iLtn+H9dyRuVU0qHj8QCW3gfa5/9hkPsysL9babxXCwAw+oDDYsx
jDD3Nr0NkNoK9qxuKLNRgGMdnvPujZPk2r1+Avr2Og8B2JpiLdnmdxYxEinYftPc
YpkRW2gAmXdEq4Ovt0jTc9XsI+rTtksBot3J1dpTfcwxXG5mlVy4+9QatvQ2XSk+
t+snUgYxoErfWcZ5xHQpwcYSzGnzmXNbFNxpTxcdGpSNUOTq6fmF27jmMM63Cx21
ALlVswVeUssEExsfKjQgV/L7hGBhiuveEzKUC8V751RAXt633WwAqLlVMIdTYBf9
gqvxjL0ICr3t3M07EGv5TgC1NNL4xkwj+kJ+3o7NanoK3d+oReuKaMIE7R6Ay8wy
8DRDQDRnbIwR7WRUHxaXWbMakCN4O4C87EQ9dhJNO7ngQFyH/wEIhCsv/AFcF+mW
3aA8mG0HCU+sPKr1lU2+uVggn9hU4A+qzNB9SMnZg3/Ooei5TAW0sid0wDXuvncd
+slOivs3938Z15Q60wvpybM9zCSueygRrys+R8InBnX55A792xUOvIA5mCwqjr3V
azc+gKI5FrFIcssNYlWDqIFCm8KVtq0LfPo+hN9ftczIVop1Thc4dtJ9M+YY9/DE
sf9n+6W0czkDDni+e7XFMWzczepm7sCJFCQtxnPE5RuP4BXi9rf5gw0AYjNJUlu4
i6mX9YJFLo2x+KujfZKDW9S5GkAMnrby/EI49YLHITAJzxD/NSpRgMD0u9o7NhRo
Ql47GMph52iGZB6vC0bRta8jF+BUCBDnVSeRCSXe8w/spkOcqxVA03cm/Peq+ehK
JmUJhoXaZwSjW3YW0/DmIYX2fDfZ0iHf4bup1dvL5uwhd/+txJWOL2Jz3XGuJSRs
Uz8P7c9TF4TD0YCYZG6HZ+HbSX8GWp7vOVyRS8Zs/txpM2tb91ZO4Qbay1KlXYOt
veA8Ad/5hWe8eO6yjgTvCJKNB3skze9dGsrVYiqiMWarUXCwOKZhfxKBdgRlVI3h
eo6tGs+JwMDJQTvkxYO6wzIJVk/Lk/LgzIpKpQNT5jHgg25KgjNvQdb7j2zIQvVc
vwXA4c0dfZtcxPfeNJFLXi9wK73Y5L608emhtG8dct33igJvf3WULko1YgQyMOM+
wq7b4IeUa17HWX/PxTtv8M4NYF3FEt5zRdYaaR4ZQjCNMsOk1EeTIahtqhtlmiwS
O0cSh/ZuOcgKNlfkU8Qz4IvmLLqHjyzWthLXxaDlp5HrYvaZkYvvIRUBYnWlbQDc
8q2n28tsYt3AN2cGMtsbt5ahx+TYlyCLx0PgfWypYKNDuFzRxGATnEGkTQjczkTA
997bp5wKQ0NlYE+1J4OPT5DnyTHwhie+hYfT5rXv0OFMItHmjVh2wTt1FLNJBBj9
6GgVfzQTPIbJ/mIJikQ3beMJFLqhgL8ljpKlkO4HSb6QJtWnh8QB7lNzKCinG4O3
94BvZ5XO7TZYuddLvjWZB16S9N5r82Uj87KSqYfXfJmTlnxwDvztvjW+lOOFQsc0
ep/K/4a2je2z9nnR8YFhvGd7YdcCShB32wCp5EokGC3zA9ICKbFVDbqUtVd5upGb
f5tUUPV9/qD5EjmoEs8CNr9UX8T8VacHqOjpcj5jl0CXupclHvMJgsHY9nqbmYcQ
++io5uW6S4zAtd+TdkvrvdjekHOEMjencW+fuTGrcosueyu+yafeqbKIz3FRNx7g
EkNpUPQJaENIpC0sh5CZH72ncwrh0eSq8PPGHwV4oRd/vGiWfJ8luKvMxG6hESpd
pZ3qe+MoZdf2KHZ9Xp7H45Xs10NdwckS3znyty54UAeizebX3XIhgW2fcuOIcqY0
S9/rgXQaOYXrwxLVkGYoH4wDy9QoWds9ZlPVxr9yUyHsZrBTp85W4MXphBHsRhEq
TTFaQSOY21GpyKC7Tt6m5ecLN80oMoYLWavUJQTA7fP93rIFFfqdb6SuIYNdZnjS
ExDbsaQXLHheZVzuLZ23Rkenvhnj2iVDfCDVoacMSGfTteeolSONZoCHgRNtj9YT
mYCnrEljJc0usr+BaasfZpadeWKfuqQyHHWqtZ+8gRdBmevj+KedxkCrRgWmoCv/
BMXkJ165LnnoGJoQWoQT+ODBud+gFK72SONS0S4Ypim1uh8fjthVD0vHQqt08uvF
UUxLYmrgJinuaeeAxV9Mmg==
--pragma protect end_data_block
--pragma protect digest_block
E+7SyZlnToQc9yWMph5nNtR32e4=
--pragma protect end_digest_block
--pragma protect end_protected
