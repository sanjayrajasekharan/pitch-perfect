-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
GYxm3Ok0FtVDsGZj9KjhY7IRI5qqNIhtOsMGlECRVaIGsVZcWVNYjxYf4tzBoXrU
20oYGyJZImBSvo03C3LZ/MBcqL6Tr1T3iUw770ZaiNRT/f79HUTLSmfUdbu4DANs
ExpdnPYgQqZkUYkurSmTAVlEaqhzCgRk1XNCiIBMOmw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 28016)
`protect data_block
Xm58iXcult4ygII/bjyxkCGt6accvBgNBi76NR2o+t0IxYMTuliq/nTyvGr4rWDU
4K8kXGmJNLQYFoSgq0DA2Pd80inI9OZwgiuAyqkfHBCZdO310wv4mXoNSbD5Ck6s
KMLrwjUuDwHF0eMGLQJ2GhGe3EPfu1miWxzSqJpR5pEpFJXYnmBTBk9WjEwytrSi
94ZQxpY6UgUXtu/tE0DeK4FHBy5p0fibhk3AKMDJx3jag7+Hm3E5XmxORx2LKOYN
yPAUbEpVQTGI3WEAdOrFI5+BMu4AS5RSEizCkHVX0AfxH2pNrwVQddQx30NS2fmw
svpiW0UB76vSwSZT0LkU7hL2Lw6TXlVxME32Vnz+8eSSnz5QviUO6HjVns1Sq78f
guEkX2P8l5/VW/azxUN43pxmxIFZb7fWuAJy6Aqpwr2KvUHi6o9j9kWpxqD9mxZs
XRgwrI/WfzA0RMhhc8vPOe7HgcABsWMg7XMhEZH2V5B8ch1H94K6C1hDtlFLP1S4
Qxb4vkocrtQXPOJIpvr//EdhdY/cPBPLSaTqF/sT/yn7avxTJ77nS6Jle6ydH0x7
1rAoxv/2xFk7GSlYCC9Jo/UWzg8joqaU+wPGw+ZQNMfHy9IncVxcWqHU0TDKoP+J
qdlTgKjTMOnhKX8a446x8XCeNdLiF1EYFbOIj3mZXQ0NCSNneD7vqZiKq7CUQqN+
CiQQxLUeTjOKCMlUTCLDUpR0JEJJdR/2GZy9Jy36766nkr9pdKoXvJj4hMPg+l1n
wnfQUje9ypjqZoiJDlHjk9zUMki9GTYe8cqhnETTSxG0HGepIHS/NGyMh5O9BJ2q
YIXvxtaAL4gTrvl/08zELcgANhdAwO4yBHIH9ThNWhnI46BT9WlYh0gQcomd6hSw
tCftm+lq1Hf4LnJ6/5Ee1LJMIY8ueq/lVuXqUscIEiWZlCqgTSzkR0JsXTNvKIAP
sFS3IHHP8Zb4HzS1YOdqfL2/YWyjye+FC1JBDoIzNG90xfI3dSpvkSBW46DyNGOw
A5LrjvyQIDxemmAOfDDlPfqyNLSgALzIlTL0jsHB7Ch9fBq5h5zTuX4GFWMrdy5W
kkNsvITraI0VARMzP/OLNA3qyGKpLcmIjobFggCC3Bqgf1Kq0MrMuwF8+V14Uu3s
/idtUwC4clQZh59Qi10G6ZpPFpFZjYxv9ck7xvXIymwh6UhSzSVnpHBjuNBoxTYe
QxQtXfBquBnwakyNtYLkukXQEvB4ydL0Dv1VtBmMvy7UbbsX5zHe/A/8eSuLgQvd
jsiFZGqkynnnUbFnaJqf2T+NRUzgXFWYduAfTU/fSI+zelfOwgqJ7YshKsFocDtB
nbvu5w/MNTOjz3hpxTtxYhVaC5/n80sVvjtv0CUIadJztKTsriV0+Bepqa8wmzGb
iquBHHAenrAVzV1ACBe65BpmbNf1nDTV53GCI6dk+VtSGbBiJkfqT1IIheI9cthu
zotD9fpgFVPr1/qO4a9UfHE4kgoUqYmuWh9hUe5MosZgZOlWqGrd25FtWyGeJuvz
pb/0B8MtHgdq6nHocj0zO6hUsCyYIWxmDIzKUXR1g3cag8QZ0AZ1+3xSSzB7j8FU
XV8X3BSRc9d01lR9Bfj1achKHrf1e/fqqk/W336F39N4olR8cIgpLvTZ1Oc1VnqD
MHWytUUYo2khU1K7eWm15A4+wTsZXR6y8UP4Ebjoy2HHFYMRz4EDU7z21Wrl6ATl
XYRPdweGiOtpYIX/TRRNN8cAJyUTjzmC4e8Z3ivmHqeNSVdPA0Q8yhYBoS+hPyLd
CNpgIMx8kX44tOz+hLxEZ3dbAoHmi/hoVmhvL6NH7aKD/pu7gOFdA5+a09ljTHNe
pyj6b+su3T7zREzQS9/J8476mN+6oYqd3JIFAzzN+gXrEs4lOLdpnb7IkGMfaY0D
x98xxAp65lgAIuf1a3oA8mzM/JG+fkMJVzBPfvssKJ6o7J2F7MFaPInhYs/lbrof
IAm1buq7BS5bfHFQ2+k5CxYYWl14hpoh1dfom+ygc2j071bMnV7lc8+go1GF7fcQ
6ElltuR0ENanhZdUDueNCBZcShF76wt32vf26Mf2dJSXxgNtI2PkF87sXeZA3tI2
1rDqxPtBZ2kt50zeDdnbfIlFQ+7xNAYd7oCOHR7Wtwp26iG4in1/iL/p+cvSCWIH
wkY/ppLd+/rQodruKdPw/RrKjXe7SKRNmpcM1AQGlUR9HcQumwyPtA9gySF0hEZV
dHHYLQYGgqr8ERWD/EnbUr2H69zi+FD0zw7d+TdBjk71hmQoqltUGHnZas4xWnof
NIhHpDIo38IDbWkTF9TUvJTg/+tDuoB++8xT93G4nHjhH4IMt9rRsF6Qp33DGO/a
9vDfGFAWIGNfbLR1alqoJ78HA6E2r8vj5r9VvIiTlLaAfiuLpe5yhVBscNFVHvaX
cSGcw7QJ0askdp/rg8JLavEMxoya0L16tFqpp5P17KIR7nMqpVh3czByLqOnVsU0
uFpSWyjyCtcxyV/j9ww5XgmKpoiDMtkFAqvkcdwO99yV7c2hF8zru6lFsMK2CDrz
LXJLJLZcCYLiqrZuzYpDCDWgJ6hzZgsZ7W6roA7g7C7JvEd8swIY2zzsWkWGF47I
+nf/V9dNg2h7HFXTIyTWFxn7gtvjRUQPeqNFX8AozFEHm8zoql5NfFNEvdTmhl5U
t0KCC+X4K4+qww2EGk6tL8pWiH7U6XduEDCK/m86BnOdTf+zNNVAMlppAEfiD2ig
adUylfKSY2I74M9z0ojLzUfAhpgIRINf7VNl1HNoMuaFpfUb57Ihzhfm9kApFTmf
xAq7PjF0SAN4ELgD1jUHZKzbsu6LHGNaUL0B7lSZ140UcqKe94xJ+v8WMre/QDaL
PEsXC8lC+4/ExBgx1m+1aKaMI5kJCRpQ9Sl2vVIdSn2sHakJVhV0RieG9dH/HR4f
+DYEVuDYYliHZyk9aWoZ7+ELeM2y2YQrq6u73GrfiV75+rCt13Sx4Vao86eXx7wp
+pQ/o54Hs7zKaLFicvERbHZwdGq/G0J0aqaVtmRWOomie8tRbT2cjC7ANIq6jmmN
XSFVuIwSuUG+9LJY+TuZ4npvtCWhAuUGwwNnlJunwKzlIx2GR6uWZEuNNNN4jMhn
7XNVqF5kcM53/DjKFfUu14cMSx+GQWe0BMWQZ2bKE3y7lBCxVspBwGkKk+Pw2OLK
q0bAvGVPm6ZzPL23GZ6ZNUHiLdKTWrsEnpbQRcLjvnn8NTv/IA02BPSLIOXqoLPF
Rbp741TSdsaZCsYLmTlGSdICUYWtducWWE/TJxpeJTcSQX0/WyIbI0m8znjf1xF/
6X0PM+LjnETpm4AMs6rTO/UFsVlc+kvWXYE5jaYy9KgK1vZTKypknNTAN2LIUilA
vWzRg4c5J8ekHPlYUbVjB4dAo6omT/w+c9nJ7ScmdU4o93RoMEoRV6UdWdkb2hgS
L9a23NCRV1AbZ2PvUHN8XYp+bb5nIlPl5mkQolta/YjGzRx1Nhj+yaho/6kqBDzH
NP4226CgwsNT4tyiKGqDI1WwCispfMS9HbDoQ+DPz4EwxYPB7h/vaJyvr3SrQJ/A
p18jvLBDNd3r3/PeMdFYIkAWyzCvTqCbeUq+/M6l8V51nQa5CDCp7UL2AYCHNqdn
fG1ASNKP8IX5Od0KA79a6gZ7/Q1DoAElt1GiUp2yxcSUPztbCbVWxy4koohp/h1R
vWxGPmJyo+ONP5xVp46+OVerFliT+OwG5D0xSmdJCW6+m/GQZKr3aKtFP+9+i4+s
3o8lvM46naviDGDWtswd3PBcYH3m8G3+9zlr5kt7uEBhexITI3Z3+fQv/iyrvDWu
72MRI0d943X5fM5cheTDZTu9fytYopDZmVmtrYKj+olXkYB+Hy0tVZTlNKpvHMdM
Hg0A1gljDfy4FDIJUqwdcZUzEX1EXPcVDwcAwOIwk6eIcqH/zMaHZy4eJh96K5e2
luxowmnefZgQkloMZ3yXBKKUXOSBPg84Q6FCSnslFwyPTKGklbP3ZVVxTyGtFUi9
mI7La31MzCSfeGy1lGhBe10sOVyCd1qRxj68d2o5GWdDFlqc989YmLTVbC8VWRIo
iKl2gsD9SB05PQ6ulmMGA9f9XE9Ont9Uu43aAKNwrpfV4HQumP9iglTOaq8hKT16
aM2hagpK0VgJWGzm7dE1+dINejlSbecwm/4gCLc8jQNoZcX1p4/2i4FFrDBiZ+q/
uDcIfHtyOd3zHFrP8ORwSWiIyQfdHreDovvKF+Lwp1rb/KqveYMprsrxIwu5eoz8
RC4nSQQL4ALX/r+GmCckVaj843A73CfPEZfgYdwNYi2/ExJL0fKqpHu3G0Finjhx
Iri1BlEYi/b/mFHGeQK3pU0UKkzQy+gNLJBexdSjeYzzttOU2xKatnTaA/b2RJHq
64iVcE/hQd2410qpfeLeBSmloZE6Rh/w0NaC+pnnlOtFIUQ07cMi+nV7svt1eGqT
c4ebaI52R9qTJCbuUKW1bsAs/zAi95mEHzARtwYxc4zHm39RBMXLH04FLJpSZabH
pIpLFBJceafkUFAP9Qtyfh8MQND7xTy9eXcOcGVfa7q3AN5XkysC4GONIoM6/UPM
YZ+N6OEZ/Aw4Iauhqha+as6/ElKvrfGBepRdkxteqO5aJ20V9OiWu77BdIKQhtZL
JBJM6Gr6Rf6ktsbwn1Hlxg4kRO1VEmjGyG6AEpkhazm/yynL74k6UdR5iCkpH8co
JlwNwjd7y0XGPr2L0w48MFVxP6EZAnruYVS5oF16AfJT8VpD32Ls+qEPKA8XfoYI
I4EUOvFN1Ww2nv7Q7KM9hLeZaRzHMr6Vx7nFTO6A2odkf2mmrxibRD0c7u21Ncdb
ILPuLjf2bY+BYQ/a7jv1nb45P0cNwr5AKBvt81aPWtNMOGpdo9NP7/+71rlasTmk
H6VeYN9873CVxwL+CBkv9UMrxjupg2oBMN2vkSCrTyJ2lyWmxGVp4B89KVkI1cX3
96RMwTmTDsf+7PO//L8J1kGgL5o8vwrInpdx2qU0LwOyLN46GYyoPiJ9TYlBeJVO
1ghhN3yGPI1t9BqCzYZmMDvW+bml8kkzztiOElZ+hwoFOwN0gsm7zsIKPGRVRLNC
ouYw0Tn/6eIk87w+07w34iLNbn82ECJSakIb07cZEavxFohPD6wqwwQWDAFejmyF
3hH8usggyi5vo5IuUMOga6/qz5RQA8Ef1jg9xMPpbEZs2pW76U0l+Vof9oiyHrMM
GGScNvVSCabTQUslxrlrsmKxQVarqd87RduS0SDlcF6XglX3MmXCucplRq8wW10U
H+TxLDK4wagA+Ehg8U2x+EfQ03f1HZo+o1/RAIjpTJ/0njkLkU4p0Oq6g74JXBt3
9IGriR5iyNBSkZxwJwF4YAQ08jINWiZMEbgIIMLf2OCZRka3JyWv8ArwBCqyN02d
TJA5/PL/G1siUBBJQ4R2YIXzT+hrnR0jofqw5NQ0pFdiwdbLtvOYt12FqUa6jCGr
GnufKL4X07LjrzjZiLoqhEJuNUg5ul3IqhqlvDbmD/eprVzO24TiGk8hm9oYZ1kq
DSIVvyTbx/x14NZIeXi7+LqI0wWR45NrXNuycuFY6ADnvM9TSKFA6HI+M6A24PLy
QuujqFgypI6vKIM1D+1CGJj6bK2hvmIHUUlVsbijDGhXWGVJ+mT8aHlEwS7m0P0k
/JZs9nlJfpUDlfSI92JxfU2uRiB4v2fd++Bf2nffXPpF2ZND5aIef4dD65lXpvTU
F6AXSJJaYjBNQkO6STeFo4F1rBebYdjJgEpB5aXtmzU5sKZalixhkT/6afSbeC51
EGb6atVaDk8p2iDjLEzzlJ+BJ3OW38IG5R3uOvS0nJItdFWNLN6HyA4H9ean5ssC
c8Gne+JEf6aAVIbXcZnP33bh37PqqesdrQwhvcn/1bvTmbkyPBN8jgkAWYUlI96c
2H20TKY0CNI8ssDgLEDUwQJzfI9rdC+m/z+NEw9LsXFZT+RQ2dG4n1WbVX2Yoi7J
UJ8HGFLr8TrFJwYNhaWr9uq9Z7FD0ehCK7FxY04IEMiZpTYcSKHbjNBNWAOLuzka
S2FdnNsYOmsBno/7VIA1mW0MQ/B2PDjLD3HPgVrLbKUkkCoCMtNBpB+Gh+xKNwwQ
O+GS396mv4lJWFd09yTuKf695RaNuLnbpxFEKGBuacEFooNLqz8wO5UBm+XHIuWH
isaRUsrRnuYVovN+nf5tO9MqPJ7B0JTCWWaOyXpZ5NrISFs0a0BSgDQ6XRoJnAuS
+99rgwSQ+bH3q8Ehl9XoZdYxuzIsDOYK33UfYsk5jscolgFUy4l9hcB/s8dkSNVv
eFyCIjCJFEBwK/kUJJJPorcmShJ9DEVFm2gs66SA7GPGLpIDWrd8vrZ5tJLzxLxK
gJGjarq5fXxKrLrHLJZrWGBfMgmm3y8iFYwnHuQNjM53pJGGt5y9uqICwgNrrP1r
i3G9YZnAIRWSZ+rcw65KKnDGLlM3oyB0TX97xxfLbrGDYxhB8UGymNhh4OfluRWf
tfkO8OuisZZC07TES+RZtMTrHJW9cToq7KvRB3METXawEbjUpBXDUgCe48XbqLmZ
OlC+6noyeAeqthoufvJ0ltYpWq/eKCqtLJecfqTvUV4prvUI7iN3WgroXo6AJMZv
z/j7glFYuRA3xhiIuH1KeNFXhiVFH9UwQX9+viQIE5N9QiIGyIMDPDOtAGx1OBYN
w8/zbIs3Wav3CJSz+NZx+hcFxo8FAOwiXBic/+lKx1aqli36UFlHbydHs05qACgW
qQqdG9zPeaS0jwM8lv8pUKWa0Ec8lMg1sA0M5jTe+rJ/NhkmxZ5hfjp9Glw71elN
M6n9tJcKVEcVSHsIJZqtc0aOfNqhsyswjVCdw2e3pMCAAv1WYDkmPhZyJnCMMmMQ
1yG346HktcS2ncbbtU76QMszlLirpAlmy1XkEMLupVIZ+879qB4NI4VJc8XiHegg
QZTCK5VVQJXJj/ejjKMTS/dU0N85BMv52jucEehlMnoLRt016wp6AldGM9i7Q13C
Ssh61sNHuf8D/5UMEBUZ2kdQRDOGGJe+GQQVfNZv+1O77HTnd7/ArCcga1LmivJY
rcgfixVJPn18ubYXEE3FU38wwxEGMXF473GsylrK35EmzlpHBULbHgW5jrPnpAOF
nJdW+KqOkgbwRaraLDli4s9bK8UizSzzVou6Wz6omfTG2EUKSp6NCmrG1s2dqDrx
wkNH/EqSDukpzVjTEpAQeEjw7BJth3S19mLh8pWJ5twz9M+S11ZHb0nRG/mybeHW
zcuQ42zLA6MWOT1uM3c1b/NPezFi4p+c3korywAACCNhv0j4tbWuyNsupUA19g17
FVb4aOFOjAnb0S/MUlO/m5e+Qs7gmcbV5Q829iYb27TakT6/UEMAwFAQNI1gS/0f
nmHeIqLJ7KxWrtptBOAonKF35acnGrrnD4bRVaqstTWWjEmBVuTJR9WaqAsYMKAo
qKNSfoSFzE5N92WQHvoWGREEKOoe0B2MQoZ55iG6ZsYH1axHxv/c/bnYH1aZEU9z
heQhfnj+burLU8spEFWkDFUdFRq8RTPrKYvM+0/3tCnV28DngcqZwaFA2GfxGMpA
aqjSqPoRnZOq4l0kEK/HYRcJSngT+LeVZFgqqKEH/VgHIAOE/ozjsnDX0lQ4Emb8
OKn4OeDshKOw2XyzB/QMbudTZj4b2AvOiRjtsYj+AhAuLeIDJWue0qjedXqP5zqG
nD3kM5A4E24UOJ4jjqLGhdI6+VIpwp52WLwC2cxPmJ3MK53KSS+ABxzpO0aNaKRy
bo/p8Vy3KhFUYwZtYRDLbzKznjMZQJk3RLfNAHvk42mtvD1niDOI3VdF33fZE0Lw
U5sebb8DLo/hZsW7eD9oAxhD/U0Gp60fbchz4rn/4AD8dEeZzCuRkRfEu74Kd0Xn
n2TubfagWRVjC8ccJes0IzjYHtYgT56ay+RpprddZWmCA8mNcTv7ifFLX1/usNlY
tJagxwR41OZTt+Aq20r38Blfe21GAiKpe7UpbdH+FZP40Y7JYEpsJ4tIEn6nJBVd
0ik/LzezxvqtQnIQU9NmfNZn5D6qQXqabz44mjrpGYmC+K5/h2mJWwvirg/cMwQA
m4rXEIsHP0Cl7l6nBPatVgojEEXqZSBVgiqnVvtFXLacZjJwvsfIGYwAOTi9djlF
Ia2YBI/n0Zo4O599aeFL3AvES5aNA20YUKIazbQfPovXRhGIylFHf/3l5a4p6gfa
ka1+siqlm7t7FnDjuPd7t1ohusSetjpFUhzB3JFUeFtpRVfvrr0qu1PJVZjImC50
PjpAWPQf+2uKrOggvX/lGgN4unwqgUBvGIGz+7ut4UMlQc4VhNBIVkn4rjTDp15w
6o2+RsAlPh76G+Z5TjztlDvS6npa/IACfNDjMrigUS9pnWsEvwc8M3Nm31uaHLFh
IkR813P9iF7dTgslztXZfyZ+TqgVPiZ9Wwx273s8ZyiN5XzX6gSvNChGSP9aZss1
uEKmW30QJg+5a5T+BPRE7lWSpHIjHCRkFukW6EeiZsdpJ9JUq8LzafO2O3NDofBP
wwFtanNRpAcfRSsPEzP2tRYe2RF28pw4zOdXxQYGS5SHAHN8BhkHjBal+vQUjj+w
jApyN72EeQBHwY5cuW6Ff/26z1UfeOC5aFzMsEzp+r1YAZ2CNoj56N7yltrVbnaP
cAcY4fo72OohifCDuZDuFD3doyzquQeCJS9s2JLhn6m5HV22zxqgiHXD51Z23hhj
43tTdrBAqbqnA8t7Tp4R23eQvq49OjgBJAaLc8Pwj6vv0vG9DqX2DvCH87Erk9uR
Zvv53hXuoTVQOHMjtbltie2HVWjXvw+LleB60b8GUsGM779y/EN136lBiVZhGdVu
NPyU1a+ADDOybPli3wupIWLXcaUgiqjMF6CHwh91pXbCSNg6oH5KCfasTTsVevKF
PVGh4mU6V55q0xV+yVoR2Voms3a+6dtP2eOFW+/fEN2d63+OpcvF2XajjmCZefyA
kjyf36MSsFilkfQgADmO0MN9FkmRO1RnxkUXSY4S19hSZDPGUQm0EgMdR5UkHOhA
0pnS0oshxs7+xbhFRAt06OSxFBKjrLvM8PLdV5QR861v7Md12mAkQiH9pylr2o8R
rzL+NJD90ygkAmvTEeD3xtVrC/Ejwg86nzYo3yMukdTOx3qHRnHvRB5R8pVmMyEO
lG8I3HRFIPe/eHm3GhFYhB0wO7AnuHYyKBOffDnttCAnKFGauIbxJZjwcz4EcfcM
fTeH5ziU1+4DRC2UAbALu7oZPz5Fq96iWRit8Qdm2+5fl3nZcDtD/ySNrmluxwm3
j3rZhx/DbkaHkZFGrrCA6rLBhZWkIU0/u29o53jsekd1mbvKz9nmXlSQ4V5V9BuO
jTINI4xXFnyR9CW4zPhUZAMB0vb4U2/mg8IaWoaCg8zdI6RgofhI+1XhBR2Eu73p
IHgF96XmWZFU/fOQ11Kx4jC/zXPO2HVXgCoCLQgOwpAos5GvuKyZ1iwvG+o3i0JJ
cC7+pDeStBAsYeceMpIBilpP7kciss4u6ko5oGLawGY8gfvxzmxm+7qQbDM1tLHR
Srnn1YzrPlWpxrzh2DU0KMgjfHfRryOMb/Kb9wfKp2jDLhtr8F0MlEowZK1Bti3t
ETfyF/rhRb2YuMuumB3CF/rOU+8gu936fll1w3wCfifyWlRn1sfvAmEiSj/5KqS5
72+fyCWE4RIZ8iKB9rc30pfkP3WEOeaZ5WzQUccyoGKuEE8xHbPeG9MJZ8UHl7Wr
Fas7eEGugh5qTIExph9UL4fy+8l5dZjCcJHPY5NgIwB57wMGQes5xQLseEkOq0YS
8xH6ZkdL3tt1CBpjvYxhflvP7dFRhsIK3HHhvDzHvZmSJ6YwwhR0EQ+lL+AXzkQ0
7XfAjo27aWlXnxp7/Mo/YM+3MCce1RHuH+VW72f7tGbldx5qg+j2BKaGfkI1n2j/
V0WHdHDLyYbkH5HWM+LTpvo2F82RuasgI3SNXjNIvoRxxHCHhMGiIFzOa0LE36wH
s/NAISQhJXPILRqgrjiu8QnlmBbB1XNLERQ3fj6RdBL/Cq9QiCFTGpKZteCOdtje
+CnDEvOCknWRpFlz9WmRQGb4/FAS5jf1ssdu6/d5gYsRj7awd7oX9gaKM81g3T7L
zOjHrtEkGBFyAiPrPH+kTTwzsuEte2GDO7lHho7LHCTh6v0pPWyLRP944+79QWpn
uU4Vd4oJBHt/vpouUknLWL8Bk0VsplBhc3LbYal0ezg21OqbMJujJJLfxQ2PK4qh
Qlu7zKx8pehml6t8IhOYJwoaYk9y+4Z9zVJOBMIYQ2s24buOjzYSgNfC63Si8W9i
4H+TAYGcwH5h2sEcPMEt2Etx2EDtliVOy+TIBqCXrrXL4+F7ayu984Z4t7PcKPGy
S8IoIRIViQfmqTampGaMAvJt/UZwzG50Ox1RpE8tEyTNGxcJ1laZ6H4XJJzs+Sow
xnZBRJQpDGcRAaUBrapTO+gCMNkwYIU6q1UJlYm+vRG3r0ZHungxUTqtRyydF6Mi
7iBSr66MFZU44RDOePzmu/sD0Dq5+Ea+jTS/P0jkKzZqUphpzy7+hvilMmR9ctfw
W7VvBlekZYmgyADZzOzTeOiAdS7jgOrEg07vRZ9hyEIkEDwgHngA/BLkH7HaTiM7
OC4xSVlYvAydTISyFRBbwTpkVU8M1iu1nLK6LP+lHUh+NC/JNFNR47qe6aKUuUmi
Z/6rygu+23b4EKyBkrPGDuGA3J/zLRRBePmy/OWnQiHVmd8mNsD99XPPo89kjmWX
0Sh3JsZwWdZd1T7wX9IXVpfPu2uaciyB5LfOcEtj+CEY7o9KRMiLI7W7wK8ZKebh
EX31mjoY8a1BShqEtJ3VjjYf0cTxjYFSpX9H6iv2oq4U6q7N3cVTU3Yn1oTqdf7X
eSbwkCgLUTigmF9QUos5WMOYWD8PHSRSD43ckpiscr1kLB2EclmKqH/qudkl6uXQ
5E+Ntf5hebW1VbaSPymPvngnV+QCa4AgE0LHqD0b+s2iT5C8LoGwrHlfKWGg1OOv
p1Epg1p7wF/8Xh+SSljiqjmvdh1TPn7/Ex4v5NrV8myzzIltA7vPOt6uQzvCVyj/
JfAKPuwZfPCIea5RYgNqAvCRwdfvcSbFgxPGhaloYGInuFqpADGBB9JPG1dxxeJw
oZ2NmTVByqC7MaqcGpVckImnvxlkydnqYpxDUjwOUO+nkvd0Cm5ZzNTUaAN3Otcj
1VNCAyTzlLs8Lr/WWOcGkwgxLe0cL0sLESkTyBvht0f1UmgCF/YDtkU4QPh/nDYN
JC7j0S5s/uzc40/KQPZhA7QMInOUZZTxDGC9CjQzjins7tdJbiynJcCJ1A269Wfv
fKUHtzs5qcf+ttTJ2hdzPCxwEVM5KNqmx47NxTF5nhDTVQt2+Cd+3XIX9qZuphmQ
s2aofM7kLVGGdFWX7JKe1+nqc3ATjq9x1vgBoE7ELZT71Dx70UYUXaYpV3SJNu0D
TNG2RYFVW5WwHs6Z1BRjzbxCFHqvzEi/li4areEdMMGWOzJbS4EedH3fGv5NIbD/
CWrHdfo4Xng2O5uAcISuFXvN0+vunNsk5k9jYUw/26m+Cnh3edOlL4ge47HbDglm
PnUe9B6ThSlTA5WT2x+5KjSCJ6uGZ2Ce/5gDReCxHeAZvzjGkcINeuyQBRYu9rmq
Hw+pRLZNrGodLsFuRgU92J+DhzGt3lCiEgoImUf+AJGMPjCrZ8ylNtPubgAT8tYW
i9YwE3yIIrmQyHW1FNPapiMajKScVUb2TKnkL19icQMVTRVKW1h/sWNWie9M2BX2
tr4yPJ8MOgEVb0uqcE25G6ywX7JP0+fxaQHT+wJ4xP083/FPW7KgErUpgGHN1pRC
h3QWefelD2Kw+LrjxXYkspZqsyZUOv2d3mzfL1z2aW8j1HeEnnj0zm3KVfrRj93R
lp6psEwxG00eWygeSFcZmHdlTG0pumJ++xBSylJ81/+W80hnxSPAv5SojS5VIVCf
4QBdmS2hTdCr/K9TIyiHiqDxKAzah5t/RZUNpR9tq4CupzZawFhlmhcwYsmLRG0T
fW+26kJpEoFaYORY3IwAZm9mojwweuEe6OPhRg5UmAnFOyx3gaRMwNTyZX20fJg4
L/w90EbprznCEO738fwk6kMs8tIFnk3cw8qbr8OgnUT6K4EoUHWqEnwccgpJMGJ4
FqCD/LQ9zCxJXTC8l1tv+M8RZJmjncCFqan4IuOVLWCRzlokSm29l9Odl4s0qnwv
fhBVN/x303BTe7PxAKr+nkIJVarMA3XA/To/H3Orpo+f+f/CET8aziSkHvcrMZdU
i0jVRlisHKvk0D0lHYOA17RhbQE1JL3aVHKMa8ae7zysgGzOYlnpJICsaTgdw+aj
tgzVTk8SHWw4lUa2j40OvZU8vTI5JUgta4MOTfTV9B7PogeTH/n8oY9VOJU+Zmyl
q1n6vC/7IEWw//K1rJMvRg5AjtBcdPfSP89R5gHjUp+f7ue9lj5RefDA+p17Eycj
DBI80iNV64ai4Ats+NILm0yySF/aD/sqG2bPKyJJtupIO+++HnaZzGWcWGzpcCKQ
r7137LElSza3UiQm/Te9fItos+A0s7iIs3M6Ow6PNOFsnPCsMIyXhtDzpBf2KYaO
ZgyOhhiWXSAotYiflUtpTTP4vBCblYlkEphKdsPbmsv5SpBtGA0HurW8YjENN+og
ZvlyCdTq2NQm3FxzGXT1sVzv93QNLNBnzihb6w2L9NwQT8TxnSUctz0VIbgV0+yC
li2xbrGjFx88pHhvjqhzhK59Cr0zW5CqY4yGl/mAoA7HryyiZVt0KQAM2FcFtXyO
VJVbZOUc4Uq4DAMh9e9mdoLPZCqo7XEK7Fk0q2aqCLVN/B/82i34C90NIJOnpRru
iHSkSuTqmhkr2nDD72FlCzdvMSvmFQNad8Kb4O4S+Y/6JssfAJZanNe1KuzQTfKJ
wwT7QzmZyV+iYdZqockAcTSMK5SBox/vhH9rDrcxSUbwrt8XD5tvXt8v3PA4zonP
qH7D9YbtwfNnbPqNNAmbSoTpjr/I8wOxo9/GEZ2fnBKHZBBCmFAPZSuG01U6vYw5
H2sfy7x2QGOZZqe/n+7ToLZZwnkYNM+mGxrPug8jwqeeSiCC15bHgFFVzSmsk5jT
P091bOfjb5u9MIJCRm/aUfOOTzNU4oKLWOSVVANCUybnHLeoI1q2VoVSXVHWkrUp
WD0qnedj4EnVFeNFvZDLEYJuUB2187kEY5lrairjqS0z/6eV1y+flE8sPU7cO17G
OvDMBxBSyoOzHLDBR7XfWmGzYw49cmSXUxi6X1lyUCSnEs1bEoR0lZeYGrw8taRZ
GtzOFxXugwHttdF1UAywKdActwfOmqU6J0Jk50Bwt3qoMezoG6NXBKdCWZACbtBr
2IV0YhtBJhVkcboclQ3WLoE2yQbyS3oXvjUjTl40gLzTpFcpSujEwmuj2Hs0z9my
tmpEIm6qwUnvK/5yknGzH4yUaVV58coYqOxay4Iw7ZOLjHb1CcpOWvFlI2Y1f8Mh
lAT2vL4LUUkcUPyVgG8OkBJNMiHMLkHk/zlKwt5FGAyzUqyMzvQA6JchdsSpvftj
Ew0DB4yYSrgxdtO9+N71thf7AJdnD84JJMtfV81uil3uRsX3wl+sNQiMh6H6A1FU
BpBVMsLhsnGkn549YhZ4NJ1fJmViqmkEXqN16yR7S4NJQADgwaMMAg0tcAgOTzUL
kb/aILh7o/bJQLo0urolKD2wlYpeuxE3WKwzpAxC7eUF4C/CDHpIT/SAP8W6+n32
norfPpeTkxiLWxt4gXJpwvzUedoHCYVhMW0/r4QpY/lM22tKOR91IpoMlAWYPZia
OKDxHq7Ey09sBQ/1/ci7/yahkDTn+dKNiFDY7enIqx50u7OLldBqqZ9Ojh/h6/Gn
NdhEhDRmkmjug9JawxpEFG+TjzV3WKQkx8vV2N46CJEgVwaHcvAPbdEbSJqcYuM/
esnOIxoGwElp7F4CMfQu2DnVLuyCxzvrcD60BhDs/VEhaqLKOMfcqzeB2IpcXRDj
ac6UDLlF2+TH5VoGXwb5NO1BuJ1gpn6UE95wpMow0wNI3wLMmUuCpx9O1P46e84J
aJis0wcBhXxqIJRHLmkIVtpN6qFiDIocSH+sTa3+1dORHGe9iS0HJPnKegtwXNDy
cdQbGQUUdATOjGhzKShESyy09XiYvvEGanAukafco9euRKQJXAutWRlFhjF+Qunt
FtA+y6kiinl9D7+0YlE+YrrOfifX9bCQQ4VsVUABlGJYVGIs0asf+2Y16OHy9zwG
vZSHCmB+XOhV11mfQY6vubWdmzSLnnwZiQyVqPpd2uCS4WLlbvunM8bka4Y+8n3y
glaRrpAdj7VnSL/2+FdqblTdSF1jbcrGEfLl2IkHDHo7VMfZFp95DYtiLU707SNo
ipJB8y9FDZ2DMrhWQ4NS8ASADEwReAF3G+UXO6bZG4SaN/QdpKCQJt7NqQvdidmQ
1USMkjTdPkP4g80U7X3bxTvhV/fiKOUqXntoda2IE3KCKuYmNzk/Heq3R5U8RMwY
81LhSwL3lyYc4Azotf7AGREXJ0Mf3nwAyVtifqHG93IyIUKyP0K0l+xqoTtK428s
ZJX2te9KSJsRl1HXWoiuSY/uzv2Jw5uMlI9eSVf+jIlMZe+rCyOLIEAD8vIscs+C
dZe3YiC8FOezZgdAbHoW+f7h7tmSxbwBn8UCUTKdx0YyMlNfd4EioOJVyElyldML
MF1ExJetQoYeu2rc7gITfVVJK3ULMiUxWWMJuoU4Jfg0hTfGyKfOUhG5XqcIPsC7
XcNPh4EE+XKYVBxuEsLiE6AabF9NffPwwvtHrqiG2mNYY+5DCosRoxA6RS9yLdb2
KE7HuY4d6yQoMlroR9PcWF7lXPk5xkdX9zQ9KveJio7trNiix6hSXYVOOUAtoHsa
CmTq33y7pdRe6pfywio26g3iWgLOKzoDNVOguL6vLxfZ8u4JaPCpDqRKuJ/jFLF4
ow8aoRk8QE3fhp6JJw9ZlmWnn9vPfH2RjBZ1qU0L12ZjbToA1mny+mD3UtNfAV8I
o84LYLQ908z6yu49511DEkCZYBjDqchH/jzjeDYdZlTY/BBBvbGpk4hPE6Y/+Px2
EjwT9iHx/L9YRBbfqIE4E7aseK5gJXQIGKvS6yVOpwkjsvDtcqDHSf5F/8f0Msbb
cQN9WchHWTqqJKHe9HQ+/RjQs5Emzqf6HSeYVvB6mopq5RpLv4y62MGNKTI1f+MC
AE+44wGeJDR1qeaehpCMMRo/swJLtgR1tZnWNW43y41guCUKipDcK7Psuf6ALbnj
BBe4d8aqbKB66pty2d6j85l5G+2RONsQJmWOQWr9A/Gi6+D8UDAGaE5mRP0VJj5B
yWndCSCz5ztQGitDSJZVz/npf2mZD7xdEOpVaDpwJD/X7nMPW5wrCviOwwAtt/K/
+2+vpt5tpnUhHsfHqrDVIJXFg9C2P41Qp5Fi3ipU7KYc6r6Ltnoy+TmzGbGDl4ug
tzQtB2UVlLtUzNno9WSUnaLkB08FaQti+52/9uXQXogeOKCz1WC1TicvZ2gAAVM3
sjxx81QqGRScWGLgH9E6m/IJeYWX9vbLaSXqMOASuM0bfy5vjuMd8RCCMlCnaJMU
VON0gDgTAt5Xzw3sDDlik2xBkT5vtMjiW2sRju0M+VKPWQ02LnMh7o5wvMxh4Oui
9bklY+hTK27IScRtDcvM/DkZ1TnUHPeDm6UcDLOr/oZXKH9VWp9QZgfz+LA9VaeQ
s2O7v/B6LiB66IwiH/sV0CAD0021C3XnMDsQ2KhOmO8pt65ugg/p7aty5fVdW49S
DcI0wKcGcvo/a6vJVXdL+W/iVb+1nBv9B/0cUvdz1GQ8oO26b/uBLBIVg1/9y49j
FrGEn0m1LMytVPO/l5VIhUwwPmISEmHVw0f9vHO65IAi0yk5446dSVk/+9HXh4vL
L74JYZ8Y9OvzYz/Cz9QPaIBuDAPsRw6UCn639v7oEjd1gxFfpx3JCfsZBWk4zo3f
qiQlAFamSFxQrYCZK+yxXDYcupGfvhYJL49o2/5+kQ5ZhOS44CZ9+N049J2oWb34
061WCN3vwx/+2OS+U0B0PgmCXkcAAyFASIM17C4In88RVsfjcVyKrK3PiqTvoq/a
mc5FUQ4SyFp+zTLc4SIJVGuAX4ypJGy4jTZQyxHEy2VG9mD65BI6SD1zbEmIFMKv
BoSKhkQZ6H5OA9WQRyBTxFSyEVtjJBEYIZAElZrYpfD3KediRpPXcy38957YDQlS
ECK7vBhNT9ui2vHoDSs6Ihkft+0q0pB1INpJ7M8REz7VT5B0ZzhPH5FL6+mgcT+M
lOQu973y2EltOG0fTImOzXzeBC+GU8bClNXVK09w/xrK8jOdIep0d0884SZTzM2h
cPrsRNBJ4+1gLEZJIGmabgHYS4F+AZ3LXVqwLjpOw9zIeOKgQbpxyVc1vDDOSPPF
J3nJYaat/HC5EiGUM7o3xKgOm2iR34nU9ZI/irdR57F90aW8JDQJrrriqPHp8Uzb
S+yh2ESxpogj75DkZz+hoEfMDTL+Nw4zMu4mrxbO/n9gwQgh3Rp7WYpKyr14jM20
QDECtDC9VOO1c4Y+mW0Mev1jKofxCqnbKXwcjtNFEfdos6qyH4ZeXI03FFBceuFd
DIPcAHF63/qbEzTe2cW22RiPgPdc5Yz/IhKuLcBqZm0xLXR3guQvrAJyvi/RL+B5
7UpcV27BhLQl8FrddhWeq/JqMSKkjeNfxOESc3SsrG6LyWg5O4EX8vaQJWoIf51H
6UXsuvXVXHDPWas1KxATbY/KFYwlBSu2sQldobi/HgeGJHz7HkDN2Vr2wvNQBUhr
Vj2AX2BySsqLQvWMJ0WjypM2gBXc6q4Zu+bbu67mWhqfHuAZg4Cs3NrwyHhCQ1p9
nhNkhw+1V03AkB95W3qTUwPa4HOQBmIt+7sXckZAxeJtm2I8ji9XyjXdQJg7Qko2
VkTMUKC6cf0cLGItF2bNqrZ9uA01MuebesHzP53ETV16bi9MZgxPUGxsO4yCaAXi
SbuUVcRVs7yA9QEclEm5gQ1sw/MghcRzlcBp4bA4GltXIq1XkPs4EVTniyxh6VBv
3hotr8V0SEAsiPyHRqUp6eG2T3NTHVzas4HGxaFfzO71NtuIDQg1G17zv7jyaOEw
z3Rz6A43CCqXw6iJrYz9kzqWyUR+35P26khDcW+ZGZbl2Ir/oEpJzoV+wyvEE72z
hp5jR1VyQQt4AopiDjI1s2GR3KTCNuWLL5t9Q7qQhlT7iBFocHIOdFsB/StGNYe3
YBGjt2ZW4VThLN4GWpjtiJWAU0k8EKxSZONA+4Fiyr5PJdifYVlqDmYBuv0p7O7q
uRJmz+70L5Bj+K3vnP7XtrgjoQceLqzW4O3OP2K7ouZLjb7KrFwGbpKHl40lhxmU
k7pr/EFGQpUjPvaZbWo7ixsJhkH9pSihMMXOwPUmaogRhCfiMhSQIfkreF/7E3Ba
O4xeHEB7zSeBzTFtsktPhJ84v7180TfVE/r4x0M5G5X/FLQf+sW9S+EpuMc5QwDO
o51m+i4HOBpGvi5N1gIb/V8mu7QqUIqcptEEEWscovJCUPIHc4sdbwt9QiSmN4xJ
j+/TzFITEmAE7KtWgc2CXEiekkd1/Ge+TVTAoE1TH6pwJDpEfnGAcA237M9Mqw4W
EcEieIFQUnlIUFcpXOSils8sfY5XLOAodC8CyDRBeF6v78ZyduolSMshpz970EXV
wbAX4Sb5z9xNSylGeRAM3sWdxrhB3aBwnsbguO8DWq9j6jwlPG0hund9zIkD1kTM
IrAiQKrKRcNUjssFVC2VUHOuiCUEWX5zEz+xseM0gW436sWvResyfHtgoKZ+rTw/
MyIEGy+K6Km1feUS9Mvedgt6DZVqrp5PKWWrlgLMV0lSPpBmOUDFfNQq74fTMCVm
WHSkIEVcV9P/ITB9J/3Q2dMZw0N9uWNm34DcI7SqdiwQGbC7tclo2jXsFDIZFrcL
d7eoHDD75Lwk4ezFDwnC8vMZFa3TGKCzfEc/PlybNhyVByCL5h0xI4scUsFxqHuR
1YnqK9P9WOQ3oZAL/7skHAMxDNpHRQBC0YzECU/CIqHBpAUL8cLFJELdb63+2ChP
0AqRuYJD2Us+m4e0LmnnJvy7oYwzPqvbS4TJnDFbhfwmN8O+dtmGIQRSaGaCBQN4
Pd6PwFTZt843CxcXKvyah8VzNA9g+339R3EIhMtv0GKQQJEq6N+ZGApzASXIleAS
eI+g+UJpUytkgyeWHWLjiB9BbWQJGGb2HsJpY5Hm/bdbMdk5dkGGH4yD8mX4hFRp
HnjQQTmXVS2gw4/qLlb/hYGAMxK4f2laqx1WZ+v5P+h4CIzPdbQCjiGxjeeQge0h
lWTPvz16qTmUwSlijWAdIGZUCnkBcHcEfhQWrgBodhvjNavFisfugkts3ismRJFA
29EfSpmLTvBOCFTpQ75/h8Z/3BmqhEkAiOkYZjOsBuwpOORg/+0asFDfldpk3hzv
iE2wARYgObmCffHyx6oZjdEHMXiLBeidSU0uoIJAGz85KN76wDzQ5hlKD06pzNzl
ESuw3up3zI8kBzGByqu/cHyulX6tV1w49gmS1U9JSfrYRqypKo6QY7mErX8X6c9i
izcXpjC8q9MIQRqMnDuG4njD0/UUlp5I4SdObMcJG1DpsCyeHmvQs8kH4xZfLKLo
qECvJ9feKte94vB7VOKe4eS48tZE1092xi7ejRTBFG9eXehGxEIVlcEZSt6ddpap
+Z3H5TeK9OjiVMYONG/NzN7/+ihjVNxKkIsgrGRkkoHT3xw1LGrUvot9xnxsfwgH
qEhpZ8ifndVYu3Xfa1pgshpMp0zf5RsjaRR9RvO50qje47OgyxyvjIt9u0rlgSge
R5/iJ7jWSdsYWHHHXWdKZFtJ8minwDbLc4omsJ4UO3VeqYbxKamU0ce+9asjeHbY
2cZPSSwGb1qj8sKaPe61NF/6tt8wsHadlx+itOf5b/5oZev7b6SfthRXR8gqQZi/
k9fYb4wnrN7bvq+5XGIRbsRgKVpEax0myWdFfzhjiLIQifqGGlZ85MTtt2//bGGs
xelotxQi4ReLIZOH3TvAT8Wcp7rTwSV+dpESP8aBoLhHK85KwLmIAs6vClyz78yQ
DE6Dryr9Jxq33AFaKuDZjXjlnMfN1kqtGvEGGSuM/x6iZMIOgP+2ko1UKHTHc4Qh
BIutPLxiRwdYjThqwgNOL3DR7QThART0T2emhKWd+RHwLcYs4JAXJdIQWcXJBqwS
c0bGtAu6MXvwyBZ/LkT/2O2LBua4PlQmwmdw5FOIUE7TyicZ2ggTlWHSwA3/VDlm
SxJe3wfFIwZaCV8tF4Do1rMppLFYqYFBiNJ8M7g3CS/fEA0jyzyPCRUquW+qK4Cg
97ypQTCfHWAwyP7s6BzR0hjclEkA6WSrgg3PvCNaK8CiHC32uolYcS8QAst12PyK
AzpyLO95r7fP6tbuKnj9oeqAVX6/Q+vthnXVTrsl72F9CDuooZWkO+8cd/n2L9pH
tVMz1Y3RA7CsCXTFnhFStx7/raZD8ydUJqDIqMBpG1kuQVd56bcy9B1miGcoe20y
BMO1bICg1YmXQz9kjZIe9hrWgsct/TXhejs3/QCgXzXMJUUHlUSlLxHMRgV21feG
ooBeMjrTkwVm6/x9reeXBQ6zY8EjP1vge2vrR3QApeJkZpKl2Zp3VCS4YoOK658p
+3/OphakyTCZHj4mYVo+7Q3XtoZsn9yFTreX6dPmpkJX8pQiMm+H4JiIku8IvelR
wViZImG7KVZ6uvR9Kd8GE2mWRrhPXNBZo6BIiwV1NhYpJ/Du7eIoN7km6/8YGphC
cfsR2x3Bddd+eUerQI3XGhiqFH+hrXAvYqKgk5yRTgF87LpLvvKENHh+wFxDOWoR
dyw5mjJ6xXphrEpc4iDbjaZ7POZNKcftNwVYwLUrsNOo77xzagXhDbDv9igj7G39
oIg9m4fE7yhYAA6bZCQ4chvRhsuRq8+cqEE09jvpYqnN4shkVGs2qBbsmvZIFQN4
VzHT8BTfdmm/PyUFKXF+cVxDstIdUMJxAF/RofxBZo6egxUuyn6Yz+qYfUxcEEwB
L52z7s8U7XvrTeMfAJqEyPOyCEWav3Kzsd6psc6eyXwXIYuxq/XyKhRszIWLNDMt
oeX1/qJWX/04Gs6aBlMuBQ3DRIquZ8qwYi3ix0t2e5ETTkSPGVumsD9lRM1eNuES
WUs68M3gxvtN23uRsSEDaOVADEAhVkx2NMqUlng6cocCDKn8CyAeom8vCZ7PVhmb
3SHN2K3FRBMPCCLXRzKUfETP/sI3agop3/FmM/LqQkJBqxK5YWcIem5X3BPm7iyu
fJwVNqV3gZCD9MSNfjbgKW4go7uTVkAZkyl+yes+sdE2UhctVutSZPJL/eoJCh/Z
FC+NhwMZYMSci/4XusBp6UMw6mHDnm1Z+sXMl5vE3NlCDq416HLDvsoa+KmXlvEG
IPLPVaAwnfG1Keekxk/Zxf9hBSQYF1md+2s6Fv4BV8alOYBKQwcVJfUtKNWAhQkZ
FgLYtXLCUshmsYpvPuqTjHqYcghZkRdg6FjFhZ6qlzvphuIJ5wHxbjXmHtEjjJZg
lUoZZf7CEvQPnpAHPQstIddFuDYdKMu7khI11vDpUBR8JNunXtPIecol8LmSIUKA
zdk6jdw7JVsy4hMt3sX+fgQKMAQ0ADogxvaxziHF/8m8QQIffgsbF3qX1Eed3M94
I9yLSvesoKaeTsUSMAXKzgn2EBxxrSL82tfTYAz07UYPjgxlaP6n36SmHAm93Mq8
zCQWvaBfUxGIoMh106wYTRdVVbgAQ5Fx9ttbetC7Is/W5oR8wZNL5yy5BzAZXvql
v7kuOGkEtvnelTnMshmP6iyzBBTB53bVXzzFDBYi88y5UcJHBSTXK5fBDAHSpYFJ
wlydr7wB5jwgK3jFE3N+RFHvkDZd9aRxkp3PZqS+397PywXIaUi49g1rf9IvQAt2
+PjvfU6m+RyIsEm4gSdHRpxm+YANceKRUM95ASNYVdHoG82Ea5C9BK3ra5FO2WOs
/Mu7VyTsovhWeAGzxOADcIAk4m4g9BYdRUHSZx5V1kgSgXsg4hFzsG7PQrZH4Xso
WGrtAg5d/ST1RbR4hAvOpjLgqQiaUsnmgEX7KNcGZuISZfqlIqy7YM3jURAQT5UN
rKUVic72fzZQ950Zs8MjiX8G4mJsZTzvyRLnCZv0TNSZ4pvAFNpvr7c5decf1AUf
Qyr0IRXPn1GSdywD3IwPo5nWcGIIAmF8EeJ0C95xcvkkzxsKaaspFKbxDknWyvZC
X82TjJLWzJkuJxhtJnpn8gBy6VpWR66JC1g0yAPfzqOl38JcCowJ09Zr5Dif3mm8
psaDHyZdNkgAzZym8lFQZ3yYrlmqTjtCrrWqRXT4QmQplI2yw/JIT9jvlJVjblQU
lW1PdnG7jTJeMYnvlSt3s7ygUEhNaIgnoOLuT75mjhvjse98aNAG3CeoBCTrBHEN
jM82bp7C6LLE3SeTVIqVYnqqEUF1U+QTziOXdiZ+gVwCDb61b4cEnPaVYtt/Od94
nugEzqbjPtvjikGewNG5mkLzdWIjrl4mSFvGLIhVTierzsueOv4hAKOaPmjYp4Yd
b+wlmjzwny6MjxKh7Y8Z6nEObGf/9HsHVRnMirn0lmWwGu/7PVQwtF0U6lFnwB1s
QopViJrXmGpF0dZ5wBHlrlsjHneSeljnzTpTuBNPthMECIaXw+S3+93Q3srHf+ZJ
lgwgO2Ic1LOOS3jWbzWryMGfO/yD9dODZEsZrDiOVg8+/VvizQjfkcnb7hxjAXuG
ehRDOu/DeaAyITU2m1WA+YSmZkJhYsNX3a3BeUyPosKcfRNPFL2ZioD5Qhswjamg
GlMwHgPf/6JPdrkdW0pN8rp1vdCz7WfSUSvOHNk2BbtHQNydpbwDC2UD8Hi9NXHi
0CS5fAsMyowONeLLu4gDowT8jS8zi0cQ+diyVSUJTPWXYxGl2Y9x6X1MUOrYiMu/
nWZVAn7H2QIAjz8pfdEuy9KPhWQEx9yhXr3x/eJSGq8cZNbcmd5P0jOBiARWqNMd
yilgNzNKHskHQCehecgdFIrEC/1x6XnToxAYM0JOjMx4X3Ti3YWgmYM7379lL80s
lhof7mhqInucUAmztvRFF7kd896PH1pBK6lqShmU3o5ukqZJ+IsF7LsoCDkWgdOE
8D2JqHvXT1lgsZTVt0tkZJfxDBvmx5gPpI0M1CIZ5arfU8D/M0dU/NS6MA3aEgjl
sRw+m4dUbaLKERJT+0Bm9/e+7tg35cceZBYqT/MPmaprZ4Ll9UEhx3l2DSGiyjRD
gE6sjWTsbJcgq0ED2uqRt2VYx9Gc15qout57NLgGarL5bNv6H1BWBmSAzc+5iYWp
i0m0/fd3jkSGHM22BKma8BWOQYbDI4VoEHiGjoC0A2iRdZAAtAa8MWE/RSundRlZ
cJ/dUaI7iGDS0xPPB5eiIEN53bPfwdsBwKvWSxpyjYD/TszySTbialJNdLc2OE/x
vnV4irKnFzq8I4MedNpORJIlEoreNPAvHFOAOn+W9iG9LLHYX2MFE4vPzQaT+eJ/
JBQhZEZVa2+axbXmKn44tJP+HOAVQi8KsFI04+JaYYPbGIxt3kl3Y2GkwWPJferj
l2xR5PFn13zOfky2Q7WAnaXZRExhjMgtdgZ7wnCUXl5OW4RfYToDu2ADvoH29Nwd
BUqae4iJAuxa28f1TIMmI57LVOIkxhr4ey3jivLyWKyswomiNrMhzXUYeRQ+8QVR
knvvljwPvCRdDylh0mQ4k1l9ubj2dhCN7tRWnbqIXOdCzibFf60J3aapWDctKcfg
b2lo9mgpVAWSQIjKq8zjLF7yJ8+uKo2pesujeJFPE+L7Hbz3w74vkSl5KFSw61Mc
O4sJD955yRmhZSFQFTAuAH0Za7z45aDJomN7oTvGr8m+XAiQRUHYd8tvj41qQOFp
zEPOqNXWCH/eGrfYmohT8La6oSCfj1p0rY3u6IyG9NrO1rLCIJJTwloQRXauy4sE
UXp635JnurtodiPl9BvXbYjZvereS21mhDhFsMlYfVaP8jcfQt9vMlZ4vNla8Bq/
z1XjIB4LO6Mn3I2KRaipqxoxRE6zEPod3EUYOj8M4v8o5zb24feAyhITPVpUGQea
XlnzDWct9CrtJvy3oIY3DrjDehu9qrR+ajgy/1uT/YSZlSxGp/AgMe/0VVx4POsX
8k35rITGVVIZi71pDE6TmwPChv11GnrlQsCBDPfePjSKw4UM8AQW4AUjNMmd/k9B
Kqa+nL60RcYMBjrIFs32iWuPEAbohXwpViqXaVojBWqa2QFD8zsZQVgfmVyJZU/O
95kgwGgopCs78Xag9yB3EgZnw0odauvTwXLXpOPAyeQ/HAhzvBH5ZCzRq//yHnNT
zNnQOJpwmUgJLRPZfp3fkURacjZSBTf9BKtkRIbz0op3OOWBtHzdaGbp3B3SrwDN
xNAXe6pZ2HJJ8eZfxNJ4znN4ngHt/iZeWHQ1s9RlNh4ElN9f9CfJ/cryhr7aaXDv
THOVg2IYOkHXD83N93q6bcH8mafPbLzc2isG8GYBH3/gK8tno3hFh1VCIcaFkUY+
ruUE0MekF0a2yCIaRVZcZS4lYYC9X1HnkkihIbwgtcSI6EJMzVNmSSvztO5zoTwE
0QxMIZBQxVvWdwNkn33iVq5hjUQh87OvQbMtedds2m3ij4NXuOFDPZjlLTG/f6K9
8/1cXQhsd3LpXcpmSHyUEkK3kmOD0K/qI7jcy7vN+ZrJo4QDbL5Pw/jDrtoBnjBb
DJ2ZEbSFXhHOoMdoGRg8aEDWzBRVQlMId/lJLd90LVQ8gmXbdgrlNxuuBGpFJRBP
cFlZv9XdGnAMLrI5Z/MLdI3nMuya7ZYMs/YCLUKx2nccrw5lQvu5lbC1Z2s80u8A
am5BffpYLNbyY6VWTlsiXVJk/o7ZPXg9uEjN0Exww538nGWhz2SSOBY1g1cGqhKU
WoQiAc04dETfR3jipkowpb4p1xxMrSHoK1+ZyiIl7LqLPbiEY+tFENIBCNgeldJA
VhMAZOYR1YZa8HQKOdW9TFV7wJz4bq5Q4vU3B2IqzEwZjnw3VfqTPxmdFWErrkR8
sKvhH4X61o+ApWDFGfSsiQQGR/io8DCo7iE106oK/+Ieh7ElzPGpzz/Bo6B4Yr+n
pK6yFU6Cr8k2bEQj9VkB7F+NKunIYPssgV1BFBZto8JFfIlKx5uClFZWpeM8iasR
kA5amnZeLZ5zGZxw6wqFETNJApZ2ajv2WNCW4qxTNnDVfOcxm3a4jwt4izxGZbtd
NiPPM9AAYQ2Z5xyr5GT1ri5rzF26g2wVHv09A0WbSPG1SeZDXSBnF08r6yQEY4IA
XcXVrxcTzSj0SytXXHJ83mQs49fMQag7xag0BvjSIJTco/dwESxi9mCsooz914Xg
AFlkyRqHpTJuUk6sJRT2sn987Zb8StheUbCvg0KrcOeFF/m+9vLWHdthcvA831CZ
s5QxMvsVXxj4O2+P4WzWcufkMAYEBF1/Sdt5Y/ARXDQ1S3DUdqnjhGVXgcNc1aBj
fwbgL/vV/Q6/c1jGoNmbOQ6nNoZNhpwJLTkSpPEyEIRPCHvkUSksiluNTxLncJp3
B+koBft2G6WIMlHgDddGM2Ic/TnBODhL1qtrV05PzopaOIEktx/WocgXiNyiXYLS
SoyAQTwU/LAkvZzxWiReq51x/ZRZo+Ci8dS7mfJLO02pT1AhF9N2pHAfxGBh3WSs
fhpv2Ch7dQ5bjfuJkrVMX04gG64xKa8rVq1VpyMa0ar6z0rr1rMmKcXra4IbSuvB
ngYhuNKHbLHiJLF6JZxWWjM6+Z0hLMMdlL3AcaId9r16WxX1fEUz2POaAj4Zzb0c
Ed01L1AL+tbqGMdQe4xKAvzbaK/+0ljIm47Ux97aLM08sZ/1qbpwhfHPthEhuOad
R+TaveFrKw1QgHM8N4hMtkcx+LSvDw9m5HEBeWt6t+7TNmkG/edBQK8TFOHylQf3
64g+pR1Cd3a0/0i26rxuRTuY+CxtsdnhtB8h8BhHjig7oojC3KV7VJpd5lgPrtyi
PQQlEskknN8rg4x957Fy+UT4YNnxPkXu4LRwDrc71ecYJDiYatmpm3vTrcY4oD98
42hznCdxEWbe8m+IMpo4yIW3RREyO+rEeDmv9m+nMHieRF1ym+BT83DhL9XoUqWj
9IMfturQWHze5seloj0p1jmr+no2WYh3Yxc9HjvH1l0rJVUj154NH3lZAmi1kG4L
lPgA1vY20OO3TeCKMqu3rcxSbfqk7ePHzTv2waGdvCtm4k5iLJYAL8miItrEYzpT
5Ltm/YANrFGduWe8XbPp0cYxpM+0AqeZZcS89asl0hjIUwsdu9V16fD+csZgHE6/
0oVRqjLrcuJTMiQMdMYtQUT9wdDf+Nsm9b470F/Yd92LizKrLtocUvVy813fE+fi
rch3iWLqIBEZbp5B/OfH2P/8xqwRjQwYFP2xCY+W0sr/1dJAYcx53DTOALtJAJUs
tjVuz38qYQeJ7WiXy1Vw8FfFSkmGsevrsCg44k8JmwYPsk1+QSzplVZ6njLLahwo
sOOPT90GlmCpgTnt8/VEAOEnnPfSwnWnfqRBoXwU16lvRgwcoiKW0pz9QO53zjGg
cQv6cBncLr5YgOeA5P80y06k62vGEfdUYFQGIw08LNv6C2MkN2rcvvswaHhvdnkZ
NfwMp4VTs5EObFSooKKR1JdbCdgfz/Ny2dh29pNHFZJm4x5W0BuCEqAK4qXHn/52
AQzSQSMAY9gy15e+eIta0gSHaDVhyeamoC5VurN3NULLJUAh4VllDKxP4Ts2p5GM
Lg+ExFB5LNNTgmQFmdWzkLl3P3R2TSYGdW4O7ovkKrCAv558OZONfAz180aEqumn
ZiZZ65aWqpCsaxao0DJPpZ7JUeOtLf32YyAwJM51bPdIuPGWFSHW7n3/9sJNT54T
xH/mP2yz3xvnFvWC755f3wLQUpj9+FeQY//v8XPJC72F5+IEoivIyEjDiNjc0wx5
wXMqkkie6lB1XMTXEems35XAkWxxNV7J+XkoPsnhnm3qKbL/Cbvx2t61UXdaNSUQ
N6cgbFu9LHibRV13KMGRQYJkEPYfaruNWnZXcR0B6+k57hYprnZa2AbVWL9EfuU8
87a1LuyxL9l6dQYLEIp8HIRKl5PnnwUXu02DXZ9gD72OFKqcvNT0Bizy7uityH3M
AhSYVt8ZE/5Jkc9HTf/JfJdEt1K7uJUCEZv+9xt6NSn+VLBh2t4YIPpCfc5zN3p+
HnpBP3dZQKol+NghtlW6mmrGIbZJGLapblCh5369w95VKbEZT/99RWjGOYXCZgJQ
Ky4BRLPKImTmTH2eQgQx73lxrNXOASr1NNDuFnVuq+gvlpEk0EhkV2xFY9OBXkeJ
SyPaQ5yLyLTrLqBkACNnFgdYVYChYs5PXq7EYg13iHS2i/D5U9rjpJV8OiFCHLU7
sEXOQ2w/JKIhTrtY++TxpApprLLo6EG7dLQuzISWC7qqFH94uqZN7ItcRURkfYNN
/+E+7k0Ly06yd0e00z/22u7IyVg1kn3zxCQ1z6XzHAqi0Q/DEA49BpBaO056wFkt
p6uBMt9myj1VLtInZBTgUVX7jEPRXa7Ld5IDGLijDfAVuf5d9rufotCGKV6Im09N
4CZvfxeoDcGWTQ0Hs/ujswjAxHPzScMxyt6ycDJmCcFHQ7gEuWnvIomgK58+B22r
Aar1DXgYnrPjkoGPtBWndz8l55BD0J92idgeaaF+EL99waG3Vzx4tSECMSIJK2jq
VjEmYjtSHetYgyoi8pcy00/1xC3nd9PH6fIng/dkghWIbW6616s8ZQrTpp2JL4nh
yiYBaRWWlBb9lSyv8JVWpQCoZd6bU3adWpKRRDsV4X1pxyLh1FpQ//BPE6wS5KZQ
Rv6KRIoz3sh72Fv8OjHj+fUdn+0LhYbGdEjPunyIT3RF7F7ev6y07D02s27f3rg0
gf15z0c7oPLAmqpL7NB80M3HmSkMBb2GdYkEC3bVyxGUjBWTwAxiDLNorqC4ZyvZ
NPx2lQoKeM6ewR6lcb+d7feqnr9HadL13d0XTSmkHCO1cEJNE5bl1VxUB2FoNfmD
E7UfMMgrh9hNsdSXRims7QxNumDt8cX7F2Vs5pSgYhvyI5km0HGS0sQbNYgnxx6z
XVMkSFnH7Pq5/kSYjAYf0/5iVdTzw0vhruHqNFhcD1pyQ1E50hXPJZhmvB79q1/9
NZM9wOlrNQkMf9kaU6rrdT+ZxscT3RaCmXw+0ZQ2VfFAqNNVYvUf9m0DoblB1R4c
YTyNF1REVlMizWbtWBrxwKUsoIwD9QqkvhKeZr5pY/PybI4JlT8H8PvIhcxyU+n5
UkSV9iKVkCUngNAMD5elcq1v5GjP8QXxq/yZoUh7nHXUx5aWdnt3stXdOjdT6wHE
JeCh8qklRL4woIBtAds+5jNNeH9g3GMjjwB9ib4xRCKnQkmkdzs4A9nXrYR1f/eY
kynMvP8EOhqw4KOwxwVF9NTnGTkiawrtjSDLhOPawTqJXRrzU41JuiCbMBcWsD8+
v8TZ1sa0O6XD1czw44nsnGM1TZQztw+zXREwXfURDuz3vGRfP1n2bT8LnvxXwC7P
CQlKtAw3gDJHhnFWwM4KvjxLp3XLMt245iuwdmmW02RLHPY3AfsZeZ8JZkdTELKA
WWghRDmF15zpxoK3z1BablzY0Nb3uMqMsRUmevlfL8Ej2oHkiyYqhdxXIoRymRJm
8CWTsbVYUOdJkf0XMMhNbTVl1rUHifJzPa/GqF1fB8z8+y0ejsebC4Uo4WcYF9AI
UwBAgH66rQeIBfWOoAToyGrc9SpN/q2WybFwq5mThoFVzU1caNWwK7yMdycpqY0p
J+akCxRQdo1DnQ8zaIDwP4mrqHGYgwuRmh0l6cv02zfXrLh+BuHFV8wcJAJuZ0Hi
n9GBw9So7sudzl5R2p4yNwIGjoX+Iv/qDao2Wzgc10z5/GXsHANryGs60k0jhtNr
npFEit2tNdiPetTH/FETBmNSNzqxSExUS+kblin391Djvx4hj81twfBF/4TQG05c
AJEKWRiWaR1VrluRPXHPOWlN/A7PRpEGDdaOQYpDFEf8kcqqVi7d87J21ZjCCOyZ
45h0B8OOBRLf9/o/1nYM/Rxs5hzJen496WXQujSjQzOprdY2j/c2yDk5zaAEwLPo
/81qcp+uXlW/M5JEFpEWOaJqU/nUidIDJlIW5t9odwwnAqS7sjq8CzriHk4JpJnE
vDfIauEE0aFYwwFfcDviNuVaG8f2ZIOIbYth1qLCBdCXZPpvZBafB78gwfHvsAEy
+dSkh4qsCd3UePNnLcAISVEl3b2jDd2RWMrllT2YZWQe7m8/SySrPyLAoa9E5w9e
347xoPDmzD61PaCXr08mMcnw2AHK2UBwgAkmBcIGphWcmyNqNOKakl0MkXKhKsvz
LjJU+Id1QLlpPvVgvUe0PV3b0adfVAPEgSzDqGPPu8GAoEbEJFYjomfKX6q2Hfes
r3hFxiOpAmvuChoImnjbQwjMfdQQSGo0nHxN9NjsCeYGCs3KY52UMLWJTVx5DXHG
d/zz/nlVHrlgMkXb/qkx/ReWnrZXOreHCDecOe0/7s/RG4e6qoPLi1oDjpm++544
PUll7ETCHUuymJhrmgmcyo9SbrHUd/q3MiznsjGL5pDpbYSqF/QdCfuPwdQIMSo2
1UZYY5NZbA4JQ4T/2bYkxaa0/31LJiUf6HMByDdmxW2uUtQrcFEDGx2WYCASDOD6
eSXHK75cc84KympgY6ZxyOHYwWjDfir53XJMFdEdiqHw1z5xxe/FHhSJ0VWI7jxN
cTNdZgBH5Svk964lt8KWtCEi2cyCLaGCqwDHTQU1Y94bH8W6Hyo/dBasaFHDcQO1
C60/Hepqsx7VZLOudFwxah8K+xzAW7KSeUiePVJPSe3NX5ZQGJeHrhOmBzF7RiGx
rYmUl71TvA9YJXAV1ZzA5VjWDkoPU0LqmhyGf16mZu72r8iS7Mu6qS7bhwx3dr8z
ohxc72TJYqAqOhEJKmRPVomIPopR25rhRYVAFJK5sZafKZ7qyA9A1awBSfRrFRdg
SBLPTpq85VpAu/cY6o/uHa1RWdlsyK1XRt2QVFeqVZc/+uaT54muN2CbeVjF3N/y
f9e8l42meESIKotyQgW6Uim8CT8PalFRqbbtq9hbfPtkY7rFsr6SY/E5jJh+FiGA
FhwgRaPp2UEu3GxP0a3mtj6wjKULqq+urhxunCGibKtXMH1lPpzcuSNHTIDwDy+u
JJsxEHRISkjgA43f44HoPiit8FejhMa/WIGplKW7jAn5twseulD+0ETpooVu/FkI
3JMf2ElQgAW2vRzqJPYK7NOfiM+5gYy9VM48wo61VMlB9K9n1LJq2XQHn+9rL1LL
EIEb5QKXrfBtL+MBsS6S4QCTuR6OI6b9mFnpOau5jtY7lKLHFD+E6vCaETfOEm84
yDJgqLvu6lxxMJhHV5GSfSE3nodcriIibe0ENFwNWECLGM5TlpUXgKmOyjShfv//
ODXUhYHurQOxwzNso+nWWzTt0DtiXdws+XrYb7gF8Y5N0HyyPJoMc61g3FRWKYqw
W7ee8OI7b8dubUgOuxMKioTvs7P+Yv74ryIdJdWa5bsmI2LCIQmhVIgW3HKe9p3I
Sc94QAYRdsd8rDnrfYIeIlJzT92nOJeZvqP+QeHtVyb8Ay2I3VagmoUkX1xSmDZY
4U7ib4D1M79SIlGpY6lp2l0t+a/1R4c7Zcjr8Ie/XXc8MP8+JpswdxLth5XdQSat
MmODXXZpRGF7KN2mQ3zxI/Pc3KC6Gk93Mp4r225dBNIPDMPKGyqx6/mHtf1FQk/Z
7ocK56BYhtLLHzsmmDPGbqp9SaDiO6bajHAh32M50QQE3/kLtdMvbUrOwPrJ6Zvn
U+CtAb2Bs5lvKcYnNQORXy18L/9ECIzRhbWOn3LoGgLFFuojbN/K9q5Tdvz3mUtk
/JAFE0JnQLpLfMywe23afmpG+IY9fJvQBRX2H73c6iEtRfmMGL0e0cKRqSjcLKLh
qRamgvXkJFuP7GlQL1cjCEISibyBgxAlTScsOYmlvIpb8GtreNIy+1ouqo3S6SHp
BC4585+i+xLu8mP3nGEtNHmRRRWh1LAR2nf9Qm0Eqr/xHBw1IF8P/dir4zZSyV9r
9igyANPd1AbkDvNinezMtZkvpntwT7e765kC2wwdnAd1YFls27hYKKTDW8GS5MHs
GJGucXk2LVl7t6bdEZx5Q+RAJoDk+NXPw/rGXoHiQPrhFQDS/Gb9H6xoZVsb7vO8
7zvw5U9uY6Llxld+dGo2oVIsCYYqgTfK31V7Gxa5WEq9OdG54jge8P/ZsCdcDiBO
hrENOMoXmhaj+dT77WowQS4FrRUvBsIZdMKPnZCvphRQOJyscFUgmH8DyK/7wo9N
JGor5gizD6EuXaYBTwM3h0Zhgg16NQUgM/Q49+PVt5VGB2X+ADnfuoruOSfV94j0
tqZJjWXIVwYYIn9ldYyzx6CSw+vZf9SkdArDXd2NfLQFY8pgZyUHHwzD+jt+tMAg
JzLjISIhiYwahR0ZVdkm9/isguChgUQ8RXNepULRy1r+IHRUVCKasRKoKr2wh31b
2zS8pum+SjuXXlpToP3uew9D6TrTEuXfRh5sgaoQ8CaFRwj9tfPZhRI9AnARPBq+
Zu/T+NW5kE+nMJQOcelSizkawYy55jfIovxepAj3nDoqtgtc0Hv7uSPLpGZMz5TE
KsxlH/f3/uC9rGznR1MKwt3+qHtuBCrxSH/nhl2iT0MB9bz0dQZ5lR3JKUZDNYv3
/gi0OcqChgFlcMxe0dbFFjteEAnclLDr7hCnhDcnrn999jpeIXuimuXvLoIWi8Df
cr1GAZSXd7rY4d6OelixFkJXyY+2mCeparuJOpFjsNXm1Rhn5nG+qEOBDUjVOS6G
xYakU7eTNR22vdOhCeh37L2kdtT4wUH/+sVWyHYZDvEEr6q2Syzs0XVNEof5L+2D
nOzNwmJTlWZ77uF3EjwHzv0lJHwteaB1WsBh6gWJmXcUgFp9jS4zaOHoLfaErDDE
1h8khF1XOR83+Qc1l2wG24R3WGukT9k1vSj9AD9ki/aWWADkP2wDz6Kt37fPVNNM
Hva/t76totjGv0jWjjOpP8CXs72x2wdsHHL6f8ozcsfIBPRQQq5eqQC9q85GsM6Z
VVFTqnCMvik6p8WWW5t0VChDv633F/SinDetqVTH9gtvdjQxRjBwAXMXHr3niIYs
r1Wz4GJPiNhsS9s8aaGSqluHkV5J6adwpbaWZLJ5Sh9ptoWvkYMMcgLzWPy6CSlV
8qJC13ZsGFu3kwHwOubZbYup5CDb5KXvMN8l9gyUBVsllOyNTvvWKTNOXLWaUX8G
kEklQ2lIuv50OiPzd3AtoyVl4kBXa55iWtbzGuADsRvVQRPKxyFJ2kFonFWEwiQd
u24hwXJNmSjvK6mWBStJbR4JRUC/FCSGbwVkkCdserubAXEdOGBDWZJHTiKu7Xdj
Cix+cYHwKNiVjCVP5MdJN7Gf+kqXvyquP4wqXrKGzi924ZLWkPDXExM2WK3CcjEK
h6vEQgCuXtkEjiaEQSSl1ui8bvqIohMucPjgqYR6MyKHXBoQb+8e4QNDVvjFz+TQ
JBk40N2Qv5w4RXU92b9ZZFbtEmuXEIXUWJWq9rznV+1xWvPdS4+ZK3eHhRHMGBv4
2lihMZAq0l0wwhUOVgaTcSgU/4dUA5K9yrJbscJtCaMrGIFuR3fUwye/1VpsC7KR
FaSzLRYF21/cRji6nY/JKekUpXGtz/AuUt2Z/nUfo2asBVFP8GPjosqoAPFYgB4g
Fwl30mnUGVSNjX0IcTyHOT+TQ+NeNs2XR6ic0MXYLkTg7NAfCHTekudQOqVCCsz0
EW2PQ88guMtrtHGfeTPOZjIyK7VYTaFO7NjuilFv6RvvaEY9UOLTWUz2NMxE6d8j
p9wHlABeMb+EKWgwQHlKwgD5XPNrIyt/eZfWoLrR3PtpPLrgglU903vloN6zeHJ0
wfsn3C0zstfeFvomZVpLP5Bf0QzkhDL+GZDY1zaYgcOdDihOTaDX+sfxReUBPZSY
A6szg4sjEa3ud03Y2v2lI2R3zMv99IOsvWjK7MVvrP2AYawMRxpYSUmbMY2k2p9/
Tok2OR8sG4uOf4JD+i0ChOtelxrY8yV5lrF52f30bhCAk9JA7JHLAQQWLwsu5nPU
MSZ7yZKQPFICIAV0Dgl9wwgjBNRaVcQkamv4O3swut1pRIzfjYgTt+oEUgdUBxGl
NFQQpLbLvpgTGE58lsPDPTWdMLNfy0V+nom2RBVFtvZ6IiUKfa8UdNz5VmBapGjW
eUgQS2DSphcGOQzWxwDzHZ4GUYgairK4Jd1gfbngmkVQXhSmKk+e6LxjfBgwXo7d
PTNnn5OriwXfmjoeEe8U7YBTYSOtm6IX2eyq7r+GcHkyMt9lfDeG7ekFTN8T8l9U
PCWd8xq0e4nlsLalUw11V+ObHOen4wlXUdMTRYC9HK2ro7IG+6dS3SfjSuJOTDdk
W1qMp2feDv9gOapqMfq1QeKZYVhwtkp93MvXSltNVeGQTEXz2aS1WMkYwJ/D7B/2
mx+uWozixd/2NRlkdCqcPpJc8AbB+1wrrVsKjK/jnaZeNO7A4FCX+zQW9AVyfZIZ
yKZd/5n/nUELIiVtZS1EIry74k3YA49rofcm4mvqPc2O54TFip9gCfC1NwK1sDnq
zhFyZ4e8E9m5zRt15d9nxNUeq4elDSsczGSQaCdeNWFbLjgPduW8N98KZhlNbhmW
K9/zr3V4trlTc/Ca0N3OGAWeg8juJI7HVrSTUPs8Al9xPO9NAzt8Ls7sqCtrITK7
MagnxHV3qFz8FucuartxyHacajJ5bRbUGnA/o4BVUOu6+qnOBiujVxs0/wvrqfU5
viYeXyoGgGNDpDiEDxttAHzrENAGkfGvgokUYwMkwZLCz95kN0kZ2cDSYYqxOwTG
1tKZKuzdcxezDysAgkTAZend2J/JuPNkqkk8IwjGL9cn9yBd5YSV7XAjwUrTXnq2
WzVFAD4B3yd5ppqY7VH82WzRVmLxbVf4ku1yRd37K2opzbOETYYNXmgaUsdOykpz
qX4zkz1v9YFf4NcyHJdkjuSSDTRlqiezO+LdtZqRoFo0d8utuX/uXTWLTEa1mU5U
W0mqeJu0zJdpwOpQ7ZjWh6s5xCQICpyBCU2iaZruhoYaqKZ5orxM9RQvh9PfppJp
Yz4Bdbz3qiPHtmVILMOH7hixQo5hDi/5fZd8QNY64z/7VxlVHZLwrNqa3GiRmMrN
8eMnCs2F6CxXVoU84Yy4KkpCBYnNGv1Oe19DPoq7beVpUbyOSOHhNkfX3AzM5e5J
dMUbwTT+c71RJg6r/wureYQZbERFVAuHdmMzLywkXViSbhGcAjNLyxg57EVLo6aw
MkpH78Jy0E58y4prtxe210tjD9MIXL6zysMf8KNvoXqXRTWJ0QwRPhJ+qzG/iCXA
mhyLKZi6XY5yH3sDPkrj03sVg4fLRNTXUVaIsikjvmbJHzQLpB/SHv0JHVr0T/Jq
aVI1YWzRitL97ok+WGBG0JiKzRutLSCGfds924NI4LECwSGkoGCbn0o+uSSIQm1A
YX1Vy5XJ276Z0iKN+fAKSiBnwd+TSICZ3Lt1ZuSL1GT3lMdWIvP9rlwBKX5EaHoS
9XthH0s7kRvr/bo5jWdwq2hEu1VYENChvV/hVn60UcTa7SVs0ZRv0VQreKoU/UN0
Dr4lcxSJof44WOCJoemMdWwWwWtDsDj2tL8orgvLPXOKwSNgAdJLtvBl2Ce6au6h
cGwHTz1Bedtxv/8LDj0dYqf8HtOXmjYyXoUppLwDwwv7TXMSwzlh4AXIJ5AbxcDp
AxwgAhq/ES6wgBlpvoL0pZHCEQDZflMTr8knKmxXJolaYUpRAXl9mUxes49CjiiT
ATWOzwKGd9peoyPEqO/0XIma1f+s+fB+5dTUYoeLZTkXpyX3Z2naU94AcfWu8+Pd
6riI5pyaAmE58EC+v1AKVnJTywR5plZzmjfRZiV3QVwaai2kK+R/Dmhs8CmQH4kS
Chake9zSlgUZGC31HfZgcF9zxrsyVy1DAkxRkkyHIxW+AkqXhIB2zgk9oye5qRZS
zO4B1Tvvaqu5agY18DeJ5g1H+C445vL1GJppT2CDIPGDrMYRS8u4VcHLAkHIEeLD
ZjHxaEJDwP5oDRTQFEBe3L61FN2nIdz9SSAhiHLt/wUWAbm9B0XCrUNndmdfjzQ0
LRBdbkn3fJZKio2BooQKJREiCenJuVDv9cO9QWYjWZXjvgDXzwi+dcd0x+rOL1lO
pfh0EtJaP+PrlO0oZZcPsNGdFoMQoXKzUhq/+Jjxz304kETN88GKMuj91cfO8chq
/SLqxTNtUe5M4CeLlQcshxaZUa6UKGdmHciNWgVGnudth1FOyuqScGUzMCyBaTMG
IP814DTQzPa7Nf7WVD01VTSTdrg/dctTNXi3A43jOEtIDu6shC2HBCuA/9FtAdBY
ihH2F0bW4sQ26c4wU/H7iCpd/xUNRGbIuKcfpJBs+vq4xvRvEnrd0t8NXW1/bVWn
UTJpA7s8hSoiJvOQajyCNTADbWUJfSOos/YXG338TOIbQFzQg0JL7tyGKDxbbwTR
+6UOkwOIaQN2gjutKqC6CHeAiAOF5LlmMqZgcW+Y3YacKGBTguwQCrqvvWrAViht
1ytdL/r0kEzgFWGSDXW/L1MEQwvl+dfMtGaLqAoq8bdqwMaC0LsPiVU1vu7TUSxL
BgZAJ/hrGDdNq0KslRFGtvIPcb1JpMzwV/YhLDyC92UoKGd9s1DLapPLhWw6KIh3
MzfkTTu8Dit2WPg5aZl/49mNpburonY2ap1HI+V4Wg3KYgtkR2eN2q2MgUNnFoqg
lOG0/Tgx2Da8n6PEX/e08p34jonRIL0aaRUz3mSjWhwhOsSBiwuF28mcRGh2uXjW
Hr6ao6L+fhqvd69ooTU63J+xO9sLscK7OhADhBEMVPdQfgd2I1iRCZgAHjlr3jAn
kxhg24tnJxv1Aixn/zUb9qSY1uOalDyfpGzOww4xRE0rWuHD0Og44Ny0ohQ5nVnM
Ge35QP1Fj5owXCBvm3utWfTAcZrHWBdc9HtgnHvEdw7O65z196St2vUljJl8jlXd
sa2Hby4mWXgdE6ZK2yISGmLZSqkKHPVRtwYNsJ5GLQcz/EiC9uh94w+1hpabmpS+
vE9uitE1BFGij6B57DTR4wlXPlhjyOYcyBDZt+YhOvGSIY0G1+82hGcx+gZImbcg
EEn4EwKZcAiy2hBe7Qq5OFKdN0VdK+pRkqZpVCDek+tsbrg+CFYwvoSnpNx8RfAs
+dXAdoUsCIq2yPdPKEMOYP7o6vRje+N4fAl0grUjWZbf6HJLp4mf1SCz04gowAQ/
fJfTsgnjblG7fvPgEYItnLKJQ9oB71qXgMupk2ZCA0JxgWEevnpQtSCTrZTMWOVf
jdWfpO4wuvD4jqtt2846H0duBrKRxfKMQb7DoaNzOePyGU9K+VWSwledktWxS3EA
CRpkF7iDYIvXTCMPqFWEC72+XseNu1RR1HYCOdxOeA0C96cZUyVPTuyAoliApB39
kgSsnPGvYFvJnGkkOZx4ZgQ0XcY5c/XULjuZ1PUM7TI9BdyEoCU0UfKAJwfPOIE1
E8lwAzWxoyiM2xkTUOwHEySU3F8sbhinta2R4WlPDaAf9WThkE00606+IVNzeNUU
eYMAHmjRg1XHEa1kbgau9LZU3f4/hcCc0BmUu6pyJA5IGLh5qBv94u7/grXySsMX
FwjJslIXSv/P+FDHV0YHEuvf0t37sRoTCet9jb8HyVPs4FavJTcmigiQ1Basf3t9
wbwaQfow/tTl6BJnUGtJt3xsekBlHGPxp421rtIl6jMcCm1FN/SX14iWM1YlJOau
IZufB5o27RMJ3yCSS4IHSL0HJxp19YxCcfpXQkuvoJCxiey5UN6koyKnIzFst/kn
TqyxverBhpbTeur4QBYrUc5dEz1q/msYRx9JWaGRC/O7kDwKVQXZSa4M+bYpYrsY
kxLWCO7ZC4Foi2p7dYT8ffjwCAstBmlDYWv4Z11imE5OU8r3bR6FmUtHNvK1+WDR
E+hdjQ1QPscRi8du+AWbUQ9C7EduOarhlCEhZOossyU/GWqssIJHg8lQrfITH+KC
PV4mSIARdAPxgWSQ37EkQEJOrDGDMAF5jdy1lOIsaa80e8+2ZO95m3YrL5gCQwJn
TzbDGysw2eN59/mreQeQCvvPnyeFwb+SrA1Y78L+V7Zw984et2U89REeaXjFTzbZ
BZbwDY0l37aqo1EBI457aC0VC+nJ3sXYEx4DfZaY6CHSDyx/O20xxAegl7OyebmQ
ZptST2rS6DKXSusHeAHcSBn1+qk4W6LJTlq8B8+b0zfZtOtC2kalmPARqywbQ26w
9mKeYUI300KhAhcTyPo0tjuu4b7e+tKSlOFMbi3oodgEx0GLUpuIrWI97WCrLbBB
+34dSPIWKCGtIrHKnBgPCQOnUrrqSjbojFwUGI+Y+CK6uyLhUQVDT3/1JsIX8B/d
6ZQQ5hP7QO38u84ZLPX85tU7Rl/lta2A43VWu+GuuEEMp6Wdw//bkOenwfeTV/Sq
bTnvd40O+DaTfqilnjO6HgZWQ7Zxy9th4sfjkPC5aUbP7PioY6FK13YuHIK+n98D
hZGak+/slkRVe11qUh4PDstqfikzsVQiaYIG6pK8Kg6fzPxLsY7NrW54dE0qeF0V
V2Cd+40/mQ4WQpiiKLcGBlS40TKoUTqx56TWiLBiKWuquvqQ2kFLWDC6AXvIj4a4
/ImOOMHVKL11RUyUHRxxM7wKmzX6ZM2mnLZsKoZ1VgzILIMtu5Mbj319L0eH6YEg
0j/ceOKnyIQUvKS0kpPYmUNabmeiwa87XnzLxKQfUv61yJUHTv8nCId09/HLfLsW
2DvqI+EqfXmlzL94lhgJ8v/ykd6+FyX0cGOimTyRHKIFbL+DrYkjhNwUUlOzc8zI
kmRs2w+T1z5BCVfDvuW+xj3QFcJouNM/C09jVJb/NwO3evUJ53N8fNvSFJpi2A3r
h0eO/v/dv1cy/Tyid69j8DzcjV0WfSP/tMz4sptoYMp9M4pXwHyHJPdvxiaiEWfF
ezWQ7ynTz1quHCq5hrCkFefmweh2JpqY2KakTlgWN42wb6Lbxiqkw8I3UfpSt3eZ
uiQka9H8WIybxFcw76M3WCKKITZe6VAdLYQoir16R1Y=
`protect end_protected
