��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki��Ы�T�￉��`����^�s=���x����<�����N|��"�����z(� ̛�	����1g-��c*ߗqT'�C�"9x��)K$�1G�e�K}�����g����A�e�����~��2!CI%�cp$-��*kj�pʶ�n}Wzg�Sޙ��j y`P��e$�	{���3��Y/����������ƴ��� 㛛p�ǃi��|e�����e�Ol1�yj�f�D�D�;r�\S .[�U�)X��͝�SI���j�-�q��6��?J��i�.K�`g�fy�f�$hI_-�;�>��iڃA���8`��w�O��s}�N1%����XkJ]�Z�z��bѨ�p|bD����y���ߌ�?�?ן� ���� �+}!ڿ��b�^C<������@�
��l��o4����0���_P0p�1�s�5� q������$ԅ���B�ibʋj���"^YG��� �t
�MJ�:�}�2�4`y��#�B�آt�˻�A_�ZU(���(�J����P��6�;��N�:~$�tM�'���S���24i}ܲ^I�T������s���]�}M�_�1d+벂IqU�_��Qm���٥��t�)�� R�0��}0�t�u�m��Mm�Z+JF��H�@?,rꨀ6lnB���;��P�����ѨT��ZN������2��
p�q6���j9�>�5�]��l�
|�Ǜ����'���~�j�� ��V�s��O	G;�!�d6��O���T�~��bK�G���@j��(���Qg-d3)��
֬��[��oe������f�aa(o�:���w�"�+�?�("��P��ۦJvX�M9� fr�z��%<O�1�{TQWƬ��nBѴ��&��;�ϑF�g����}�[���,XV�-@"�N��3�����Yp���}?\Z����j>�R�7o�%3�������P��Z�`(��$J��ggt:�)�Ww�g�o�8� �������̣�B�!|��M��]EO�,�����|��F�;�X�ɠ<�s���O�����Ԥ��G"ٖ��C1v�^��֬0[�7E�[��g*��G�W\�Q�l:��yw��֒��P�AX��1�{bt}Q"M�8!aA��:qw�B���aթ9_��� �^([V(���*����wi�j���-�$V/bB��p�3�dX�xO����j��I�b=���A��i��A]��ί+�^s\E�7�BІ��	��br�d#�tG��}Q����R� ���.�{<�dK)I5r�2��T��E��Є?�h��iM�U�k�U��y���� B�x�T���a�	oxjLhE���˺G�E��2�Q�O�qgR�* >˙���Mq��ɖ��4J��xm�΍h7*����`�k���nC�D;���� V�J����F�4�F���,��)�(.���zq)R��w2��kUH�{���#MM�w�� �����A�]F�����ꗼ�ܞ�F����n����·`g���3Xs9|kh�-M6-g"�t~��~�f����Q�L���3�	�E�4ݤ����c/�T���n�C�ٺ�v<�-%v���DE]_(�R���&
�Âz酴!B���%��ƨ2�@�gA���*�b��e�*D��P�f����~�V2(eV-D�f������hMbM��-���T;��q>��!��]�>�d..֫BBͿ�1xZ�|	����g��ag=�[?��>*1!G����FʬG��7��W��ّ��8�1p�L�0[O�M����g;t}U�1�@��JɊ�� W�T����{�e�5�$�<h�T�t$�+G=5QJr0�I�]Uf.�q?P��Z(%��ЋUV�1���3D|�x�;�씓(��5�cT橍�n�Mew��)�i%j��D�E�	��֍�h�yc�K�a���V<��D��!�?��s������d���1iHDɦs
���-�Y�4�Jby˾����A��uXL b�8��q�Xk����q��'n$�2��fie��Y��J��������'��wt��1���zm,'j�����=���{�q`�1�]-��/��doT*/��W��P���2R��`�Ȱ��OЉ�.�۵\��;h�/ϔ΀ޗ�!]}x���_-����g��>�:�,���?��Y�"�<Bm>�\�Ab��N��sxfUU�^�ވ�3�� ���n}�at�
|E����쑰;΍n\*@ogkn��Ǒ/j����+(���)�9O��g�
vr��Zͭ�Wv�x�ߐ�j�C���yj�6��j^�;�<��d���=;h?�Rzj���Wz��]�__�9��4�����g�e%K��W�nQ8�A�>&���EV����Tk]�Y[V%����wZ����ڸehf�d��;�W,A�<�-EU�^��oL�F��X.�tIYҁ5;���:����E�y@F�]8n㊋+�,�5\�A�<���r��D���ص��N�է%%��{��޸+���I
��P֏�W�l�ʩ%��.�BG,R �}�p�/��?b��2�'��	<�����j����p��0�{y%]��#��<�j����*�ڳ�|a�P��@Q���ژ���g���1QW2���H4,�7z�Eu�_�3/���|!���>1��(��)�k?�T���5GA�+�c��s��j��U��
��ݳ���"��G�Tz�7y�/Ʊ4�_�1%�z)�L��V�� 
e\RfR�h:��4�!'�� �����ϥ��� y� \/\ȗ9Q4/��#��+L��k�ΞP�OwV�N{����3�T1�w)�YM�Y㘆z�1�L�]d"����+o����jʆ�tը�6ll)8��c�鴈o(b��:��$SM�<�6�ng�壬��(6�4H�Md�|���2׶L=T$3/d�v�(���V������k!S�̣��`����{2ZRAd���>��a���f�O���π��`��" �����R��U7��Q��=ό��D#�DR ��̪��A��i�$��dY<����7X�"�i�>.f(o�DJ�
*�#T��;�?X�*�1@���ii�6�Y4[u9��<�6:����u��)���P�<�֜D������vXR	����ڃ"�f�[���i�|A�"����U�gh���LF�X��˩]��C���൹A�$�Ym��/�kI���Y�ƶ
_5����[�����f-�nF3����2�i06��z�[)�5|����.a��6�hEH��(�.�\��$`f�쉘�Lf� #h@����{��2f�\�t��$"�H�Mɂ87<Nj��7�X �����W� b�O��S� ���cY]�y,=�O�MJԻ��a"&]>��C%���2t�Ճ�8��)�8u�Ʊ���=������n�"�X��$��{�V�vF�ЊU�j����{�N���Y�>{�T�)��;��Q�D��m�l���<���ݔ��4Bøg܃E�D�a?<X�6�)�dl���P����R�	:2�M��qܡ����De7l�d�h � R��L� hD1�ڋY[�֕˔�D��ر�b�7�mg�U��/z����7C=;H&��TM	љ�Zt��k꺰��'SŎ�	ubX#V%�DQ��<Њ�13<a�60'��Q�C��e΃��S(K������3/��)�*d��0\D﯉��n��(��S�8����I�>���!����	�_Ҿo�,<��\Z����`��R������1��6�����[ ,�3߹�aN
.��l9�� ݿ)	3g�-D�jP�ht� ��*�A��jzవG��7���>��8�ٔI�s*N&.�X6�<���� ��79�u�rE����7NR�l��m����R7���`�
~�\���2�d1�о�p�~�ϏO�8#a�/�PUC�#��	��>�R%U��aC0��&��p�mX�O��?L�eF��؂�!`5����J�_�"�m^��G��8e�D��^Jkv�'�A��vxb��!���6*S�ys��д���:�Q�`	ѯ! RC3��Q=;���?�gA'�3��;�ʀ�J���c�Z�ۭ���[���^��^�!��*��+ҁ��h{C�<��S���*��Dl:F�O�=!���QVO��+�.���7�a-E�"��Ur�l}���X_�� L��<�t+$K�.�l-�gC���l(V��x�º��d���=.��׌̮�Q�ɐ{���O�*s�j�?��3�L�x`l�"]
��Q_��sQ��?|�"2���3�q�4t��05�u���g�&�2t�I|]�6�6&+O��wW��^HL���y�܈Ŷh�$�4`0��{uu���=��0]�rZ��4O�el�~孄c_�L�϶w�a�J�棨�,�R>�:�c/�-��0�0�"����⫮\=���Z-E�g�~�><�隦6?��KŤ�=��Ռ"�W����#o/�v�&٦Y����-�bZr�ջz�>ߋ����O1%��xWMA9/�)Z���⪓�^�J�ˊ�_���"i=a��l���*X!����i[��e������~��6Z	fPE�$7��B�$f�e��M��*q�5�@"��9���['n��5��_\�)A�XD#��i�|7|��Xwo�@bF�ϭ�!�tY��J`�6 ��`��Z9��4� \���Rİ���u�s3���r�\>��lC�لf� �u#qV�q�u��SX	|b��X���dxcx��kD�L���5p���u{�9�ǭ�)0��L��~�C:S_�H�+����>�ڏt~n�)t%�p+�j���Uݢ+	��$�M|l'������@�H�a?V�.��q�k�3��\��So:/�6�%�ӥ���O�	m�Sj��h�,D���R0Fќ�M��ڇ��8�
�ٿ'9�
�3��>�Q�Z�85�Vv����=\(s3y�@H\ �1\�~F���m�3N�T�w���z�=�SzO<�7JVɛ�Fj�s�W��.�Ck�K��	0o���%V�r���s��g��tIf����',K<
ܘ��"Ұ�UP�r�Кm�;�),3MH���I; ���L7�Wި�3r�-bѮr>����֥q4��W:�]
�ۉw�����I#�*�@>��ml�}qQ���V��t�G�����-z��6tn����O�Q�;�{Rl�b)o����أ8���������+�eak�)<�JO]��|����B�7�p��{-�����pJ01����/*F0�wb謪v'���G�ꖐF�e^9�!�@kU�}�B	;46�������[���b�`�y�k����t����I�[�i��sլ�%�l�%�C�u���Z��cQ�m��Xpz��|��n��̱L��r<<O�"K$�E�4RB�)����t���QzC�"n%z��Ҟ�p�0����C0E�)DN�o�`5O�q�a0���\R�̓�gsU�3���u=��W�&�V�cţ���$(2gX��fM��ɱ~��\��=�}�|ĝ*lx�z��uwH��i�S΂��4�Nv1(q���e�c��~�p��؋~�*/�D��QW�?�͆J��x���6�r���b2CiF�ͦ��>Y�e�su����b����82�_\�B���}�3�w{����
��<@��C�粌U�Ii��'��Ш�цh�%�m��唓�13�pil��6;���h�[qHN���1�� �=QZ�8$4[��I�e���Z:'^LW8�z�.*x�C ��AN��M[���Y}�d���7�
�<odR�%P��D+8`{��9�}2^�M�4Xx>���N�0���gN��O��cՊ'MS;�%֦�0�|�d��2��<D|��6�x��o�Vp!3S����_�W1'M���wk~��9Sv�8I���.�LJ�5�`ٳ֘�l���4���>q���U�@�L�Z���F�LD�x?[5q�{͚uS�>)?�p癿Kp��Z���E���m���yo6G%���r�4^I�2�;�x�=V�[���ʚ�Oo��es���g�Cޞ�0�����m]�E�Eh0���>�$:V����)�%��Iy*ۋ�݂;�k�o�d�~����cE�/�XAF�,p��E4�8؎�|l���ɃB�3B�-2�b灖<��ۉ�J���=~�ԯhéu~k��T�H����bO{�����ѰMX��5�ӟ�ʥؗ"b?��'��
�������
�^`�����?���M�7adծ9*�@sH�8m�����v�I�O<*9�x���I��Rn;Y�v�ܚ�+���a9�F+�Ǆ�y��"6�y"���H�c�a�U�)���/�>-�H�ț��'E���[�#}�������!v�.v����1�7�U?@[���=m!+9}�$*�ДU�9�<�;��5y����C�-!3�Y�H�ד|��ј����)��d��a�v��ڨ.�]��)(�D�[��'�>9�,�cԅkC?��`�La���G�K^�E�q��G�qڢC��5ܰ�d�B3�p�"�@k!����:ڇ\�	��Ѕké�,��f��w�GF#J,寵lD�3��g&,���`P�I��b��2]kX�gwB����4u�/X�j�m��J�����mj�(���1;1�3��V�`�:;����&h����?M��y�v) �N�*����2|J��
�n�t�˪�T�:�+�����6�o,�u����+�a���0e�̸��B�+q�;R]�{{+�%���bVI�A�Ԑ�\�T󓡕i �:�f4#�ڋ�X��y��z�t����/a�MBRV,�|��������.Zx�|�G+:�B�G	��4B��7P|�۸�_��,���k܊�W1����n3�Pw� ��%_y���p�C��D����)�@R#tx��}�B���Y o\����ʖ��z�+��T���<�wB�0%�R��U�w��E���1��9N8=ۆ���܍��$�*{�2�gjS]q����,��J�ii�����]nN�T�$��L��U�(�Մ����+�a��#�Qmm%vn2�WHDӴUH� ޑ�G��$vz�#_�]w��Y~�_�2�Y	^�?�^�6��0�=c;%�S�9�.�T呁�-�z�5�#g��<Z�7r�@��Gv��5�������e���3�%�!��G�Q�ݧ�H!i�bMѢ>�'�Ҳ*^�G���N`��s\�U����5�R��v��/�`N�>����P%�6i��>Tҝ���(�>������#,����Z��)��6�s��Fxؾ�h�S?�6�u�&�����A�����8O(�F�#���D��H����oX/,F�!s���{����oa=Cy�J��.��tv��d��0�j0J�Cvq��t��]k^��'�;[���D3�a=��<�|�JH*R�����_�������b��O��س�������J�G2� �Ǭe��gV۞q^.�KP�D�K.2�B4Ri�d~6�.����4�0�cU�ϟ�"z���ԏ�A�+
N/��qR^m� ��ފ�+Q��-�[�����给�Q�?�Yk]���7�y�n	_ ݆��Ϲ5��(5+J` ���3��4�@��ҕ��z����7H��5���.X�@&����S�%z��T�iE�-�QF}tY���	�\�RV�ji��"#�b�	 ����:�4�'�q��+�^��n�Nq�8�L<�𛖩���/���PAk���t�w|��Sw �F&CL�6$�Sߊ�{
wTĪ˩%R-��ym_¹�ݗ���!��a�����&�N@MKA�i���q�I�p�現�f��/<���G79�ox���l[I�M�}�CC�%UT˯"�$�cAC�%ӂ�w.z� Z}�W���x��h��$�0�����u���+��BΊ�x���bB,]�=B+ I�R
�j��3��X��@���Ц��X�x�LA��N���(��_V��'�1�����F��`j7�8�#��Ӆ����
��kS��ӕb���#�垳+m��6@̢�sb'Vk�������35�� U;�����<q���a)��%� �.��aF�.�О��_Sa���I'���q�!��K�Y�C^�.��%�;-�~�����K�Ɖ�@l��IM�sW�@���
�ځ9^N�A��FtU
D�=�tN��_?]��Y6K�$J�R`P��a��8�%'F� ,�|L�,��*�
Kdq/y�b�<X`��rQ��b���͚ �)Y���OGn�Ǖ�}��0�����fM�u<��\�c-�̎n�܂���'��؅i���������̓G��=� �40��6,��YZS������ׅJDr�i��	V~-&+�t��=^=�({�U�P�z?R��9� =b�'�N��r���P5�MB{�����6�.�Y�_��\}�΍�ˤ���e��������X,��z=�{t�7��c�� ����,3��ur��b�����Z�+?98b8Z����˲<<i��xj��X�ӈlC���j���#@���U\�U����B-���L�F��v�8M��d�n$��F���b;��iT�ѯ]�ajv+�h���Gg��z����
��̀�k�Z�/ޒ��M..E���GT��噦h;L�WA����O���2LK%3�4���Z�.EUP�@�T��BW�$}r�����N�"O��Z�Q�j�މ:b�a���;?��w�!�Ǡ��#���I3bZa&�����������r��1��C^�f��p�kt��0��c&���ɯ<H�i@��"J�hTՠ.pG��	}�@�����%4lG�#h��|��( ���
�L�ù0�=v���6ʂj�T��N��> �����B���n�,�S�,�Y>������ie�?��W,��@,���f�-/� a��-��괫tڴJXVE�Hg�ߢEoL���I4a���1.g�y1�_�v�Y�.��R3��@�݇L=���Ru�.�D�l8V�	J��J��$�́&5����U��L3k�<�ˤ��ߟ8�џ�r� E~�c���ǉ��n d�-�E"�,�q3`�|�5��W��E]`�1���(����A����ܒ|yt�o�n+���F�{���ģN����I���́zV��ܾ��{��#�yi�j�X�Q���p2���!��7��.��
��b<�7�C�H��}�vk�C#m�̾����Q�����g�h_�+a��4O/�%��Mjo�d5K�;�1�<2&r�۱fY
��*-~���v0����ͽ6Ixu u^�k���O0����S!�⨠���j���s�7Z����H"��[�h�������?��-�xJs�%�����N�������e�"?�M��Q�b������a/W
�p��ټ��\H�"����S/�g��x�+@J�~,��j��U�!I���_�#γ�m��o ��
��A}���j}�2���5�Zz%���uZ��j��珔�;����U E�ᐪKq�<g��w�Q��9��J !E7�T���E�~�q��~%���~���wa���?BM��)�X=�;U/�7�g7(N�k��CZ��7@��+E��?pPFuwn7�6vb�M�;�ð�
BV��Q��c{ypM+����`�3 ���,Ґ�!U�|3v�[����L�rF4S]�7)
Sd���a2��B6x,�*g��� ut�\����U��?*������d|���]�ޅ�[d~{�����������8Ѿ���O��u�|.&��'leG��n���Tv=~�	�h���H�)Y�0�um.w�XS=1��q��8,^D�D ��7q��& Q1h�m)4¡��0�p�&Q;���Ol��d���$*�އ���#��3�
��wH��I��X3R޼᯷'��w��nOn*����:~G���"q�|~oհm_�2�J��oWֽ>�ȂO�P���e���/���=����N���l2�#��MĐ��3?��Ǟ����f���(���99��n�p-C�=< �Q���簅�;���ׄ'9}߿�$}�FQHL����9�x@n@H����I�Ϣu�5L.P�
<��Z��D���a���BQ�-]�j���gp{q%��B��0}���}Q�;�@�Z���s��!�K��#{]���wP��������q�@�:�,n�z Ff;�{l�I�1b�z�}q��j�0(�!yÌƕ�:�4�F�eqơ����H����Ex��Đ)~=��1��]˘�E:����*ó�(�F~��`�d�`����a,�<��D$e���=Yeú>����9�I}�ZgG�7���~�u*�aJ]6i�Ao��P�7 %r`�c�{�)��ӌ����^����%c����%���E�B��Er�@X���4�$���2�ޮ�G|��G�7+1��6�t��f:֜�&��K��X�1Eӑ.K���R&�o����5$�X�<�m��:�
9�e"�F#R�b���s��?�g�|^�JM�v�L��`!^�]�ȍ߭i��G_������?O��߬�����r'X;t.��σϜ�g��7(�C�y�� l�������1����w�)m�P�R�'���|��'���M��pm=����s��n�,���z�Hea���+�D�d	��E=KzX۫�Ȫ��:��+'��q������v����$�%�<�L��&�U>�tι�aPH&H6��ogȫ|R���,G)�@���!��G��9z\J�X�J$�!�0l]��b8�J%����t���JcH{$w�.͇�~a>�x�ѭhr�N���Rv� �P����'�:�G��tE/�gҢ�g|Щ�Z�Qn��߽q�����29(�QD�.��B�-�HgF�����`2a�2�2"�)��a��R����$03�A���@TWc�z@�w�E3X��B�J}�X�U���N���f�7�ڙ��f�ڞ���H~�҈�A���Q�!�Z���<����$���g�S���]��X�nw�.87�s��7䳤"��7|l�����bK�H��b��h60�g�1��k��Z�z5��q	���sE+I���q:�%���%%K���L�-,܁e��$���w�3�|���ᇠm�H�>��IP]8z�d�,2/��"\��fH���i#񜣃k���5���nuIz���V�h-2�-Ŷs��������d��FO����J��>���q��2k�g���$��%�<�]�F9�<��v;�;pn̯�ޝ�4QgbS�)����������v|h]L$g4_���3qe<؋�1D �_�14HB�81`*�H�i�߽u�iޖ�vȈ0г���L܈�����k��v��dCW���Y����������������4?��U&S�/�������<��w)1���r}{���/_Ю�tO_=�R�� �IW|>f%������O����%I�,a+�����<;�uJ��P���mK�( tj�6�&�x�Ml�1|�k�
�'8��[!���Tj�<��.#��^Dt|ꡨ���'�d�~� ����só������Rt�N�O4@�;nSo�P)e����RU��?��JMՕ��.Q a���{!%_|������&���Y���HFL'�)��f���p��Ҡ�IX�b�Ԉ{z$��8�����|4n���qs�H��g�a��5_+k�	�C#e�i�_�j}�W��Q�@���:r�Zk�t]d\Ņ�C0^��_խ�9�|`��"����>;��?��_=�WuKL�SO�ަCT����f`(oh=`tUƮ%�:�$j�)�v@w�k&o�t{���?�UQu3G7&>�.��$�?4����x��zm!�"��3pʹy��@�i>A����R����r�b<L=QnS%!�+����K7^��x0L?�\Oμ{Rl[�vd��*�(�
�����؁Su)����ğ°Lb�BZ����d�8�L�A3�ހc|6�ϗ����@9E�/'&}��rs��?����>��$�h��(v9�ݢ����Ɩ����}ƣ���0_av
��y���Å0�J26Œ�l���H�F�?&a�ܭ��4�ӫbV3
s�aI�`���8��W��3�b��}R��F.~,�uͶ	-��l��]N��>0��VU��6�`Iޭ^� .A���:�D��&��m�O�չ�J�^Wހ7?���Ø9:���
����(�L��`�0_�S$�md�!r�WɶN��91=>˜ð.8���ʇ"P�Ѳk�
 I�b-���!.��P�B&V֕۽&�6׸�"$����[Gb�(�Ϙ���*?�̋��$_QKޢ��i
;���O]m�jJ��A��p��e�v��0Fޡ��1}I$���R�?/ܫsd���L�k��� p@o2ג�PMc*�axj.����T�� ����/�h���J�q���(�Q]��p�RB8�p,�͛��~k�)�]�i;�ť�7���,p�C#U-��B��Y=D�k9��$c��N��P!�q�٧Y��� 
G�����C��gx��1
�=�B�m�W����R���40  i��K��Z�8��£��dY���~`w�iI&�{�[�țU��r[�� ��-W�t�Ҕ���䪨������zR�Mו��'��t��f�"{	�X�qvC��T�ƗO`��{Uϩ,�&9;�팣�r��@��eŋe	�sm�Aͧ�IQO����v�_sD�G���a�.g��V��}�i��j�$x���Hx��:G�P�dW! =ubE�g8*�7�C41�bbz�ʜ��o��	8�hN0�Y�K�-�
��"֐�@a�*Hj@���{��C�k'��^�E+�"8����s�?�m��;kt�
k�!�_~,��A�b~FQ`4��^�wL}��TRHr��w��<}�����	�&��\�ﯪ�q�(�8�p�r���1���_����KC�h���TG�R��<��'z����g{���0�R+XU��Gp`(ӯ:�G�\�$�!L����έ�0q�E�p��;�� ���[Gk�/S�I���1�W�P�`������&֌���٥����������(�1�ﭳ�o�)\�PՋ���Ҭ�Wk.�@2���x�A��..�Yc ��w)%+[���6�6*�y���n\$P��ev��^َ r�Ao��(�V���Ys����j����@}:k��8!�}+��&���fe��ZT61���1�pr�\k
�8r˚^j6�%������q�:�C��ҟ�×�����8&���L��3u��^mfpമ�l|�A�^T<ڭ��sެJ�}�m�uW���×2�)hT��gfg��zQx��2wKZ��9�j�-!�~�TG:}� +]��p�˽:����%������cV�8E�M���6i)����u��g�j�R�zFl,���NL�#���; ��="�C��vrsC�B����ER*���Y��L�z��ұ�[ʫa�	D�$��kb�/�_�z����t���&���@!c;�3:�䖢��5/�Q!y�2Ŵ�GTD3Ɓ�'䈤\�]�l���p`�����F��e��yVT�gk�
����]�܋�fō>ѥ*Al^L�/_Z�ζ���}�������c|���?���{����6ߎJ���zo;	��Y,(3�����K��+�/H+�n��d�����#usRof����y_حnJo
z��$Ϡs�D<�.��j�%n�t�o��\6���T8��ڬ�����?��e��/~���mo��!��~![D����&i���.y�(s0ZRȏk�nJbV�N�ͱ*�%x0Iy��ߧ��L������@���]ժ!�҅MG�G�3��TR�y����#���:��K���M[)�.��\��VoíW����yUZ�+���v,هj�Иp|m���v%	�#:�K�O�T��^�1��UK �k�
��j�.q���&}��Փ/����x�D��׏^��;�R��� ǳ�qUtr��G�03��,�#d��^��4r�jW�p��'�q0LR+�N��nP�h��ۧ/HtޛG�:DC՛ȫ,'�L��šR��EO�7~h|���,�,�ԒS��"IՍ����[�qi�g��i�S�m� 6�{F�k��W; ��@ە��&�J(�M�b����o:�b�o��@i����GW7��k�q5�f�D����δ0��s���"�5![��!��%͒-��4��ݔˤ�{�~
���霈C�E�MK�#��]����p� �C./V �M	�J���?ra3(��~G�	�x.%E���51Cc?2��,h�JtөsunE��#]YH ����`Y"�/Q,ߏaY,F�C��b�$���u��T'n|	�W��@���'���u�=M7�l<^���{�B��U��)G��d����̝ W"�'�kϫ��KK:����Mǈ�Fж�^������pC*�s��p���+��6u�ԝj�T`B�V�#\㵣J)�k�V�mB��+�����	���,�
��a���'���� �r}�|�z4����=X�]��L��Җ�Dn^��ߓ �qPy�ƶn���@"zE���l_��7����l|�;0�ErH��!�vW�GpH(b@�ʢ�%=8A	w׬q:'2���q�yR��xRj8�P�,�y��j:��-��h{I�Ǧ�o�������R�(9?S��)�Ge�+'�����z���n��7Z�!D;M���Z{9�D[)^�=h:���šP� 
��^��/��U���SaF�Xd$�a��۷�9�2�N����n�d�VJ��b�C�V	��i�Cݎ��rg�&�～C9��@ȅҫIJ�a��s�]��p_t���=*Dƨ��wLi`Ϲ�u�W��Z$������2��?��>1�{��wt.�{vX�k2�3ݕ�S*�iXq�$��v�gYӤ��/�:�A8C��Z~	�r����0L����_-ݗ�؊i��z|�C�?�@���<�ֺ��1��I��~��:R����a�?U5�w�K�na�a�T�;��MX�����t@շ��]H��Ҥ�ɰ��"<�TY��KR�l���  �*��	)M�*}���_	�s%�q�}�ZJ���-�nO�2��$��2O�K9�c]ͥ�rISrY���Y	[�1��{��rJ�sF8>OE��ڸ �����Ъ�%�	�ٟ�xʢ2b� e�TU#��G+��%��b��x�O�3l��j{���ݒ���m)�Ígí
V�H��W�J`�z��v�(ߺ�X,ޠE���Fzi]��s��а��uW�ۃ`�:�T��Lz��޴�����񝛬Fbav߲�����3r�@�u\��Q�khUZjtڹ�����5�^%i�۞�4���^>!��!���uR��f���S�]�@�8Hy��hQ ��%��z���%��Pnk�2�q��!�WR;|��F�����$;A��	P�Cݞ��t��^�0��<���O����m=DMH��w��K��N�؀=���I2�_g��2��-
�B�ݲ����>[K�|���[h�h�V�>��_���ػ���ߛ0����U,���#�jT�j"�GZ� �߮����;+Igw/Bj�|s�g�b0��e(�B��
.�MZw�G#i�����q@!�C���9kƌl3�-5#?$����}eX���1���v�QЍ�>�et(���o|�l�Ǳ�%I��w�O�y_�
�۩��Ϫo�	�鴰�ģ��]��q���OR�B�v Oי���U��s_	�;W���B<H��
B�Ao���B�7���9������o�n�)�� �kd�x����� �F���jDdKɾ���n�~���xT���뻺�)�B��ϖ����K����ֶ���Q�S����L��#������I;��~va
��P�"�ޗ뻧;�K����́&-��b���"tC"�*�@�!f(��}1h�{�m�Ụ�+D�8|�Ӡ���+�	Jw\����������kQ������ �]�H���LߙL���ƻMLA͟�9yF?"d\)a�51�'���Nd	u�&i禌0,{���d�4a��c�0hzMY�ю���|X`��`�������:�ԛQ뢿���B[܎`��` Vu���-q]m���ÑV����F2 �M���+{�y����A>��͗XW�����Yù����u�P�|R�2Tb>�~:#:���k=Z!�C��L{?6�^BZ�uv�&�bW��I�{`j�G3Q�����aY"\��Dږ�a��f��нW&n�E�A������@���_�
re X��'�=0����r5�y*���La�C�>>���|�(�נV_� ��P	�ɷժ��:���]�m��^ff*|N|�D�m���m�m�#$^^�q�XԄ��s�!�l4�7��o�1�E��H'�t��VU� A�{�۷0���3�B&�{C@i�8���מ����TSS'��&Q���?ƓQ���>��a���P��,��}D�����-Ǵ p8F��ӣ���ɣa�����X\������z�Mt�b_2�4����ɀ&6�3�%��'�*t�u/#����{�O�����=Ѹ�ZL���V�͉D���ɬug�͋WX�߮x/uk�b�?�.��
���r^�}+���sύ��4� W"����C���eX�[�	4Ng��<7�<݄?vo�>{Dۺ�z��&>|�g�p,��e��xWN>1��+2�,`�_�g�qru��%����6x�;E�qM������,⵹���-Ȝ���>"������ǥ		��
����oe2Yx����?+����wx�J�ժv>�ސr���%���ծW��h.��c��@�9x���)k!������������x9I�j���v��(��SY��dB
Y��.����Y|'�\�p-���xيkJ��ɍ��@M�}���% f��D3���6�z�d�F�5`��u\)��/��ƲMlkQD8�ȩ�﫝�Un��?Y)�At#ˉ��ny��Fߥ���JR<�����r�'&o �L��]��Uֽ�����u�sa�"�
��|�j��h`�$�����l< ��R�DTvS؈]3B8��F����M'D�#��{k��=3m�Ã4�a���F�M�X*t����6��Q��=�'MWL�!f�!��RѰ�vWdۈIfn��%9EN�����}��[=�_z��	d1�؃�q������|��B�{d��V��L�n<��{7_�; ��j�};��V�f�WX�}�Gǰ�t��3��#3')`�0[QDP���:�i��n/�����I粈Ъ��A�l�`"��1L�6~{0&��>e�%.(@���KH���̊W��H<��c?�n��ۓy6i���sdmv����-�8L���5�G `Gr6�A�̇�EU"wD:kx��(��X�-�|?۳k�~�Ga�aW��A�n0a��/����'J��1x���/�>���Z���[��R9XJ���U��f*Z{��P��\7���L����bP�fs�^ԧO�\ؖ�������*�-(�4��!�DMKݼ�m1���h	�f7��u`���)��R��V�Sb�Ӥ���uNMAjNc2Ԧ'o-T����ɒbX��U�7Y�˗[��A�+38˥�V��tn��ýO;N�I�"}UR��:��������*9�c��>�#��=h���BB�&�3�p�� w4JG�
�f��)�^>J��� ��սxrs�{�6<��7Nx�',�@#�q�9GO��8�|��s�CQ�'�)e�[�r�iV�H?�w��z[$QӻJ�ogVc�')��%�̂���o�&>v��e�g
�^ee�uW'��1X�|����ʲ�k]trˏ�śo^�$��
�e�z\��,�`���_glDΫ�'�fꀽ�����r�2}�5�5ҷ��y4
��� \$!�~,@�!�!�� �v��Ѡ�ң�?;=`�L�F�y���v��`�i��Tu�[Z�tu�'sװ�Xe��.K0[�T�T��0[���!l��UJaa9Z�^Ȇ>+�l���.��Vi�D���`�7.S�g�
NUQ/�t<��:m��b�xk#�(fe'F�bԑ�Q�<�'@�B�2K���o��<Cٯ�F���KV����
�}ZT�l�I�8^%\<�G��N������,�s��A�K
<G�!}��kS4UҠ�	�,��!�5y:L��6{c��CG�HDz8�ė��+��i�p�S��ϳE�ce�*�j9����/�������K�^���<%���b��&I|ρ�*"Y�W���2 P�cś:'��@�.����MUX"8��ấ���B��mG_�.����*t��:�Q�� ��a��+�D{�~��OaH�7�����i���O}�D�x��k.0!���h���x�ݙ��\��Wu��X�ϗo���Y��8�_�D.���82Y����JX�#a��&�ݒa�H�XE�{C�j�1��太ߺ(����8����B˖�@�BBF+�YC�n��Pt�_���oIqM�Ƭ=#k���Q��i4�e"R �Xoϰ��-�������hP�G0��l����K��9r12B	�hfW-e���uAj�J�!}|��K��w(�S&�6{W��`�I����QnFs`2@�����0<xPu�/��)�7�Y��V���R>D(wZw�An�m���:��EYi5��`�e��:���r�y�F��'Il0�48����->�M�cC����$��CR2����&$��N�P�r�"�aX�����V��&^!�Z��������\X}ڥ�=>d����Ɲ%KN� N����?W���X ch"<�	/*���U���M�B�((r�X�À��'9���'��y���mV⟍�ˤ�C��F�R�0E���M,�0Dm?���sK���">��S�rj�!���k��>��O�T1��c6�}�m3��(�RnU
�ޡ3D-Q� �89�\���Hn���JNwJ��Lʱ�N����X����Ew����E�  �
�G��8�׽؋��<�w��!��)�k[��#�0^;�ZV����#��[�>n+QR��0�����,ᣜ{����ϼ��~ƒb�:��l5p���R��s��9�(s�="�Ɓ�ȉ\sz�\#0-E[>��XmD.ӌWX��[�:cg�{��԰N�s,�N�Бbd��`SaQ��ie7��V���s�����Ֆ��i(݌
8$�7x��)���	ٖ+6% <�ȅ�Ű3�#dġ<�������h��=td�@!)8���nS�T�82��2F	�*�Y����V6���pz��hʓ�A���ٰn�̍�����#�vf�xl�}
�6��1�V͓�!����N�1�ܹ�s�K�9��49��,;���?.I�.T�S�V��Du�嬇[C�N��D[8��$4���	Uk3��b^N�;
hZ����f "�);�jhV�����v&`��Z�ȡzu�)x���eUC �޿�0~�2�u����<sW;0?�(X�]nI���
������6����ѡ̯ۘS
�SF �t~'h����O=R���\frݟ���W�wD�O}3��n� ��Dy��{�7Z]�QnR�j�Ye�+6)M@��=����-����*!���g��6�Y�)m$�}��g���׿�1]���y�Q�8��4��Ž�d�Tп��_=�'���i
�R���R�Q&Ң*|X&?��=-��{�Z�O�!B�E|f���H�D�o�F��������k$T`�g
�צ�w/p���h��.��[±�fb��ȧW�����G֫)b��oe��8Ep��5%��É����a���4qݜ�鼃���(�8+ n�I�p�O��;Z�p�x�
5
jS�m�U��YV�q,�]QY�=���Bb�0�Ej��-�QO*e�]^a,�f���?���0�.��Do6G-�>� X4�7�O�>������,]��Jg�Zf�Y�/�6H�_H�m�n�}-*�<�j]��ds�wmw�1h�����mvf2 �s%�6	=s�6��;]S�G �R*��N�b�krP7�c���i����T
�#V���.K9��$NNqn�C�g�?�_��[�7Ƅzn�s�肢˪&�T�^���@�:,��{��W�evο��ە�����/��N��`�C����u�s���y-����ZM�H��M?+�U���P�;�˚�����뒬��C�.���}��MCϡN��&"�K���t�K�o�*�jlD��կ)�8�ye��4'!h��� ���^4J�㕝��]����]�YP�ȳ\�6��hP�i�%�[a�Dɿ'��r�o�gG4�r�sk�ֻV�~o��gvD]��L����D�]��p�`E�%v�\�Ll)R�'�'����rP���RpЀ�iz���6J9��R��BY�%=?�a��Q	��,�q�Mx��'=R����1(����(j��C�  �-��E�i�f�|���e���	�I��R^)�J����y9Ă2Q����4P.=^�;t��]xE�1ڨ�l����y�|����J#���c�3��J�Ț[� ��t�Y)�N)�5Z���eZ�y�dC&���{�U���c� %��AH���(�ԹcM�a��i
�PV������F��]&�����-�=���o����k�u�;�U���0y��O+W�3.�r�!c>n���𢣪��j���
V���#w��Rη7c�0��փ����	�t#���N䐐�hVYlPI�AF��ĉu_-xN|�� ݿI�*�2���BK�8���ٿ�Sj�b������mC��t	�IG@���H��(NL�	M�k�R�l����{�4N�e���-�I}k�KSqG�e�$�6n���m��, 1�����أ�*�SS̖Y�Vgl�3��%�?
�w<�R*ߜ:�fL�9�����>`ƙ �s5FA��7����Wv�%�%?Z��iz5#	`cq	��ǻ��L��k4z��iKt`�&���Q��7E!p�c����a-L�n�.�:�Πu3CdC��
3�
ш�Ē�a�j��Ц��T�د�:�WBr�(�2�z,���;'�����+_L�YNHRx���*6A�f��(+��iA	W;��1-H���Ѹ�{�Ƞ��,�TT���߂��aF��H�5}z�*��+]6s"�Q�������u���,���a"��À%7m�}C��g��$öe�K�a'r�Z��Q;>����6�D���[��-ukf�g�K {e�} ���:�)��A�R�Z��Ir}�ŮîNk� Lh����"���-[��y�>L���Ɣ�U����L��bfߨg�t���c�hs�۾Ѵ�ny��h���w���>1|F����*��`�e��/�Xv�/�b�E�V��壘��t}u0e�G �U�&\21W�`����{�a�y���:K���{}�BL��_]JS׷�W2�'c�Eh_{lL��ї|y l�[��x� ����x��_FZ ���y;K�{@%������6��v����8V�������*��z|q���H�t�i<��̜��������`�F�T�t=��0枏���s��+�1h�1���!UEV�����4���+�D�zZr����e�]\������F��wNa��'�J,�g����%������ e����ʛq���B�����]��P젾V?OOcA���������z\���ۖS����!C�}�l��(��Qc��>�5:���e���s6]����|n!a��@�Nn�__T���bv��j���B��ٛʉ� ����|N��Ŗ����*�� x~��6��	��^']_��	�'�=�`,��.x��W�������U$��f��/��thV_z"�3�y�ާL�s:�Xp��;ߙV<�0T�h5{��D�0���)�g��7��nN�m���d�z�y����D������ׅ�w����`���R]"���05QV�2%�˫CI�K��Q�E�
�k��-�-��1;�0��[(KPe/#6t�?��c�\6�߷�Y�_+�h��L�i����Y�H��Ώ(nG����̊����/�}dZ�]�6�����Ry�����cl�0s������dc
%<��2G��K'tU^�zRo���Z�?M��o��91}޺�=`e�*��MU�%�V�N0@~s���YH(�S���PB_hW�����������8�8��9�+�q�z�(h�$o�D�����Mf�j�Ս4^�~�+c�??�Y�./ �7�ۆ`OY�0�'��̻v8��S�-'������m�u����^�,b�'����Z�M�1�F
rC��Э&� ��]4©A�܈�;�J�!�2*�Z�\�k�����{��EM/)����;�[br�%<
s�n�]��,�1��F�Y-ՙ�� םӢ]� 6H]�Rw�N�0������G��u-�3������+��p㣪�PQ���J
u�#�iL�:o1M�A+���[q�̌=2I���ƀKN�~6����^w�A�
k��o�Rڙ������癫��
(���OD���J������%�4(�m5�`X�T��m��~zG���Z����4�l�lb��tM~�|VHH�	9u��!�d��2�?f���]�
���4r2�ft��^ηa��*�\�r�|:�G�|��)#ĜW����E(`��W6H4#��?��#)Am��������g��r{��)�M��\6�",9������;�L��.�we�g� ��;�.�4�	��H�����x�㬶u�����{y�,��}�D4�uc�dR�����Q���l����:j��?� ��8�m�R\ :/�ToGy�H7��q�������,���`x��-W6Q�F��㪌´{����%nᡔ�z���|��2�-Z�F��K���@xk5�&ҭ��7G	�f�`�,��>J�貮�&E0$� j��,ŀX|d���e��̽�ւB��.�'Yλ3�۲6*�k���JB��o&��c��8���!���q�lƝ�l�ڡ�=t�=�$z�jߠ��&4����R�/�d:�X�S�
ZipGݥ�BK������4���N,P�e�[_mU�Ζ|�