-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
f0dqzlbdBlI2MvdXutgWv38jHKoQXeSG6c+gskqpVRhs7ryw3BsjyaAOAZmByjlm
PQRo6ygeE7vaT0sFYh1Si4VNgdrrxvBGX5ZoupsphHIwXksNOx2MI9QEKlzcxIjP
9Q2xEZE7DtAIjxoKjNCRRhafle5RB5+5zq84Ww4uxOk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 2944)
`protect data_block
PxiHA5UuNFjMWEb6inMRvROQGqntsE3AwsbHF6GT/ntel7Wj98PtGj9zY75oQgmy
bfMHPgWQnRXnSkiCnZagpFaTIQIlFZR1yUKXzD3h7L2hYtxMyJi7Y+d0TJ5X8zb4
vUzlJfVFz8bITYDy7El03TF7dZwvx57XGiItpWbgGr+Sy74JSbY884tGVj09yX6P
9qq8lauya6S9WOhqPhUMKhVmlMgoprQ+1tRmNVIOEPv+3smRTAWl3obGaV8W67rL
bCYkKEFhTsKA8f5km/W58YIkLCR221VQUDGX/3IrTtS9vhz6ozqi6s4ikOLQLoL4
TjfDi6t+Y6GWLZo/pu76h8ZXrqkccziUIVJ7GHPlSHAsuOIfo7IcC6KYh67TrDJU
sswnyab5COFaDNDZNYaA/dPPjQYxkbVFqCavF8Z/ce5sQ6LZ+t+WDRuCnuWTYWSb
fgOT6t9Xn2Gny4i6pqdCyxoW4j3hVc16yZotyQK76sfFiJAxdtbScNcJEnvgImfa
aF5bZXcyS7nA48WOXK9qBv+m0cLo6asPMqsvhlf2sJEJ9O40B1FRDbMbybLhqL/S
ByNvhrQSt9vbXTLK2P6IzmhLtk1F4mmRwVBzzYsWIjGTUbVbves5zzJI2mQwRye1
byL/V/RQr7ZfvPzdn0iOr+ITE+N4ifTFWIshtr16YsIKvF2NULuxYyBNAbIxHlsn
CCz5cde1LWWbDri5evCwyMYXEMQkG+BP3wKEIlgUSaOF22SSwPpNmBvn8ZcQ864f
ppvRm1PBiJgsLYAELpziZVBUdX+HQX/D08qrjEXgjqRLVAbnIDHJ6FF2/T5vSBgX
MN2oZuqMSpKet0Lq8xXizewuD4azOhKYO/BELrbG7J4e/aFPpXKcpKHxIcwW8y0t
wfO+k/Ny/6ZSahGKwNPzFVuBXo3UywhtsSJJ0E0Yd3ZOD+b59fHEgtF48bA67zUS
ITC/V2vhkuSdYGlIbgsCR1SgDK5zJJslXtv8RMR6n0NlwnlQ1wPugzFOoD9sBjrs
8jlb1VURRKqSzXQipUzvzgE1EwXC7yYrr1ZHoqdQ9ABKkEzD09Ssg8Ngv2M0eGzs
s7UnThRofe7Y/xGaDfEm4TKXxq8z752Zho08o5vCMHsvKEzhRIndinie8GgxuLLk
k4X9c+mVziUolkW17fXZsuW8XFbW7M2PT/IkD1o9vfj8PcQ0GhhkMU6rAv8Is1vn
DAKzBvkQ2An41rDdQfH+chs4gzAwirrmPzf9p7HlkOtr2hiGm0lmHNZSn+urCBuB
PMZIW6MFJ3dcO6tF8s8Gc2iKoFR5/GUp/epSxR78Ofvdu4usb0UCUTbHcTFq1ZGu
jtahclJegfNNOzmRjXnmvk9rxmGdJ4xjmNV2RLWnR+u7GUnGZVwsC7ps/YjP6Twu
xx7mk+S7mZyhMP9aFJQlem8FXzyUAT4xUrg/kxwX5U3j8UATJI6HQSCmnSFxNZBN
ZLAk4+VKwdTJlmZ0zqRi+0WtblQfSkcaeKPvlvw1OJDhKYCDUG91GChxiflZ9Vtf
e+oJZ+UDEVQkIFzxr1Wldt+19k8lvkW37ELiRGz1M8QJZT9JYA7EGKT3Lge9Orjv
MIRzN0WK44hcAdmSQ2r/wSuPi74Uaqn0tFtAjHWLqfDKo90QUeHtAm39PiiOp2Fp
MjZTrxayo5pNusX5XcP30IIGb5S2Bgbelzs4byRkGWltQL5v+qfnTBwUQ0wtRW5h
pxHLVOZhajYdOXEXi8Y2HQcsl6whcH04uYulNXM4qwY9L7VBOVkUW0CPidymCWAS
+Ig8pOvCYwvEJXF7/W65FPznmMB/eJirOTCFxGy43SWBBQTAhBj5IN2ffCX44d5g
Bzub1Woo61Hi96lOlWARZ7z6iWE2NcjDiErcMTWnSEngm2jwEYg62ZXEJ8QvKyi1
Z+4eRu+oujZ8uGRROd4hnb/td4EFZipHtB3NaeR/7/oQ/x961jsuzU3x5GCrwz1V
tuzasd5sX2UROIpyDA6Enl1CQosHlcWwgmqtYl4zmQWe24KnzrSy4bAUOK7a7iI/
CCxFzHX8VB+UXgDWnIU4LzIrmO2R/8VXPG92sFTIcExvXCRktAPImQ3VblNKK40c
4ThNnQv9Prvip7q8XcCrhIyjatOKZAGyZuX59L8dalr6l1hW6bq9vLXfRqFPn+ug
SBD08xHeEwHfeFObiewxxcxD8earMia0oS7u479EXFZG6la57dXBLVpXFJrwkrru
bzTgkIo5Vx5r8EsoQRli8HypL1f1cEx3fMGJJZB4OK8ZO3BmYc5vDzt6pPsMeBlE
rifOhV8XPhuC3NNTWV5XzTcODZVLtX9NroPRL87GKTW76i51zOjHH1wmfRzji21u
PABD0eeYUEaG75Gd6RDFMWjPE7m3iMiwqWVn6k//Rc2s0dpNLgMGN2fAkP5LIRjk
cR3iT0jBXgr7yJ7cEs/e+swkfkzMWDT0cYcX9bvW2FaIDa+erfRD/E2N8bBJzMNV
J+AoLCEaK/5a9CSyr/rN+wmTuDKw1NfrVffo8+AaPwuvChK1A6KHqrYDmGT5adHF
YcAf+6GgQntlyiUkGL8q4TdaAtX8nAd4udBed7LmcB/6p/utdQ0H0DeHc4TS+Kdu
oLXDe7osZ+RSK5dfyeQO7nEP5xzYoIvwjNX7bMOZf+zSukd88uLqAdrIbshCGn1v
cZMjEijmi/9M+nFClwxG8UFwsJL8eQFYAMalrkgC47iZwHLazbLAhbOdBy8HuUeb
29JioZ2Q03hH1NSHoaaj0QkHCyoHXUV+WEKJU6KLOfU0zP8Wh4XVLsoaxzW8NFwJ
36zERU5YbBSpfA8loPCK75CzrbV88b629GmS+7wgkgEy0A1+vLDXyk6k79hQQvu0
lAHGmRv/Uy619e2v4PbH0u+nVHFKlFuEo8y1gjnbkR4dikosLdl2QKWFCKoKCMFw
qY30EIQZ3uwDkfmd+MBC/GE+Mp9SaIIsvgbgNPO0fqI29gnSke3K1C7ek02T3t3T
22aYMCai+t3PSfXhbrF+l9rEeitYqMrqbTwcBRdU+xwwbv0Eqe+N9BwHgMMmfyuz
KjW9lsMO2HEO/XsFwrqbgyinrIstWemT6IlmWTQW5I/AzkquITtbekdhgql+9DIe
Pntz4grWfn/kBzmQjVMeJ3gaWuU4GhZxrglkxuiZGJqlWg/AvI/OZ7FbVjWIV7bw
ouaj2R2cI7rYXf9QdfZH1DNAp3tn3i10YZON0yf2Kv5gg5SO2ePANMYKP41Q5ok8
AER2TsT3UYJl4xEkfag1M0z9vqWiRJn7JbRHaVjNVwzgE0N+qMl/2AGzv0Iz1zUW
kwYH6jUUTfIyN5vliW+KJzGsQEvDmFRu1S+bJBP0cJqc0BIOmSJ/+T3KvzQA8DeS
aJjRyi2zNPT+1+2jPnzgGfvXSvTWEdQV1mAf3VSKKj3gRWZKhnn/5kgDhsnzaQbF
fVJcIcXtdOcA6d3lOHzv0V6kqZ5d75sF+/67S452DcmbbmVIgcje0+ziebcaCuXD
Ab7Y1gWGtjDsuhcRIpZngzmFHg8fuuN/Nj8yvdqiFmTOHDQjqsYeLdhs5kATtmFI
GjrQdWctzY6Q4+9s6567x8TW1Zg8YnRoSbtTsbnrT/tLrTn9Xn55l/R+O/cG+ZtT
XRMy4JsLBO9LU/Hh6eVer4ATEJ7JR5aN8SL6K8nkzRHdaMvoXbK755Kr4eeiCQGZ
R/rJKsGT8+wu4yAtmq9uiuaSm2QQDN0M+stqU4MeCMbo85OqP0blZK1jTiMT5ORD
puiwIHJw54JUOuZ+gWzLkAhzdpoTz9IZD5dl3X/lEALkesvyEu2LWwY/AOUtehLc
G5q7zZYn6bhPBwHfcWq85/5m0TmlHVN9eJMLorV7HQDEg0lwj0tsjTfnpDyiLH4D
aGs1xMDvTYawCoWS2UYs3g==
`protect end_protected
