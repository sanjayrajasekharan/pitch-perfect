-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Kx6k+aOAQ6L6NBncCzpkVoYbl+V1Npqkt94/s4bLEbB5t0o+U8HaadAkHXq6AuDz
F1XP61vxlCErxiMjkSDQCq5gwZYYsvIYridFRS7WMbOhi4RCSB3Aed/DbEdcvC6x
oOTcooRDWK+34GOE6d5GoHLdasdzaB4bpm2C2WSrfBg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10048)
`protect data_block
SUMdW/tVqRvhWG7waIweEqhcQpqBhpg1yzWhwVRqdKpZtD8NpoqW/sLZIYU8qYj7
nvAG94Z9aeoN//KbgYnUwx+UsFkRiRcWiDhFHqMx9+7Pe741RHshOimFCSKV4/TG
vV7TYHdafUEOhNZgBmEFS7lia3eiQPLleUOEkczAvS0wBxq0NG0Llb1NusBt5KQJ
pQmNmFNP0WO0W/GZQonkqr4+RAPmWgvh27sjYoR3Hp5uTILDT33TXFx3CO1QJ6eX
r16t2SPZo/jW1dP7Deqvt/L7x4STWmV34yqWYoEP9cT1EEi21XvXMEnM6nNCbr1g
edIMpL4VZGOdfR2mLnOzbVONmrFp6u25PMnWnxLoyGgKixcFBtuzj+EJxdMyuc+F
bQ2b+cgkQAa/HFvH5GD2pwgZfbo4l5wUHXEwjvWSjRZl6eZ6R5/VrsydX4kZ2GTP
X2lkD12k1e72WDB767QjZ++mMK2HUtNRpp1E/HtzYiKdclFOVHeyOwFK2A3pn1jl
brUy7G/ToGja4fvc/D+tqcEIvwS0z1veRiPJFDkJwxwFvmMq9O/T+DBfQeWYpZ9k
tF3SmVOUP+RmOyqhK8NivI9WcO3uI6/0zQZ1d5uvmGOiJohA+P1EHFAYQ3y7410w
WX/wbUQ61chBYqXkXoQ6y9sPkNl1juoTFlHRNQ3tbwrcmVy1aHVN3SRBjsM1PVO/
IG2uaqWkw0x20yax3PSf1dkXOfhJ+ct/BfQpvoLgRsHzfLxIdkTZCjwEqweNF0ze
JPl+cPFqCkyIz4HmtQktu1K5kYCdw+Uf16sO1VroULCPYSnpAt66ef4dPeYzhmCS
DcyWxkQyv5cDad1BRY9YoyewBhNhEAyI0LSa4Zf1MqEdKFGGP0IZHvq8RB7hJ8MS
gAKO/KaRfNwkf9rzKvzIoJHTH4OFuOJrAP/Vbxhtebc1znA2KCJFeh0GOFfGs2e8
yM0RNvUyiNOm5rozUYhZTZgp6TeSQkFDOxEsH6jykSQbBbZz316tQz04uD33sV7A
LspMTAjn1wk4oHqHo+XGLf/QrE/geHT0X52FK5CByWRSWxinVpakKFoGBtrnUPo9
7SfDVMmVdSDDnu1ZqscoY4HudSbOSswxH8VJ8LKt9sPg1EdsRp3v0Dn0NZsxcNY+
PvhDG4dgdMl6U7lMhn9zm0KKAJuiF6jIvX74t6WLUyOYtewa/zIj0/YeczcfIvwk
N9ybcVm+r/B8+SpNxMJyPZxa3lNH9VWYIp9Op0/tqdQYorpIZrubdvICEjEZr0Sz
3i0CCbWdixTxXreaB5Q+uO0ozrHJzgjjLRFtNLFiKo0Ax0139M30myOqtVc7t+Cn
24ecZe28Z45nEHTKMl2O8bDGvmoReAOnXYdpNyHM1aJkiYuXS5AN9MBUShysCk6o
ST/Obi8KV4VHD35Fg/+UzthtaErrTpnOdfXKhnuSarwIqZy0OGulmSpGc5kaVIvU
A+PHeoWfJyOlJai6rnruS7++66QxqPP8DOZltIwVRfNsXEy29F4hafrZBYHBcJag
kHZpIQWY2JDQk5hOJ/HaecAP/V/UapeCsfBus8F/qOD1LiHxBmVDwvumvnn4qPid
GXmbatLrmcPegGgGdsOI+Q9QHI74fEK2FqqsqzbkzlPvicMDWW6d+DIju2Gz+oOV
+W6x2lAAdnR3NZ/iUWrJ34SEiqrVVxgzbPyWzuCguxwZxmpfE5GY6Qoenk5irxYU
4GwwTOlfPYUaT8UM+Ze9F0mkIgwSxrNJT3u/Iaqlyo45IA9GqDsUpNUf6MPoiOvS
97zNa7oFBNGCXViSweBwpd6uSnk57n1P2elzvDfCHjbOqzIvs38xj3FxrhJljuuF
mBYObUC8Uh8gNs7nGY6OeNMlLE8zZAanhUcYi7sBSXdUcGdrAFd19Dyw8gZ58STQ
n7BRR8+fHYMe0JbSeLOOOX3ofhbvjsr57OoQXcJh5DswWGdOIZEo6OFersgcdYiz
Fv8NKS4UhUzx8qpn1hf8l0AuShQHrwxeeod4b9HwrUX7NagnnbEveD5QjDcHZ68p
KsuZQz8pjh0LDByTMa569wxbJhKEWhw+SkqFRgo3w4r/AFZs8YsyB1SSD+65rzdr
UHtQS+EmDAXrixILSbSwGFNVdXJ320Xxyh/Zqx0Q8zIVjlZvk4cDJMvTZQBB77ZP
d91kmjJgyExNxzU+LCR9t/OlSmXzKbkIni/GfyzNOAH+KJEkPtNxOlGE9EYhoQNr
EMBXm8K4emI+lQG3KMI/GVV8FEb4WXLqzMwNRM2BDUN3X9dQWr7x9HoXm6mr4JWf
Wftn/bwqxThBzt700hn/gFAtd6z+jrvONl54pqKfdcXQUexE18m1qi5y88UjiINC
+FdWjXweonsXZrz8HCN8p1pynacTywLF879y5yWRstmHGyJ84vdmFHyrdKWCAdoX
isWd5E2g7zgccujePKFd5avxxtL2L8HSE+CHUz0VkorZgnnDyXW3ZO5pD2EgmMrZ
NbHzk550vTW6aBxU5XB7u1lmScC3EWIsSNwYwYl3i8OreSZsTGqgsbYSQR8Xl7yJ
yI38JeqMcXSF0G12ZvqrGWmdB1yq3fVi8iSEHZkoJ00IEUQKqaaV1/CMmr11APS0
+qwhx828SdkqNSo2BHJSNIcvXJ+oq2PUq6u3cBkfd7/kVCjWXM3IRTmCYOkb5S4P
rQkdp/USpSQzjcCzg7VG5prDUQz/eGaNelysS1zQUQyJgqQB8+mHeyULlg7PzbUW
ovToKOYS86VE0zPBqMYqiYz4MnyBQGRxlJYAEaE+rv97GrCT2LbdFaJg/fvBi0n7
I1YKgBEpU/LKOYNjLB8ks+NNU/lSAPbazuuQULau1NKfnEoLtDNc8NDF6ReptDYz
TIlLQkkMfL5DyfmaAW1XHll+HRh9qQPIH39pVRPHug6aIAGbCGVp8fkPudwTwhVW
vqyLm1wUeINf0wEr1eGIj6awCNQw2IWrdmLFSEEG71bHRPxRoEuVKlhpN/xrkkDq
EbeQ8VPkZy65GkcdcBa+RjBF3rBeTS2OGpugXi/EY5C1P8ev+imgSHPHKYuk9Kwm
/+bfy9rrfSndqISVry0zu1F8aokdkQ4Qzl0PUNTd1z7Gw23GhmK6o62qN18WCTj3
3MXtyDIR+QKnQEIey03400cI6Wctl5bTt7IHJFtuP2ldnDQ5TnriZyecZWM9zyij
1Jw4BduMlkFdZ3UrsgplSoE5Op6jiorkF9Rg6+Eiq0zNKpwvoHVip5QVGPvVzGcI
hE9S82W1zd76Xa+AFff3BRUzI+avyZv2OCqsgKUJbNT9XfcXpOf4cfVYFDJI6tPE
KvqCSg8DdQV+hPNQhxzP2JZ/WWAYGgAlJyFMfZL0n2G3pb7BDCcniNqLrDqgs6s8
3/il0o3aK/tmt1bg+R+T6AIdRElLwt+ffA4Xc6coyCeRJ3mX2bssFn4/2iw7OHFy
022F2N4vclIpHiTHXkWOOPCJ2cuSZ8CklCYjNO/2DWsq/KhwqDFLdNoCe73jtfyi
ZItZyoh/oBbc4IwIV1o0N2Zl0AM9NJxRGgCaU1gq0YMEd8jYL7KhWtU2vdujWEpV
4+WMO6kQzV+KOQaQLuDw2SwkH7kB2LeySAffkOqVKprEFqPVoLZ5ukgPQ1l0sAuR
1UnwQ/fYXKHHlfZP5cYqao2Zn7tbcYluOHQk1jq64rcbnFHpWYasLfvVsoKjXVT4
DK5OYubkD1w9eJci7FVUOcMRaXWFvXTKs7qnZqc2SIswB0pqfKJMVVjYTssRbvek
qoyiEQynXEWkDjRc7dN8nEB1EUAZwetn1ITBOSeg6MXehTFrnOXUdQZbh+4pJMWv
VRjzsEBgzICCLXR9C6+2nwszRwWfLo1YVv0b1gzEIO6knsyDr/hP8q2uOkXR/3Wl
ylasSStQ/yYPU2Y8JnAC4dtv4hsgRIaRIMWSYGnSImuCqoqu5jtZign4evrKBSvd
9zGokFz3qzqYQpDvi751INxYfFf2yrZqLu8mVrxpMaK3lHOKGFFk9atEje7m9nim
x44CsMpo+6oE9x2QEob8F3R5Mx4EF/dmpMMkR5+eMOBSVw0PXRW6bodNj3qIXVfD
+oS/tPb07T85F0Hqtmia7XbB0rC1L8rz5nWEAPUy6NhLBqzVViS+xRUZh882+NG8
ijRVXOn4Jot69Kzct8qIqc1J0srvflvAJWuU19C652Bx9Qh1JeD8woUdPSOZDH3k
WtsSnjneATs21Iqa4DSbBt5l5D4a3x8e8KohXRS7YptBzx9q3y0QOqrjdQvvxm4h
xs4NrBHDXeC6dX+exqM6Pel6THBgqHAZK+mn1QyemBox1A5P/Iir73csrWbqNbra
IKz0OkUpx2Nq19htnDFWuCSoWfspgGqNiaKuK7OFT7xVaOz0Ge4p/fSBpY6G+flw
EAPzfpSL+pwt41cXtYV3wbZONBg2FvOvB+UvkGRE7CGbAkp9z537+LikSZQNhxzo
bkIVbVRL19/AOLBB9Os6N+uFnVBEr6uQHyvgovpbf5f1lXPAIjk2tDoUDxDrSWZ3
cZSz+y1XbCGK9j6BqbirHKMtUTcDWuCX0pHGZNWOgA49wjjDKq9Q9PT/EyAl4xls
2va/oo1Gs8JrQTiOi7S/IhKAlZBR4YXKJyf+y94i1Nsbm3ZAHWkRMjeydSFoQkUy
y3EHHp5Mewv2cSww/Cy2KAU06p/QA+GBCH5WdUnAZTvxWk0fWp77Wr30s6ZnrwGG
46ju1hbnftweHp9Vzy/I0Chl+guhrxcLTuuprCpvNgWBzzcKaUyJcJW+IcDMMy9P
ZlTdQ1SL15G3peOPysghFlK3aW2S21RGd7tTiFs1I9KCiGFcD2WYa/qjhYhKhT03
iWPeOdGzXmQPX0lc1W1XL9aWA7GvlGy+CBW0yYhkeV+JoWaGWkXqMw1G+NNXXvK8
jxnsJqzZ4L2JAEutmIULkA3BrmKH/XThhopi0otUqxc1vCHq9NnqVlbg0H8ZCSxR
bTvGWAe04es7Puj2Os6laYgMs0KCt2exW8anUrOUP3lscLPA4euQpdlwJWPP0n9h
S9+8JEkGmXGF0zGdITljYWIZPH5JvvxdGr+Qv6xW+L0dnRMpsUDatqr2kz26UcBj
SQQPlQNPgEOqO0dsmYoXgWylrKqr1HpB9a2Jtyj+oOnDWGe2rR9uzC9Qeut6M4iM
pZaKprc8l1ygJ/P7qgTVzSgJTQDJ/AUnDKlrTaPUTY2ZUB08KI8GFFEnf0+b/CIz
PfkM4boiz2IVgIFlRe94am7MtQ1GZd4zOrH9Wc5jqpfK1GuyKn+8D5LiOqbM7sfv
B48qGP2iyqLL8XjHZM7u4ATTxlb+4jc0/mLp6XrHtyXKl+8YLaNQv+MAczymt/7Z
3aSa1Tbe5EYtjVEsOhiBn9adt8orYqSPV7azvWff9ZeeFyR0Fzl8wJcIEqVkxqBi
kIyDSv9yJXwFYEj0+oe0maVA+LIAPg4+vOfzFKf2AIT91EA+y566BeI3ERjVLas8
d9UDl2tNI2tl78GMf0v0f8Jfk9axNX7RuyJ/mP9RYfiwYJNmHVfbjjW4YdI+A3ml
FfQUNCFMh0f78EwL8iHUQ3TIbqFX50KE9LceXpGBUmMXWz47FmTRyumpLgtpAxsS
pU4s03VtJTd38FT4KQ0LD9BQIKRqk4sRR5dKxohvNGgg5XHeSWMNL1EiKQiVNU2K
g+/TSLtdy20MfzUH40kFiRlPKGMBM9VJyuusxl9nd2/8IUvCH49QcF0FvJ3l82gB
YB9I9o6fSrHSb7kSYe8F0rT/6cbQJjpxsg9lQeEsfrzLPy1JFXwVgonNL1VLRqvb
gidoq7deD0r/wlIsE/IE2+5ATWKbT6Bt0V8MnA/LSIgDJa+KfdQDOFaezu7KlMeN
vJ3RmRA5hMcFkNAtqmDkv+wGTzqE8F2pRFuFlYu8qn268xyd7RA4ozcnU4GhgFuQ
S0JqQ+im8MBYubg+kqcXwn/88R680MBvkm1yUFtxwcCOf0i2iasJt4DEroMp/fNd
MElnveKvW6gKa4OcKLA5uimBQ99r5vlozJsUSNtcvGQAPYSjNpbyffDCThx81jjI
4CAHRIFQw886+zOfj1c482DS86f/mDVD+h07nFigR9jaP6S/OjMnYOozEN4gH+lf
qoSNwSe9VOeqzfRChrTo+Q7TdMkk2ilhO1b5d8gCU6rT8fu2NxjKYXMdIXyzR/pM
KvSj7qTxmOkcHrvRq1GHdtlLEQxHvpBjEXMB9bWKXQjbVchnQsRF3vdXzOGUo5c/
MRApT2jwUiuOqqVdHwNLD4Ic3+Kd3N5snkP1aExS8vfASy38yvjjieRgcpaDnUWm
nMvtwcTiX7gWE4IXmO1uH3vRR3+GVo/aiirqwg4xot6Si1zlxWHAu+oqCQxcWWnQ
dA3Pdi2hV+kc10LOqK97IdBxWlde9tj9OZcSttvp5HateJwaeYXOYKmIl4eeMVyP
UuPRL6DM2QZpPgcPv9h6wh3aMSSr6GfGY2q4BUf6Rew/ekLzqxRiYjfQu4gs3bby
sWT0PAS+SmuiL7topeKIj1ZQgIuthmfyO7AYccr3hj/fMnASRdxbN/MBZbEGHR1V
bvevAOWNvIdzOv8G6K4et0FqrVNlMRaIsUbXb48th2awlMcYtImLq7/RQfKoh5CQ
k7vXbRy4cRCYTtZw/AYxviB4IKdlATf80BzCC2C7RZ732qQnBXULYIw0BEx8aEis
kbSZghvbGkmqNhQos4UJEnIWICcTiminq3TgfCkfpp/3gUDA9bftsJvnFASaccB9
qfjhw2wtYHxti2UGwHPltRgiM/iS+ehzKOe7Dq1LV2qyN/DI0jpUpgG/Q8Osci5Y
laq/DZPjgsj94WrBgarOY++gMdW2BgqEOMa3akupEc9S17bFugene9ZlYnVFthhr
1nc02WkuBMcx8+e3YS95ZUXTtR+4ubxK5tX9Es6mWuZjZZ2XLYAS5paRRUpj2L/8
UG290uAT1AiBuH+N5JyOsjN/50RdQ2vS5a0M2Au7lZswfsV9a7xUAxgqhuFFmBMH
XhGoIdz+MfgaL0Ej888uhI1HtJwH/fUyYtpH0nYmUMokoHyOY9l9AOmnoKTNHABx
TnDk9GB28buNR+J/HZ8a9UIboKB3Y/a3GecoM8uALOt3gJya+tUllCk8EX7lABa8
PG/bvYzFTnevNA96X+3s9ZrJiwy6FN6I5l14N7Fb+unc6uAI5x0HjrfUBRzYYmPK
NZxYMr1rLG83n3QFnlpAuvdNBD9SuS4Bctw7tk4rN8ud5A3DLT//eoK2X51pkk/d
i3gXtss048CIeTqr/4gFoE6eqv/SLGaacB3mP64JfY5fOvFK5GoqWS46vFxXLf20
slG/DRpQ0YKz5Vb4C7hF/I0YcEW1y/zPAXmQhUBVEewvOLRcobjdmHPEaNrIYNON
XxhOvhVIQZE4SEju/q5kL35BYqbYVAgF7Z3zu2FNwzV5k0S3aBcR0A4zpyqe4faT
QMTk7U/zv3llihRxIz/ijgSx55Q0/Ai8JV73ZMmvqLknOKlq3T/9PzyOrnDkipS9
r51cxoFVxkKiDUFQbzP+W4qnAc9H8bKJn6+Azc+ZRkRSwtp5FH2M9lCFOs282pDh
/+pmnFKACGRXdyjojAbUJZmt9S1bOKkCPxBFLeEjN8psRsUb9jFT8Q1MjGPNj+JS
ySrTAiGnAkGREjEexShBa10osrgCy3Kda4Uem3bNuEinKCUJtZr8bDD1pB7CH2KS
tNsxAWMPvkIKdYeK44uyQu0tgvNTWLtqyAdwV+wXpgtB8kqFYLs0elvZOTiSVGFZ
2BQNZLtAmZEwcccagBa2gS06LKenDt/oNXkXMIQLQRcLqm9K27K0VL9I+6Rmenc4
SyVFviTXcGEt2UrFou2p7YL7RJEcZlH8Q6NOdiooIbVd8QD27oDig3dT9ftsrZpY
7zq+s3S8WqE2PnvRtZsQqkAYNAj3MGw1Le8nL5YhbXopAY3TpY9No2kt/vy3t8L6
GkAVzVTZiCvMaz9mPqC0K6xkY7joSQHV5R5gH4xW/eZavG+gp3ZGxZEjCRbczLq9
pN/Oa11z9d/mF+vy2aUFpfwVXYdZaK0SlvVdusm4iJEtGk7VIqHtNUMf0/JOT/qT
7w5udlUT+0pCYHDhrihHVqV/GUZgK1wfj4Yo3E9YaxoiLVs4+BIPi5DhAiZ3wGCn
NGudvo/PtVjQ7Be3rNfoeRnp61+oNHcgfEQbEmny+9535YQnYm6hUmCKCXFhaFQs
XJ+BAu4Ic3bt60psFW6K0cV1z2n1x3rm0SPLCJU9oZJSHFUxu2m5qMlNCo3pBKhg
rvFUgUG4tk5iuTzxeGpSqRM75mvLewyTPCfW8dbtWlVHVUd810Y3/CLMoq6uvuTK
CdfK2pz59fTFuu0VB1isR9I3aJUqwWgDo6FjbTt73zI29oZWNS6LpRMXoU9XbRga
aGgSOhCuiIquvh2u2F5oFmQ8g+Z+yu8YVIRkMhSigGhOQvFrG8ErPRBYKQqDplml
ODG2wkbSeLwv7Kd07E/UU/pv5XjzurABmET8jko+kQDdoE450RoBGzuwbOTvND02
jhGRR4YqACbOCl/mVPvnQVcS1XRixiEZyn2n58un9aCkVYvLO5kHo/+Gbb5U0inq
GBugJ9wjMQL/2smXXAEz9RZl53skoYufzTDrtrzFOZBRqSApTonqzSh2kklAhl80
ZvvqCgi3vgmhjwEiiRGtFipDnVrrFvW8F2D1udtDMC7LQJRUTwZLo8CZ95OluGtt
YOiTRBfZ97bnkH1ialtSHxu77NztUVBsCcHkp8/hmOU0lYvooBeXfnQ0Tidw9TAi
rf6KMPhIHLdIPoENwi8AtqR4gEyeWZv2fjw2+9kgoxHP1VBedxML8CKut5nnpXsj
1a1/OYBzg/RJ8aC3ktBJEyBmldO2RGzm6ffgAPsUNhFrD6mr4SS3SiODV4N6844F
WqkcvGwrf3UzZePN2YlR5pQ7T9Pg2d4pno3PDsvJGcwdXYhuw7WThMOP35wUxzjc
AcOCg5WexmGFadwrepra1zbWv4TWaB0RyxycVABlvG5XO1muQ5XwrvHl+Zr/Pnug
zi2yqF/9gELpuuMTt4QQ+vVxU94m/b3OU4zyL5zMJUaueKBDsSiFLaDKzi3qHzcr
hWKUhkKcs5V6Ftkr3/wZ5nIJv+j4VLIpZwja9IpVsKEBSOhaZKUV9NM3BGk+77oh
IJWI54VYQUySpxyxhhjiCFZlYrL1VR+QE00wai/R4YkL9GSp5K/5obGt7XaFNbF4
2rsWgmlFYPlYgyHhQDxGVryjcP7fiWefVuaxe+fSvI+zV5/EfbXbeXgBtICxHW2C
r13m/oojlPWOUA6gaPIfxudXGnPdZ5NJpn9e7+4SevmFij7+vz+FC3bdu/Y+IQtc
/XLI15OL6I9Ld8Jisn+PKjkqxN8/RLF/0wTXiqejTCarlykqLUgfTPH7Uav9dGeF
/u6UtawKaDeYS8xQdt5ESPJIdBBxIjRpc9U8R5dz+zQvykXIvZwsmjIz6Zu9S8Ku
xyn9GiwcDjr8v7OoPOvhmTUYasv/NufdCjn2ft6Ao/nXarpXkCyVDRuNJu6z0lkH
hFerIhQH+hfBygsQAm8XQ/SyZ93BiJW1R0P7Rbtxb7SGJLj7W/8e+9mrdSgeXIBM
yTkIXTJtcQ9WcUQSmk/l6spC37NWcZZvbNlMfdpW8h9W1uwjCB82KF/mWSxKb3SY
2VCMlufYWKfBC8bz2rIdyX8+nH8PfkyrXop2Jf2WqKI64fupozLwuxXf2xf9Cj0A
BxYXI9WNWVyvHfaGXK09ryGBAUcz6P1EObUlXhirSxjqvX4lVClvTgQYB9MVO2dF
zKVs+xmbc70aXGmywIL8sqZsg9P5TzHfmWjrKPlElOjbXblze5ct1YMk6lRn+sTG
GBK3AZzig6WAkX6e4ggBnjqzjPxUEQz3cEWHp+dH16kevGZDCcv66kRyO6e/dh2x
fHkBUVjnT9Kv/pAysGkQLZAK4GJ77iSgSNlaFWaq4IdPvFY09QO9kSxWTL/dtf+M
n5qU4CtFyk7cmGgTJjMRktpvRruH/HT6ivsWlxwq7ngiPj+3EZxV8T4R7V8VANWz
5e1YC7iQcfWpx+k3pnb58wsRax7B8VmGayEfjfwlgG92mdEZ+Gn1EeT2RmYHCqUi
fqsXR/NPMGv0Y9mKyMw1tkNAaPWf75tyEpAHbF+iwISlkGZbTgp2SM+vIbnepyoy
zmQRORqoy/7MbE0MwRHfioWQ+zu20JlcBqI2gViRuKhJ6dt5tjD4hytoicOnplwM
RjzzBYziNU1hzicNW5KeCBG90fmpajWcVu3vkEy+Z8HcCWn9XHavjvgtym77fhCV
Zq/EXSprv5TXh4i2gEUn7eP2KgYmUT6n1MGsdMwpvBSjbZXB5WfJdLpwDPk7c1m0
jFf4jSSEXDLnNjzklpQhjCcQM1Tkg2YUgm76dKdVeh1zWolLRkrKYnlLMc+Q0RK0
s0eVpHtxl6RYgFZOR29ML80F8whUUEyqc6Fou0cXtiNOmw8bEqB1BCImhEThzUFY
5lwspD1jqokdHSztEa230HYhMa4W64yS1dC6acPHSg+oy3A78byXr5jsofAzFIwt
1JoV/oHVSvYiC2ubu49cuMZ8aXEYcqBoW3Z9bUhkyuUbGuzCiDokxjH0n7HZQEtM
8TbdCoys7wRL/GQMSUbVMCUmY7gx1q+vt49rG3/09sZYdFRR7MKOVatlx1X95FeO
qyjvq24PYhPGWWeE/xRnZrCpPahNT4N7Iln8pZqCgBCYDR5sWHXZz1XOUYfCi2zN
5MmdQIyZC8TEo3AZxzdSAxkp8pcA9KXo+KbRD4dsZMUEyfFu94kZj1p9lTQwdm03
U2YPZNoe4THiggViBq8MDkiO/LYSRa2K/qUeW9yJmDhJESa4epu3DfZWfC3nN2wY
Oxi9HXzaj4V/k1NT9rWjB01BisrvVY9FrReX5c4I+khIlhmbgMD3ao56iuZcGvrY
/J65Lmr1dJsg1HfB7S+tMy90VYO1hVVda941+Em8C0LcV+FKQ9f0ediIDkbKeaf3
ZC0JSxE7LovJmtqPxML6Jdmvw1cQRxGmu4rHM8yerU9lx/mKPq6sP6aEUF9glGqJ
TLPAPtRlbUyZ22k8VCgAmOtJMAW94P2P13fd8UvmCKNnP8G+P37Go+tvVGIUai9E
xtbpSj+dA/lw3R/NezwLxXHnGgcuSkSlhodHCSIL0DWrnyxuUS9jASb2Q32tRTRr
H/yzibpQ8/JiMRub/qd6EkJUeU3PyIJoynGNWocaUmICme+qjOaHoSuBGolMJYgU
/YhOpRqEOEy0BRAOd24LkOAuVhsHInMbuRqo9iYesF3QF5qb1xqpChSt3h9QyfIH
4SD90BDcWX1tifFfm0+exTllZBgEwO7qL/G2wxxm2m8PQIELLBzDlEYxV47ml48n
NFb1gCqtO3tr2Lqqg45DHbMoOmf+fgx+9UrQHC/Q6nfEeMvbOJM2eP6VZM8FMsM6
uO7ycivcxwpWULStTbLojb4qOgeczT/TOmMTQYPF0YGBjBJWwwS/6Blp1NF0N8DQ
UfUcCcSZ7XKCD8aOd2LH+oiFEFpyiufgjTNA/quXt96TGDeWgcufm4ON3WKpFQ4Z
BCIpVLYhFeTelQlXlnoQb6/2xSw/zmGZEt/qeFWN030jgWVSImUTRuJdwTYY2kZi
xa1rhHqJXb0t2LnnijoL4ors1nx0/RtbEhKeubTqAp+B7XA9/pfu77woVPYWGzrX
cqSJsycZ7nzHN8rRwa+zNLprhPiW17nVTWZvzHI/8TrctulO+cifLcDL7Z79R6ln
aNrv/uU3kvBDZz3bapD9/xLw6NfNXsI9T9s8oeP6uhNO1QS1QxIawF2FXaFfMPUo
e7/14vP95zm14YLTnsXx1qvkXDV1IlsR6sqCLXp8r9r2ArrdD066fXTGrcUxww9t
eHhovK5rQ3Q0WscLzbkMoGb0nOH5A7COH6hlqJsr8BQRxiE5pa7K7p8iKA/8S8Vk
TcSzx5jM+/t0GPDWu+s2p66UIdGpiNo9SIi0POZmyvnDyRE5EGHsISaROxbJQhBt
BS6U9qMrVdzwJWXLX+0wPbUvkMACd4Ns/E9PboePxc81gIIGZemI5taZXDoy9Rk4
W152gxIpzss6iwIjFLscD/Mr89GGzY6iYhpvyLJA27LZQCCgBdzIKDH/3RqlTMsP
v5GYkwjXs4/0jO1B4dq7qrFP39v6wI81C3M9BMsM51UGLbdHFnmFfyAZI6Mts9Ec
oF3HFJaMXWoWNyuanTfk1AoBwRto+LLlLhnNmMS+bukJMe4Pl7OjchEg0RGnrvYf
WeOJkYcDLkB6Te5dNMbJALA/3hqENeH8DaOoZINQYCeXjnpS7mewbYEd1cmFd8If
21XtntBfl4e0fBnZedgAP88+4H+MxHZ5m7Ie+6Zhj8zlSTmbw7lixXETACxaZ+T1
+OgGfNWxuq+AaNZ+r6lYVr2hrJTD/Rc0CdNR1CkaDdIhOiizmmx/6B3qt3IDLMu9
DkGuF9nYLUJwoWkrefHV6wTTcggDdX8f0pEK0Rk8B7PujBXhmFWAXG4QnWRsL6+Q
wSASuOvwA64jmgx712wCfvTQ5m/5/Xp2E1gi8tosJ2CHh/CUJwXC4LsAipOMvC/2
hNIhsDkatZ6VKaEPZwrzZUvEeDldqG4qHXZsgamE9YsjY3XUKawG1qNOMQpPJEkQ
lNKvJwGnN0PUjoo3UWI/wRcyVUIvS4tz/dN011qVYrUlVduFtcwaasBr7s7txvEW
Da500hXK3I7uuJ3j252dbraKJp1DfVDmAHPvbQf0TNcrvHlLFMGZ0WteUBT8TaJS
svW3TNBbH3X6wRMdZvIU+9FYJxa+tbFz8Xq3O4Y/yImePtQekrQinCJ48lzDmUR5
UxkUas81RgkCcTH4acgzgPNxa2iEbE8gQ0C1H+FVnNuF2j2oJKNQH9zPfsMf8Y2M
EKLkGpiHYL6wSoYG15h7gqYvjRMCpvOQBIwcJV0GEWlpaBpX8/8XRK4UNsoqaY0s
oO2ALHX2reyP4fZ4H7NbX9J4YFL+gWptkupSRZ0g9SmHB/bzf6kLFd6ot7vteOYd
a3Rs/V5g0kUlKIj/dfDsI+0+FUN/wLzJKWFXFZyVku9cmC8SV/aljPGYv9oxN66Q
DD3P3X+3WU9CjRwgz6JVEQdb/ah9ATYzIpqIMX19Y9bOoHxAYzZYht1iIPIhOEi7
GUpXwpxqyo0ry+zyUivQYsjQgOwP+n2L0Tj1//84GufQ9p5PfiARu/xrAzCifoDK
H2Tz+Ez5CrAM85KCiWtTTOJ5RLzpEelRFTBBSoAJ7H1xM2UfU7tKijd5Fxt+Kuwg
GgSPKR2LLWHWdCfbdeY5kA==
`protect end_protected
