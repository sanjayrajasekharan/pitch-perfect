��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki"jLU�RH?�|
a;~�ek��3"X���!>�����f1e��9����oe��tX{3X�� лi�׀?�T~J.�T��}/���F��A ����5i��I��� �1�gt��;8���τ����S�[�C�7�x��t�}�1,aa ��]�����
!�0�1�-�����\E�[{��	z��ܓP����:�����x7�'b&�HP]��Eʁ �/ ��}/$vfN�h���@hk~ӂ�*f�i�:TW�q����M�9�Չ]0> ���隲�=R��8��'�S�ߒ�����,��/�F%{}"�?R��dB�B0֩� ���kn;��������o��Y����)�%-�k���l�@�݄	���8ġgY ��G����pU����D��.� ¢D<5�T�qŎ����ҘD|Y��)�V4�L"@oU�%�Y@+?��E�@_6n�K���tB���R���*a;�Y�l��:ɇl
�qi�"`D9��h[�a�c��Hx_b�B��#�_gfRv�`�\��T�}����P���aJ��9���W�h`Ã�� �k:}۫����8h(��< �K�v�dЭ����B���w��nG��C�{��!]N�쉘Qh�
�ON9��:���$;�������B4n$��P��R��ßl�Z=$���:]���$���0<Zb�C��;]w�I��Z3�9��ʀ�1��m�I�>X{�&�t.�1ᥖ����|y���?����W�����*a��dv:�"5K\��&�����f8c�6"&cF�]��p�bD���?��8��v�m��C�nO
����[�3 !/d�ln���K�Ւ�Z����Y\��I^L��E����j�l@; MXs��z�pϿ�Y�9�9;<ʺ�ʟ�x�pl��&�F�?{oS}i
���UrMg-�o��A�ȥ��oE�'���8hi��WJ�o9�@\�6�[ݣ���t�:�n�]���\��Ma��y%OԔ������K�I��}��:�H��1��Z����E/���-ء�~t5޻������Ʉ Z��P���7�#q2w�&�c2y��Ma��N�3+\��8�����eS�[����:t������(!��B��4Q��д���Z��_i�m���Y���D!�c�"��Kh���φ����r��-0���~+�0��3`��V��|S�~�p��^�*�{���J2��߱��D5�ll44�����^nc�mϓ3�4O4�L�90l�%��v�%\dS�o��O�Ű��7�����_�3|������!:/#�9�f���[��0T���KT��L��լh���������@�&��w_���i�4?��C�fw��!�k�2e�н2�e�x�7��R���E¿3�=�@j!1�6�@w�����0�3]v�a4V<��':&.y�����!�qAϋ)iu��%W$;�5�
p�13x�[��9���k?��.��Sϐt�V�(���ϚBgaBN?�T�K�
��>v<*C�U�ᏻJ��� ��w0�̢�o�����ܻLA����t�Ol���\��f8��䛏��:���+�(���
�y_a�0��c�_l�x
�E�V�Is�&��\�;�>(�u�����[���X�Iy!3Ra�RM�	L�G>�Јi�UPp��(�9��L�g�l]A�O��j�L��:;m��C7�"�>�ƕ%�9�Ɉy�n&5���l=��C�x�����`!��tH��G���\�o? �,�'��!;A��l�a؀�dGx���X��4�
��J㨳���H<�أ����Rd��+;�f�{��8�l7�R=u��#��\b��p�1�/n�s��c:dn��ր@Ҵ(�Y�Y��D-�	���+!w�1���A3�H�T�����o�}�ɻ�锊ٖP۪�ϰ���������V�|����ͼ� �]�O�b
���D��"(�R�����	d^	�������|jz���'����Β�C�Ox��Wj�*]8 Ϩ�Dv:�`�e>=eםG�hr-���,�|�#��ޟp�
�
<'��^�l�	�<T��-�V��6�&�%�U��.֪���+�蜖-��G �L8q ���N� eX�J@`��$�9%���&M��tC�f��ﮗ�j_��H�-2㥐F^���c
W`�	�@���, �u-F�������h�tz�	K�s��X!�F n}Ji���� }��_i��j/o�����`n9弁o���v:���A��Tm%ۋ6�����D�9Pt��"�/�<�L6*�i��dvE�S�j�6�� c�V��s�Ղ@�sQT�0���)��o߻/�J�5^���OQ���N"t��Ve�3^F���C>'�r����vu"�*�wV�ܶ&"�6��*���Ư��!>�$tkS7UBˊ�o��Rc�����[GpK�mE���z}����|	��A>�S���5t��n�qPt� ���Z���B�����$��vA'���"��۝�rv���G���x�پutV�Z���Lxq ��ag�r��4ǉ����l��_ E�����)S�&��A�T7"�ǖ�:�:�eI��J���JeJ�&L�n>��a�5�9&_Vq��\q]v�aE��'�Z7��i�MŴHڥ*��L�/�>h����_%�3B���$'�H��Clvh�`'�N���K$�Tl�eЙjJ��q�OWg0R��h�1��Z��U��y����<m��O	QfiD!u4&{oe�yE�Rn(ſ}1T��@iw��R�
=�6�~{�TX�r��#�{��x�h��t��x��:��Pz��%߷� }J ��9#5���|�lh�B��vm٦C�X`A� h+�BL���.�O^zn#�u�&_�d�>��	�-�h����uj��D�����@���>���d5*��XD0[3#:i�*~'��U_x�����}؂T����_ײ��m8�:{ˑOg�����a�;�1��خ)�.y�^�n�@��9gZ��6ӯ�q���\%�0_��Ϲ�8�*�2UB\�Eܶ�'�R���L9)A��:X��H���Bk:a�Z����ڥe4 K���<NXex0��z扯�h}��b�|�E��oTuI��\�j�=_����[�1l��>�/V���ttg U{��~[��x�Q�fgۿb�6(S/�Ya���Dc��<��$��o�����w����	��֫��m<F�\�v%n�[����0ƒ�5[�����X������ˊ���8߶Dz����Їs�( u��{���#|����w&r,N� �QMT��)�y� �RX#H��� ���A�3l�*��2U�eG��S�� ���V;���A�)Ԩ.^CЂ]�AHR�9��_�q۴�V�_�v�?B3K)���|z���ژ���8�p�s��4�iy���KG������oٍ�@jJ���e�jуnd�c��y1�^���St�M�������="���/��W�NN�c^d�h��IK���h�	Y������`�Y��cbG�=(���o��t���AZk�x������&���D��_k"���'.7?)���9I�g��ʝ{ *��9�z6؏��<�\a[?~lxÞ�L�bfd���	��������B=�h{<7���uC�q�刑�0���T��@;���q�¤"���C��P�3�~S2����Xy�SZ�~n3΅q�B��.8&ғ���F�m��=?�@�4���y"l�
����f���JC����=7qE��"k'C�Z��)7ſ�7��4f�o��k?�#(C\����{�C~E0Ñ� %Ξ(��| F��壶���Y`(���S_l���-��ݪ��>�ߵ��΍��*�X8�����B慄mTkֶ�1ҵG����R�  ^�j�S���kIM�sT�9�˨�0q~��%2k�9֟��R&C�vp
�^�$�4QYM����~��>�z�[]�@�tC4���'��M��:.��~W����.Ս��3Q��U�e��n��*�	v���	�͜y���ƉRw���e���C)�@LV!�Ǳ�&�9�-�Yt���<�����C��H��VT�uh|�l��Q�����VȧGQDa6�ӸR�J�<%��/@	��Y}��1�1��E�w�i<�L5�[�eCkp�fs���2��D&��F��1��}�G��/	�y�1�V�yXpq*m|e��@+߼rJ�?�u�㋾�3�.�5����h�-�ޢ��@kϙ������վ�Eh՞�kaV���F,@b@��m�qw������-�`14N>8c�'(��=�� ș��ӿ�s��& ��wD�A12���R�(�Y:{xY+ӿDu��:R�GٗH#4=��MX7�rB�v����j�����i ��o����Oǹ�s���,m�]�0 ��})Z^H�pX��^��o�砧BK�6�ˆ�g��.4}���.a )�j�XF�0Ѝ��->@Q�
,,aO��bwi���\�	��g��,ώ�DiMVYUש
$��%6Uw��V����_�8��[�_b�1}�������v^s�@�&�s��NaX�	�0}ph5���kG@W]t����2��D@�ߝR��DU��jz���u���(�����L���Й�J�q��z�J�N�̤Ed�"��J�l�`&����OZ֛( X��;##���J	�V��qm��69�Ȁ�����zj�]b_����s���oa.Z_�勪����e�V���_#���"���ۼ���ys�L3����+��h��ɸ*�d�N6��hT�k66��=�J�c���� c�MFj՝'���Y��]ZB��ބ��zW
Y���"��R��x-=|�q��G�d-E;�s��t��\�����]e���D�q:W�����)]�7v��
�I��+fI[N�d�ڿla2"+z�܍l�M���i��� =���;�WW��s;OP"�۞�O��ɳh�Rl5ӌ����,Z��{Q &G�s	;1l��2����t�;i�����׶�\v6�.jM[�7+� +c�>\�����Ԩ��l�z��6��]�f��	��T�H��$8��2qX)�1�sPz�������Z���l\�����I<��|	�x��֢��Ie����-.T�,,�X��4 �ċJgC��2���4�ύ�H]�I��ܵ�̂o�ҁ�"8%�;1�=N��#�?[����n�`���v-�K�eZ�>�IR���!�Z{
�<c���vd��।'����#�ғ�@�a�#���0�*l7C]&�.3��:�}��##�J��2�����燝ڙ�썵�t���R��ǁ9"�)���Vb�"�j�;#V�dI�wv�\9ޞSrG�-�-�m��L4[8�_�.|:����:�"w7�p�-���Mr���]�R9h@�U�T?n�C����h��N�G��k�}�F�\VoI㏓���qi[U�����I�?x�s���fc,'i��v���Ȫj����r����<��)S��u�(sz 0lk�(�ɶ�j�h
!@�
ǽ_������(����uob���Q>�V�G�V�������Ƒ���������@a:4'�߇�1����@i��̑픺�~�C"Ìܲ��D��w����88C�*�����?�մ�Q��W��nq�pDϼ���z�4_��|:�+�[)[y��)��)���U]�2.�E��C�J�݅��<�F]V�\����7yO䓝`�
xhɸ�z�i0h��x�����U�e���t���7t��Z��&zq���XXiiSs�������J7cE��\~�� UsB\RC?���gt���[�����K��m�� Ξ��qA0Y�Gb�vF7l��3�K�8������YO{]��y�5�ot@�AA������K�0E��|G_ᑃ�2�Cǂ�����d��y	O��I"��;�MU{�"n8�w')uI��w�M
��[ikI�����HY2��Zq{���M�p�5�������P"��t�t;Z�k�~��=N1�[p���E�����Ja��X�2nW>f�2]5sbv�g,�jp���í�H�|�L2T^��E�|��9o��',���� �7�@��?ິ��ns��d��(��z�nc�����C��]�:a��������1�~��+[���I�#:贋��M߄�L�*��z���Ot��Q��<(�]g �EA� &�|�N�&��:���M�ⱏ"����-l�����]*J�˚�'Q�`s81;�_y���ğ�?x��H�}�y}�o������櫸b�q�YW���x �gv����	�zQ��i/�8����t��arCQ����K���S'�ҳJ��.R-f�fR,yAR���&GF�r�*��"Ȗ1�Cp]���n�H?�L�mS��t�$x���OM�򉼄���䌧��(��`��_-]�$��1�5����cxE,�}�?�Eh�H�C�~�fB��8QL��A��P��|��r)�S0A����0���Y���w�}F�5���+�G�X���"���d��K� F��Ysh<��?���jz3z��N�����A�էI���{лXM'��]�1���Zƙ5bM��^���S��%�6��@?8�� ~���(��?�r�0�Sf��{� '�`��O������\
"���D�J�ŵ�`�1r���5 7���~М�Ĥ��,j��.��C=�rd��aE���u%R�����u��Wc�_њ�ɐ�H,Ë��霙��r#��a!�0<i4NAu���ѥ^�;�'�ê���-����黲��aX�~;/�S2<�6� /���H%���!�+]HPŗ ��K�>G�=�wc��3/1���=�d����͐�-�z���6�n>�(�5��w� �'��7�+U7]B��@2s��³�@�^�8%�9�d��B��;�P'z�o����S������
��L��d-�B���~?`s)/6�J�_ͦ�Ӧ��Yԙ��h�3�FCR�!]��V*{�n�i0��Uˬ.��	�~�v�sm��^�顮�S+��s��|������<%�w#ܢ�S,�l�C��D�H�:4 �ޕ�s�25�G{K�fI�&s��q/��>Dc}���Hsu �%KS�^�+~y�o��zF�> Rҿ ��~��:w��/�Λ���b�g��~�J�z�T)�o����^o��6�͟!3�f��~E�U����΢:=�l����`���ηT|�숶��QȌ�7WEq�;��h� T6�7m\0� �ߢ��w�q�-�#���>���OY��J������sD���P�]�� ���X�#̩.Ë0���mk�\�k�O�_5�ln���:"b���b����l��~?ט<�:�3U�O�Jm��=^�i��I��4�l�a���Z���4cg"M'�������+�]965U��s���i��G�� ��Uny�������b�#��&o8+]݌lx7�l$s�Q�����N<��j�8Y��	��vyO���׆���V���p�ft%�.��x����|�I��"��a�X����cz��Kfj.�;A��B,SL��2_��tz�~�p����VG���"m�`LX�	mU��!�-������</���j��]%a�iu��k�e�?y�����V��P��ȶ&j*sb�0���#햛�}���8���9^.K"9�|Q?�u��eL��n׏�V�[Mh⹐`N���~=_����&<g�|���Xxn"�2�F��u'%������K��.Fsv��*�����P0&�D�+7Y2& �;��즫����r�z����Ig�������|@�.k��ĉ�HX�L������٣�М���C���X�7��V��׳oko����CQ[��x�O��/��7�[R_F�Q'tbX���J���������b��^�잍�.(��	����J�^�ENh̪�0���G��F�h3��Io��QA�bv��ï��\�U%��]�̏�lE'�ǵ��[�*�db�rz�Ԥ�I�^?�N�&����u���칉o�������Qwi�s9��F8�8��>�_�ZL�/�z���M��+�煑=6���%M��`5�
��>�dQ�rH�l�^�k7�N�j�ݼ_˓��j����Ι�R�J�!:Y�����ӂ��ޖ�-����b�+�3&��rkTf������A�S�R��w��r�6w��{�N�ߵ��A=s;�t>�'�A'"]���_�F�1�G����B<�.0�f���o�<�$�d�w4�\����G�~�4R�Nx8����0�GR]|�|g�����&��Kr��_%� _W
�}!�4ޑU5��|��|�����V��l$=�'3n.���԰����qI����[�� ���(V(�L+O�<F`��t8֤V�kYC���O+#��#�����~�N���沠c���:��H�}Ƥ�O�t�*��m�k����>�m>!KV���F���ʳ>�i���&2�����q|w)�#���j��TKNo,�����]��J�Le h��5���{��T��t��K ��_Ҟ��ѳ�@9�q>+�\<�}�� ���K�kFh_�%ik��͛)�xP���q`l����g�W�X��VeY|����cS',��@P�|O�����*����j�:�x力"c?툎�̦&�O�
�)9^��jJ�iqk>G�21S,�i*�Jl�:ீ�R�;H	�M4l�Ll}�sy�v3��J<v�X-�#п��o6����_�p�W��Y�;���dB�´^m!Qd$_0�.@7��ʹ	f�4§�}&�x���a�h�����ՏB$1�0SA�2�A�5���n�q�
?Q�}���(���>�2�\4ǝ�(;0lB����x��L���>�z��ί�߬�Gx&�K<E�|�[P���c=g�	�e�s���A���fw�rώiʍ;���(-ӗ9ÊͩI�����_I��f��Y���C9��|}u�-��y|a� ?al�Кl��@6�]�q,at^ѝ�t'b�d��I�u$<�_�ۢy��h�)�B-���ɒ���� �$��q���['L	
��M�q]3A=�\���4>��e�� �b�	�R�}����4�C��/��Y,F��K�f�v�WO+*���X��?����X
���#�����l�0#���Iz�n��b{�^X���R��B[ǽ7�J�'r�uf.j�C��O�N��8��yg��)�bV���t��%,���@�Y���!���˙�$�1���E}h�R�瓘w	��ķ�Gծ`?"�veK2����<�z��d['xz��uqG\RPw�?��;�ִ�(��fiÞO���`�w��D���D�]��-*��=e~��w�1	E��jg���E���&:����b��sәNg8����Y<� *�f��/d��]�Đ�,�����}�����ۭ:=�5�X����Xm#�㍽i����&�U����uUP����\8���t��`S\�c�x�H�'l�� ���05�?OfY���E*_e��%�W<t��r�� �0q<�Q��0A�ڱB(���R���?uOh �Y�q
��ّ�S�=��������}���-��
@n>����-.�wEq/�LO�A��<�$������sK@*�޶�s�8��u�͒�<��p��pأ������JGc@2��~� ���~���`ͩ@�\gv���"��*;\������Ӂ��K�a	��ehy��� /Y`��j��0�5�����mk<7����]��U�,�]ݟ�*�S֍]� �%��I]��,��/�^Z����D�x��i��Oi�g��Ο�z�6jKj ��FӘ���&��q���Fg��&�����qZ�oяzQ�����-Unv,�_�S~�� ,�+د����z/�|��;�5�B����#hm������-�=ȼ��$�>��jQO����ˎ9w��10ݟ��fj��W���>J�X��3!ٌ�_IN8,�R�gU�eE�'s\5@^��;��"�ӝ�5�꧚�&񚵪�����R�yw�U�i���=����Tq��"�z��P���^�E{�zT:� [Y0�����<�,#y��'U4B\�;�i�H�:�~�?s���A�p.Da�ֺ��K���B���/Q����V��HȊ]���)��B����_�.���HP�J�My������4&�?��8�{�W�f�ɘ/�cl;����ȉ�\��t�3��1�,/W`�Fї�h��`���u�${���q�PQ���a�(<i(`����pN��_�՘��n|˴���s�z���� �i�΅i��Ɣia�C�2�V�I�U蝳���S��J��Q0��f��h�o���k����ʯl~+JvdjU�(�c�Lu�Q^�����<�����	�xN��x�z]�q[�1�6�1���Δ�jµ����p��¯w��7
O	���r���c�5zm3��)D�P���K$�[h��sn���όg�-�����#����6�Z1dO���r	?_�[�������z�<�.�1�
u����;{�*�����=ҥ+�7e9\@]��}����@㋒��J�/dio����vE��u�/8 iǞi�y���T��5(�|/�27H����K���12�=}��~�̿w��9���+�M7s^.wej�i}����D�(���rK�p'?t�8Κ�n��r�j�Et�K��L�9L[#ڢ+2�Q2�'�-�6���%����qO�o&)5C\�K޾�Wur�d���8�e���;7|3uW��;/M�?�uS��G��8� �Ӧ�s�m�8#g���x���Y{�����-�j��Ƽ�$6)U��gr>�W񥋧i7Jp�e��F3Jξ�e�*�\�q�4F��k13h3�D��|�J�)Ü��������}p���ț^���\�������p*�\|� �I̍H'��x+}�H��~X�� �JtX���P���`�[O���K���A��NBqrc�lX��V�%�q��u.Y���	:�W���}u_��\��LASě�Kg��S���������>��Ĺ3��Ӑ�ߋ/�6s���F�.x��z2�Y%̲%y�X�+ɨ~���;v��*�%G�)R�P����k0dycs�zp�5"�Q��+�Q�?�R��$�fø>  J%K���5N^aƺ��E=V���$C�H�H�'�Fg��,���(ǵ�&h�FU�T�
���^�t>�������| '��y]'�t=�ФK��]�V�`����h�QOd��hD�)M�����c��<��B9I>6ѼI@��t���[�e�N�8�8��IX���1V��=�8�X�b
Tn 2�29��A�T����U	�_�W�@��-�Κ׵>;;c�����RjHT�qc����ue:�eW����,�� �e�{�0L6fȰbmFAV"�I��9/�@������t��ҝ9\D�Fs��C�7��N�������ܲO�Q-��,.vsp|�R)6���?#�4>���2�����9�.?�9�kI��ygY�X�������I0�^:?�,˞�{D�����c���d��_���$ANI�Z�|Ot�oR:S����3��d��4��9��YJ,����*ւ+��G*�7pȊW\������^�O�̓0?���DÒI;9�;�9j�M�������6�8�t@h���ښSI���l�����}q���xI����!����ORѭ2�T�/�և)����ke2%j�)����#96����XI��B��u⅚~?�F� ,]��ahm�7`�'r&:w�"v3J��<)za�E�ꑾ4��{dW�r�0���?�~�����J���} �9^Q�2�<I����1������D{z�w��a�O��
R _��'�[;���g���H5�]���B,7�Uǹ����iF��T��3�h������ ����9󲧹�c�n_�WH�~�S˷憾�'#�S[���5}�� r%%O�{x�t������c`�I��H*�A%ܨ�&X;����,G���BO^>;����^����K�2?���1�y�vݽ6����l��ߦ��h^]���v�4��$�O�3���s='F��,�6���R�w=�Ydo��U�Aݵxpb ��ȶ ?�F3\x�d?�B�5����yL�҄eҡqU/r#w�����D4�iq8D�ѷu��_�O�����	Ax��������
�y�W���T{;�hlT7���{����7K��l�BX/��Ld,Z]�t�롎�+�B�j5�m���sJ��Wr�A�>�t-��5�ui\tZL).��\ޡ5D���P�9�����/.dA�����f�>���vz!ܦ�Q�nD�n�Z�޶:�(���H]n��
Z?�RĴ2!�@�9<鿰�ow�xX1��~G�7�G�3��Q�={�Q���m�ۑ�]W�(��a��j���L�����О^��wB����"���� �u�P���ؚ,�^�a��0�*;iX7)�Y��{�YP-v��7��m��Y�K���"�������yo\u]P\���l&��.�������iQ�5D�[�*��*�(~�7��A���<�ԧ����K'Ĭ��Jm���	���r��K&p������� 8@�/<&(�*�@�2_Ҙ�0ۍK�N�2"B��yݻ�X��~�ٗ����ű���7gA{.�9VN",,��w����3O����rS�	��,���/x>	��#u'�|ry�[�X�+%G��E��0Bf�9J ��O"%9�)�x��0ԉ�VV���8D�[?)��f��ZjzI�N�t�~J���I��[��=��\��96���8��:J�ɠ�?�����
��!a��H�QZş�rB�]�J����\�T#�m�4%X�+�aT��ؐQ��]���vIg(@g����S�S����͜��7�}	|���xu�$�
,�b�q��,������:�����XD��h��5���W�J^]�ٰA�큔|����l�[��e�If�_���.�R�Ʉ�&�v�R蹏��d���f�D�V�!EdW��L˜�n�����Y����c)�8+# HHn�"�>t�k���R+��몼A�� o@Jͽ������yh���hw���6��n�@7�{��@������=_��/�KF�[t���|T'A��y#�baR�#����X�s0�C0يy�R��u���=�5 ���eJ��V]'^W(N�4��9�:�-�Fܐ�eT���¨PI>��]�8M�$�H���ӦOTΆ_�^�~@�����
��=[lxϕ=+T&��d�M���X!{��#.FXBȣ�.���������@7'��Z'�
A�y[�p?n4 �{���4�ׇ��v`�/W�kn���<�O�P��YP5[�T�c`k�ةJ��w��
r�$y��}�֓��nKy/��Q&�{P�p@m�l�p(�t�����3 UoY���ܑI=��/(�=��n��!I������x�1��
w��,�,(����rBy��kN��U�/i��՘"�`��AA��;?����܀�GBek��dE�@�h�?�,w���{j|ǔ��=dH�a��#Oq��ZXt��lr�hz�e(�}P�g�?��yV0ܫѿIv~
Lu�{N���,�?�vT������YNC���T�p�q�kA�6�ӥ�2oM�g�E�('�$���7��|�O����ώ���#P��=HT���#���e�A{3ZDe5�v��z�J��u�ں��E��Z���/�T}�8�+��A��$o��^��o0�N<"\�3��߾!�o�e��ŝ��O%>��Td�S����Pi�C�;,�Ҟ?����Wz��|�4Y؁&���k�9��_�V�]��?k^�g �y-JM=�6.�-e�P
b�نŃ�O"XĸL~��S0��-�9L�^�6�c� �hRX�B��^���owz�����z��� �H�h<sU���^���!�	�)�������
��C	���$UTQ,n��-�*>���{uL�*����j�OiV/����A�����F�3�	�v�9*ድ���g�TEr8�{F�[�3�*��c9��_G����G�i�,���H7+zKB>9π!���M\A�`E45ľ=���1Gu��]C�ج� <M\`�I�]����U������P�q�ɶ$���Gv���I3��9�w9�D�K_��n���ӝ�� �7�d�^���z�ď�H����Pf=i�~&\KB�!%;�@�\g�*����X�7��AEc���竰쫴"�Mg:%ˊ�ʏӐՒ��M�����|���V�>�������U�Rd	�m�\�EV�.ᴓ��*��Ry[�MjP)-fE�<ۻ�*����A�m�u7��+E��yQ���!�
=}�[�u욶:��l�w^��ۨGU����΢@K�O��~8k��`�Ο�u��=��
��}(��X�vY�����=�>'�Ͽ+fG���e����p<�ܠ�#L��m���5���)��qy�ٵ�'���0"L�����[=px9�Be�%h�H��%]��Ԝ��'��������8�Ɗ�'`Q�q�~�d�"�J�h������[\E����*(o��S˼Q��@N��p��3���"	|������em,�k��>�U!�/��owp#Վ�X��4���]��%l@���ϳH�\�+#���5�o�%I����:&a��?��/wqQ��l�8ⷢţ�d��^���'X�K��p�31��D熒Gq�"v�}xs��]��|��)*h`ʸ�REmʁ݊&!]���OS�Z&�"x���l��}�QOg5� ��C܁ĦT���88��ɴ����IY|��5���)+�QH^��_K?`2���$�r���PZ��F*�5���A��>Hk"y�Imh[�� דP ���c�9==}�F�w�U���Hp�h�Y��<8�$V3
��=t/�ѩ���=����I��/lM ��U
R)���rh�����KT-�aRt�3��?���Lɋ����aC�!�bY�R�W��bœ�9k��<�TܗׇU.G=�Eѭ��	*��_~�sX���m�"�
c�V� �ܸ��l(�eFg���A�������ԁ�I�9�vMu�w�7w���}H��T)T/�V�tz(���m7�����[��ۍ9��~�Q�-���w�!k$��B~�j�U�ٔ"#���2!8e{z������@��E�.�f��K�/�G-~50_|�: O��r�>���{rZc)����kK������A0��5��[:�K�&�f����y�l�S����\(��|�L�]�?=64Q+�a�u��.�?��ںߠ5���C�7;�\�̴Z�;Ǭ�)�Ɲ��j!��c�fg���[/�߈�xF$r�c�q��P��?~_�2�Uǉ�cbn�m32�&'�'[�[zCv�k*�

'"t����SM6O<�+ā�L%���m6$���t�j��˛��&�p�-����"(�kd�P L���T/"9�z�)�vc1~pB�!r^Ax@���0w��+�|ܹ�1ꓑy�E׊!���³7�5\���4*ގ����E��5��d�4WwF�P(� Q����N��r�J@q;��R��w4w����i�O�ڡ����h.O�yЯ�.��2>��E}Y����V��b�X�NQ��T��yCR�PiG{U���il��Ah�zu���-�:Fv'��_k�-E��w2��	ר��̲��n��"b�(�9U��3G��=W��ܜů��Ǭu�H2���_8��ʒ�TQz���p��q��X���p��'�ty�l،�oު��^6!`)������A�	�p���=��~lƪF�H�U��~~���H�x��M�C�?nI� ��3P��kσ�fb*C}(�pF�=��}�/�Q]�K_�z�8�QX��t%Ҙ!�����5��.#���-C�bPMbV>��>Tf���є�)�`���;<Y[����2�!�'��1!*:+8���6���T���M�ԍ��)<AעO�,��5��d�_[(��GY }���;�-�_�b��=�a��>([�pD�3�y��Ye$p]��Q5ݎ��}����%x*P6��)��[c�!���������[��%��A��
�d�<�v5-d��� P���GG)�f�)���` )w�#�;yV-�����r��;\ȔJ��aBh	�^A��7�*���$-�gׇF����<f;�ID���L��<؄ M>l<ϋ#�i޻�����
��U�h�W��R�+P�趟�i=ԓG쾭�+By`�%=�E�G7X?��|�����3ׄ��{;�=��B�1R��|,ҽK+G~�(%�)��9Ќ�_��K��pRqw8�l��%���UZ�.rшP�1���Xi�>�:��_�p����K�2΍%�>mZ�}W�6���ŒI�X
��[ihJ�l�"�V�F�V����0v7"�Y��5�J鬦1��#�-�qg��1 ����k�f�d�YJ
-��B���j`��M]05?��ky��Ľ�"��������E�Q�:��c	]	��x hP�t:��o�}X7�!��`���o�<�p꧎�o��LV�Q�j�����8����Z�i�&0�7��VA��G��(���m:q3^»a�
��CE���I$��o�=J�=0�`��<��yǚC��f�2E�!��Ȝ4��j/������>`�����dii�+�G+�T����͜��)y�h��
.�P��<���"�$�<�r��T�0Sc�������@��hɝ`BY��n"^����`��bh3[� �Mb�t