-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Jghjhx30sE9OdrH5jrcNBHxsYYvRcVcHLDDNKUXz7zwc3AWFmJ7Qwt1tanL3Fi91w345L8qwJor4
jKiV5ciXeSlUjYkAk/Dfxi5h+fmctex2dnTICXoKji6zpefHLvk4v2pqUhhDRXRUrrEqStBOYPtH
xUwFQNksOkmHfL+D/sYWJioXUtx99N+FUrON4z38zyWQI7W02FJPWS9OTtYeNDA8y9B2ix68C0KU
qjXLYLns97uFCBZcJu1ZThp8y5y9bmEJfMXyD3jsyXIfVGdQKTX01rvB3xwrbQCuXzgXB50IFdIQ
XuWcojJ8E1aWGboNv54IyqZk+/6vDgK/9Uw7iA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24112)
`protect data_block
an58lWuL2mnr5GL7AoWOlDSgAgoWlWUqRpnXc/Dln9FXstybfWhSWlQGagdhbv0Ml9Kn3nwK6ESU
raN1um9QCrAaXJzKphBlB3XQU494xd7QkBFzNawhhMOuZY0tOMEE6Q6bQ1wAp0UYEZwMJFvnSluN
eTvKpiNmTQ1tmp5LnKGC+4/daVN2aqddGufyplao3Eg1nlTihD3t6/bIn6lELfkCTzwJOCXpEv9N
WUY0Ddbm9t8BKOXsewDfC2qSbCexqq+qHyC04pHnw876LujPsFPtial5usOIm0cQdvDgShjYAoAr
wb6ofpyw31WM7aooaPcAKAgLiFrsatoIg0idUcc5xuCw1FXta9/ZLWB5Xu5MZ9ms6kvLF9VA3wnL
te9CYMHz5qUNJxb/Q7JJviuC91PYFtWvPGLrruXFJ2mjNJou32NBhMYlcn7c9nj6UCl+H2qQWEpY
r6PBWarVztD373atDQw91wm0GcJUr1BplHOrbwUYCBltkfsEEUGLsH/GHcoehhyh6vIwtBPXM/kS
sYsp617ydJUPFmqowPkYmpmf5EvnLo/RPD1BXLuQJfTyOYgp8/EChperw8WjMPxzuAbLhXq6ByYM
2JcJoayAz6br2BVqf+gHghlddvIonKy4VYLIez34wRh0Nb0fNIijwvvRgecOkGWTWA4JlCow5FvC
ALhnPQXoLAQ4gC0jwbHof8ST4VkSkp3ZJthZgc0ljQh2bQWtMCakJGbBFqCfiBL06sZhby6fHb1M
OZZLLKyTu0R9gqHmph2VeWMBGNH4RdJaagLm+yD4fX+zsy6HttJ9kJQN0eRsZGBhYdrC8gl1qLUr
EtyA/spiF5KMY9QUsbTyy07pQUfiMteHqJ31yBmFofV0PP9G0wiFjdtNEfBoktVfoI/2buqo+j9v
hbfEKhBDJaWxJsKKpvJw9XvsfZviyKrPzA3j+rYJowDzKxSJVJPZu1/x0eBHNjNOkc/aW+Mvl9/r
KZT2SF+eHQODAzc1Qbn3pSGLf7UtFRQXpyijY8tJzXpLPw3KYK7J+vAUYcEl2M3zRQCuVgNNzzzl
LzonppqKCHnyWz5VWMZgoEIIO2dFZ7PmkBfP4E+fLp9eolns7lLxLOQ30ZJW6wxI2LV5+hil42kX
PngRQU2k3zM2M6YX+6aT6cIdqJvbyqGh7NeeA7NWcaychvj7NSlnfyqN0TQqCGQxzuxMmqYmqVIx
NQF8oBCYLoDNbQDnAUzi4ueqYB5mx0EOlOG8OdN8Fias5dqjSDRubsfSc95IQGNLho88D2jbzFDc
6NYkqfTk+imW+ZRXSgkno9GYeaMUNNGLQGcKwkREqw3yzF1ntBopkGDyrkshJc/T7PRANEB/NYRJ
C12Foafxp1NyI+ca/44/qGxDdKy/gn1Hyta+GstTATwhKqr/wZwd1ChXggDpr6HEjVvUsrWsRMgT
aMtQ2R/xlD0djS3qGPzZsMVDP6468HgbKucegVCaLDshESXvUFsgVCeFfOkEq+/cDW6b7fwobX2B
eZu3vJiAVirncOrBqCbaIBT7SQPGWa5E7/9vFrzsA+WB1tj4VcSpyw0/3xDalqGOgew3BULluMYn
xb0At3FOTlAKaUQCEjsJBOlg6ErY9JEtxM8VAmWTuIcNZiLcxGObBO0JFz3VHWZnljGVFHWBmiLC
FfuuwGYVfRThApdvSSZtCypTe5t1aKYHBtCYn9q2KEyagdNAk0BuIqQmMxRlU5k21odYuCjFDK2L
7/ISb1NXjoMnB1BBmd8lzYHVtkb0UBHakO8KtRtlmp7PvKiwRXAMp6Pjcy56Xt3hf/Ch8IMe+5n/
jECf/Dz8NhoYYAsOFkYhn0Ex+LGLElQIfdLZbF8eqivj+qRTl/ANMMnxDoqRqAKV+9Up9YB8W84g
O4yBC2FIwBIBGcaduqPmDkBmPmE9x/ecvhDnq9wG/RbsHkQqlUDtG/Yr3RuFLn5c4vOfWvsh2TWB
trb573k8sZT3b71FUEZ5mpRgkK51xNR6dKHRfpt/aJx8HZtSf179zwhbfZkw/q4BvNmcwbBNv3fK
II4Xnt4CZpc5fB73f6u+GHGaI5GvGjixajFMZGva+iRn3IkaK2etiCrg1qCjlrc+d8zLGTqqog0W
DMf1FIVJWe7rin010H/lSWd4FdsPwi9IYs21TuJBu+h0e2CNgs4M1HASX8M27NMB2xfo7MpAtoPF
I6bgmUZdVQfWOKBSlQio66n17ahoJpBMgHVb9bjsTvhNYF0mqkpHieX+Hwc1x/yARwP3h4H+pjMc
YUlK75LK0d3BClVYWfNIATIqSeaclwhEf5+RJmg3/YF9E7ziG9VZvgBHtxhyiTRej+6DZsUF6JMH
K6hUCFh9vP9PV6RnsLvhKrO/Y2Lrmq2CPb0oA0sEsJUsPD1ZGXh6Gucg3Eqts0vqUq5Mj7mQadQ9
INAD3oCQWA67FRJA/4jYn0t+tFmOmdivFKw3bVsyHRClGxpFZy3lwFib12r/OhnT5J3YekCkcVku
mBaukwP1g8IKNlWcFSH0v39SKIqQDWnmBgxbjg9dpXgLg4SPHTV8HUZ9FWTyM0xVQ6c+lLuKiGTj
0a3MWo+ibYA0FZlD6Hcr6eWaUPA7DbKXkkmmKdy0fh/vUMRF3tj5EkxQqnhw0ax3+MvuJ7ZJl1c9
XXTbXycxL7/Ien0tcFMJHWANsqlYGJ4vzyozhdkB2LB42OVW2MAK2VwK2c1O2b+us8aik9SIzbDj
Xtp/zrfF5DF+OvRT6E7R0MjbhMDUu9il8xZSWDYrCtWh5KFS2YyUgKut8SOk87cvEjKm4uHrxpba
g2IT9ZAAxl0xIEUZo9T1w2aVuYcSeXrwR3kCGZgGxSXfhVu4YmvlqSR2Z+91bsq9COxrwOk57Jwt
SE8Irft45JK7SsniQB3MmZzcz85x1KVeL3DAyyQPSX5VVjl5VcV9bTHH2fcv/+smTTW31rvx7nAf
4Se9p3LR4UWl3g2AOrDIbLSa8DPQUmDJvtK1yB11NwyUQou8lYSk+CHTgX8PBrFwoFq72L5TyDIl
c1WOqGA5i9mM4xHLuCgXJWC4esPk8NEPmnkK2hQx53gQgj0cnwRdt7Eu0TiF8G3pyOh7HGJJRhAL
FKZy8bikNXRxvfDoRw65g8DjuKqTshePwWc7wUb0TbHauSqqiwIPy+bu/o5t/CzUSy1i6WvDvmXF
9nMqSU8WpSXy9s0uQ/q1lgNefcqR/GuMMmFD3YY2h5Kpu0fIa/uelNQYjQlD3liNxSCYiefq0Db+
cwiuSXCWgIcjAS/dzhHwfe2fc6WFEL6INuByEcput7qKV5hr8C06w6Hit2AUxUUBLonq4jyzr9VU
mI5hx7vciSh3FRpuYPDnmIpo+OoIQ+VGCNX/l1RY4pIe+CoGfuFWwkFSv56aHhxBMHCwi7HgEI1j
CjhbQj7XMco6Tj44mLZi6mPxgD6vjZ0npitrUMkbyxQnPQmSLte/P4AVuIio4e9IswaARX1yFMho
L5rodgiDLuAxyZ+syky3Q3alFvs9lf8/HvottLb5Hw+NQmKWa9Sozi4gEfk8Izq0VbiHBV2wnHxf
lNL6I/9PYxrgr2iWEGGOpGN43onQY01bvJFDw7dPNieCsn9sDx3C5QPFgp5CR1nTrhUXe/b1aSo/
WwkeFoi8oLnj5GAqMmzBjk8R9ignUyBQhYMkijq2zhkgrJBqb/ucs7OEzSJ/LuoXnz2o3JrJ22vp
IdRT/anbIa9wtHYrjy/jnc+OUDWxeDz94qUvE59iIfx1QEKKjvJK22jMC4dfYI4r7iA/zY5niRmR
59sPMcUVwFfi24mGx7Z58iU0xt4v6MHfCjzIrZuQaZkRFPzB0S94wSHd1CA7OjbomdJmVXXgeEqr
5fB95hd4K5cb2/yoD604D7NQoC1xmTQ8TpfyNRHllk3i6tboDAruR+DBlNtOOUFDDxY+QWdMTI/w
mIjagbdUJDDowABCHb85QQumk5HMU3BdMYDkESTVNoMHdcJIWzPRtWQxvdbGTUMaHdXCuvWsJxXs
aRKyT8dE3A4Q6mlbXUfqm075jPFermcr6rTVifspWIE3jAc0m7WqSh32+w1M3wreQA+J3Ls2rxAY
gEHZRJ04FbtYj5UshPVxO40voSOmTRpPeTYqzmca8Q4EQ+JeBrVZALx4X3GRsdsiRVsi/GNdeU+E
cJRlqgI/gM5jodNi7UH0PwzQ7jd66rq8hdk55qu2ZRLbm5f7AJW78xHVdFOOFq2uF/62ZaWmT02d
rQ8ZuQ8BA/yVpAzQ8mMVJjaEaK5KQNdEeHMZMwVv8rGo9nqi1WZDCjeQ+itldyBVtre34PVNZgIJ
0/NGwDMQ3AP8p62wiVcNyu9bHGsI93ZFeW8W2++IOWRRxWeqPkpYBuarena32khMlaFpZf0kOj//
krR6FHU8ojEBCYMxdTU6FEYas9UovmUomgQGve7b1PYAieZhCVmoONZ3tBgzRgv/FT8ZgzlWSeYt
DLXptUe4QhWpBWBR/O6INUIEJFH6nzQ4WctA4VX6MfbxfafGJ7Aw+1HcZXUXStK18mFDT9qnCr0R
lYBiExQ7nCjNb9Hv2HS80joNfMDMQSjajLMfH4qlGZ6irURgT3eDc8JHplwlafLKcnUVNTfeL3N+
zbFc9t4N5UgzxyHjeBjc4ygsdjr3pbtO8AuvzpnQa+bWay1Or4yv2UYmFDW40o+rM+o1WJe2vI1s
BeIsMmFnhu2UOXFaPPcsuBJL9/H1MJxgKBdasADapwgBJbeI5x5i82RD7Cf+86U+/wrY7I+qnPzl
fsOdH1GVRaPlevUjmuLxNoZNb/XRQLHDBHXZ7Om+CmhqbPWikAW2pnjN5VH8DAEnNzaoO/EPh0SI
LdEXxxGlp4sXBrx7a5ePUpZECgutTP9xS9a7afCPxRoAT4IfJcAy5/ZCYoDWSGrBHf3wEJGo/w12
IjiiUTufujIKmuJhMPnuudUYCIfNxmDkXWbJE+0l22U4QqI/MSEU3pSXNyA3gGTuZPxIqzVxLt0R
7bbgdLewM2+Ui06v3QMjotsrnyqQVnuhOeZWgYlXPd9Xnq9BPhWvO/WeYPBL+B1UV2LBfj4dHMit
aQaCrUkz20bDUocZ8kfQHJIs0O+b2yalUWBIezxv2KKFbBLxrg0bGHqyBKE0qirc/m1cYbN21Vjy
RmPodRQtLSlOhbTb0eDjrhmleA/0ybMQzpKH6fhaggAhYJoO4y7k5U0Y3TDtZOsjNPw6V3QvdVUp
P74veoJKGR02uOPXKwdhRmbdr/u7m/mzE+NiW6yxiQ5gGY5U92oDn9keicwIhz5xv8RD39WdTU9d
6T+8kbTF7OsghVxGZMoB1k+rSdrikaiTNbDrF61bnrWJw0TNzbAlPMzW+cZON6oPIlDng+CltM1i
OgM4yilUzei9wQZR0c2nVgXuH4f1gx04/b9lS/X6DXTcoo+JW1Jntl+2BM1ZC5QE0O5LiXIFgEPo
5f5UA3m/N2L74FTmHedo5IJo6f6WcTdDMvA73SRXsIiqqTNgyuAsHTaL2TEsnpwqVBIDGgh3cN2N
nACJEKjan5iPXSjSVRENdaTEKS/hlJdQnII+P83WIUSu4KPTvfrVidEwuoos+m6nVk4Hn8ocwB4p
gapuDEvODOfiIzBndHaPM5UQbLEywa1Suegyr6rqe14Zn+BaJ7/P8Lz8uMpAGVWWYVd5hqU4eb12
7R4WvZ2RiTm1OHE7K3LIfwf1fftJ34YJx3d5RneHczaYeVc98+IpuXKEDf5xf42EzkboiRK2cK50
TBYcmh8rFj2F8NfttecGaKjfcf4btrKhM9h4qmYL/hUHF8BxEV52bzIn0bagLanNFB3tGsRYxOKh
bJ2cNjRKmZ0QnFxFWW4kQ3irkkOK6TOTvZaJuH8FW7wbGLjkR84MYHooH5SCZ/0kp1J7nYxtNiK1
Gj0KCLGGiA+rJLfavm2cgSLrASQGT5TRUk/z3x0H6ruM++/I9eMZGqR6ETFQUpRd6B5ewQBQQVIf
vlMDJWoLY7KVyZkPa4KyjsSe+pFIYLqnkuhOiq5sxEuc/3FxK3cBXzvPPNyF+4cgN7Lx2dhBWLzS
h1nLbpi724hjtKMxw+NKufyoK6Iu23pk6pffeLpAQAHpkGNGe7QVR56t9R9yYDjOhNUfA83zY0b7
RQvwK2beYs+HQwFFUyxuJjZ7kN/uwVNvkOnFz0Yb9PlYSeoJGAWniTUjFG7Ge+xPYlb2Iujpk1e5
WsJFmsqL7haARUto03fGKL5Y2I5fZJ2Ysrdc8ww1ryh7ME9Ne9DWGW++iMzB3krvYqsymdmz3dcY
Xa2DUfunD7Y7tgB2og00rzoP9AWpR/N/tHr2fgBXKU9ajV3yjPxQR7qDfaD40hoOsC76b6m/YX7A
LqQIt11USSeMgGcqjD0LH9jCEy1xLvDZm88iccrlvrlLY4nkpfP/n0CIyH7s//3F6nXTXiRpmjfg
3mQ8ehgGLkGMNuVJZuwigOjbfRmWqqDnNYEEEZKYc91kHZnaAdeNFWf6HZ1DlOIvvKNklQF0qa9u
PabgJIaa9sJ8i16ILY+mSKD+v+xciTxR5NmsoghzwHxfU8gGuNDMIpvNs+ahpJfuTKh0JYs8nbNi
FvwZW8Nz9QQcDQAvV8tVbEQxTH6OlrzgpmeXZ7nZuy344AWM/d9chlqukE8ddEzCUvEzpkyuYz8T
zEdDOUYstY8/vpRwc6h1J5xSpLKUCNiS+Oo+m3+CgNqg2ryeLomkKFI0KnxIvjZAqPZgc0jZ2OWF
+qCR/N0mWM0iGOTRFrmlt6l6fmuFdsbHoHEHHG/Dohmg1WeL+iiRoyz6QbcpgdRm/g7os5Qgk0IY
k9R9kMBHQzaBIpEMmAX6XT9/DlcLyGnT4LBmZuxp1PnXV0527h4JpVu8cvCluz5pDpFR/mnx9mFQ
Zx4wU2cQCWFadPlfqGc3I8QRbScBO1eSYrBS07tRMYo+3XwgcAdOYTqlOMGPwFz9G6uG2SOT3w1G
8jXGyRO2ShbQuqncn/WagmZ10K7bUU3oo3ud4f1u6vvdHZVocdVlUxLeh8BHJEVVFuwGgw2/7Kdv
7gYaf4h4JTXYHbupccdWin+CmT8sAc1TflihEE0C5ATz7UIkrvAiMsrzojL2hhgIbTXzW5xdCOPc
qPQbs3N4+NvSk3F6LWvf2HsR/JeXJyUBBYSLMVIHqm41JPIDfXEUWqmk0b19fYqYrDtxXmTrQsjC
o0utkiPDngWhg6IzxycXu8VbtufofAulTWHf3+iN9imhkyMN0m2yC4zTtFZ7TPbn2fUbsnZuNmpx
/BumnAW2eB6kTPPkSBgcVHhebeiD9HrWT0fxy1JNGK3fClM5XgRad5eoAqH4IkmPmc4Alw1n4MN4
KqmITYbmVT64vabGOHxu7P/iwkW+AVdy+ePgntqGEMYTivE3ubHaFPM2FeuOiDCM1B+80zK6i5Xh
/zs+R49iItUYBsT/EXZJ/jCuL6z9R1LaUrUnDVcGv93fNDXEoSiZUXEyOTPIxNKIzqjJ7Y74/8NL
SxjGN7G/D4ghGnw2KNSMi/6RVtpj394a8A9edUGoVWAFPYLxMWV0R50Vh5VQuKENBK2/Qab/qT8g
K/Tk9T9y9+sg4ZCVUkk8LMS9ikMuoVBrjtnl6ugMuOA3a1LOtZcIuUT0vFHaH/8wyeAWruELp0px
xItOJoMVkudn2yah3BIoYgnRilYKmFdow+OfIecUAhmlEehAua/p3OhkzECzuwDwAJreRG/3cFnc
sxy5+RAYPIDsH5qOpqEeua9Ez/F1R8m2cUVlbXJ9HBD+SvsEIMJosIziGKKJHv5OJ+4s5Yvocq6H
/vTmQDG78ImaoPwKK1m8g+v5gt4qkuTtNqFs3jcndrr1RsenEb/H9Jh7gOdpdN7ZR3BWjJla338Q
pyChtkprf+aDqXjFC/Ob6qX7/Zm739YL0YOOmh9hJbQwhK4FB3fhBgnDeNL6zjFRnFgBAkk/6Wsu
evKphlufPJJQywv9lY9lYhvveMyLQzu0hS29WvsMeT6/3URfdmb+IwQ3UsKG9mGsm8CE7B+m/mYK
fLVXBrpfm8CKLhOkhoDVwfOFkqjwgRig2Aem0P+2HwUxAE7au9P7JCA1ldcWWTc/o99OZw/QPa/a
CcL/puLaPqR5MrcegAe7+TcFSIO94E0oxrDOF71YWLl2ZxSgv6bPUTX6kAm15JdnSp0c28a807RB
+ObAqabOhTLXqzYSDmipBPheiCYXNLSbsgObAnXnZmY/Kx/mG1+W/9s0GHySs3Kf+v0rUHdfEo6x
moRX3lyOwVPb+VEMBqKwaxyY5AsOC1MMy+rYnuaB9KLExfUoomM10TgUyijqCvA0HCfLud/6lwoV
VNmaUUoqLsJCjBr5aEJ7qPXxF9BpfyCEz9ECfbWJJ5CxABl16pUO5c72B/dTrTNsNt8aVlrBQDNU
pCucM9H/abMZFzdEyPOOwe8dZX3LVD/hZpAO2t3P4n7FfiTbm1PfZNjg52b6BNHeCzxnpMf2IsvM
iHwpxJgR0gc+CmyJk4yw0LEm/7aFTBKYA14ftqAqjum9dKK3TqvX4d5aYdNFMVac3pIS9qicfFs7
a4FDURgn8TIlwJcgoJIPhstyAonVrDFPkpu7D8uYbKfj73rule/DjN5qg5e8QwbmlgWTUsV97Mtn
BjSzwPzRZ5yHgK2ihGBB7sRFFdmK5HxbuniBHMugaAQVTr34O1S6VdDpDKGaBQBEutyUcSR1H31H
cdGuPBjku8sah5w0J903VsaENeG4QcLnWwet+20oSPRC6EIHGKL5PtXtSF/EKkqaURmw7jQK+3gZ
KO1vbeEwDzpVqahg9MovZ3Dmn0vrq0GR36uuXte+1d5Jd5xbufccrKC4kTrJ9ey198b5YuXP3DBy
VHImk4Jufs/hjZ9tvaiTtuouQGOMinHk7W69jFloh+q7yTUqM9Yuc4UmHb+laGoOn2+IkYHZqLt8
la5bJeKsr8QjUVdb/N6hAFiwOcmDkeXhsmkmJRFubzIyfc7FIRYENBsScrYY8Hp15zyfVc+eVO3K
4dPwo+p/GV4QL2KxzvpkEk+qxNjgtUU1/2QjxyPAwDRm9W/npqdsehFKvhH8odWgipnWJUnTCT+3
Am1I1wA6Ibdgf6I8Dco2C30hyPnOm2u5opa7ZTH7AeFC9I7vinIEle3mCgizFTx5m352St7ULoXJ
RSj7pnAXu9h+AqxTFzpnmJMoHkRMJKAD29pP0lGoG/HeAmCSvjUJ6R68q5kmGSUkkZLey87xcsei
OQumT+LleqrbveUBqfBQdOFUalcOM3N/7PebzzFUCd33zwaVy+TlunPvWda35vsZFzDQ6Cjo5hYO
D3uYdNwJae2b3hB3Y05Du7AS1cSqBDTAUFag9JsxmF3I8tTcVM9ClSaGujgOPtdJQvrqz+kjgo73
+rkrcG18VvhnCqwGw3bZsjQEO4ypv4qONeaR/WjKx/UkNgMVEKmNZm2oI9OOLM0m0sMA4cBIWIQ6
VqLruyq7QunE/Chgi5fq7aqekfvXbD/lllSkaO/VUcFa+skK1njLVaQV2Ip4W6fBGiG0XyO39NJ7
9bIjGh6f/2isYELgxxnV33R0rg8c+3DbNvEZ8EP+LxheaXov2F5KOEkgsThIvwuer+m32yIwleK6
LzFGXVaFtnM0cY5xaD58NiD86PImHQty8WLv/gyGWu71EC3nvTduOx7I3eJ0ZZlRUfSPVZlKKaIi
xsKAwvOtYJo0RDqIUqJrmLNS3o2i5YMNxVBJMDSXwjYrEzgfzJtkEFIyCrooF91KklN+0/UHI4j8
KeXYUQZDfTQm4bX9d2wKgg9y1uF6ENSWYN+7blLR1tkE2viZv46iw5xS6GMJIYPWiOiPbwI7rdy6
ZxAZC9O8Dp+B6H6zfGzvwk1UhSBgu2uAF4D6mjGBgfxP1fIz0jyC0YdtAYCsPIBfBzwwR52i0A+U
8c2KJzwBFMMhTknMFH9ai9+osMcduKkaBw5EsU8rWS9LLN08JB9/0xo5JAuyD7UNOITlq4KYiEIG
KHcHoX+4/98eyxT2Uvzc33366qLutstK2NRYqdQwnZ6DNqM+kedhpbir+rcWzsE03xnFi3BKP3Rv
owF4JHos2GqXX/8j6Rd3wOScaPj9i/SOLwPE6fee4lIBKyG9eLUmdZ7jj1Hu8qBGX9bMWWRgFHWn
E9UiDZ7vmWj/keeGBZP348LBNQwDk9bsAxoDhXSZ13qA5BlAyEtLxZNLeo4a9swMHsGMBPNkEJUI
Xd7GwiMQzFiHbLG6rj9ZuoHqraKEem1Nq+6uQRZxcjO+UO9fzUavFL3zJf1KZontrhfBcQdTg6J5
5HljP2OLwcxWc2srm2/HcsStl3YSMYxI0jMvj8Z//cABiQwzhqlj7O11YrQ5L2UdVZYBIFVlLG/w
P9+61l1veR4hxbBpTPU1FG3Fi1l9qHJ0yfA0lK9CGALFdWXj54rTqqpoC9XRDxKlyg/4C/ErNRVW
lp9laLTxmp1hPiSu/WfAZm6763OSFh8ghikOFWnhYXZDLJUTgamkJPFtegtw4IMeVXpfSAK0b47s
y8i5soETei7JNUZ+m8G2XuA8nsDow6qNuIYM5JrwgjxeERPm/y9Jf0k+uEutDL8dgWa9pKSjkmXD
u69GEbMFqXD7FRPeqAENYEiKfoyo2/lr9zKqmeMzU1KpVCNvcbgcNkMS/LPQLGhdO7DDt8NTrON0
4DCKjvpUcTtINHK+IyvKD5THzfZBLOxb+F+2q70V0hm4y8btAU46YuLhGJoBqxBFjF/l8C6J3/Zk
VQhr6dXnWh1m6tHd6Qe9aaFI3wnkfyu89UVXAUsuYwCrPol1vfi6rFKXPgC5dBseYqJfh6BAyR0l
E0e3N9PjMkBHh/CSxTAyqT9by/p4APgkOREtDGm1vZQcGJqJ56RkaXyqgC5gH7kod9Qr/HrJiz1X
wJ8OTi3tE306BQeIrFAbsWEtVc9FW7C8H7zdsJyc7SMGQA13Wv0ZOuw1u6ur/2CS75tVv+kxGoEb
pWCGhRdFCwaHjv/bCtARXbxdUToKjTWvvXWmjguub55QY/VQ26wvzSZypXHgLlReoXw0lM/DVJsz
Dj4vWAVaO+YhQrMPaAuM4pTym22tQZwRvVkkFZzCpFenUERbeSXJBCHz0eCO3IFb1KSSCN0yQbll
sujvF7CXGGVCUZhbHn9WRKlGtBSDO4C/uJgL0tzi+GkRTGORNC4mFqx03V2wJKOXc+51hiwCI0C+
oziVJLZyuG1Fw4NhrJB5qDBD3VEPYWQvZkRU+8ks8dlznnx9lsWW1TrUKfmM+BL2aHjHWNVyrgKj
666BKGcLALftmWiUbu4kdsv0WcvQTlRM9f74lhYkz3Kg2JkoRHTIwhhNnt0wZEOAJe2DRDVZG+d4
Fk4G4N9JEdOiB8jNyH/C0w70U18yYBMb6IIUdkgqSl1wooyK00CF1ElTA9WAFVqc9t3PZqdtN4+f
wpvppqirDBrceUPJJfkAskZSttIG9/Knw+ESODyWpH84QEkTu/H1ZGgPwDJ1NGDNwAY+z0E+2WtN
S+wAIMIezFNoMwFiBGTRyHqseLEVC6jVAkThs+eXMU/swVTvduJLxZtm5C2ZxN2ORt8dUfzxWccZ
rI0h796IB+Gj4LOpMduWNFqphjCHD5BnxudkhC3PEJJY93P2t+fdovYSUnhWLdZ+wqSKgrxxP0IS
rsnT73O8nk/oGC4dJYdmusKiQOhepEi4qlS9BqiQoK1K8+yxrydWj6PiMfRDvEM52OhHIALWOY+Z
kPd4lf6kS1LYjLXwV17scfQrNR0BmPKCsSgelyY4/60MUkkVGLsKPYhqdw67zqXFgmcJMkRcrBWv
vvQLGP60H2zVBtf6wt7UgZzJ4xiOfYwv3rIiNLz3swCdVylATFIVjFYRE+v1rIRKOkQIHJI+6ZHD
tMlXW3zBdReslgX9CxYFORJbbi3p2Z8kk/vgVWfsOCs18RTo0W4vNXXWCEcM2E3mxHA92PyfJ1kh
xrSRVt+ksY2JOdh3v3685+aGP7wIr4vXEAXX3GFWAGDXXQmhmsAn0ffuYDJ2gi6ZFyTXd92ttLvB
5aPlMZV1BFm6Po6WZdwkq2L9BEaF9hACpTewsTNeOVGQHH5hKoVrNUY31aQzyEr6CkhFuFE4AtNi
ETEiEFIDebZN9FR0jQNjQb2uzQ2HQqpgBK4k3/4FAXGNd0l43UYpuHhS8sMIx/uxNFxmluW5I8qb
uabQxzu20ZQzMOTUvJGrMuqgXmPkjyIe+gmrlv4AKobH81BKPwHDM0ZlubhaZPhNMiILHJUt1HjX
bsagQnbCiwanb9RVZGQ7N9PiPIuKs8LQfZ7rEJ00ILUGvVJkV1DTHGq6T5MZMIKnBhMwG1QEQGo+
sI5WXcM3fxqvtwC+aIngvudALwSJw5w+94nhD/RcLVNFSQ9TyAR5OqOZ6uNOUj2PDsYPrgN5wn9O
t1ke2N5StUPeCxOx3Kr+QrKmvPYW3P3J7zL/XsY8L2uFgz13AtFaxgjVMJVcqbzIewtl1jdabsS0
cC6bg9BOTMn26vx5rdKzlynex5NksgPu1FOzBgshNQRTtSR0DuJOh4qsu9yJdSjzaLXir2k/xUVG
DZuPOCllDkkWQc1RCACE7xhO7g+K6gisT6M7WJ6Og/Dxgb4CeGO4PkQ0ODT4OHMeKZbND99WMRjV
Xe5xdA7l4C/ixfvV54VX355MGfDQ4dwqYSxLGWbiF8vOiFK7Bdj7WmZ5uc7pIIOkfZq2hc66C5NI
Ks8vhf62tqxhF4VVNtCoeWokUehggOWDmx2k3VoGH1/U2fAYhghHXPbMSHZcP88vswHxjPxgxhoc
Gw5W6exqbD+A1zWQvOAFRoaLJvaJO9xwkvfi7busWXF6aeIBg8xeHkwYpyR2lregbk0rZTQAQSN5
2Hw8NKt72E7C2TrcRS90fK/quTcaiGUJVEj2A9FrJtR0C1haSWKv6SzKzJMHyvO5jHfJGHoEUC6P
Seri91M1utlEQsTH4bkTa9F8eRmJBTH+rDaXjj+aUdp05iR7cFIX9Z3eL7RnLth7KWJJbIr2RD3Q
ywFX79aeim9itom803JMNVtSHjQDJn7NSFEC1JqHWdM4HfN/HB3vtXXMlItkxmhndKqS9pkt587t
8OQW1IhlDJSq1Bp82Vtezd43Mp6UsVvWm8O/sUkTGw/TbiPwUtiaQ8lShMyxk/rEC5fL+0bzDBnX
bdIEYp7/cyTRR3sXNzBCoieg2B0oII2FOazJtIkEFXb8pwa+DHj5a0tcVOJGOY9XOsTZu5YHp5zC
dpJMCIaMlTi+FC2fEInvmgl/XCu8KKF0fjyxdKgsKuEIUcJFYXTtsIT18Ar1eHicHFXlIXwwNLrG
JPCnyzlOQaidJDdumBfxF10GKpNBcrCTqF/uTOudmii8JHJSN2bF/XpGNrTBG5UNNyoPmqlfT5Mz
av9g0ITmvUA0RDTLIdmo1+uSbPQU8kbKSVm++Rc8/d6X/diAZu8WhGGaTZg7mPn+lJYNxpfH7gdn
q55iu6bTTKJpRVEA1WUEFZFIStV164DZ3CyWd+buzzNKkaMDxvcSND0qNtcjm24wnkaTVfTRQxm2
GMyzzA8/fwNZPZatDpcFwk7vMqK5aOjs79ZeXbsKKaRjRre9rp7BU+vOZrR6xrPycrJWGljJkN6D
72xwYlNIUuY8KyM3RsGLn08ej2pK6wiTTOrJLWoAoxis3oywNuFBFsiHFocRLKkj3CJqmCkjQc6z
THcdbsyFXIPH2byDDl0FR+IMrRk4UzFjI4d03zjIvwO9WmDcOgaUvFDiH2GxcFCV13Gp6RzIp67o
hUfjiDKMM5baDuxwLwost1BrDRTG9eIqAVONxZTitBwrNWiTCg23LH+fJSt1aaK6FNh7xFqnd9+7
/fvoqdJuC95rHNmKq+OSi8ihP95M+Zno6IwKv/bb7mZO0T0RhsodveSuU9pJVpTkxrR0p2jvLAUQ
9Bw2V/DrDXAF855OYt2/DnX36VWlZcEidNlOaUIjrlIAIfwURxkwHpoF5DvtxDdfqi4YgX8rCjDh
mWWNZP+yWWHPxOgDg34HWDJm4evfEVWpl+ecVJdP3vX8mZxDSnB3eFKt5SbZ1QJq9n7ZGP86FkYx
y6iagboHcacwS5jaLIclzULmzFTH+pEOcJQ2dbZLNO0gejnQNYq4byE72a0FWIK+Bxw7TXORGEhv
TosfyLyxmgm2c5m7KyhT+GUqCHDCyu9CFcY+6xPXhIxziqpfBtoVfwBAC6ZhZN5ovWeqU6KZB3VF
mDo7IyJw9Mc/pj1UMnjEvpnayG2ZIlquAuqbmxJgnYiANCxiIGO2Vs+Pysxe+5F8jZkod8LnwY4o
qxtevsa2Q8TaXJfYkMCdAjP+TZSc9qzXXwIM8zkemRlz43dmf4eliiEaZ474f3j7w+qC7yWotmb5
ZdE3hnWj+eQovpJM3sLYjmV5LU87eDIvPqD2CTW100QmUZQJEGHPNaw6lWEcKIQ8o+Vp7O4WikB3
EvZNcdH2qbEyJz6PJX5xcx6qmnREZcbf73UpKHSwoVs+432Y2iFqYBHRGNRwUUgM3edWgPdc2U5Q
9ts7mKG+lql6u8F7y4G9AFI4eL/exgc58T13zHWN163z5NcFRL1kQVBDJaR6WGDr7rKr1kFfjEg6
wfewJFRHKEnsIF0hSZ7TZ1ab4oHpp/NjpIBnNi6LRE5cAWfqFJGKgNbOdJCfuuZOGx9Qnnb3m5Fr
/qCaR38vithddzUO9I32z7OGKTKI4iE0lhWIYSmmzVoAVThlkvrYT4h7Sj30u9v/WHpz4BozVadh
D7fsMjIP/JraceRGwcMrBPPIBXI/ZK6nm3Pb8+H2ohiWGN5BGIPxFFwbzNTTnYfbuUMqVPVgdWWw
HWyqCBPu6KExc/iI2veLTVRakSeT+KDzL1x4FLaZIJhRLCOMFkJwfkFyeCt9HxAcfWULVb7WC8QL
dLn7GOsFkRvEiHOESb43YC9JScOP6Q3sBNDpgTFAebuZdKpz/tJJiVTsDGmtTEHKSfyz8rec7a8j
qEFiBD9VU/ODqePwh9kfk9s5fj8zJHYqctEwXaUX+xz1hSDf3Ph95zQ+nGOK9xrO7g+UlGDLI6YP
fMNsS55zNBHqQ9/2WreudYRh0zfuuveIWtplGrvEZle4MO4KaAikntQMy5OzcUqnoqwBgLuWi/pH
Xkv9MOtH7PGxk+8K2NsgxHlYyI5Hbp75cO/+mPvUPwD2U+1qdOhp1VKKmf6WJyvJCk/b7aiNBxl4
JqxkEFLWfbaEn4FswBl2JC2047fpB2WgVh30lHw7B/VzaiHDwbhLYScWk8QrY/XP9oRF4O/p1KaA
703yJ3u3PHGMNnDf5pYHaQ1WbgNs9C990hVPQr5Def+oECjlVi8yy/9gCWyQIeYdIk/EPB4mdrgp
4nd9kSroje2LBprcseWTlqk/ZdOM08ynNSxuiSJMEjiDwOJJCtwyIqbIMQ3n6O3or5P3c+4rpW9V
XgWy1wjYlyFQh45iAFW786JEOapHtXTWkC1pzdkQ8pQ28I74KcCo98iOpULac6CRtLOFdab+eJg+
30Ztxi8evzmVfu1DP4NTG/vvC/wURrtNLWyO3df4s/VxRfwlXg6MnT726tVT1m8zkVTcEnAia0j8
H4yVvFG43qB2A3Qayz8aVxnm60uDXoSPTRByqOGrsY00elNrNuIAcA2G784ES0iWLYwQb5GeX7tL
pOW9UVchlOKMIdiRFypr0iglkgIOys7ycAh7yRgNStXSMfNhW2cGdL1Z7C12MhehubpsX9FDBlNp
dsNJlFgLcaTzJpgRiwuExwNrdvkdtMuGSjhN/Z9BksZ3g9liadvX9sBGv8d6RbhDD218TeP7Dntq
WodfibGWEb/5xR7jWih/sBn8OtgkFOhE+VkX/3LSU/+9anxU75SXk+T8lzjl15pcbHH8qygW6vT8
wGun+becOq/+kuTFTigS2IA8nslW+8AqlzIrNzrfZPFQARjL4mjV8Dy2uQlYim5e6zzRKnIFk3WS
1o6VXoLhX7Des6xJ8EnOLFYXCktUEMebvoGq7LZIUCnzUGlI3+HEPITqF7U8lS0UvJnrEOWSN55A
RKD+0vuKUPHQzqQL5gmGAaHKE5YSTwzyrpcjUJyquRuHgGMF1ZQhJ7gauhM7JsC0kLzDnX3iCGt9
bTVNN3vxBF/g2mETF7h//qLR9m65hXNju3JhzrPbFcMxVefK30TBs2P73jF1Bbm9lkqg4JJdi8wv
yEUuaIAoetykunpDakGR8bLABGRKjBtXPZBxhY/cJ4gKE076t7uyldZTjqBa2sPtrDdvTsA+6KhW
vE9idHqssSh+BxctQzV31LJ32e4amzfGZL/Xmxt4sEM821uPAio5KI9SMk1iCEbRHmH6fSo0tJmb
/B6Hj1TN4DLlST/QvmKx3nn74gkdr0bWEfeO4oywkZ8Fjxyl8jiIDgqxS+wWpk61ap7e0nc9cnWi
dFpMqeFVopSqs9QXkec+J4nHA+mTLK0TI9pAlco8nAo1YKMF2lX8eg5wve4nKuFmJ1RWATOXoWrU
mTk4p2eKiHu1IG3giP1o+LWf32dIhhQ2WFwB0tj/SkpNiCIOAuGleCodsz91C4MZB7psoYPAHDow
/hJ5oA7CFfVuZ4ZtfRB2yX0txwtmox7HlOQErGyGPJPUikoczdB/PnxZa/u8ElwMv1DF1g5F8ESZ
7g8DSzjOtL6dfgSCLxikITWALMY/pgji1FOwabknoJ0CZcIWi/NE3K80ukryTPASGwSPJ6sowJDr
QVNrfBhpFlw4T70Q6OmzF3KGDA23oE0oxwekaNzZSDZIg3db4iMNJwgSCtmQ10nQGVA8yM54XCdM
jWjvyzFepj2eMZsGQVeUeWqAFWNj7IFYM9IKPXpr9yaSsbKRjag16eczGOReeRQDhc6jOfm9/AnD
dL/uidPErMZ64uAXbxtz3y/ZQDD2IIvqdcRRszlnGjEqix9Aba26slxMH9gqbwKT1Zdi7Nf2+mR6
mLg/aX/5KLSH6LRfHxzNn3Kqs4vkHC8rMcTGnMb2fK1Z/JifkRb3RGscSkri028+3EdzaQc7yaup
79Xvem6uGVNP35UjuhB8gZxu+IlV5Pq4CVTx+4rIEswrLdOQ3vCxxVByQKNMUwH8KSeL65hIaNeh
gOreDCwE2nzBeHu8Gk0OZkpdeuBcTf1wWzxvKTZDNW0gYRL5S8jXUfdZ/wp4FAYdz5dXK+IdOttS
90NYUWoteI0OobMbrdVQZ7BteakHee5NcnC6PCOBpBbdvNjZ1wMYvQSHkQbslzl/mjqULzZNe9lM
TkNZW0D6HPcyLLeQXW9jwDodlDjcVtQta/DXxHnFEAP66j8d5Na+1CBuxsbIvWHmFz/TVPB8twAl
bt+p4BEzlSnZGkrUqlmQ1mkucDoAx/lJasNucv0XIPzJDqLMdI/ujT8miBxaUMwAngajk4yfMqNV
XSzIURcQvYCkMPx2XDOiuknN7EoTvXwMw/HF8Xaf0Vhupv1F86dW7RFG9VkM/o5suVajgNlDpNrp
vDiPmBwnnew6NNh0e9+qQEOXZDtVrBiz2n+vgQAByoB25K5pR8jVaSR3jAlqAaxMul/K8ZuDeM54
E6xTkuNFACTh0oeZ08Ba2JKxw7AJuVJibzdmPAh164tS/jUgKTbWNfApdUyl7BYpBfkSKq42tLG6
Su+RILSrw3OCZKGYBfP4g3bcK001L8tOW+uUs1sq05bw5/s/ZFdPevm6bk6sQkTafRaEgFG74yxr
ZIlnAYc9pVRwOvk3UChV5IL1nynCBb0NkaRVUdF7ZnCH1YG8uZwIJLTjdYoi1/Gp8IxmNfbZscfA
UEqtoG1tSs8xMD34/I2uu3zFPGJpKSTphmX0nHIbK56RrMwhEjMRiZ5/YFd4z91fZui7v2LXMy/x
otyySNBKKx99PvhvDmvQhhaubmeOYttiM/kePfAKfdcHzUUOuu9HxHtmANkUl/EOtKMtE2CBcMGU
btxOSaeqW3CQ/Inz7+bPTa7zbhq5ojEDm74w0Wnwm5fGL6gAKLS7znp+Ix2AUWSuRJezULYjoHB/
EZSDD3BW5TQ6K4oBOir7sSjAfOnr4b70mMBOrPe08IT8LiYRkXvsygfdDkyW4kDd10WHNU8lCM+h
iZi7fD2fJlV8JMHdMUQfwEXl6QvRVU7Z4Z21I2wvGfH+Q3RUAGz2wySF0FO7NC9wglJEBC4GXKai
g5JW5kgL9id858YhnISnqBYY9bntmoHeWeF8Gt5wySnC9OAywGei3S+tezZbnav9evyBo0/efDon
pbZD9M79vG6QKLP2xkr7nLhNpnYqOPAmJlRGcw55tacgv8gjHNRBxT7TWBjzt/xq2WHH7d+1/R2D
uD9nc5lS3Ql598OJLOo4xEmKM4fJ/YCE0tc2cAtza2mIIJTdNoCxtuxA6jgZ6PsCApi6o0zWHR7r
OUJn6n6BdWyHivIY/1CIlq1rC6TOxfmua6oG+PkJRIXsGpu5rUWC2lu6JNDEIBZjr8vzUzxzI5h8
/4Lm+BOBlM839Vtk5x3pZb2tIJBqjRs4d1MpCI61NXF7kjlml6low52vU7/LBw7Sh2M42Me+rbl8
yclgIH05kxp+DsRKjKa8waWIcFTvIE2Hlkcs9AgqKoULWcRURz2DD291xp2Fz2+C8m3aniYp7gLu
AR/n7OtJFovSqY0Sis7tznLADoo24TEtmrvtx6BmBONeEGvSdQeKaB0nNaZxQEFUKS6GZn67w3SR
fVBB8T58X6qtCTjy9pCzpcXZEte4zNF+/OMLOMDixKIr+CoowKKNd39jldF1a7jw7/NZvWq6+981
9ELKWkhC/UNtAGvEWxekHw6tmexNyrmo+J5hKbluxsoXjfz31HaTY5Tuavk33axmFq+A/oIC/Kcc
hBYqTgYoCykvHkuXcQ//OpGwmI9MF8eox0RAVg7HzFAHTiWwjdyEXiZa18g9MwkkmUjHm+wJOSqE
URjEffXmApp8uBwimFAZfpPYX9shvoQP9roEjZev0EXMrf1VG+Gk1pUYqWjjJiwt1Dk0ilFauKHH
qBNCXUjJQVkDrZuVIcRix6UMjmLCayDr9rq3nB+jvWfJjNTcq57RxOB1nEv24bwQhNilsdtDOnFp
gDEzH22XsYL6S/Bh9mu3FImUuAGOf4CP7h8wmChRlRM7jQ4+gbaLnrU8QLaUZz2yflSkFRdAfBC1
Ywng8xqaeOciNFQHZew5o3vI4uV2PftEH41o3qBpqihKdWG0qJVzh701EikH7rT7P+2HudzP+PYS
PhnurG27M1fEq2ZYLo6KbdzyXQjXCcO5ob5MpTXcak6IjrnxCTHcO4MGeQGBNWZ6hV/txmvI6B6m
ThNOp9gOj5h03PDnBzhgiyaV2NOj3Jn3spx/7oPwKx7w1PGqvyh2NHOKZawZzeTKRJioyzZ7eCtJ
VnCG8xCFc/lDvLVbB3b0GyH5Le62Y69mPziUGohdbSq6F46J5wUQjs/pM8QDDuKdUE9fYSZNTjne
0oa2eHunnXHsBPRR1YvCAm7gQQc+o15d/Ok3GFpqdvfycTDZ8U6m17EPmyvgcMMq25ljdoH0XSlq
cU1pfryGYe+4OXQwDsLKl4zPu8XgZKtlzpl8lJxbjpJE1/K6IKkRuJKcPhioKgSp5fYkr2QjpKEs
DysKGR6TsBhkJDBvBJPz3HS5pOZcCNmW+bV0Uddtcu/HyfK43l9WZMQm+Go6F5HzB5bfefLWLTih
Cmm64CaZFWnQrPzm/5sCOz6vxYF8NpLc13XzNk5nEhkzV6MdHGeuLk/VXOvYRK9Ks5LedMNbYOsn
fAaJJ+FEzfU5K0tBZSuNOx8VZxXCLZPOuQtKYShpfzDmxqermW0ZYBjtb0oHAX7jq67CWS6irmec
4EA1tY9SI+JW3V5zjKRjZvh2N/aLWVcupqRz28l3q5alb7faFhnzo8W9/wBIFtsj3K3yhQ8qBcMC
Sb4vOZcqTpOCLpBOj0XJUX/kdl5cB+qc9kslUpsNoBeXt3wkkgA75ID8hIwfvhRYuVvvE47oTAu2
Ila3jHAf+5+3eW37ntlwXecEeTph2ImpneXT0iuyYpDbaPUAu7WACQwCjUEYYU2v3ll5rBXGwVfx
OIsteSEpZclGoXzCCgKl34hxm2P41Plk/kKRKxXZOfY9mydwqWTX1h+BIo7aBLaM55hvYGQSjuVl
acwCLGkz9oZSlI3HV2t6c9hRhyncCPkHFHItzzrngvpswgrPadvVU/VDOM9MATo0x91ks4IicIKC
dN/RoI39Dy7oiusCbo9A9rNzNdW81RRphaILdVbfCo9Yx9rqXBU6G+KeOSRkaBpspoqJDXGhv5A0
lQoMJR520zu85ja0QT06xB6v24e7CVj8dpb6DLlTSgg7RcmHaIQ7X/wIAmaYVCS+EJncEWXviQxr
S51B/clrA5xsL9VuDgpqpbCtXu8UUk9/rE/GFx32pV8UyorE5enK/8zQcDQSQ8g7e1zmPo81+ibu
aPLInIX3tHi4v/+UWOT4v57SqH180mJK/ZSJ29NRWodTICXLPG6tAUFS6YHFbkwezRQNwgz4zX1F
BnCH3LLSWO9dJFxdsC7KXmlCiGDJdvBE7CHYBjfqcYzArThGHK2d14hKtSdZqUqYkC4NAFPRf6Ei
/R21eWMN8A7Jjm5gTozeOh3CiFLmdsHvhfLWlzV25GxlkSx88h+HK9tjTK3914KWmKl8WkF/ODRs
y0P5TGilLdTgvw3Lua1s+FfW1HwBIlrsXlCvyzoSy7chfFeQesWqnYtI7jooHqAg8fmjOXVC3a2y
VcIgzIYq+QLAka8wk+BpHRKMrrmiwdl9PsI+QwrDfCYNbWifsdhM+LbNGfP+FUlISXvEhHb+/fP7
HYKZ6b99FGJk8yCXhLu+myMhF4iURppAVUfyEtRDI/zU5g7f1MIXv4VXfz2AMyT2+45xR1L/cDc7
b/gDxR0U3KKLGdYv9l4ueM64kZSvJdqLp4JVdEuI/yRYPi54y7k78fxtCdMG2oBDuWMjICEZSQX9
0lcRLceiceNw+TKC4QVRbtH2+PDUkumjFD3FDDnyVywF+KZC2+MGY4bmvPXnEkrJDS1wTbHDp/i6
d8u1yt4hyWOLe4DgiP20GyKEx6BKneN87X1H5lH1WSHoUi+QHneHIHCi8ESaLgH+0zXFY9Vk2zPL
He9JEBY+fTxZLEWs4QQSHJTue60A0Aa05RmylpPO4wgWytuuJS59oNP7AmoCaJVywln/bwCSXBDp
ZDt8DzzK0aWRuQKcTsF8JO/9xWEUHYZvcizo1EJfgXLNSA6+eC+Efseo5cRrX2aK+qM78z4hvVtx
UoLhdqA/HGLBGv7+70GXM9TMsU2RyuQT5mZD3jOBA9IDAyXPMn0Ytu8tvg5lZnpBdgMmnN7iKPL+
zVkvsGPaIr/krXmZB/XQNJYDgy3SotEqfU+ZcC7/wIWaHbaGjToP023J0k8BFJGogCGjeFHBT25j
bJyN8xso5Oa8e24haX0FyeLbrynk9gQEHWNEIwCRaKuteYEwfTp1quWaV6nBryzWbwkd6H75vMtd
uKc+uEI8dQnrSFHk3VEukP3T5LaLvny/CcivGsj4I8V5MYzvWCQnBMYNrgcsQdzX5fYyN8P9OzQN
Zf4Cj6NFN4A1ZEhODj9kbGJ76OGy1j9gJ4NQ6LGdPtEKbRLelH/1jqPjsHYA7sDKlcFgZsralzgY
tzBeZLoAT2c+346GfYCIemjrJNLz0Ea4X4BVEUE18CfZ629mIjmCBHJZJuOAOiBMUrADRbA7ZApx
lSqSlsr7RrN4P3g+mEaNbNjxsy3iTzvVFbstG8A7Gkrf/BYMDL3wtDa5knlhCtD2ZoGAkj1rLTqg
H+MUiAYN/hLHgRFT2rgvk0w1jGI7kIz4Qt5AWMeL+DXI3sjKTigs+EJnWDFdtjNh9jWtiD9bQK1t
xrrgFGYkpGgh9lU+CiQXWIQteoVW2sTwgpS2NTvQC47kEdOz2D1T4zXDdJFX2EOYDOE6Thcqoo1K
/fgjoh+Jl2pXgZL3Wsexcm+trz2IUMYS9XFLKzZ6WTxsZg8ddiNeR2Hg9ynbr6yvDPrHY4tjWuf0
JiYmhQN+dnw3/5jabwJzLUyZdvKMPZlcBLF1ARYjbfEvibpQgQDyk28DLAbx8kW5pZlNQQLM/Wa3
TI5my/JNQ/VmrNhq+JK78Xc3+GvUhUdlPFlpRLKSYHhqrEEqootuEqvlqNZsRlMsvNlyVV39CpAO
iAwXjX4VkceA7BrZ7AapqGMWDbsY5h3L8Zq+LnIwpuXWdyVZq0BKvbaLCdJp/Kmf6oaD0waAfH9p
z+6LE9rgoMp4LQAEZxM1jsAtBdhMXLi/k0c6nJPWpiDZNnYrpttYH/J2t0hZtqrMkTbW9SMH7iF0
r+bc2ywxyIWTzQEUxeufoRbMReSc9YzPO+fZi/hMNVoBE9/5kFj/px0k50484em6b/fWjs+a/8Gc
arUxUMuf/0a5wKO8QiFf7LThWbHBh81e0c9Nnt6jCrT8wdXS3g95dar40XwEHRTuuDwYolvZJ7jw
2q3Dj4Xh2gg/+MxFRIvx9cj/UUWtNiCw4BtEf65bJI+TJqd2ekvg0UlaSQuUtApnYTg0vuRRG6kC
hx/cHDC4Q5l15LsAp06VM02SGpF4VaOf1O5AsYOypU4A2V8cc7Ny02ue822lCK78KcgpOd3iy8FD
w7ZcIbpZQw+cv4xRsV2nf9JNl/1lYvJgy69nZz7ucoY3pQ+J4v9kiVrW+GTJC7p6aCp4FtmtF6mL
CmS2HrC9poXTJsCaG0h7efkT2D94aNBFXSBzQU08vXn+wWxVmOMmeH/iBXRZXAa2c3Yv0PgWWeRq
eRiEviw1oLQafoRsAplO0QUOEirDjZ6Rsqaq2pQfKDlplgqMqSocC3jHcPxTddKNIqz7E8M7L196
C8UoDxaAwZbWqfO6C2nay9VSpd0BOFJz73z7h9VnP/3Gnhj9Yal8OSCTT8Y4Am7WzhBIk6s8JcGE
hxIC+b2phke2JQAfGS7+iQu+kmm9Vqm/wUxTN8EVlDFvyT9ReTHsYymk4vVuDzGGGfuSn0tQjYVq
aHS/anvbYHfTcUPSZxWj/q0IElPLhHY2pw+kHPJMdWptVrDr4AzNlLBA65sOE6aVvglGcPSryylD
E+ED4GV46ThuG62ekMMx1Vh1daSrAP30VACbEk2nHO9EXz64hRrOQ67ORYbZtRfoX0OJ7CZKL5lH
rTP1UDdeK3Wxbkjs/ZqV86MgqLKkY3JUhu4Z7FUg+tQUyV3JQw9yF+1dsTEc7rh7TIR0v34m2cno
cCc0KAQAElKzbwtNJs9kWePE7lPKMUw0tM+chmJ+f3qWXKazD4RBhFB/A9xLMjzDwjl7WIRf0ED3
WmFYPc5b0VdqD9MdeI24ndpzlmpxcuRg6TtBdFb2iyLV2b5CkgPRq8yBXahk5CuDC2qyujcT3ts/
nNrx7kE7NAUH1yEaBIoTHIqQT/tYPdu1FWNhoEYM0C65pNRNxXh+mevp67XPoMZxhTDYzu8v/YeH
2sz0QTaXELonc+iKW3rdWKPPeG6oBDZmZSvjC/Cjwv6qn3XhmuOcBYdjESRw+BrgBRJIf3EYXYH4
/lKijdgDeHA9vRFYZlr1MSIyKeLuGe2Bosd7HTCkfm7DDxMcfnz+xVTvXABNLBrl1Xs9+ENeN+S3
Pf7h17mAie3v5bVb3M3fhNgMtIxButOiBu/jYRiRS4ibZbP9dnre7shoZ24ycdX5XCtoEihKL+nF
5KacXQqaQkWZlvwRZhVo7IRIlcrk3/Vs14WGAWCIHR1Cw7fhcRkf93XPHdKLKUpKBAvwKzCrWJ1v
od8T8lQRBmRLXGiF2i/sl6XJfRLOTN9NIb8GOXxLkkJtb4RxDkJ3th2/VN5DHPKsv+SY8CmMnANO
PEo5ipESDB6Rk5lpkBNXuqPUO6PKu95hph0JfIK2GgfywvhEF3qE6gV8LEZV0dSyq4w0Q5m66O7v
c5BshRguErz/pD0W5W1n0cKhHt4wMxpXADTpr1kGOctp7YUvgPWk6543soZnG3UEo6demB/QWumP
hjj7IjzF1y7mQUJTF39Ru2yZ7eg3KTs3kKg/n9pGg7Gju46YN2yiTD84LIKfQR3qqB8eJUbstwcr
CA8FFVn3cgGJiaNt5KcI4Mlzct9/XpX5xXxzxwYvwq9Di5J8dtBe7duW9Boirpex0M5lPoYKQvPz
qF1rEygMUsZFkBqixBGUaIgKch/a46vqDM4jqTwrY/Ljx+8kWoomVUmjPF4HLd2To7anhZAKjS3+
N9XPOdf9TWkrl08It8V3YNJrymeYQaEdVmPopNQZx0pu3FmsipOig497AjUZh8rXbFs3H7g9BVDI
4e6Ov/hz73fqKE7j18N0wDszQAR3Kgh/xMttnNmjcHNhNgJ+ywbbklZQvtnbNTn+BbBw8Eu38za6
DTWuWQEvZAgS7kc24mKFTfvcV/DinDMlmTqVC2NG3+rOJXBhRs6dCGvQuUGuH1JH++cJP/1rSNZS
pDz2DMFZ4RtXKMr1MHWrH7HuGSwJpu2kmaHk4F7Ll8S1B0CK38c7WX32YmsUrdGdYJvAejg10LiF
npaA1p4JCB2r2LaHB3ROF6wSGuTEFwBfvMw+OUmI7FKYb7Di+MaPUWd1aLSreymYBRAXt4zlXcR4
FI/uWv+k3qXlbZTANSm31nSzrB4sN/bzzgGdAm2bJN3fR8TZ5aCzeEtCIms8EM/1sucvDD76Doi2
p5OCv2wnaqHTtWYLS05MUVcM/M4fnnrbFVv7McVHt2R4XwaJeO4YasU8WHe9jGBjV/H0TTm/tO3W
Hlx12vTXnwgZsoy6ZxLRlrz/02e3TTc1wZFueSUP+Auj/aAh9GFvl+eObooPttq7I/aJaM6Tid3B
Y/MLzY8PzELpntS8NdkcAI1sFHDsvn5c55q5f8W9dUZOYNduyskqLE0vqjm2DayW3UgbpBwwdog3
iLwe7iUxsH8ioA6ZYN4Nq1R8Y6E5StvmE5FuPl0/gXyP9ZxVNyWbIr0ZbNUZx/PHUSAqiZOQWWoz
y5TEo/9Qzi+UkTb41ItHNtMSiRujOKGNwx1DDgKA5sWvTrGwqPMPQqYQP8A5tC5a9VDwKjHx70YG
7++qPwsdcuQWIJZgkvAdMypTZpM1lZl14Px1S5Tpx0U3DTrF/VQDo02ckbdRCZY3b0B27XTKUcFS
uBB3/AthWDhMqlEtez0NIfUYhFRLc2378W2o0JIP8obOcVnpmS3RwHwxwv+aOlaaQ3U9P+R1mZ4g
eTyf9FhRY0Wul5b+D5dN3ii/E+qclPW0ZSHYsritAeIdtfzfQgDq2MiXMRPbxzvZ9qfD6e42vfEq
uqseDKstCXOuaZqDvCK3G5rZiTDJcxLh5w6Ym3srQJ8CwsR1MhSTL0Fu7mrg5bYL50iQFCtxUssg
J/InDPyelG4ZeL5ArJj+aJVTdkaPU3/+f/bpMDZNJnBMUZT8WX/fFrDcZGDOR82QrvBvdQBMSZgv
kehVUVrjG9u1lOHRjVegg24RME8XyTpBXeg5a3u2/UEd7mrD9mEAvsUJpciA66SRyu/l68fVAYwJ
PvNSQxKzYXuvSLDkZFZAw7RujslXi2FdAUP3IPndoosR4iL3GNeAoQerdBxZEW+aPatPN2SJ9h5S
ff0czfHFCHAHqWDseppnkwL+DNwPCGcgEnCiHMlCBX/8DV2i4z3w11BkmKBfbUrwezjW3KOKEvKx
wcUbx8ktkJ6fSn9/0g25wUq43RhyQAAqHefdafVFiBLDrPXvsc6wxtpDEZN4GwjSN87iF83kMlaY
0MxdHlFW/JwEKS7IwHWH2CBfD6xg9Yw4kZXSUdJHUNOVmNKqqekJBppW2yg17V+g2WBwCqex5M/1
UnkNElaj+MokOE75xx3D9y9RcrhLsQuA6ybT7dWkziKlKA833TfFBDb4edtLUt2LWmDqmbSH585G
aJvmQ77nTU2u1QhiBYUyOsFU4Obpi9madphAyqveoF+T37rZbtsvY99qqIRSZo70oIQiIW4YHDw6
GSdELL6zoTInPK/TPq/n5QLgyGryoaIAJ8vp+3t4XYu8aSadDkJoIUMUEMztSj7MSY4hcrOxB3gn
YzbgZQVKAMbtZRJzJwmuCxwjqy8fYiCzVGwzALWc4jYc8kvpkZf/cry0shn5m77igI1rltvCKDee
j0AZI3T45Sixog12rJTOibO7sxiiQKDRdkIoOfuAy9uR4udALdJuJKQaLQHnZpBmngGl6+1tiXIB
8n/ZexGSZ4KE5MEC6Ms+2viuytfgTmeHecryyaALCPbAiUufU+E4jBsLrSblzwwhpO22qXl3EmBA
+n7ZCXU0WWyp/a4u9uU+zrAJcJ0SrgrYz4NAdqmKBXKG+9oj4BMSscnl1H4cwxrlVMgpDN8AGnsh
wEL0DWN9Eb14EaZf61q1h/3pvflCFzLMgqcFucj7MOWtVLZet3F+5mh2aFhY8m7C5jhD9qPw32F8
30aKzU/2mHcLt+QMbnNpBWmxLKHo7ozaK/H+pAGfcwhBm5lLD6pyB/3HZugc9qKvqxligojH4kqt
Jb8nlXctPo1PR/NXpL7+0CuaevJVD0eizg+Wv7fzjYEn9MHNz17s8LvT7DOKp19tMbdwh0nOyuwN
YBIH2nBbTO/NDIol9ARO84dJQt0/vN4pZL3gWCnxh0C8yqr5GjZVn9Q2vxc6oEvI9rRuNjn+WMds
iWOY5BGrXeN+r8jQCYJfKnzPUDZxmN5VpmO8IrYPGdk6Bwy9z7ZsReEo8Zwz2A5PuOtbdx44oaPy
GLKm3h7H1S9N2hOUiTpQZYtYgdL6i/o9Tx0tpEVKd2HcloMLfo6mo9d/BrHFL/m7P+N4oTeXs3pH
k7whcAHqPgpX4SKn4wxpnMsm5tcPGzRrazbaEu5TgSimpoLKQ5TJjhS2cNJhUs/EDznSbjNYJjPC
oF/vjn1aK/KfoadcLqlk8YYpy/9J0SEVefDYQ22W3ZnkpNL2LrKwuaXvx2DhPB2HwmR3tYvK8pPq
1fmV8Dk0SbMuPsra+7GD0DOv7JN2k+Igm0vGD7Kyz9fSqq0h2GBRoE8wYuZtzB/0DNmL2jeBxfnB
P+F/29OytZnF0ZdnDNAbsQ6cgLQC6XO2X4a0biVazdSu3MGXC9o0hhIit6KFtlX3kEPRp2FiFwDE
eKKJEzT0RjHFKeR0ZtcCSh3Ffcvb/1dS5tqmTX8hNhdZkrFpGvdSYOE6EzJIxCLykSJvS7mHoyil
gmCtNwsCi9b28Wj+M0QNmb0RvMiK7UTH5wbbQhhqJCzuSaZ+49O8OkCbk3lYSLgpe3ibHXOjQ7wV
VhoFr7DGkv/zocP7NJdV0lqBj888vijcjZUZ+qRrc/DfZxnw81oSfHgx74/QF0U/7xb9Iyi7wBAV
u65SXj8Khb4Ij73cjU+t0Lb8hdyTzsW81yrVAQbBSa+j5BglH+Q6pXMzzOU2KwbkH7Xzkwfz9uow
hz4404rtwWREk/vIz9W0kKqlb8B1Dgo6v7pcrCQh8bnKQLbTN4U0RBh0gCoYKSLdcUygzeuNi44c
Mm13tdvDwvXz1sKdu5IdxCMgl4FD1NIH5+UVGahz4vuBnS6ugqmaeSBUrDThG6abP2rNS6ldqs7v
/5Zed98K09DBtgvkskxjJ85nkyY6rz9GsfVEYuyXmsT/Headp8nI+v0zbZ4NUZMolynW1VjOKdds
EFXfjYMqowe4MtnMDURUnHBKWVyacSl5v0/4b46N2MDRj3S2J6zKBSohqvYIzH96vcvVQwChvjSG
Ai5sbyvFprnrudkKXbyfAyimEk0yyvsB1/cFJaVggra0CCRcslA/ffBP0vlz5/sGzOQ6o3PHLO8+
6gkGG2zmdGvTXUvmubbmz5smNa7NOeAtwghL8uY1aIePVXpIiYQyiD0E2giJC6QobHvDSXNzf3NA
poV6wA8GB1LGUwaZvpGi5AsD7xnCQOr2dyIn6Zw3xXfDdGyZsK6xJkYE8NW62jJ/jXo7dJIDfybc
ldTXpenDdUjHLuJR64KlmJ4gFJBH9Dvy8sMV5hP49lDTCM/m5tOeVFB9pSSeQjo8+V408ei/mC9O
GQyqQbvkX8qGwLjO1ps6Ur6ubadsZfNdfdendlDKTWmV6LSJ5h+mOLhe6aaGE6gSBrfjBSNj09tN
BBDf4WFzaCytKumSHmqZk0Q80qNXdFLb2dJZShW1PtXr5FUNLn5BE5Y2/UWeeeYSPs24BrZvtMTX
KnzTRjLhMSVmr/KJeCJZ4U2CT8QDgm1TP52ui4IY4J78+hZ+SHqjz36aS/7jWItHqKhceESFJkne
mMDmFwwR+Lu3gYxcw8ML9Cr4X+AJdUyQ7MU5UCMtUAJFuBuE4TYUhCe2UGZZ7EUbzSinzj1hbL+M
xySS78zDFJW6fWNTMsMJrGblNfKv1R0YQI32Y5b0HqCJbytUXA5OOY/KRRSn2tAfTIxV4a9WZM5I
jwqIHBNRWu09WOFDVhIIJSYFKySrsZDJfpTQOQ2AOjdZlRqnCoHUC+qmqkKwNFl8sebVyZTINpz3
SeLAC7JL6vIQIy9gXTKQQMZ8KezmUxjWX0izPbVKoLCXent1HaBfbQJ1gZV0CxGifSmHUzHLDY45
54xAnYXoxf8V1mu9BM6cXE43q1+l6NsMG58c0tL4FH6VVNYLYmRmbAXOfmaVaOu0y8zOLiKK3u9n
1kk4Ko3vNSc/nDCV0N3nwVhswwRtui6b0PaercpYPo9zy0m0wDA4C1VSWtxvECGTlFjEuSf/V+sQ
rtrNm9slBrYqiHBXAb83Q9YtPuKqaoB4ML7OusCuR8JC4vWSI10H8sTz/nNgLZDYgXU6WhJ5J7El
Jgr91wSBtPdFtFweW/hp93KcALHw/OkiEdRQWEJcUOfn7DmBfuRDf8jb5PV3S0/QTOn0+wkLWfxI
1ZWIGYnEhkGVKLurk6ZJ5u/ngfOFO2C74OXxs78g0b6x+A48B2Uy/I4hpshtEB8+6owfSIrgodvd
q/oKLaPGLkmtBq425msdkQiy+b8UqLN0G2N2KOdeJvuQ5PxSZZG87oCjQzMfok174jD9ocoikndW
nV4r8A5+mz+tkqDbYXRRopurlmpNFc/Wc2lhLBv9RUUCZCbRVwIlhUeC4LZ2fqy1ghkdWS45pw4K
65ab4drkSjAbIHV9evxAz61RwNF12Y6ezvlelydmZXQTujFAUd5w1FMRmD5r3gV+i7MLBuFbVFNV
ey3S9Vu+q9BGWHYMO7hdk7I3H24e1nqaToZyQhZXNfgOdMgqrmonkv6Fa46rb4n0E9sQMNxSeGi7
hkjW1Bc4lZvlsBuQ9/JlyMmlhxAX3jtFT7gMha82OhgkLJ/82qch/vwg+yHbWkbeSXLqTWK2Q4N6
eOOW3+PYPHJbEwclI+gD0JMrfBq9Y+8rXIoQ7b+Mrxz7Y4Z5E8OaU9ByLzTXG/v8xs0cJPf7y/T3
VM1eM/u1XXGt+JKIfsxpKiAqe6piMFTd05Sm8UDn3vsYksI3HirpNB978jdsxqCRcvTvxqsE/58L
mpHOnrja1f32zpmmOO/CtLgI05qOnj/FoRJANOF1YhEQdGYZSSoRFpW0g5+2aD+Il9dfkbggLvjz
K/irFUmvtqcUb5nE5zadFSnu4tkrpam23vqCXaMhWC/zinMypsdSzw7NY+VWzwRnLcq1DkeAiVY+
EfHBuUnsVMIw7czpPyJn9O/mS5uxZxSPgUH5mvDY92XgS7CwPPpzkrrDxh5IIQezy6EwNGk4Pmq0
+2y2X07a+e6/nX3cdCtHK90+y0jXjkjQCAOJCwSGYecwILzEuEapZhgmQUoSBtyFyTTPGzJV8oOk
l72F8sfzbw4UFmKGO29sr6Si53C2FTgstoMZAm9TyW9Tyo0rxcbSZEDf6kZHrV0BrdPpW1MfUxJI
tXJSJJQPgpjFoJRlPVBJFlkWU/0l4BrmAHyCEUpfKTvnHu6Esn7ptu7ciwBXR783yjsvG23Snr/q
oSalvOkzTMWlt9I2rhaXh9Dcyw5bsoHBwbh7IN3c8vt5IuY4+f2SFekrgH8Qn1lGy0p+cGlS0mdY
L9rL5zjnQNJaV7oCkcq9f75odBGHD2qTlLdcVTD+jovIXhS4dyks5TxItFn1j42iJck9ggY8eBZD
xO06fqTMZMuKyPVIvPeCTRl/mTl8sTvk48NtCxjjMjokv6+8Zfy/Loktlk+My/9k/FVPELH+VcmF
z4cYvmuFUAomjwv5cmRLNiBLwFqvwAqr47KTvK+LlLBZcAlO3o+eNssT0pSsd8m9Ga8UYDzGuMS6
Rp2mN4GE2rr+TKwXiA1ZPpGaE3Ja/wdqnwbI3o8gLhqEFr+5rdCyC5HARKUGI49+2UZzcD7OrpO6
2eJogF9YSEuTuzP9k++V0cOcXYG/0m42gEMNJXfFivzfftq5pYwNT8NNDcTYRVZyQEd+wM50XfDI
gI060upEns+yzmeCz9GSMvCaFtU7NLK7fdUUamWOfY5HIWoeDLQBAyJphKc5D7FahNlWAuLSs2qo
L5dt8KnBFSYorRbp88HVo7iLChyzsj5ZY0vMgVp5b2LG9RH49ftB5hwJO++SOPjtvuC72Y+FNsb0
NmA4NAz8VbsRwCOjpAapJkSsPQY1Q0uEh5Ca8npbZPN5ONvYU2zWkXtUE/gU+yEvhTf1xFc7zGDc
svTPGCYEaQF526IVGZs73WSHyTeVtlduTT5wPH0xuubSBrbcEnATAX6WuC/grFXFKV7QnnXtzIdL
cdckUI14m/+hNKraRBeKuARI7ihG7mTd+wQmXa2mBLG0PTrwLVZhYwCzHevVLMfuL79Dwrq+Cj4W
s5zs1Q16nqkNYbtuQ2APBzeqG1s6naSntKIoQoOsKRBVJjLTlUXK1Hg+L2WV8+BGyeTl2uHKLgjp
ue07IOtyflg8wy+Nc86rswXA4pj8vcrh4KCEhoVGHcwuybzgTloxa0RKK0Y27HBqzTeawpIKwgJO
/Nk24mEgVweEAjxpuvKQSh0gz03auNIn8P2ctUGmkLXjEh9wJZdkoOkN2Im21Fs6PVBQcI/Hd9fm
94czVLkfq4uTq9RcISIOhu/RECaonMXAVJ+1x6W0JXhBK97u7NYwA3dgjdyLSpZyCuMeRvC6YaiT
dvfy5sXUGb2/T4+fggPrIpfy27WC/V/KqMtjAU4bB68xDO0+se/F+e2yYsWshh0CQqD5Um/lT2RZ
cg2H1JBgC9Atkw5sKtEjrMCSdx7i6iwsIayIZ20F3TOPPB9vZu3fhkWpqyI5BUc0KPfEuRo0gwbd
qdQjDrenfff/FN7X9grSV+0XhSQnU9oSLn+uFkqtrM+oL8vJzUnElBwEkilmTUS86roGGgAijS3a
DRU43VH4JDKUfjrdz4AyWxGpz0wQCFEbHhLD5CquWHRFPGLu0eZeRpRMP3L4wZrvUMshKxZAWhNG
FDdaGJ0JkNdFcOVGpQGcItjBst4hT8wyWN+lhjB6oTa4Mzf+o1MMzDjzI9Vst1hV8OUSdzQfHOdF
Ao4PBRxsdPMXLj/nePiA7JrX6HtR8KxzZHvb/vJG/A+/YRC4kL0bAdAPpR4NSmn7k+mp9V9wgMzk
JvtkLEU5BfXcNcn/4Ju/+inCqKLTuJtsn0dso/oHpK+sbmL9CQ+1ztioWEwKbYjGzTHKX62J63di
U/0QrzcKGsAm1djZoia3xYQPzgF1ZtdZyEu0ILK8zzxMNt6UXt4z4rPcwpqHSWYCM51W67ABRDQ2
I1UhYH97W5F+nxMJ+ovvqGtsJHdr+h5/MzFUMgoE3Pel9/3HEKmmNAJe85ZGA3xSfrL3u14BrFWQ
PfQ9PBUH5FyHtCjNSQI0V7oa8CDVWrJ32fB46wYLrHSZDRbMkTaIzP1Bu1R5VdYIUhmyeUU33vhd
Raop+pariNhLOlO5JjSN6vOU/wAOFdxrGsxzcujA8kI9NEw4mhTeMweaxKuhnKqz3vAiC8FNqW6X
SvhqfLvWvSEICm6KJojQ5cjyRDBtcWTb/xfeGRo7xPrCpqzvEGYWsDkKaihkZYXNKbPuK9weRAqd
czViBeVYM24B+WgpaPsZcUovOUpVm/QUms28/o6s4VRyjMDI3EXti3jCUJHiuLh2xm3eFYpnJzeq
gQ==
`protect end_protected
