��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x�O�=w�����v��z��I�=nQ��t��S������C*Ё~_"W�3�3���,�r�J�?��D���_vއ�j%�ձ{Io@����YU^��A��J"��(m�)#r]�����N�W��G^�)��O��}Ȣ��C`�����]� �޵��o��GK�b{8�����`�A*Y�>�ec&�e�Y�����gu���	����2�:ǼW�}.��%�B�C�{_�ޕ>�|�Uv6\����8�[�Pyv֦�
Xí{��rNƶs7�0����z�j�]�p��S��3`��������$}̢�.
˷�+m����8_��p�K�6���,۞�$2Vg(�wf�{�ht�੔$���T�X�o��}��'G�G,ӽ����|Lޝ.X����d��'dб	q�ee��h]�T]�VQЃ�a9Rpb����<��'��=L�a3
�6��C[5H�#v��b͝��W��w`|cpfo�m���������(�~��!�z����o��RZJ������d2L��F�&�}���b=O��O�Ku��e(
Hؚt��������4�Z�"���y��gH$�b���i��y6e0<Wt֩�1oo�!>��:���_[W5� ?��󕬙��H@!˝�N="�@�]p��pQ#�'<�"h�Z�Ȕ\%mhO;� � �x�Ltރ�5y
��4ߊ?W=,��\���1�#aw���v��V����#?��+�5|�I��:c�`cC� z�џ�=t��
nE�a�}{cd7Z<+�>#(aB����?	
#�Ei�"����E���E� �wFDn]���]I���{�q�.AX�?Y��yܻӖ�%{㐇����?�9Y9��؈�P�9X_aЀP1�����M�E'VJ��Syt����D(��mU�4�9�"��28��d
o}T;G֝���K4U��1f���}}�n��^�"�	4�2�&a^�c����nv�sڛ�faJз�d���3�a�Gv@?*�k!�=�#��FJ�ֹ�7牊�&
q�?^ր�O羬?��O$>���^�iݱk"a2WeVhj�H�~բJ��\q���L�oH�^����A���`�B=\���ȇ���k��(���d��+D��c��ю����AYJ�Z�7�%�缀V�+�a��uk��OC��6��G��N��`'����V�cATka���@}ǚ�z��l-1�-�0��������~)n�弖�ΗU��H��_,�%3��\�����iExA��uE��9�4����s��W�7V�����h���w��C�����X��U�2VVv?�.�?(_9Tv`±�{�ɐ^�i���!~��m�Y#݇������1PXI�u�ɪ��(��-Wf}ө�A�a7���P�������է��3ߪ����bpP�~��%
t��O\u����4vޜR:�� �0��0��_��}�T.a��[TP���cu�b��8�Bl��B�{��Ġb��e����Ǒ�E�;���5���B���_d���4��"Ǟ(��*ա��(#=8��G�*�JJi5������pȇx:��3�Y��oϟq��D����0����2�^�h��	�=�Y0��v�lc��9��+n�	̊h�"��b�2���j:T�.��a�l��2�Xyo�������3A�i%�����57Q8C&�M6�h_R�}��6|t
�]S��Ԉh���n\)_��S�*c,�G���� �[��2�Cf?f@����ck��"�>�'�u�˜�(����K�Z���R�����8iO=�1D⽂�P�?�XV�ss���8��?��P[��-��j����I�D��Gm�N��+\
֤_� �8h�Q�+v�Ж7���D����!S@�/�_=S,�i�%�eV�E�O6��w�#��QP�F�{=V;�6������:���I�.���C�_oQ�(�A/��)i����$l�����4V��[�6�%pz�M{!�W�=��҅�ئ�2���u������b�N�j��=��?�x���=zٷ�ŦEB��DGY�_�]7�Qy^כ#��,��oǓ�Z5;F� w��|o��G�S���~� q��}2�u