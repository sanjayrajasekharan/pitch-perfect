-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1b2FhHEPaJe1BSnuS8as53ZBhamVoBm65LmJ83du2PxTd5PlfI1Drcd0FU/eReGwMdqYlWTRDxSE
7F1WW9e+ZcIzVJUxw64msaC6lAI1RTqbas9uuwAzLb3VjZJG5Qg3YGoFKP1TjinH6PH611o6yPUW
AfY5BNLBrKtK8KcyIFu5HBrkXF8UDseAB3f7SoozYtk81arwAuKlfCYOc873k97cE9oLhG8z+eq7
kZ24NklK90TT9VB2R7ly99pQ5yNqRK3eyGkvEFHXHkEGcoH1JsVw9VPVfkmF5ApTKc35JdjeFY5m
UWiNHY8v5jgbr8TmkjYudpvddOJaqJZtFe3jkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6080)
`protect data_block
lgesFqCEoQqcTP54/ZVXU/hInibkyRR05QzcboHOsz+nBAYCC8KPxlw6LOxGWGKpQX1FyCeTESEI
tmxttEWatH50XTuXQMDK9330EkX6Kjp1pp83kC6knAW+94XKRHVHRH2bFngGFOaOvwl8aylbJ59C
YTfslwZjmF5Zz1mshdBNNiTu5TSigfk37Jna5OLILUQWT7eLfmG2ai8Fsn1KqOB8VceZY3FPL+TH
2CvVdynGfdnGRAgfNLDrE6E0WZfOh9CHkmDkA1CrTK5rFGJgwZCshdYnbNZswymVfVT3H+oweEZC
WXP5r+bfPrL1MfQSq7DzUcCINF66xW/CKNCesQc54rXpdMeJdLDNx40U65q3782yjohOOnr9Vjfg
XqxY6PNexplerBJIerNtGPGd20YSRQDb0dYKfyRjxhzogCuVyqnc7uiVW404C2cqKBfmAsxw5vC5
smYk0DUlxY5ddQtN+znks2rhle/ldg/n6U2FtWJyGAZvo8M3emdqWX6OPcQ7Ec1BGs22UnsCddSy
fC9Bvc6q7o2o0gi4JaWHo+jwblxvdrx1zQkJ00y+KVTT8fehu0bYxEKTB56Qy5ZARKeRCpbKpcUE
O5jO+D/vipB7x0MBVvC+kJhFJDKrb3HgITu7e5rNBxhFByxbO5AqYrWk45re1/hop5IaGTtSLd78
5D4hDuCsXab/IwehpBN62OsJpusm5qVZ/kRmG8tmjH+LhhVPLjnrEdeq2frbEy7FF7SROTqHq4YO
5KpF0TlsVHt0kFhD1THRWYcIXBsoGDV6GbbjZowtTi8mFoT4ah483RENAFXLugOY69UFvfMPzKK0
y6ibGNGsZUFlwLSytMvrOYIWZ80ZSjyXsIj/8EwuDFFsE2aglVjj0obILIvu3TVj/24O6CAJxRdI
ZqEcJXawITma+jJRl9+LQgVlwOXGfX4ZUSa5hpQDKBE+XEAmNVZ59+mmtzX/7KJYz/2C+5QCJqQs
NBdLXFzSCIv8Qp3bRATiIIv8VDSg9j+flh6dhVczholyEOg6fyh0/kwkYYDKFUic17xwGlslYKxs
XD3us+52UBdAVaIOsxFLfAPHhq1IzaDYJDf2ukVyom3pv04u9dV59Tg+g9g/BI9c6xu2BGjbWo6U
oZAEVCQkmDQrNXbGQpscebOn/N5MSnL0oCeqYaECZQvfclWRCPi1aKC2TdqWaWpiqfgF0k9b54h3
kbx0Kc+P1snM+ww4tRSqf9z9s1cFTiyYR9e7VGg1yI9HdAq/l+N1dVQfyhfg3urxfgveCM/ib8nq
MlrV0Kao5BKC+X25zRVb9jz3WGMqTRFwH4flcNS+V4NZe7wcyYGJmkrpJ+H86MpmG1OIdOi6+fNt
gnn70SxtUvxp5wYv1N33Sl6yyzgizRvgl3Oj9Dc6tusInANPkCK1cgQQByqLNbqf65nAOpLtdtkb
U6MccBaONz95nIFaQGPH4GrxS5doItFhU9EhwcR1EQuN744Lu+xbMJwAbDNxYx1RdTdAf9VNZQ2J
ipnudCYD16WlFselUVQnw8ArfserZvDbSyJWABWIYFTltfnKGDAzbyoXv55yJiUcfMTB0Nl4QEBP
Tb6xOPvFGPvq6oRfSaL1SCG9N/7w2zbbu+d278vmwDN5qUFLPS2xS/dg52H5YpCBivj8ll+Qs2aZ
Zpkt5xo1OE8FDo1b4sc23WHts8Q8yS+AyNVCEuVj7ZL6QftwEhKlpsnMISOhxZZ+0ZCtyePMYwCs
gU7dWf7Ne+jn4d6i2QspT/algus4P7mngFhfEp+l7NaFL09Vw/5VCnk0RHTloOPJwGSI/blY0S1w
FzCLltMYzCXKhFYzb/fU3uXa8au8LWq1++5wiIjJW01k01xiDsfeGrYsM2NkFsLl520ZQ++jM2cs
fHPk05PFeUNnRMymo26SclyZXxmRaRWbKQQBgokN5COr29yYWTz1DMGVMmYEaFbg3rTJ0eUxxWQZ
6+2WArXBhXa0nCHGstnY8ekT5kG3nxyONnL1fdi9asOGNIOXy4UVJtNxOXl2nCcCe5DBmyyX5wjG
PrgRW9DLo7MOzHT9mWU5RD+TkOcpsu+8lDlHpXgG9zaMWoqriqLt6dD+wg4d0EbZLrYQxk0cUxJE
4c5P18IjU9i3tjiXA92L6OkzXo/T8YcOTtXF4fv3YSkXo8DSITXtQyP7IFxOWQpFIgb2+8wcedUq
SCDLvt1EjZbbwFhN/3Nt7Q1fc43meZ1AGSFjq7HXMEuDs38ulq778G5juzJk3Aopo5a1zWnNNLlj
hxfU56e5g9riOfQGNOu85ZeL9AQ5D/0AXNMjbKfiJORQ/eir3kP8YlJR4loC/IxSS1CSbsw/+zd2
V0H2ARPCRfyG0WNShELprK2ziwc5255G6ZViGfksLne5V60wHPrslWUgshDi9FMAZzITr6zNoH4R
tZzkmVOy6TCwGciOjPBnp514dzkSXMo/jJq1kgbV01oWXk/cBzHbblK+arDHTiLMjq/lFw+dZrrR
Bc/ulYOrQC2sUoLZ5bQ5BGsq00f+WYEYh4IXv6j2pXc8qMvURHL0fQRMfxQGx485lbXDJVBC/B9e
Jenan+/8LuQJ38Aq+0b4ZCgsF7HxCGBbjFHnTz85oq5tZ76mdUbhbPHX3zF+rPcK+JDYMLP1ovHQ
1Tw5JV2a0acfvoDwi68UW5lvNmLhS0J38nDk71NJ24CWocPm33f/LTvvbKyuimUQ4WoQuC/u7Atv
VBQBC0fgg1n3gGAW3PAFiCKl/Qibg0KQ/6+w/wVUcFk4HqqVuqu1jL67qTxzrXwZBAthxeEayjXn
uFPUkBM0+JbtNogl8K9tZXzK/ffvVXatwc8zLfAL0YQyyokpsBdXUd1vsl3aTB5i8juMYSWhi0Yc
M9az8z8hMA2wUb0hcM5NxHY92W/JQxJMgX5gBwro8M3uHpmBm5jQAnrNxZjq5K/p+IEW8ynqNceT
dTd9hCyiTu8LA0Pf72DzHqajYGTneT4qyD4AXdjA7xN0P2nKBHRpj7rXKA3BPHZJQvRijHNL+wDP
HnVa/V63BYKVoBOOF8das9JI92G94Uls5Yj5nb5tgBXFLmqiHCimjTAHGQQctGPXoT9EGhHqI9Lc
mRpM0q2Cg6BAulkcU1uKk8J1IX6xI3Dm9cVu7MKqBauE9ogwSARhs4edlV6ARdYcg50fSTqBtf4b
Kf+X7MGjseUT4RnfOqNSZaLQLFyStTZGEWU71/epQWaLm4jE8O9FnO4XbA4PJuCVYeFU7woL6qCt
J6uBLbrVj9p7N0ANMdF+jitfWKJi1+xLWIqscjKe9OYOuKrj+fNYSAVpDtHiWtzlI962xfOGS+nW
7mTQ63ONXOxtVHZxWpzk73Ujh2O+F6kVXItDmQCuDnfV3Bvy4KSwjufL5+nsGncUSGbNsq5VW/fn
ZQyT0Cg485LiwNJek7CwKCYqbP2KVuo6uzcSu3DmaDOVB1mICdFlJalkW/VcMnLX7YiUu6IouAkG
8OeTqzavEDRjPJ7zFWJnqYldu8a8uAD83xiEQItG+s0HRkxAAALYKgCqWyzuiJwIxnFQseJs69nN
zi5FldG/2CjSoZMOLTyrVDeIBPjWDeYPUMl0ES9hyDFydZ0O0nbf94l87tXsL21gcYbrgLTRWBAa
Z6i5nEX7kApAo47na/Ylhq74bqlI7tkz1wRJZ1I5iqmdCFLNWDzliHnm4nmwMScVEl3wnK7ARJr7
ecn4ufIYCY9xqU7XOYhoG0dq46oHzX+WpnQARtdHkFj+p284TSgY6kfuc8NibRZX8zayHTctGxeU
i9TULfxCGq6jdn/D27zosU1AcEGQL6mpOsfZfpKg5q/on+nOy8TsmcmToDpOBtD9lRBrdVrapZOB
WnIutuPSMDf6PUYH9xFvKSun5esdB5cMYGZa5esBNAwWqqYC1PUuF/Yzz5kNHut1QuUbe/L+halg
42iPxEsU3bvGxJGsRoRZAFvQM6ETYBplvbrx7vHoq8ZN9HsNvOpLH5UcnyS/cJbVU159r1EOMS43
BIjRgRjSANNEtGmRxfKzqlBcrbUzUkIHzIa1mAEl9f5r3SiXay0dZX5QiKSNJ2uqkCe5nOn96GgH
dPhoRRNm6Am+6UY5mVmT4zthaZHZC9s5mQXlgKOPn4E9nDxpIm0YfZX+7wVb7+gAAFiOfdbdlbBK
fiP+VPpm5KFUxwXNElmGhXXYVumBB642JfPl1neNx4XKsCofcZ11GpOXBdxADqN92HvqntXT8DII
fIxZB6/r1039nwHbK+foit8DLf5Q0xFRuu4mc+ZFNXVKTUU/c2sFLD8vaJPbjybPpvfgxDj2Pv+J
wdJpD3kmXv3LaPuANu39+DuOLuaSTdltliACnFweh6lEMlJyOTCj7gcgDElgDE22pkHS40THrXMJ
Xhxnd3WnSZ32JrG8OB21JrNMuJsgXGvisOWhJsjg3XsqM+xMnShl+xf9CuVDRVMFJiRPOmE3gacN
KQJr5i4wkNJ1Yh305o+/IN7FZSCggQJisGaLOHtDT9OzjpP8lzVD8kN6d608fYXqWLJ6srHbWhbY
uUQ+TH+Nxyuzs3afLwVrw3m4iRr30nVWRuqEfvN0g8oolppM2cFgs/AQX4awiSStmi62KWcPhBRU
K1EeLlOFK80rU9cIWwejb7xhgTSHBEsUdPhOr0hTlsOko+JMsgQUS/9votxOyEbF+WtCbe/awVXX
8teoYlYsklnJxBefXt9m3K7J6twYvOSGIVR5HHny/9NOM3Jwrzt90U95sVPsEAU2wzNxXr5CgObB
8lvRAXUUXB2dgCecu9VyklZIHVRXsoEsNz0u2bMrzUgIC+LKlGKxTdDzr/Kt+ii1/gvs4ym8YMc3
W9LPhlpnRACRjkjIPrExF2CtkPfaiQGnyP+AeTy/ezWQuyWAW3EXHkzp+YyV3IqZGvBgKOGaPKf2
iPA1pee+Ji+wJQvld1e7DzgrCH4HQl51kmbKJXt8Ynwm4zAWEenRBCnZMxCj4nfHyQPFVpt6FQLP
gsM2S5htJmEeFSXgkZMMUJasjwChBDM76PTH/Wi3gu5CdLZ7Eoiyc4gdF1CHUUCDecRoqdaqgy7a
VX3R9ZIg9vjvfrdCH8Iq4r9Zp2j3z8HtScEf3LdXKwGnQVEQrDwmTA+idrif1Ou+XJZQnTdYrz/k
7PzwZ7nSHzrxvyyqmeBh1gERhDiZUcEfZGCVwWmwwiD2heJyrtYNpYpeK2HXvrmKzgABksUqdyQx
Oa3lEaSBeVeDQaEa/XtS7TcFcSHYFcMnzYpj6KjbxTZhTOumBqpMFghaOuRdB5/UOmlVGt6BZ9mZ
FS+rhk84hlSwu1i32yylW2VCEhMAo8i3AAwGqrJOuwohvhI3vN3C0mpy+QaCB+FEC0SMfBhg9iO1
6/mZ8YGd9d4FRQr6/LmoGPU2nGOIKzmVrY53WWSWBuyH7OVSVcvTX51N+f/6vBeUt002tjHgx1Gy
kdkNBU9WF7WTgrSz1sjOV36q5H7WGLDTn/bXHGeJCPac9fiE/SB35ny5PMUDM/uUJQqE3rMptMpB
UdPhBP1X2dwQcR60xEt/RFNJM6dakkEWTXu0UGm03zFN7ApJBd9NQbtxoc6c8jaRKW8TQKepo4YS
drbZSNLmmiVVrhfcolhSzybzr/GjlyQEhZsaShy10ci/5Dz+tHlkNBjFeAeMR+zkITEYokKNOHcP
LvztrvYFou3bjFSWuIbrHxDiVf/B/DeEc3/yzYcGbbNdKwJ38/egW+uiu/6LG/BMgQgARg5b+TaY
nBkg7pk1HeN4irJdl3fJ3KQyo74A2sGBc+sJrUfBDg3YEP0/djs8zGQ+kbozzZyxvoNSyElk+Gyc
Ne7J2jSa6Z49F4PYwCQ7TDWu7Zvdy5wWeTGnn8VWnhPlsZeQGf0XalrxLAYHMmlkT3j14nN0ij0J
cbdgir/iiLPN3PL1Mp0ONJkRJKVtfUp9XxuLzn/c24bDUJ6gH/pqNvaZXUFA9raggISIkBv5elUq
TgdwZy9lIFqj3Qn0YBYXqOnMK2/2ONtpzs7FpEN75d0v0ch1hfv7aWLKTbX6caMJq5Hz1XOwyJ2M
gPf/cEm7ruvCrymmNkVSxLHXQgnS/N/Slbq3nTM7ISmcR+l5kXXoLHZfPpPDshA0LzkpNEgAqEkP
GQORcXRZyAh7t7oxWevjcZYQP7Hj28aUB5/r/yagOYcT+/N53DFEgHwCcoiJn6r73/NnWYnOKcO5
XOIQjuIwNAcCI9MUzkc5ovKS8ZHyUyJy1ik5iHkSr5adp1XhQv27rf4qT/uWe8CL5VMyXfWrYzFX
WjQ891OHTytZsHitRsyJ5sWRP/M5l7PCM7lwMwB9zO6rymMIewBnAk13kiJWuurjqBy1bjbDyCdF
E1dhO0bGOEejQLJUAX81T4l0dYFsCuK/NWu2HWnR/tkbj1QuZKst1vTw5YiAxHHqe3SSjKxZq3CU
nNqE+8VfGG8kd9I/7KR+m0xXceeeBzBIk6o6mdHI5UfR/CpGdywy4AlPPRWfaSrkPJTTQBE8tZNh
h+VbgZUHRIUKzd/UgcBeubidSQGPVqOu07rNVLKepXzDBifvZ+yQ4YCdu5eTHMKVFR76oyd8kE0N
jLJwkj750rHX/GLnTx6VZ0Eh1purTkV6BFPEBlT0TfwpICe0saQOicKBYBZiAeCInOnXPhzFDqS4
66wi89j9B2dhFNkCs1j5cVOBhq+Fm9tLc7Lh969iWimlSP0HH55LfxPNG/P2+OqjcRxuO+19T9hK
BMsPPNQlMZ1nG0TCscvgXDTbPOrnuXwV7kcgaPj3RsI1KGBos/FORwn/DFFlekPL4s5ad6zjMEXc
6jiQbLhSx3cgMrrBKFMHWYnkZS1Xh2Y76rxscLp1dEiZV0WxRQcFwM1t9mB3y/7TkJgpA6BUqlFm
67+7FSRGEr32ErnR5rtW1zuvYA/1BAteTDpUuPeATtHN8r9J+ZW5zIqB7kT2GbFeg+GBuUzAZr16
dyNz0hzpHat9bVYJjzgfUlg3b4nH97A+1ZtK8I1cBGBH/QAI0ar9r6pe0jfyC2wTitLICY0faGVU
XUmWlrA3RlfrygyhXDHVsj2ocBaFexm5DvTe/6eag+9nEOC58BmUO3gV5l3T6pIJ6FHoJS9Bfzc0
Qq7YbryBfBxy35FlzRWfEsROJOXJfoGSfMZRfGmRVmPIKr5+ty9/kUmeG+AOqtnWuJU8MTL/ex7f
NNs9BFcfeJBHa2HddtLw3Dy4QV62kGn514aJHo9miUzskV7jfZ+T/hhzV0xcCQA9RsbKfh4JgfxU
1zbBeU+aMP6llzI8Sux4qI5pQy3Qoc9YjSwO9v4KWhd6zaxIa0I6Epbfqhf8zwuYaRW6gcETqlkT
RM5/xZFkVIX0SJ8Kdo849/JqLVpQxSZ/xNEIg4kOJ2XXR7Lj4eqp9nGIijVulkV+7RJnbbU7UeUX
FY5rx/rqi4sCnGvxGcm8wRDkeixF1Fsyo/CULUqTXyUP1c8/Z4I9Kp0ulORTlSy4mDwcPi+aPSvG
r0fcuwGX7ERBUmhtqFky/vHmCSOK9T8qPTOXMBMMB2Fw/W28Pd7WEbIwDZ5vjkNBAUxTWQWyE5/l
uCYQAecCsBPvwFM6+H1cY6No8o//iu6z7d4I8W2/hamc/y66cxAVkoMzzbLToQgkunvIY0RsDdC6
pr+U2wOzUeUaWQqHvrdZrjrh8BcJL/hdJdFIs4cKLRCnx81nFUD4qARAE7yl9XqSg71FGcdA8QKu
XNbnS0D7Jf6e3oPK4rTUoZjO3qlInIzAVrp1O7dc/7AJTi5nm6i4M5MrhUum2KIuIYIGuRf6byGO
+96HTot2EArCVebMdQEibzZF9CBGL+daWp250TuV3+WRb2YH4Mj3Uev0rwqIe7nzAx2DAjBq18AM
hOyJ9Ma4AQPQeh8cEMCRY9ENil1DmWjf1MgakKBV9Jv6tuWt4czFBvdBo21yUivKs/SjqZFQ4Wi4
hgFKd7V4WCu9ubbyoTjxZCMOBDX+VSeIfrnVz4/CoG39bftfi4vzQe983Z+CcRt48DLwgFd7jxsC
UPYlC5NG2NtAjzDXAc+VJLGCZanlxkjwHeZYxRn60azptSlYX5k=
`protect end_protected
