-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
JhQ2OgTCfwXDXgtCLSI6r93d15t2sgMZvrLp7tPl6Bu4qmgf/ZXPsoPTmi13Sjhk
SPlqBALb/7zM2o9yfG54kupEoUbLWppsZ3AYefJdj6WFVSLwJK25t3C4iy/K2bWg
h0iOxwllBcJfXDzO7ktpBd7CGgbaA9aiPNAVVlx+aQU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 12077)

`protect DATA_BLOCK
FULDpq77SRshmTwF84WuzcOTJp3CmiijBsqhOqWBXF1kDFZ0CnihaVDnxjX98Gdl
8skRQ2iLsrMSzkG33vHjv45KnDxYicPvkybSnTIXOnZmIgCvVIsOWjTMbHYOeNjs
1zqwFhR++UzGs5SRss1ZBOJQZSivPZ6vbwxawJRH+AuOolZunPXSTCljJR/6rY8R
xrhpwhOfVdKiU4B8JhP6woVLOH76jInHP7twSNeSWln65dpiBGLVF2Laf6UtmlJ5
U6bOWREle/FxBHMNe93Ruw2R28ilGn6JvraFrf48mypaEQs+CyhwanUQERSIxsCB
sv4ZeTyX6sS1otZqRkm/TTCWW8Sj3ZiJCX/M4iy4hyX4ylqXjMlDZsD9Tjp/z8ag
CM3XsV7rP4W3Xo5YsLW7YagSCRn7HMy62HeooN6hwhKMw6GDsky7PbHsJcVhadai
p2UUf8o9UoO/P3X3sWcroCFi84bubbo0YkXPCCVY4yZMVd24JejhdG/+K+k31KCG
rv9D+oSK7ic9bCrMsL/wzTZrUZA2x+DR0uvzIF+E1LEcuaNxPMyiLq18hOb4ddfm
qMCGovJ3xp73pissYR1BAN4ZGZwkWbBd4AQP3+xxWI3VHvpJvWU+dRIeN2HfegRO
M0fDb7y0pXr1BuYPqVP42ZbQq90IrWtvNYatNPh8exIU3gCpanrDdNZnDm09Pd6A
IGTUa6lspK/RuqBMZCkyvqmpTHElnya+a+QCSB2GuBe/Rz3LnM4OOzqSXkUZFrzT
cWQWf9RbRnir1KMeBszrZMOrN4Eq/yHRUg9h6OQHF9MXlB6Z8ipy9V/VlJoZ6rat
wUHHDkOgKidrvJbiGEX84+KZp5nXNXGWIpnHFShmuQRk8M0FXfSPGYUPP11YgLx6
fyILUlqAZEexq5IG9DRBWs/Lij5cFsHeM8PU/P7C96tCQWv2u7U6U0GIUJCAo9lm
RoXPf6LehudkUgvHc5z8AUVH58PNuYeAGyO4Vaq+AV/tcTZ3mqaIlpGmiKD6mKr6
87dyME+ssrCbAlEUMyARaXxIR+YukVXyyuMSUGfiR1cCa3WafUwXpbLbP9WN/sZK
QB95KB0ccpK32pxAAZXGbJj3wWQSa5JAa0s59vrI67CNnHJr2V5QZSNgjb2lLxTQ
QUG8phFrjJLCwsw918y/moXD7ipahjwBIpigmbfvki2Ij1kLAQKARNu1X0l2b6rd
9H4+5uE61SjNlmbZqgYCG3n/6o7U1qxX0CIzSzegQ6mbfcNHOCRK/Zi8BDdzgz6h
sm2nexmnqBL1EkdzLN5wZSnWP07XOwjpyhr9qcohBd5TvfOWA0VQk6nfuiEW87a9
4CaiYph5UI+xXo5Unnk56wFc/I0Mvws2tR5gB0ZzyGmPc/OI91EMZHpUrgRQWZY8
98AZv9Q2zjTzPcZDDBhXQTGThG0YRToihwrTIgzZoP0+wF0JzCinSMYV/cECFR23
Gnf0+P8bQuywcAlTaV/DlY8Ijv2VXgvP4/B922XKu6cguUyGmUOu/EUZRzid+Buf
0Nq20zBo0MlfE0/t+ldcGlnfr9b56xdYrWA689gbFICAy2GTAqDHC5gmNCg/Tynf
QAptNVBp/P0XdbxL9MMMNPeQRRUSIL788jHqk2Z1xhCxhgQ2y/900eZqNGFc6YgQ
3sHKM+8tJwnEI7/Itz0fQjnfTmDZ0NN8JrQkdYWgC4/lRtgYn5qCrPThHx7vvRyT
KzSbY5cXSBQW/NP3H4QkgwaSPMVoKjymn7+sp8cDjjr91l1W/RINvgLejLQruo+L
tlzsLVEVd5o9qAFXbG/y4GLRmn1Xkhh6Ttf7MZ1ZU/oXAsW4sKTFwYZznzNP4peR
465dIXg3Uc20aBGT/SsFfH86dfhHvt4e+iD1M9MeJdd8Wndb+uFbz2U9uVzVFUfa
IGkavLfDDT3WQwxHo5oX1cSsOSTWMy8xPlBiHLywuNUNN1oTcgVy/WGzCWhDW24l
21RBiKyUk8C7tdkOUhwQj+PB6xjqsjOIsa6LEJU2Lne6DLN7QcAHmpAJz+EtQYKx
OaBG+HvSDwh+BZMkEHlloCn7Yu6ZOC2W4h8oSCbRC5dlFys971Jc6zZHm86wyFWD
xpf/u9dwf2jik1L5YIleXk7mChGiLzNQVsPie0DCjBJFdoddYegkInR+LSn+b/A2
yqVmG6/tJbk7TMp6wnZ6JrEKIkaBgx5wsnBKhNia3n/eydewV5/6Zx5VWaecKSac
VbFsbPEZj+bhUfoLdCa8O1ctu4iO/w4S7PbL2MICbqHHLl6NEux5/YZcn3rlXuo1
w7nJnKKR8/eMgJ6YCCDMV5XKxbS5zf1Gl5GoxodNUZ7U9HnpSU9D1XGdgw4CyqGY
85cegc5QZv3zygg1GvFLYqZsS43Fu7/RlJaDjp8H/8JWFQfrbxqPI27G0ntM+TUV
PDdwobK5OIugiE3Sz/NzTFTx8PwwVtbIbGYrd6GZGUb5rcWtJQB1iLOGeZJbrbkq
LgL8u2lvikDdSyZ/i3jFvYqSM7zsMsH4aqbkcC2g/l3LExQzC53dawKnEvTA/jnF
vkXTwPyfhKhGf6/Gv8plDIRmAIXhBlioTzusOyj1LrYOilFRTehdj9S9fiOsV8IZ
Q45gqWq8K9eJMjtCly76/IG15pBVKVFsXathMQI4o54K6cY4Onn0Q7+i2Xjfoxen
cfMFLGbSnKyWUC8Elzi5VKDgMW1fzZp6rH3oF1Aziw+R/3PfcQ0pJf95JRvp8XMJ
svmIvAzt+L8RpMEtBgbPRKOIHLgAcJOcEXnpo/KMKhMKMiuqvysBBn1gYUKKljqh
CRpz10CS9zoSnse2F6yMhxl2LJlSxd2kJD/6pXX/GGfoQdfpHVX7o/rzW727fOMr
j+xTKc2paNTPKLcqk0GI8pOef1xpeU4eeWVJJOBq8tLlEZo2Q8MSyckrOVvhM1Fa
WJrlW7ChxxT1PUqU1QOiOEud0KyYo/76KWhf9DwTXE4GM7+pFWJOXPpcnBUzvgW6
v1YDfeHFnhSb9i7OalWW0eT8Ijrp3Ux9y+IMraImZ/DDZv1ST2682zuyKZ/hrOM3
U1T0c3lg2BI1zWTRr2rrJ1TeGG4yNvRAnJL5S5bPgdCcr8mwURFugnlqa4ahAOYK
8LotEmF1m+iOrM58hO2sBJFe9USkz09f6MgATNh2OLOzLrUJ+Vouaf4S0vBvgjwL
ODd1IF0CcJGZchQJbv5GwrTXbw4S+UFbmDLv4JxAmvxBlUyssW7NBVJ8t5kBnWlt
KrrOUqWl0Z40EUC92+DIJK31gCC1iCvdVAGEkY+oomMnaNlrglc1J9Uqf8RVVb+y
7lJxmDFpnKGRlo5LwVqBpLZmY21LGbYYPfwaBftDBiWLypAPnVJEEBctUaBdc3yo
33xEubqzcAj1Tpj1vQLZ6SLjZOzTx5ewRNa1EgkZ2iQFfjfZ91n7UZZIPs0ABlyo
7LUNXGlwjcJwM2VrUUR7Ab8Hy8cI9u4Y4hvlBeL0kbIe/XGoTIhYfSdXsvqghPcY
kec2Rckf9PccYxYYutDkV5rUqu7cvJJgrhCz8kpi1fbc//CIODYXtvIG53pWICWk
tOZ8rR9Zjf5egksvNjDMTHYL3nrPIotoU/HYBREDpoPgqES1IUhIMGK5GL72WZE2
fmDa+ByWl117x+Kd1ekoChVm1qLureO5WgJsk3FLu5b3/bFLKXDiXb/NE7qZt0Wh
4amNY7a7uJi5mtBUmaIcmlxZD0NZ3srDcIgUwIOyVDQDfSplF8hs/hpRhUqxKySj
LEpjSSn7o7smAhFueMfhGjkjk/VlOaYWuITcRHe2bl27faKFlc4zHYlvzXOo+bpZ
DV/O0AK7lkXEA7tvsNvBnMA1PZJ/WlvOEOthiAdZbSX9hlRTJr/rXVlD9v+7lqT7
7B3tU346ocrB+sGAS6N3Ds9sWS7tzIj31P4qooK/vecElYGcgxkW4ipkI+x6/PpD
k3SJBCowGdI3Ltvy3EOHPMJ/kcSTbDD1yfyMAlQFtp9rYLLCNbvrPwuXt7KSeWg/
TpDlueTuy5TzbmWvRTsrrMoDd8o6kdi76XKE7fnxCq1alcACxA7p1Rw0np3rIte2
q6xWsZ6dC55aatHUhhh/C1w6/KoRUBjxQ7MXBAQZ3lgFI8KWPE9MgXyyyvKtkom2
p3rAegL3c4ueV0Vb5rmDlHtHslHqhZ+S3QYkHZ1NyADHGiE/EdzdslE/hj8z4Aq6
Q2WEli/MJ9lgBVe1afjgQqGQZ6LmVwmMBj6Lyu1niDI+umJziYGpPkqmHNjViXHk
qw8y/+30tyjjmTSccETpJRYVZtm5Fh2Mniw0+dlzIvxyutkwIhQI2vgvt3amgU9n
hykSVJkDhnF1mwJDLct0hOJ091drlqXV5HlUl3AsNIUJ8oznawVvktF8DRcB46cg
FxqxzoFk4HtQ2lpJCOkP1KYnWyxMNmOKlJRWAm/aDabAvf53aMz2BiVp3xlufgTX
LspG4NgCIj9JnEndcw2d5BJbAZHotRGeGiaLYEotpzix6toOxyVtWhQB8s/fy1Yx
xuiCs+6xJHmZCdLVcTxg+kCPJI5CRXapR4dfyujfKRyAnpLw/Btsd1tUbqPVS97L
ZaMlf30H3ERyXQbEuXj+EWmlz9xRInxFneeOLuXavbuegfXh5/hkv2YCJnFSzv7x
yLm1JOQecVDFm0/PuZPx3ty+kSJcDm1Mp+Gh8in0d1yDE+atmqAwSU3Gnp9indF6
36QBQPYgmxDg18iRK0Ic40txkdiS0PVNvIHbXLzIsRXXOYZ/1r/rWgoSJBQPy+kQ
E0TNFMbyP2038cYhYg6yKE2utoeNR/ISWjHbrxwqtIkX5LEKC/oymfngRb0mRXaB
Rkw2T9bSxkGANgl65W08EFPgI/1K4I0xUgrhpXCbdeb+0MrcoZkCBQjhEXQD7B/k
MRWX3a93XJxO2lGTvECWP38obLoVclgDKq1Hxp/bIB7DvZgjHP95vLat6XlKteun
7YQGxHeTyZ6ZTdIUNwZ19OAppv7sOkKh5fNCkqCmyfBRNkP96en7J20i0PLMkmQ9
WGwXBO3eUQWDDqWLMYMl4JavZXb9AQW0oSu+azJEO6+QhjicZupDPa8gwMY+1VJk
BHtKwl/uPFx5qM16flX6rtff8QGMk8FYeU3beLIYfwUzPbUy9AZ5DLIQbhKt/RAq
coqv9kD8ek8MHqPZS6sCg5ECBereLhGW3X4jYpEBwgNqIvvyQzOwRgb52dTTnsai
ebBl1E5nSAZ3ypP3Uj7Itu6gGKR5i2qMFhXuwFrbYTrMHI6il/4u6aqdBuYVHHdU
MCoZ1BPUkcyihZWxEMVUVu68xA4b9vqHqpnMieuUGDIDMkGVKw0AUOPWoOFWimsX
OB2JI73MocLzcpJ146af6seYKFiVqKQDEF1aP9LsEiT9uFBOoy+TgSydsLrWIqsu
vy/b/qj/ZS9xO9ohyLUUJCl2ZspLhrl0gXG7JmrwT59nc2E+8AyTubsShkx6SPvP
os6n0eLEhspBAHciQ2+LOO89w+PWy5Rp8GUqgEdOKd5GsqpIBiFNkQeVHIvabFNW
FLE3+d1mBYspWcpOM92RwNOOmmPInk2mYGKHTc/c1T2LqDkFtynbRzek/B5CNnSv
BfG6T8OWcYxrTEwyQga77gsC+5dP7Cbw9qbP+GkIX27zunjmesRM4uwGs7e6Ea16
PpSrFeGUTXBSNBzUaZMnearmICvHGcAohetuq31PguC+xKUivVMXHwt3+sv5gq7M
KLrKLILu8rBEJ3G4K66AIwxZVSLjSRceul/bUdksvX+eApXYtQxs0Co1m7OS+WUD
E5xqlVk5E171v78pXL/PZLYgYBsCGnpQ4krT/2RRaYR8JOABSTk9IvxKHOevJYun
ODnoprLRT4osAx9jI7Mjm5x7+7aueJN5VJC0XRYCUXfSxD0s5p9oOD1rGmekP+VL
nyD0YlUD/MKnRlLJcMMf0N6CAnkf0knf5SJjHb/gmw2NrpXyBmBB6dYFzWxwjfxF
jNaAb0BZfb1SX86SzmDhPbib0Makbq9y/q8cqkbGKwozyD3maOuTirgXeguCLdLZ
F9fdNLg60B9ZJCZrbvWmalkHwH6CtnxmDABcNJOF8GhMAWYXDThJEEzcvlzU5o8l
wYm0khLhUAAlzbKwirBT5Is0eqWVLhZ1BKOzmgwOW+JekCY9f4hCJJyN6LBmzg+s
OI4XrfXE+Y6TDC32go9SknIz5c34Kdd8iVjMQrIRGIlNodhBVuUMTNh5s7kLsgq8
Vopy5N2Bd4mWTJyeYjUqn3l8XzCHCP1w6yGNljZFvpupXUBShHgEsMtvL7N0XNEU
m2H+LMbnSaHF+HuEbanHAHNQFgfe3dt5j7hWfJRnUrihNu3XUTlzxGPcFZXmp0qs
wgoHUMFYJ3t6ZaIWFQ1UzvP7hjWf64kBwSxVHZ15Pal7v2JrGwa4aTGuxlgA5PUA
ycRk1pPEtA5eCCX1x5TdQ5tbHEHnfRrMJaw0U1h60I9pz5tkrLLnlveTYr7ZqUv+
y8YKtN/LiIGh1if2pECokhIq16NC8C0adv0O96myw3iizmRoA2YTROmO2HGdPkiy
Szt3Tfs9lT9i94zUBBIDUMeiK+pDr8zIsVVNKrl147+6JCky2UiRhSOk+MXIlDuJ
maeygXcBdAx5vjx3Z0hxg9+wU2FKkOVwA0GBQajLlPbfQt2gTbDsB6V+XkPpejni
H52LxYuT9RCU2YZdDrGq3TikRlYpZWB1Jl8TU9R+nbHAerom1gkcEhw7CpqUPpRB
R/EN3YsY3yxXB4FS+NpS6K67Orbsb4TtOrP5TN3UOwubKnBITw49+L269gT8lXYj
kutLT2PWGKzZWi6yJmseWRPaotKDtFVoviv4Z+VxcwS4E3pG2JwBmm9JB84n2mnR
CuE7c5jswr6Rm9k1THVOQ7zbHQ9YaG4IzF+hB4vwirsebg4iYatu9t+TAkzlxAg4
ueNT94DwZdN+KUAG/msgB2ZKenCeoVYCOhE6pHHBakBGKr4FtXsGEHBqlVXOyp61
PexO5tvF3RCka4I5W5CfyrDMh2XgDRHjrQTvBmSTZx4G886dK2qcSD3D0sb/vNvB
WGd/EK4WXIxx6szUnyKnrOGj8Q4+tgN+IYf81ATPDEIC0G5PKh/n/cb3WAPwcWAL
nZf3mzfbCjDhdBxadIW/NHGlODgyrUouvfT4IMkD6Zll1LDBI0SoQIVGLs907Ntb
jFlafuAYHDlj1rXb/je/ujV88iPb4pDVvbQeqJmnM6uNJ2+mVSoI0lfr/UwB7+l9
C10/oBmgHzKI9DvRm9NJ94LmIDu1fW5svZp+EYNVNxaSdPjYepwvg3vo2jwisyyF
DT0yGnA0OyRV3uNfEqW2EdGBNvDDNmTf7P+g0PCEcrmfAd5lm2EcGtFmBQajHG68
5wL5HTzvDX8iOeM/9e3VrRdzWE7RJ5hpC6hX3P6bOY2aCBljY3y5RXjh58nbuRbW
V/iic25hUKVsO1/o/y5VcY0SOVSjB9DI5Oxt0hM0+RYMZB8KerFTtABINkJfeTV1
gkJl3MkcDtSpbt2xUpqk8yhJtaKy1i2xtXKq8ne/iD7V3RHBZE4pbpf3Y58DcYD2
BUPqlfXjeF7DuxgmNsqbuqXO6cwiRApqxrfw6YAUAYs7FSA9guTXi5r25kF1skWy
lQwng0NlORkYCij+x/H4H5zdd+/TlCEdkMm3nvRD+YjR+rRyjBIkcg9+zCgkeA8u
EQtp09svU+cE7LypckRZSTJOtZ9mmd9QETRfTMxjSCuI1MVNTwBMpo2iyQ9ctDcJ
vNvrANm+jSmySUPoJ/x1VsBSTYwUDFW+FQ9ApdRcx5eRrPOPK3hhqX805YlHRhML
V8mLLAozdF2t2h27JyTtP+S/2onzTWu3JPkrPyTwzbAZXV6kcVYiINo1wiUzYPx7
mD++hDIhYaFIL/H3NbNXJ0WhHUUAHhGmN5hp7rTINIno73t2MSkreAwzOlMznSVa
cLEktODCpP44RxyX8sJhcNX9VWn/GhQlL87jUiJMNMeUYmWba/lkUXIRgCL21Lzn
Ej2nLJlodZEhpxTq3dOp1kyE0o3+am6W9LBMfutcVReXmOOAUoBb175TxaaW1JO6
TNdZ3jTrLMyetkOl2qK56k+krrEPbDcn/p+lUS+GX81jlnlt4AlW66FhJ8ilCTnf
g626uGZZZO3JQn2j9gK4+c8Ihqo8VGrdP9q17JkoUhvNtwtDlUaHcYSM+KDGb8zl
ynXYWrM3V7T1JpT/sXGU+TENn1Xs4s34pNB152l/LZv1Z6kKmgWwULyo6s3neaJi
tAzkHli649p63hFsu4yUu7qYwXvcoxa5eL/hAW1IoITkdEM/6QEKwhq9wn04HVUC
QufO6ltBCu69+nlKS8rJHO1cFzamRPMw0yOYTmtxv5cX2+AC4Muqc1hqnkULJEkh
1C9QrJyxvVhJYGZpmc16nGxJ+iPALxH/aehUWwOhW17OjEKN5gLsMVG63vLVcW8v
AZaaJhToA4EP1emkRqQ6ufP9VLRirxGsrpSODmC/C9y5YssUiEJgt43QWx9rjQGx
isOb5S4RMWe7vvRGQN/5JklZwhIdTCfAEokFFg8kyb8Zfu/LhVtZ55LdvNk1O1O4
ou54+FO35ajVIwmZvf4bc9FldAdkL7BUvzVpUpolJ+8NPr1JF5JauuXnxnLN/psM
0pfV68C3m8vcuh3FOgMuFJQbN/n+jyNMkm64feYDJIIxrfa0/7xbKzOV5+V+7b/N
qZBg+cpLb+Iuy2GErhaj4JxEuLf/VgkhLfzMylY9GwnZNa69pJfzhsoCSLGzMHKr
BjaexAEprGlSo42EXfEJrjgSEFfv1HAFPQDkZ7cciOgh6894//9uU4faccJM21XJ
F9jQalDt6QXvgbEBLdEwHz5pA1ebnoBT5bRBUZt4O2K4Tp5cohbV3OWQ8fRr3eCp
hM+G8eS2OKYE9Ln1U6jyql0C+WwD/ed4EgqQGy+CATT0Z8jK+MMsWCnSJBpz13uY
jpDellw4NIEr2fgQZ/NIReO/jLis6/OXrlLD/LyF7hBa4LUx3FGixzXP+11lpRE+
gIWziSCzRJwE0nVvxSygbewMN6TcqFDPKvpKl7fHtszIP9QW9jtYpuvmnFz+nrFA
4WarLCasxovDPNxmvYzeWC/CCdak+vu/oEON2zDilAtphBVT9Tnmdg4FgkkTRKWW
SmcEftjlTL+t0hGM1Vw0WuWpTFrT8YajnZp2TO/hdgDflp3udnav9Kp6c9qU6Vmk
a2wiqJ4N/ZePtnPy3sLE6CsESPzPgcAFIW4vVybXish8fkPXFBgmn2wzxnH50H1j
iV7CcAv6G6+f7V9xMwZWDkOEXVw5GIdHbMJIEDEUYZTGE5N1MwmzHy3DpVFfXDpS
7hkJnkQ8j5Xtv32RYTNx3iC5s6ZYpJrckfR+ueMK2JrZsLvSE+hJd+VGp+HHCOQ1
kWwwurqnyrVB0auINX2ng6HpIJivm9wOqQW6UGZeMUqI45/NmUekVfpwQxCXUPQa
20yU/8kcWXGD58+4Cnlx8WrFxFIsQezC2m9CwtuU5K3KdNNOn/bDpa+DvGUsq9g6
1eBUnE2uALrMytpLU4dyeKFlIznJo+Bk2LwoP3e+zRtMTsig/5SIPYtPX64b3yrX
dIu9TcQBNY70WAyy4OgHsr7ddnFxEpBaJC/7QfgLbI8aXqOaeZGy5DV8b0BNHacQ
a/PRwwMp8jHbH+D1bd8cFa1PzCycQrLZE+9zyX0HtZArcWjpHDCPAHh7u8xo5bwj
NDgTcXocZlMAjqx1eQW3IofyOIsNHHq7f/UspN+LGVD/LpW8ZQpZ6OKEnBwj2tix
JB8ZuugYFvfeAizWYeDH2KtME+8e71u8I4ZHmuvkqxtQrRBjBnH4NLB0K7sGMMyD
f4Iz8Uweef4jKHB8dcKcFi0IlBrfIYhYKJ4gP3uKihWJ49CZbg+BuqHO4EzW8JMO
99l5mm5OZyr1NqYaaQXRmlcN7shfgI02jte0qnyEkNCn6/sq8Pl3rGZUcCSLnyP4
aDhcjAw7KsOWoX1X/LlDSPIznCzrzn1HYNRtHpmP5A2AWaTPoP6vFw+POrCruAg9
aqNDjUjKFckMqw59LDKY2QFgeFcrcIw14pgDWNHXzf58boVT5cqmQrbjfl4CFsuz
hxhWwlfAY9YpWlD4AnC4rsYm969g9gnEnqAoYXXFnPbTIu7jcQLzGCxk+7TPfZ49
/xR326bJIRI7k1eRtE1VanPUCxSYp39eBbMEzHBN1A0InGg9k3Ebp1dizholqcV3
RSxGIbGsKZEcmx2C8jcP174yPm3CkJdtv3rHaYRwa887RHHoW8MtUpH/0hIhXuue
aXao9ADA3A+7ouLicu04/CH4P/Wx6uRGWizlzn24P1Iaema/ExX7uLn7+n+4aZpS
CRHo6IvtlMbOvoMr24fHMzDePik2JEJfhFsRU7+lvEXfZ87Av1mR7v53tN1y+vQL
W6wD5+v8NU635l/1E7bzim5lW3HUOT6Orpp/EtcFsx2NXYlJ4gSKA9So1IXYmun/
UD5C/Nf5bdv5VNcbkE9Gu0Pv/cCe91413pZWcl2sAjC3Xa/Bsew3TZ+bmDv1rwTr
rZYAyZvycJqZwZ3F8zuBxE/4u12g9BKRq6cBgLbuHBE0/x7TK4tCb8xLqBxZq6FA
GvSBWUn3FFrnkRESxTCRheUNw9qox3tWXSsbIzENW4lBGo/hDC9lkHAoCak3CP8P
DYbBjFMxBpP04XI+HWpIjYcNoXXYvOveD4QUgeM+9LjyQweTgejNM8m1iSIMRPrH
MbST8icCYpu+lS21b0Pv1keNpnjuBsPR+vpZhNYbPPjJYCrolQHIo/f2whv6ZzM0
E69iWRhYLtd8hurdRdQm4q/2CWLRxXbuPmco5Bdigl4d1XWz7a6fdDXnDXHlt8vz
QrulJckml185fqCmsM5DmPdsNDO12MxxVGasz9w8kHYMPYGCv+OiKJPBiJ3/7PFA
7ehA8XPssBD30/XJ8yQkzdQHKbUfU6doX1Awti/i53N9l/KjyTN5cnRZyStQ0AAl
pQu4vleHjwsbwcRXl4cHM5b0cM6i2SWj4qPUNgYfVyJlJmHE88uQyCUbV/anAirg
DCyVvy+25A0AFkLUQkSpNMSDXIwvFNmT+Ub4lqcsBuXHPM9e3nu/LU/ZcFZ5MR6l
QMUZlxvtp1KZUDK29kuXfOoLMyCKWcumzyn3CxwhyHeDXW2Vshj18z9fSbPahL8M
K7B64ZGpJLdvjJebpPJYbDowVb87ZeFEATTKcWauDBD6rotYbMzKaLJB/rPhvma4
T1AY34FnIH+Nu/+/5NRuYX9dTLs1gDL5BPCoc0C38XM9/+blrghsGoTckUpM8Qf3
b4yZKPlXFIk73hM8nlkwatv+h/sJe3i6OAfNVSlstbOgdEAEuZB72P+UgPfElToY
Og9i2UhTUt9JB1BGZFiA9LC4HHvZHY8vJZA+l62KY/QN5a0eKcv/NYPml28G30RB
f6GMGHEtOGbYJQy0S6nAnTIz5T5zZN+ETRWR0RW5bJmR5/PVWtPbSkTiArnAwjfl
A2pSJAR4rUxPTXUQ47BhuVu3M080LeYO0XerpaEnRhqq5uLuaWxGirWerWTWTxqM
dTGnrjKGd5SONplUYFjXy3LbM3OvPDKaLVE+7WldWtEYfAnXMS0O7NT4CjR7KF+h
6kcrzdNnP2W0m1oLY+I0V1ejU8c2r04nZPkHOtrgTUmHLHkmHXdhEtcWKQnFuB3S
h18w7kkdgRMy2tngnExKq5ubZc6taTDpqEofOHkKLT87EXnOrJ8uwqub4I0FTHfX
Ev/X2aKywAsfGOCOTd8EfKdzyxDQjAVzzqJlojljGxy4Pms1rghBh4+rbCajgI6V
Vz5R8fuOt4WYmZmYEGInDz4IhcAJz2W9GY052fK1ea80aaaMK1ttkEqcPrd5Mjky
5ygS6GVa4sVlE8I0tjpruKUk0COQ0tAjBaENFjNmhZDzO+UYfSVeKD1S+Gm+BSQH
iOB63DarxAHSZoNIsMkfyKVvXa4mRKp+ECLfGwjB2itl7AJmFqQVhvKBA8ZnF0Xo
eLzlZ81jqWbaGP5ysWyyQAaSQiBUEOKXu5INlUHT5LfBIutww9bWb7TbhAmekLQb
PUo82IjsPLtvifnLQTNiGUbv8DEBQtIqipVAeouPDQazQ3KzPiIwlOYCXgTv/1Lx
UIHpwf3NyNI2IG/PaPtXolBBtyIJSbtVXpEGMk91vM/9rA8ElzFvrs5ufX08JmjB
3MLcdQNXbwsjOp4RbCohjOIPH0v+tobSekwQmPrYNC3y2vBTQOAnAf7HXebvD4XZ
R9AGfxikpGVAuJ/84/6osWMy1loxy7nKXgHrfPUwea5j3R/KGgqBrIj+82Jh7jcG
/8XEovfZmcNHm0WDBmOVl5woEZyTXQ7LrxyuQR15fYpfPsMXZNJSeva19O/WgT5S
lBlLYfSNXz1gT/OkiU43KgE+4XMmL/CZ8gzCoKFyxiuE8Ymg6Rv/cFuipqkV+GMU
UtH/2dUZ7zALSqGVuL7gHDLIh6Mosuj7IcXftj1EHppDu1x9eC4W+ePBxGnQZht0
Uunb0mo2g+YHOf0/NHu9iHCwxzI8uJ4+3rEd3ouPiavoVbuX2zajOUtjt8iCzm4a
bePICuf9VUxPSHyVe4cblYdFHbEwpG/hT53MWT9QWmee9RNWPxhNYLrI5z15Hcjv
16btugoCux/vnfFsJl4+Y/R6PTH+UbAk+xM2Ql24Qn4UlxlIKh3bQvme8IEUJ++D
xjYsOCCe3QnCyGJro4dzLNrEKw3Mkg8Qh4ND8pa8H/uEkY4GLCKwWNEAOgHnhJP5
wFplatlGLYMULAIx8PMMWiq1a6l+3DFaOMTA8x1yn7maBdQmIFX1V600ApR7zUD2
PGKmtjYbzfxhw4BanbjTD6G7nCTgjzQYWGcQkCpF8ziJB8l4tdGTOma7X2mo8lj+
//1wMyY/9xX5rqAKG/fun/rUnlR7cJiKWkdLCd5pmV8aL7Jx/GWDnl5xVsxXnsez
/dcvsZp4MkDpah7aullT9qrYlV+p4/c4BCPmsNvgPJJtOKKP4ZeqXg2dw1uf0q52
/dkHCc1BRarwjAaPbQ3R9N30oK6X0xLXgaPj4wXBDJxvScWBoMxNv4Z6Yfby3HoI
YyT7ZhWrWoyZYV04m+v97dDa7UtfODgpxwfCoxalu3bFfot9KV6MNjBIu+UTwsat
iJPo9vs0KJgs14nhBkzTywHbr7e18CB2CUAWxa6jDu9TDS9z6I2MdXQEbWiIJEwE
qCQ5799HyNhCPBHPqC+3Ui7bKnoUxTnH87cmI4mAu/+RAh/ucxZjwZQZunQZfjNo
zq4/sniEP4u13Jwz/WtoMf/kdDVMw7e52lZHIGS52Jr31u+8/mDe25oiCcPR1xGr
N/t+QLaMi+AjJUCIm/oi9dZcwJ8uXkeZOgj8hbliSRgzfIF1YsEY7JKj2u9IcDHh
Kx+LE5gfhbSGgdtiz2pKu1Tq7qQZtrJ+6KiewL5keeOG/W9R7m5EjFFBivcTU+9Q
0/fqioaekT4F5CgW4Y3RrjHF368YUS11zLR+gPUMLQ/ooN2IE1heSVlYPRF2++Xf
FQdImAu4oJ78i46DALjizZOzzANHQ7sk+ZA6dlndTIxdI3/YHeqtuGlGQT577SGd
nvc5BdCoRj5DZh6fjckMBOS0zhNSmun7m7rv5OXvwfSvDEsEhHYWYLFbgLeLiKfB
XJ+fsyQ2Up9DJDTpu++FjiamDt3C2B2JB//xrmB+HSAdmfMbPbR9NytQmDlBd5d/
lHyTnJ5i1LqyBLUBsBj4fGpLXwGf/ZHmNkbxdZAtaxzsOVlij+9BoaZUs85cl51V
hKa0UHJOa/2oigF0cBSi02mcxbs3Ro3SPBbe7Wg9CebdL6In9M3Z4diD8wtta79I
xr5aU3SR6gkPlqSDDFBp8onqkfv0kXSYdAGt2xpKna3a6Pthsw38KNq0Chqf7GAC
NKZQjXylN4rcXARG2ftZRuoWCCIfs71ezoXuPq7rzm+/3062MxxsgGkG+HXtqGj0
0zvRGz2qbYRDR3OQHQ0rIO3s/CLA3fR7OpC3l1DTDfMIeJn7/2+X71+4KpwOYGBi
hjnITsYwKO3XRewe1LBphdq8nfY+EFZC4zEY+mu+CFgczO33kUqbjoVFZB0xNUf3
paYo9FkAoADhMmbeW2/UHK8Xs6cZ9Oorb6ZUsXocHgglA/qGMAf9pXYnQ+7ZYX9P
LP7BGLqRuPJpc40NA3u92mF2yDJhIl2Kbc2OtAeKlLHnxdSfG0IxBzVDfjHBIuxZ
gcVjzqRssuKAiXZNpx/rTcJUYaOTlnj1C1R7S5niehBUkEms4w+gjNr0n/ZxyCiR
c789ELGemRDFzZUzp3QNDIAC1Yl3UVKeutEvqosSuiyMeE8R4NwP/AAvQCncfzDu
gvAPjyB8k165P2Q9A5+bBhp7jumyEqwcyaJs/HzLvTUzmsOuD91LkLZ/QSZBD8P2
fIfWnKcAp+U38E6B4GZ2IHVC9N3VZcr29qfs3HUKuppuNxpL4RcDiA0JLxiR+J17
CVhr2bD01zl+KaSWIajCnsby+Jqzd4M+0XORI95ur1fqPn/bV4hOeSndYSJYutmh
bEJoW0MnZcv3moUZGpNm/i/D3jRyYzlr/hNQhdqsFl9PZZlng5wCEKqs+EaHLZFw
xMl1r+KC4SjuhtbN6LZpxbMfFOYll10hyBny0Zbxk1RURbWCYxNDV2ySBcbttPWQ
RIEYX4um2B8loladm4s6O0J3XOa2MjCrkfJ1GKUMcGCcWQjoaRvBQYXKuZkqruKp
erYfOHUGLnMvzm/sZblRQmroIKR6/8jaMrF+kxuxaAvgXxpS08z786RHDS2GlViA
fM6E1JuEH3PryHL7xUywIm05bhc49v5gwgNo4nN9sDyTJ2NBpFTKlTlX3VwSE0hg
26nuz4h/wkLbP8pC8VMF97oKxf6AMAKwrRDFOYEGyutv+/b1kEhVXtQaHrxPGMAL
Sv3yVkM2z3NAr+YGnBfDxs9Rt85btVeWQoJIokOUtmdNEvuFKsZlncqTyEYGLLoM
bktF9k38/TvkDEzZtMr8/AbrWFSE+wWLGuTLeplZDvqvV3sdFsVJu2oOVtUx6dtR
pUGB136ojLnzlUGQbhXSuo/LAJIAGlscILWXsc1mBq53oRNwfBwoBqAN+wXImvOZ
rGSK2f3FSxK/EclLMqN1wtdC9LQxO04Sgbil1NzRP0LZWqYXsEVQfAlHNSAFwZpG
qyJ2NhaUBQk/3Dp53CkhXa4PTanV6jDYK1evRzfcyVloOitKU5JeS5sTIENmpPZY
rvbikxZX49LRbwDY0LgZQbqAyNj8SIfX1PL3c53WoHQ4/70UO98oLsbbKQ9+xysH
/kla2hvCrNU4I2YPmJEL/SFwEmum4Zd26JswxknX3HJ3XgAg+B3Vhrj8CRGOXSw1
6B7ZeLCHC2NNgPzIeQgaYeeqoy/9YDcZki3cym59oU1pypds4HhF1Df//VaozaKO
ZEW1QPJOmsdMuloxGSzIVy+LEXQ4f1ZMRcjtr22izZa8bLpMR6ljQWMHR9B9EZRQ
HOcDLH1pBedXDSucx/sccxRK5U7rNWYcd+JahInQgJBuQJWc2IpmIWA+S4qveb1u
REtPlcyqBB2Rc5M8X3y6Fj3DIHkbw9yd9uc9ZK8/yyp0ECNckFw9miIEhY5B4lJu
WTYiinIoYammV1jTnlmT0kHqkFDbm8N6gp7+Bs8NHSaFkEVDlq8WBliLfeVWO0tm
wrqLYDyOhGayHGj5RffTpJJ9Ijrz4RpsEKfAlTOx9KtZSrj/Rl8kRHHIVj86+htG
nbrRcT5fQIuNf898ZviNbYdlLz7Npfq3PYnKgpWnx4a71Nwb9jrzCUjb1WT+MtOi
m7SxZ7VNwip3/biBfzVcIuZUQEQOEXeP1WnLs28nDZP3URTMyOt9sCyNDa74W45k
GNW4pd5xZf9aZtmtP2nSMImwyJN/5VBvW25djGYBo200IiIEfuOGZGIUZOlr+u9a
JBXRyXJqdxxi4cZCdpN+v0JGLaaDCrUCrMyDl5P7I4UFzuS6W+emD1gWqCcfhbuj
`protect END_PROTECTED