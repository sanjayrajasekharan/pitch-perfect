��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki=/�U���cJ�>C�P������,WDǨ.���kYԥ]�ˉ�#0kz��W<0�-���$@��3p����~�U�0gQ� a��a��T��8W���~Pƴ�$�k�L�����U˕�H��܊Ȗ�_�*\��Cf�|������M|;|�ݑ�'�f�&"B-��a6�R�Vz�B:��
��H"	㺇{(cX�{�C�Ք�1gv}�YB &wnw@��0Um&M�����ŬHN���������tb��rK�B�_V2�*`�O�F���M�ϻ��p��6�uE,�=z��Ⴐ����
����a��L�7�%g�F�9Վ77��J����21i���� z��߽�?ק����B�8}ęt4O�� p9|P�юl:y|�$��]���������|����<�G�����:��o��i���7�[=����z��A���Z��D����v�k%�$=��1׬��ӣ@�P�$J!��pk���$Jo��թ	Q��M�	���'�?�T�bJՆw\66Z�N����uD̊p0����|z������BxZV�r���旽�PԹ���\����D^�r�1 b��>�U�!d���{�����bT���<�
�Tp�Q�=�<p�ciEī�C�ⳅ�9�Df���O�����Å}pzl�8�P��+�Z� ��J�"|��(aݜ׀�P���.if���E���{�!Q��Cl�!�6N��H��/�P0��m�Js�T�̸�I���bf�!���UK�jR�&wN��E}���Kp
�9�g�?/�L���M�a���X�����L�㚠�"luP��'���� 蜶f� .'&F�l��;��=x�cƃ�����{D�O�#�|�?TIY/~["q�A�w:5}Ds�̰za �r�������d�14W*#j�r[]��9����
�	u��H�ss�hk25�z���� �o�"0��k�P�V�[=U��{o4~��@�'u�s	���e��dW m��dO�噀(F��Ɲ3s	nS�%X�
w�*̸�t�=~)�4�To�e[�	����Ǖ �ݵc&_��y1�Z�E	�{AR��p�o֞�ir���y�d�8��
�&��T����K*l�eE�1{�����<,o!Ͽ������="�,_cirl��-��{�����Y�������I�Acg3^c�� v�����'����1i�a��Y��Mg/����������ۦ�?�����U(��U����Gۄ�k��1����i�k�֦���e������d!=x� �nj*�J�Z��=���3��uu��S	6aɅ�D�=5���x�Kj�|��5L�-J��-�������RÖ�=�~� ��2¢_�f�>X�U���QW��I�Tws仵M�1e�u�V�cb?�&r�����c�z�ЈJ��oH�/�SE�x�C|��:k�Q����5�L�;���A�J��Z��Ԡ'Q�2�M�!��,aM�L�x�1�t���"��Q
��}Y��j��Pʤ%o���D-����>-��sU FԪn�(��@J��^��� <k�<`��@��/�3A�B���"��g�h�%"� C:��C,�����6$���#N:䧫����R��)gJ_����7�2�8��$������/�t����esp�'��f�� �S}[(���Iر��ǲ���6g�,/�G�^�Qk�x�����1.)�2_,��OdZ�Wv���\����������}�i1J;��݄���M/$u��m�!��7�T#1kY�r��ɬ��,n���B����u��=ټ.�mЖU��?�g<XN�P�y.�_22B�����؆�%��I%����T�R
�|����oa���Y������Ap
!udF���q<*�c>#%?@�և����P>�r�z)":���F�q���;B�i���K'�Y+�h��<EI2 t�#P���mc�הLJ�W�ʿ:�dl���΂��`�|���Ii�֕��}_�/���(@+�����w�V�����Ԕ+Et��U�?�gI���_�P�5�w\͞Y���@�A������=���xE��w�v˾�#c���M'7?�3A%ƽ�s�)@b˹�������+�,�����<��jRNP��.�m��3�>V��ڻ�R� ��x��kb��0	���������'Ұ�-首�k+�4���?K�3n�d)4��W��߯��&=Y��cq(]��c�a�s�E�����޾�.��@M���I�vv�i�h)���E_�1���B�E�k<!?3q��o��!3�ᘳRcErx$��\u�3VB����}n.7���A������W�C����*"�?{04�qI�b�v�A[8�cO^��I,�|�,Y:���`+n���Q�h��7�t�-]2
�����3����&%��a���Bm�q�"X���*`�~��d�jo٤��S�B�7���2s�P[�[۟�#{s��)P=gs'�1���PC��zGmGI
��6b�yZ�݃:J�SZTx~Lj��v�@v��Ԓ�EA�<������^��ɯ0�R���b�Vz�;��!���FM����}M��6�Ն���*�)�y �D`R��Q�g����Z�J�b_:�{�O��v�񢂤e�Ia�ZD����,��.�����&�<��8�`����XEiD����U$�"����
�n����D6�'�����8�P���H�������A�m�t��*�aߵN
�҈�c�h�@1�߁�&��>n�'�H�M܊� �}H~���qP�~�G�Bȣ�����;�܇���.�`:�ʤ]
)<G[d_���E,��86��ڰ<�	$�sG�?���`C(=f�����������<��ϪU���r���uo��Zèû�0��J}�^�����	zV�L��A���Z�YpP�f5��}+�j�u���I��v!�@�]�:yI�.���7���,�?����7?���,�$dD@�ۢX��ׯwd�|�&Fʓ��!q�g�5�v�)��ۆ�o��.l�x0� �{=�	���@e�l�w�ܻ$vm��J�}uu����f3��H���.:���iQ';���o(}�@R=�rV��
���̜C�>�#�#�uV��ق�B�����NRɜ����ײ�ep7H0�M�)Z�݃���
R���J���GS������#��RzJ.w*%�MSq�eg-�\awEw �	,L;p���g/�cZ��hm�}�Aj8�`��$yY�m�s�N�Y�J,/�}���HR����1A�f�A�m85K�Ci��GϷ1���ن�iDt���W�����3~�� 1�5�z|FK�JH?