-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
WwUA30TrBNaEDGDbV6pxpOWWUnwoWAI/Q/lg+xSpHyW4QxLVEts/7yI0yGOF0Ffi
RBXQmduL6bAqKigLAImRh+9toEx1VN7n4xJ9smAb85fnJDDFMYuEnOqmJx8vF5CA
WzKb66YFuckOqbzqHC5MIcxlnN1Km22E/kkPnzQ5N7A=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13034)

`protect DATA_BLOCK
VTjy+as3XybWekmbf5ZR3cJ+nc/kL9z6RYtqF9p56k1lH/ZYVKzHfMtkLBr/RQuR
NQHtKmDFZ4CsQkJ2/CZ44aQ1NuYnRv+Ix3GejgUuOQ6Up59PP4p1rmnnQLuyrSpi
LuQhrXXemsZbBshr/CqlVGt7BWYrnojiwSIOMoiJZ9TVu1KqP5dfmxlYtz3Utu4S
k2c9yCxLgVBCgvUdG45I1f+paMfK/pj+rOL+ndUG7LC99YtvajQMrIkJNhcLaelx
OwS/8HP1pCWx91CFqtrJDjTBC/YSDaRtRpMM92oq7UohC28LWXmSCHr2hFxscYfm
h+ApnoGh+/f2xqGvRLaeAhDxupi42xVYrUgNnD6d7YrcNB6K7F5XMbUN6YIBbyD7
QMVwZlMkMqJR3nZ7ilB2Rnnsk7d85xmz9LTzgPfxhp1W7bLNLOtCLjgl1+F9Ohh0
QF5Hoq/OSGU3EgBDG6okq/qH5FBaYYEY7Bw+jpsfiC0lGxOaobvGoa4ea5PzEqfx
Tj8iEtYdL7jRpmmipKNetKnsaVx1j16jm+ySWmnRxS677Qgk5M4FhXq14lKG7Jhe
SKtiV3RNV8uPEsGvLnx2p69gnCIrvn6nam+ASXIQHlI86pU5x55YT7ooXjc/iYtj
9uwaaJKwF6uVoxuociF29sNXbLi+e5dkMC5cJC5QAqPuel1K1K4ksYDTbCv+YfbA
FWbwL4GSpXR76h4yzySlwPskD651rpP5xVyQkWAlrAODDfFLTwb8Zbkf3lhh9TUR
gA3c43N1dw3IR6juXLngmbdO+w6MPAEMZcB6bPDo9YGDxQzvLgk2wauq30xivsx0
PKUhmROTAQzCLOewcYeMr+4TAR5IfX0hNvFmrtQ058x0PDJEsPoWvhkHdViPD/H5
ejIb5rkgKpAZAOJjfSeNgaUdLP1DtONdRroqb41du7CBIHsyn/o/lPQjzVI1I/nd
XNzGxhP/kMlBGalc4CMeID6v+apeCgTo+9hYRJ9t2MCBMb/yq/bR2ba4A5yl7sIe
HYT3yBnG1gFe+V7FrmPkxfADXQotKqWil32pmi6+ifERPd9JrnF4UieDB/5hJcFj
4jdmxgtRMdaPQNUQKJuwSCvMqdnSTEtISz+P/ytFnaPIe86PdQYxlYWXylsJgsQv
3j8c6+bY+3RWOajL/JaUT/4+fd7aeqBOa/OFvjL4uirgVN1DkDcvJ+wm19lu80ML
qpAN5r4Z3ktA8+zhMAWh6Pk+gK3yCRoTxvAnx7fQAyMd31RKC/ggj+ktP5O0qQ8/
LhnCNoN4Madsw+Bhq4mu+vZ49gci6HhGQRS6MunyFIxde1W53t/0NH/sfcfIVlmx
tAyuYIx/btsgIc0/6gbXi82ip1/AXtMlRZfoYw1fSfULYAZlNFYBw4/uCyM4HJX+
CIMJ091e0AlecH89ugEngw5xHjZ7jycDl1bfEll9I6OVkWMyBPZ3y09S6EgC6Zug
EvbvR7yxE8JrJBKOPJ7rbPYAK5WqMzBgHmcl27lfF6gdGmZfwspEXYP2WAa7PX65
GZMH3P84j0ps4bxySw2w+cBTYXDSjlmsCUO2/OwJx7tJcaevocndtUtQkv52/6gU
mRK5V/UtTRCUGr+6MORWINIrBr69q7ZmDqNMmAYmMIOvTcfbEdLa2q5cQaDI6ywf
A1IK5ht4aWsstL1QGuZszhqIinOIxmI2fFgr6GSL2rPNm3yZijH1k4kcJp+jcLGg
AF8OSjRsKbcJbTAGeNiyOlKISl2qAQy5vnKV3ShQric6UMz/FwrcyPPaXTExj3ye
DmCEveHnjlMIwWhtzY86fuo1aU9oe08TQONtBu6Sol6IsQX4Dokwh+ahZfsIeMO5
YCT+M8ABqpUQv3e5N5RiO/QPCnyp+M90jRyO03CJPI6l83WqTIqpSy1mRW1gh3pM
q4UxucDH83yw23Tt5zUsv21qbKqRnywPLnK5khm2DyHZKNs0MvoehXmftO2UnUV7
jxETnMXJTtLhP8nkpOZWe2WsPvGUI1l1nuCcKwIwT9HT8PHgguS0J23Uijp4NLpd
O0C540M4ZmYz+lHiqleqfqJXhuYvVla2tKRgC+Uv/cgH/8w5c52lxiVwzOOTNEa6
MpTn8OZRE06v1UGJsmxWDeN9YQLpjkWRwu4xJBl1PHEAJ7StLrmvzQVlY5jLmapy
MtP+ZHYnv/VRJaRaJBwLCoI6Z/jxyQvRwfVAKb4pJIOwB2LmUQ58GZsp6c3f+rWv
Dz2h77DZQmA4/CM6n4JYw7RoGnQCjVAR8db1Bixiyl/Uj+RRyAvRXwAgh6+wLoRu
hjU83WXril/JMqAqFSZTk64PmgWRny0xkgHyQarm2Gm1kFr1I4QZzEHnN77RtOIH
Zs7g4Y0DwkLU34S1jBoPCoRvCA06iQomcpBjzBLhLo8ZTMGYixEBGn71dMXZuXw6
2ZnktRYzwgFnBv5WwB0Vu6v9zgLPqBIB8Ta8XU3BRdGoWCjaU4QySjHdQxy78USS
TgdtymgkHvknCV0zlAHRpZExiQV2/Zdhwxy4Ov1U9E6WJI03+fuoMV0bLNo7K0Wr
c5gDjVb/lLCWZTHA2sap8bU1QNM6fkFY5T8yEfLdj8Eh2X1EIEBA6ZRNDwEE5W0h
BGn8H2QtkhKsos+cirexC3/q8Kp1R0/BhHCoxxuHb1SBkzmVNIY30vi/IoBdEErc
HzI/T9UMRj9YW7Stuu1NbLc1FK+88VIf9Jmv4MPqKYkYg6J5bgWEN7i/t+nHMDfr
z6kw7VKLTzeSsQzHpmCwfOyP9SIJGE8xI6hZEQObA+JNGmkGuyzxKn4qpD0HB2P2
uODTJDXk+1MpYDy8bELr51DbbqT/kHOvu2qP1ongnEq7hUbmoKmWso6MgCVJY8X5
7g5ciCrNIQ1mA2O4TPi1e9gNH4BLslqwW7FfZRnK0670IcDWWzR9papVcrKUbPPh
9tpaU8gBLpDWk5F9ZfyvW9uY17/SP/hD67NieqUzupHToBVzttkNhFJg8pFylHMz
AhZrX4tmIOVkKPWK9EgRvATvx6YTsnjQw34lA5p5S3GDyszQvSYuO+aktkSZIrOc
JnT4uXqvY1RCwPvstOBDygq5B/P8EyeWSvmTFGkgwe1YETJPOTy1aiNZ5DumuQng
3Lk7T/JeKLRQcA3ey481Q+frzjWVApQBngMzPINFPK1jQVGpOKyjuGd2/2CmAap3
RJXDhqIv6ROsYLDzjC9xQ427Xz6iscYQHoUPhuxWaQ6g1EhztwcGmw6Q88t3/ZI6
XPxLwO8jTHNTb7he1TjqCk+DceDuV6my4far4XYjeNYv27a18NZxxCvLh3cxGBuP
Y2CDIDSb0nKFP5FBg2XSt0zK2AgdzZbDZaVM2BdDUsdlCrJO6HeCKx+E5wg/lEzF
cXxmzKV/PzGd1qX+ZJNu0v7OkSds5vIvlkcIkOjLXRw9h32Gqnljk0saSZBLVabv
bWyLfr9lNzzQ9HR6Cpa7kVKtwIBSHHpTdyKJSwUbWUXl5AHRlCQvyzcgUeRsDKam
GuLVf06q4dHBMDDTTABewjy3KTOHszQzKj4ALxNaFcMi4h9vkQES76OPNOkJ1BXu
E45acL1165Tnto2fbepfrVHLQUiM08qUR/j2h+/MLauzSM3888QDiYAxG7brdI2o
WImP/5Nh35Y6YKaEbXX7fRagYEwWYrv5wO9TJrSeROYL4BBjyQCEaKG3pAdpqKiX
CGcEkS0ULWv7uIyE+pcSjOih5teizxtCYNrnfUbA51Av1YMggEjXlz9J1uC7RraT
jNZqifp8LMXMTrtMgHlInuFKFeEPntNTyoIherRoMNqsBbZhhI2eOt9fZziEleuh
qoDgG2vANtwiyqk+9Ae9+hVgTf0TGC0R5fKC0SRt+74PYegiB2BFyDLBlOjqpWD3
TKpEb4c0ki9OSXrHjU+dXeqMnI5N2lgodmYM5toxDy33bz41LkjYgNvtLSW9jAL0
OFemfMXF8ZOy8cf3MFsYCGI7Tpnw02bQG+ylaeI5hOxztN07uNductbDywYTviIv
QiVhy4k8nj1ndx2rJDGjL+13s5MaASs/BGlUSyNpMbLVOz2jMNSA7opsVeg/q/EJ
kl8F2QCUx8PjADayr6CsTtY8R2u9EK74WCJeEL0kqGJz30wym1VGyiz++WxcTG71
1xtHEKEE/DsnzJceacX8W8zq44qwoM4w3lpdLFUSb00W4ieKO96QiEU+DqX5VFUG
r/G7ycHlCE5suUwbatrf3GihMy6VQKdphTNZEkIsi2hOKeTfym1RfiFfx19bdbC7
nGYiq7STIS62GczUMf17zQ7IhwXSh6H4WgKqNrVkoAV5NgG1NgFqERlDfIoGIjEp
KH63qx8sbO5fjxtKeb6pVjaqxkGlE068OTx6ZFX5Nj/xyFKX7rSf40Kng51BtzMT
tDCLjPrPOVNQj6Nc4bU4YZcTU5w6MZNCeMz6D3mSfDh6IcLU/T9/nmzR5zmdFrxF
wpowBd2b7iQxBZZed8HkkU2nt0E8I23l55ztYbKLyEiFOk6HALd/59uZLKvb8WXv
/nFf/7LYLwKM4lfQ/fPIYcgAh3xpkxUieSs6uAXbQeT1RLP5fKlWbrtt7+0A4+7l
Ba57KjKsWBFKjaIfcuVRevU06EYs87Kdr6ihsNlVNBG0sNioyd/8lEZ6G886hO5L
lz6Y1Nndb/JpUByqUMYxSB6YWkRl1wBjb9e5aIj3mjCTidCj9Tln4zOMgIIzMvcG
v+Z6tBR0/DPWdX+r+FYrXUcLL43zCc1f0X4j4OCUIkW5PUAu/KRfF+caSNW6aa7K
hJb3prWRcWsfR8lnBVpY2saOrjG3tCHo92k0Op5JesBrkgy8tAvGBEV7D3yCobfY
+DkdQfuEQ3b3E/rdIkVA8jLjGM4CKIsIqRoAcjVE2gL4eAG90UiGApT9VfkDcCJF
GWd/dAz88gkqMhZ+C0jmdmukgR8zbc/nAuX9HNlOEXEgEt/sggdSqyP0+IKnzN+f
5jDxOE6bVUO1RTRxsZJgpgYEMunIFCtYO4bXd2uo2ZpgKtRBUBXzLykKSXO3ymVn
7Jy6w1pn+ein15byEuJLZaHBs3TLEwVG7026IT720MO9mF79RfyFdvQM2z/+oPR1
1pA0KERNJrJfBrS1iNBBu2gdAy+ZwwrRG+mcJTBzyAAvXFc9VSI98vLQ0+43LSmF
iqVDPsYGiMPaWT7SC9g3VRKKnm7HZ8NS6rvzAxI7rwG9w+U+K8+oK2LkYFJWegvZ
UciddXNNS2afkNemX9th9NCUP5Nbs92XFZ2Y414bWyVkkM6pz+zWGOFiqpVtLTjZ
KAxuG/W3d0X2vDZOOVBy2hrUOU/fmSaNF8tH8vtQWH4xt8MZwN0DAo1/FVINqjbK
yBFwxr9uug8JiKcQ56GME6/jbqqcs37wUyRGMT5DeD97jS4Y6rAy9s03Tsg7n0l/
7kI7fW5bbRWmYLiDFKaVPMjQwQbH6eR/QvMJnHmZLGpvPlO0etTiO9jSzm4mhhSB
hlcnGBoC2KggcSfs0779AhISw/ElotiyTQZlE+YHzAT+xBXLET/gV6KO1ST9Ze9C
yLX008/HPTHCuWm+2L+aFvQuyrTPkFewaaLPTfg+ombGKCsAQz/XDWsv0cqcCOFr
n1AYc2OCIdaiHTfTzYlPbC/cknLW+GmeUS9j/H7WU9VfY6VGOelCFSYBdWTPYfK/
1FKqZYCWcSP8p0+lhbZoCgQvusZekJXFVSH1lM9oqIJ9GJf3Wy7I5m067QY+X8Cy
HbTFDDqlYc0nth36FmD2WjOWTd8Wa18xRbHOuDSDHF9sqOcRC58JcRfqNf/gx7vb
CN0nNoIUwAa+9zjWo4Cb5fXJJMM43Upw5USwDGGKY6s4wxeWknxTX2uo81CulyFO
ZGogh439A2ZOdyj6fuoOIOB/c9LRXhdacrr5J0Ie1kQ9MqoO1eyw6hM+3jaaYIWm
Cr1p4xsf7h+Qpx4dRmizvcZk37W3MDJHiQyFKpL+v8eCMtAQFKV2gxgkBOO/M4kh
Ub5sdqgUfJkIOjyoKoXyjX6uOIB5W6Ab/7k3WYfhJ6/eiL+pVICBHBoJUfa32EMO
vV3yACBs/tBRdUf1fpXXiGoQYNbzUJ9LyBOTA5G4t7Wd9ZTh9U/DHjHBtGvhj74P
IOWqWRQH1NsnHg2hLeLIUDQ+jj9jireOfDQJ9FrxSELiiMKKzLJAlXzCxTOHhG2N
H/nt/gAzdvvimulZWHQuZJSTJu1X6V4LU3orDdcnJIIEVTafRHR5ftCA6NLhZ4Ez
oGvsMcxRDKeDkAorsF8rLttQXe5FYFqxjpM3bjN5RNq5h9Jy48lPK5cQIFfw+/v9
Xolv/RJVaAimpjJOB6cm0GggkVy2BT5ph1B0w4YSOvgihTuJm+mmLMnJWP01bVFb
5RmVdxRmt/VRoMplPzK6uUfyZ9CejE0qZ66i4Slwcv6D5+bXkdJN55VIXepRdb2r
pq9A1onRo7ZsXA59eEWESJjKvpfCAuolWpXCrlVxRcjwQpkfqhXP+gj0s8UlffF2
t+bzVZHofwOE55V7AV0TgWDwlbcJR6uzz9krzcZ14XnBMhaM6TNw1mNZaR54qThU
LAnl3dDrWhWCq5aHuEphYl67Z9JiIcKT1j7BBVt58oUW4KQJG0h86mONIk6Q0sSu
X4PLBUFWznmYGwHAUrs//SOy7dV7ef/1l6xWnX641iWdcWli9F+gmmXeyr6/sjoh
m2T5BRHZOmaMOIRv3oIFxGHeBGdQm+I2WupS5YlthAEiB8ui3+22UF88EqIRQBHA
ifgGMxXQLx3RqSaaOGHNzcq3wIonrNyQ7w/2jr9cdBrOujA6sHNSAgUQ9gXaZqsH
SIQ189L1uSmOgheRbO3WOZ5/97ubFmRep+ZKlqYV5FGUm1sNm0th75Sjp/r4ajRy
M2TPxv8cgD5g1WRYpB84x6TQh94sDxVetu+Rg3LL8IxluRucddRPmfAE0HI+XjHF
7fksisWjTzCdgzMPI7KEh6KBp4XKPE6+4NDqts7+hBw4LKHLfdyvUYIYDn2m+T+E
mzvXMMrNhfWWMCPHYb3FdIUnKrwcK8fAGEhW7LIc8PPi7oJZcre0SXxewBygf3RQ
vjt0oiboFvsYvScb/dXmVnxfS3JYMEuFab3UfhkyurnbCD9o9QOutWoUmTmVGYdJ
YiUIu1KIPLlBHXTKd13A3aKg1J9D5cMa4Yrs9nnANB9wk+wgP9xRqtRIH8MhbxW+
YvRGRzDiR1zQ1IRU3jbT9j/GLryP9uXCviDZMZeapv3LcvawaksySspu3oek4n2U
6t9GHgEczmKHzcvG7RA8mbun5erCCbyTui2vgXxejW4Yoa5u0GLkU/nwPUOPdyQo
I6aWG1+E+u9meRnSlg0VbleDYBBr828YFmlPbwn3WPJoVEc0QnyN6ueEGQenQfQu
JS+mvwlcwqcXK9NIwgWwrmMLekwLURVEDubxFhomw6YbCI3gigTfTc/49DlBojrm
cInJwt154kAhZYwYA7+ePjIEHuH8MFjHn4/Z9iPlqxebC7rypWkN2YPQH9tpYRAh
xIsXW9/aBcR1hfEfUIyacLuP8jLaBvl+EvRmxBVtxY8NwAAM0n49tGLp8NmBvOq3
SU7dosQXMTOTxRwWNpZzaQ+RbJnhUmCYWhJSy4auz7wy6WK3snYLIHjlpeP9Q6DB
L7Fn9H6s2q9kzgZ/Ik/gEwBa4KFrBKAwtLpYKoxBEbMUu7Q2ZsLP/WWK4+LJC7zE
9rgR0pbXEzCZR2ydc6KtB8XHnqCx7lroGAZV1+MwBF6DZlqR03+LaF5EraBM7Eqc
fs6ytqRSFoMfSdwoBG37OKYodmJkYhn31pG+xm/jnOdJ8fzeeC401q/kPhwr5iQo
JsydANj93b45TMbaAjEX35ZO1qTcUgFdV5tiVToeYYIVsiJppZo0O0GxpQvhCy/1
UJYBp5xIY++sprioCYTgIy4A06YzSY9f8Gi6zcuCh2Xo3KkU5zEy+p8RH+kKz2EI
9sAdN4Fq6/5hq9+mMq1z5tQGjZaPku3QIcM0bPGGnWdvH+uMoi9ILbVY2AytWNhn
mgpByi4SDldYbQmIUFZo2ds+gNwRaG+1mvV1x9K71cFWwxeV0P4q9WRERdEh5Ho1
g9Y8o74+uROZ8yZGHU2ew+YySmwE8bkathFNPNTSVQ+1palKq9pDwJEiquVY6LYL
0thx7P9FbfzytW1Orss8yh+52I9xxDWDQvTIa+/eX/KUJ+wBZg06y3RctIDIIBQZ
iRGYZjIMN125HriebVE82oWxQFoBo0VaLU1XELqg/k+2vcSW3JE+yTHVBZZ29hy3
sOCiC+Z/Xa4dN9QxLgKrRfU7ReovPmEad1zzPoMvfB/m7dcZIUnlweM3S+8cIFf1
Gbqmj5ap7tIXOcSMHSC8C9E9/85Ku5uH03agbCpsvfa4RDrWEFFLk9Ua6Ue48Z38
un/tUuyds7mjIGKm3H0hK98eG6OlpIfFCZkIrcqSARmxKAJf1l5UGjiS9GUM/gd7
2DLL5fOCOcO/15v6jA0UKwX0ohQ0vrARCQi2ahPO1DUKaLmibH1eCYzxAf6K/XyX
GXeCx2IQVrNKzDKdf013geZEEn8ZWd8J2JO+4Wkbo772DGI7mlwvKucZE2D6avyC
txNWSpmjMmzS53sfy2g4MvRPtQMzullq/evpf7KDyYGFrOPZtuqB141t9aTGg+wT
v5J1UkCqrjfJSn5K01uHy+bKV5eWemq4ckmkxQF6V8bzui1FPHtQkb+n5sLtiibh
9Y0ai1L9HhHUgFjhmpqZNxhajYRNFyQwt9GeW6MJaa7UDPC+xEoqQGEsS4UfZ/WT
J38JQ1YohaWutGH8M6ao0NuZxUabo8LKxJWX6KDVwJehV6N6yDALzZ7Ahk4tEdA+
HXBfT23LBL21gmsoy07PDPK0sIJu+lYLAVH9NToW9ZTqtHgqYsxdStogaBOqlP9E
/x4BptW/zgld2I5qaXKQv1nrar/RvgBrJGP9fjmqSe5wLkhpC43+ZRTB0A6GFKha
5KMuBfgq6CKk+PJ24GFfV3Quy2blcRYNeQBZr2RcZziPMjroMXs2daOKFUYI+mQd
Z6jSL92ub6gJdycv/8dJZQZZiJ9x6xswN7Sy0uDfa4LISlL2fIVG5z2fAedSuOFc
uO+HZ3dwE2vYMZp+nv17q67FVwfpdrd0CEWpkWzoJsL8Qdqxq2HA10o7SujYBfEP
QNSkoVik2TpUy5ffS2gWZeKkvXqxeJ/35hjy5iyoquDLR3hJzVnwYV/5UlC1mX4j
OySJuFtZvnT1AzU3C3efoVmzNf8nc8/mfOErG61/SO4M85Ki/28gqvKU22tcAUTo
/VzpWyNd0FCGj3WRZfJ2OadsOgENpvgvX495o1nhK/LpRrgs620TlXN0rANHKVgz
BZ0M3JMY0Miq90cie6HuLVI2dM8GyRescLHZkdrrCG/uBkcKE6ewUlOnrs3iwvRB
l8wTEtCy64JbrAdS2bMk7/GUqHV4Ys8usp9LwWXHzyBwhDotxWVa3ELvoNthwBti
bOj719HWm59z9eNqOWL2N9SrzVpyOHexpsTV/OriTdG7EhhyMDdKX+TDY4JgmuEr
BBEd6+baqTYe4Wiw57HZRZtrjXzHLVKj1ZCXv73Sct791ymSrfo4wc+HFcD3Y6gR
gRUD4tMPWW5OLlQiNxDaZK2VCWFWtl2JrZoppcRdk56CojQC7GIHEdI2bu87Aj4e
19aHzFOqOK0JU3QSGrXzs2grdrIu7poTjb7YHtOJB/Q1qT4yQ9zA3AqshP7D8LID
VzGr/KVVZv9PTNw+Q4F6ohANe4DBYyBHk+gUIrQXN7Ada8qzvi1hMeyLOlAv2Fic
m5U7xNkf7VRNzbWfwwCJbchDt8eAT/hDp6dsP9C9G0tfMUNX+DYlS8MMQG5PznHY
lQ6wPJ10aSTGT41PITPRhF0JW19FA05pFSAF0H8Tf9XodGgLSwhjiDARPZwCFau5
Lc7dt8smzm4Pm8fGKsKwBgOQ0aUV21MJSpc9hwM7PsxSwDDvyShuMqquflCqfb1M
poAdsRiHykKgeGZ5dSMxxk8B7/0QmKaabC3yK1SR8unruynLatwvMCZ4C+jFPvZt
H6Lwxl48HxUbeUVkpbIGpPQPz1lQxXFI1E7lBc6oRuyNw9YIcUu4g4ozMQCASa7/
6mHcNjorgHIDUbSWOvNJiofwWJTaWAgmGtLi/Ntvv9Es/A28LGM0S9UB1DaYrOCg
0JWkGgOXUs6N4lA/7bbwTmSxd/6HofmU0mwUK8Q2h3TZamSzXRsanPsCF9j0iK7b
uyscVka/9XCcA8HUdYq62CUJHjo4LDFYGBpSuk7cmTKx5fwCRE6zgCkMf4AKrZGs
FxKmA8XLK2kvTBCN2PuXgIVveLfk0wemtQKSL+jRzl3Ru3Uwlyi3tLtHZeakYKJT
NBpe60bkC4WqyCpz5xKOYUB/6fL8dBX3pK30Qf1T8vH6kRLFnmiaZ2SOtrHOAOL4
+vVrw+pmjvQvTQXOh8AMT3JuP6jnOB70G5NkAjUYTJQO0qzRX9tipjzNGeBCWtzb
fgia554eXdZt95etLKTD3zJnkS/tzzxCsM6hYn3Vafu+nvsAch67/WUIV9g5iwrk
mZLadCElMGX6Kl8TwRniBGKcmJIBbsb2yLqBsXVNWBvBmCHasdGkSxy7EOwENllm
Wqn2O6jmyWdqHgFNmx2X+trkrbjlD1mK1IgWmqPE0579F4wsNwqxzKww5vbYBd/b
hoyyI65RTJs2B8MBIi68XQ5/ItJDyU0pMPScdA9c5dSP+H3ANlm3a+JTZmVwnFOO
MSgdHeqATs6JtEYgyeI1b/I4jJA9ri1M/GTM3o1WXgDPVEIkaQILApa7pSJfdU04
SAJMjtJvQCwhx+tKse4W09kps3OOQBb8yMcNsRIqZDfOBPPHKjmn9DZuluZLAtnR
WvVMTpmz/sW4azTwD7ohYn0Zfo0HHiaQjjrYuWbZHZzJPc+OmCAmcri9S4KSvPuQ
1T076pbKuqLWNdz6WtK5o8xCfUHQiIIhQUriGX9w7lgrILtaDDYZdkGqwdOlWpDX
7PO4jbChybKb82gBuFpv+h3cA+x2BZqJdQdAQcJ10QNvMtfts0rOr87Z2H0wyzXM
+9JsiTGvVI4B4XcYsYGzlOnOuStL2aRzrNKUlC3jR+Sf/1Ae1gkCu++F237Gs8nW
KCWLw998xlc6lgUUKZtsnhxbqgpPq1LBWXQZC6vWPndcwxxPlmYwkCq4mbgGL+Rz
vlkigneh4KTDU9oM2cxYlTLBLIT5g4UwYdvX+q/W9M9ggtu6ZUauCVVP11u7Gpbh
EMOsIzSj4/Mmi1lPOz/2x+Bnghawhjg8nRlK130ORXZwgk002DNqW3J+Eh1a/+c3
hMsjPmKPVOcJkOwzPHtJPeAVFhAeOk2jem9eFeNs8z9jkdJRROZPJBMHcumeqYaL
q1et3lMp23dJ2FvM70zNDMeRTLJfIgGgwauO6zLId5O/CSG5cEXFQ+WUDUlVtgcg
IoLaXuVLYedOmbqUIZlVLs2ACgmPVu0kZ7++GfXjtHpGfV2nEs031seRq/FJWwqZ
zVi8hbr4BdbQvwTgjVyzQooUkFh2WRwsEwWki6RNVb3U242ySt6NpK7xzABEwg6e
Kie7L1SKadDys6Ipwa33+yN+Kiq/JMEV1yVbG0AUWEeYS6oivRRKZj5gQ96OFYPo
fdTwDwYI2+vm+fRXXKXCENbweWZCGy08eFR90FVnxOaad42udBADIAjweRHMb2AV
qhkbp+GfNy5T4Ipyc2PpmZHH3DWqwx61yo2QBIANkyN3RHw4J1etIw59qdtiiwWS
TniZ7WODwMFUHlHUo9LOtUFLdKPRuwyoNMSraYg6iJySZqd7Xm47Y2JWMYVT06pW
5ixDVGBuNtJmhrmOagISGbqlLi3aLd0GG52lyd2n7mVq6LbDhFI3quEuFhjbI5ez
ZT0y4rc5ApJQzb03UiOo89NIlslxLC9TVAlkLfq7h9FYLTn/BayCVKuiHa24osMM
PjtLEwew3nQp2fKkIElOB+7NjcXsz3E3H9N+d86pLT8+1vG0nY4aF4jpAiAp0Q19
DrwxiRU9MzCD2PfTAn5GutAvFo3ZhiesLqWYDzMHvkHz8QhTvoSGSvEln0i0pJDm
rcIampOULnpu9mWlnidwVMO2SDDVhErrFgh5p0+IGFFBTfj2KBUsqur13xHRtYo5
K0swts3TdsFeqBXo358YwA2q3K67CLetBSB2IsT/GSfGF+dHD1KB+/+lrhJa8euY
B0XqlY/CVU8KAkaIicgcgZpQWRqadWVM0E6JvIA2PJ/qMuXjmM5NeqtEs8oRnM+M
wcxNNc5CMea+K/9KSlV99+MduCNxatkZtOnOADmwObB0XN9npGiSa7vYB6LCaLWD
L2oDzWNw0gu75dv5MuGmSujGU12lcSQj4Uoh4MCalVRuT98cUiIrySvhZDLUACfE
aW0GE6AXiWZVjv1fQNQwjVZKfxvkrmP14OI50l+bqxWYatTok7PqplKp8fogbDb8
tyRII6vbLihaI5iixjiCaOuxUgO4vjJeWge2DGkRYJnPPuvw1DVuvm+RSHQnjKF4
htbvwFjoQ+DbFJB8lAiJVFgnnG/3pjD7ILI1rM+2Pzu9WB5oPR9AlUBlBLKExoK+
pDGIchFsGGQSPLX1vViAx2dvLUL0GQy+7FL8Y6Pn6tYS/FKJVI6mHKv10a/HehHj
FdaglwzsXhNl6Urn8rqbXIl2ObXg8qF7ZPl5BCwEcEcp+Vir7dlywLj757kBiJzw
CYPGJk1gxMa0dIxCCWSucDNxjEznhZIvwBLNicAzdv35o1tohiS2Znt1cQsKkdJj
DY6mu/5U3vNe5/io+wENJtGDrDhem1e0WyfxqmlXA1IaV+5wNzEzyj/leKlyhgOA
o/w+BkAX8jOUl90dH6XUCvRcB36CkAcmV+UtXDPGOil1YTSObdBhOGxmg6WTA2RR
ra1w/Ku82ZfgkIGMQpw02ohBYLZ2J8DPjjdUPmsUNFjlObtSl8dLSV9CS6dn0BcJ
ucJc44FpKQddqNkzkOKKU96rGPcVEefjIMbtA42+Qq1msr6hUC5Qo/q/efuvPnxK
yzWYEMAcBcsiUO8H6EjucBo7YyN02O9/zZp4/+6IuIaObcK8irT1u3Mgd3HScZ1z
ATcZhP02YYcYby0w5uvKzgFMToh3sMSjue9nKR6eeaXpPshsELZfRwiWABNjZvyp
uorhRpIXvFOe+zjsZcv8I/WcwGD5pXaUKyOupavEbhK/EF2mA8D0B/uYWx7J0sK4
Lmy97nJZ17DKzpkuT9qn9DIUhlgEAYbIdQKFS34a13a8qDETloGRlwNZ9i/bCp3q
h5vWlBUREa2jGZDqVJTRnKmd3ySrYpjvFFWufAHImNfzH8CAwd6whYGCslLjOtG/
Ep9v8bskn81egv8h1PLPdNaA8S72J/AT/P9DsA5kWEdpUk2bY0DYbNJIST/N5Qk6
isRkaEBBZt/B1oPV/7+3lsEl9HhmtlCIMi+QznyCzJe/opDa4iqAYk33rrHBNusQ
tASRvi/anCyBbATPSplEe4FJwvhO0KnuH2tM7tJ68VXVP3rSQ1C2b7wRqwC6JIfI
p0WXczmq9hGetwzFP+uRNlwmFdMVqkHtG9mom0wlNxAwOz8mj8PHkwSBxyvDC2k7
poKtzsRCnUurQHfWBTKvgR1TCrzUTzVJ1q4ugBf/kJYacOTF7qn+niXouprjNys4
Aah5C6zsR0oiVjJt33AUOYxfCZBDSNGIfrPRIkS+D9gCaogchjwQIoHN/UmnV2ia
dajzqNooPAWPO53NQ8otvCaBQWpmlVfSl8s0SLC7nxJoKhg0xmDgRoZt7hTJ0jbt
KG4OQ3O3KfDe4jfCwo29xhde31m6Mde5sscYjw9YeOi42x5jHER6lDMs2K28lccx
34shJ7btwjP/4tm7sfZ047JQUhAE9kAEBNothXJD6J6MiJcFqudX79LR/MDhwgSB
ropJ+0iINSxbKff2y93aO8UgMRuECYnT4fLogjN9ZXALOk8yJNk0iaQJVucZ7i7e
eC4pq9OSdvDve/HRAYuVpxAiKbAmFuMHQpPeN+pj9YCFAGJV9b8oo9oN34RQvbCF
mPr5C52E7AiltfsCmy6yEULsAuUqohPV5dqaPUyPDgXWko8xhYbVSpIDR/iVhcG1
NTkfO8orErQ5WInZH3Z1uiTRIKCCA/sicyAuzYmLp69Ngx1BWNMjSBKT1toruTb/
6oidbhFNzBBCEPsLT2OQF4zqYqd31x4wRzr3FGa9ck9rnmwEWnghOkiYZacvPz3T
0sS64fKyTc6/gNdofpyCQvJv30dBN4xSV/DMrU1D1mgleNJJjIBsWotbi4tVGp3F
WkPBn5WGpmkJ2JqcY50pKH1AyKLTRr2MU6rQLJLGFkfvZO6ogBvjCeBwG2jWmqq4
THTK3BEOk1Jn9weSA5YzNOUuoyK9id8dbhRHa1Vhex529wngEBoRGJrNeLckOTSF
Lw+k77KHSCtdGa5BfaUOx7yGI6q0f0BHUxlvdQozm+VQAPwylR2GZ/2S9haWVzPR
TbGojeWkm2TZ+zLcGnRLb+BIv5Lxx5MZhbCICFg7H/6mJVZK4zh4Jsr3ztexE3dM
bWs9zNnwWdC7Mo8hWMw7rWj3FU/WlpJha4G6Z3ALum/Py9JB9Y12KXdJNrGxePZT
tF2Gzjl+YQRtPJgXtn9+dactJzCKcUbuU/5sybLIMyRk1jmSyf28nB2k02c1KsQp
Mqi8f3ZIsbuOVntiKa4FdGKA4j+og5AcQpiBEUqCGfn9XsZUJogd/SPXu71u/zKl
FW6TLzytY9gQn5BiUvOu0p17+HgYPyShG6d8DtZFkcmilsodLyVQFeTC08L0VsGR
myU3URyfJRRKucYD6zqNsHZal+JZeA+Ix4qEIh/9gnHmLS6jtX2bmizV0OqNrFzA
opzii2y79QetV5UqfWoMnCBLjTt/d9Uhmlx/NWo8HSWObiyJtLsQq8SOYR/7x1G5
5q9RYjE6XYTD0Qg40PQd6i4uZvV49XIxvfpP/IFcu3LmFdJw2lBOADerG3GfQ8r5
W7BEcJGH/v0zpCaAcWq1+/5/AEJJrFFwdrnk2NEAsXHipmye9wKHzWjxOGCenmnu
IPo5ZKf2P9ABlQvS5R7Vm2ZNitQB/ayKJkHg3TpucdLvI4sgbu076irc6fye4zXP
T2gujttfmOZSpWhBxGKzszBlZMcYldTVzy9QbvnGayMcLo7BP4bQ+Ptk/+qcEXbW
Lm8dy3DXV5GZX4oR2C1YusdIgRirM7TgUv9aKABZrNMwrQOJO3eRUmkLMRBI4QV1
YxzU6J5xG2UHNXJ24eTYMNa8+ZrGzKJMBzePHvdB9PWvmLC2qcl39TmrQWKOS9lJ
ssY0wGRY6X6hYG1MIPuBNiNm5ncS7g0UtvEU5R49gqv1xm5T3ttDPgXtiTWXo+aa
YRmllpTM2l/QJy8t3NsCKVsG9WyLuXuqilRfwkQ9ekM0teUEVP54gwGKHewYULL3
zfhlzwf8ZO70hBD/urvEFM0HRValmab1hUxUAWhzlEFQR/JANl0chCCP9qIiOat0
qHdFTGTb6vUiDoHL40Bu1iJrlF8gffurUtGNgJrsPUlysWk2OCSPyF2jXmwWW1pD
2Yk9bpj7y/ydMTzhLRswSosrZ2zPmOxmqkpwg3Ob26APiFeO9mUes0dZxtCr80gr
3Ro/4uaQsiY8HAaJvuBoOMwrnZIuSsCDCpLSFZ5kSqsxuXlEngjbnEyNHvXB8gHO
ecfQe/YuJemCCzw/c4nKx1ViJGPLGPUAmcxBwUP/X50031H5u2hIlVEql77HEAYh
uGJRS5ctqSTWwKcgzLcd0zLa+ibUCU95dDXqldVk7YdpOzLr9K47B9N7ALbtPOmS
sPR59qOJ4THkCNX0u8WEMwDJjQmovou9JS/SMQeWPCWrQcU4qfSq1r2hPVUZmqaU
0JAV/My7qcMmWJOE8RWms0tuR1HnBEiPsWaWm58OnpeiWE9QggDDrhiDxYS0+GHv
xzhV+lJzlNCho43nM7f9EYr4ewwQ0js+regdvYH6L296aCijodY3+E8/OZFU5pBI
fAJ0Skoc31DJw62RN0V5yvH1BTFaPLhRnzSzn4wSMSN2gDN4I41TELL2ck7jvQ32
sq4cZMObvGb4f0jrsTChmcpwwbJOFi8JtgzGpoagHijyW2/CHeyWpUKI4ldSIx9R
gAlijKlY/pzhNMgG1ggiFsqhzlqoZGfBiRluHqS3uXWkgHt3Jv/6wxC9ESwQRQcR
8ZDuL96miwdsBIdam5VQTBT2zJz/ygwHX8LOUx+pnhja6IU3HvF0uMzEy3Qv5G1T
bQiGuQAoe3bouU8O7k6DGmPEQqnGQWRHMh9G1hY+8IDVjB/D0aDLLivlQC8z4XCJ
wWKtsiza3LR6InmTtmyLXNDrDgo2FNsB5XapPzUbFxohVi9aLV08Za2Lr3Ls5Oqd
yjmFsXrDmSGXlpw4uo5vx5xOBpK6ywsJMn5fpbiIfUIefAeRUQtT1NMcE3nKolCE
TFMC71mJlioYJsW2jLfkBQz0uMRa7GMSzgXEX3LxwcCWp7l0LY8frtR5edQ+wTCH
Kmcm+rfquBZQYCRAUEedsL9BRiQUhS5Q59Jj3pUGIrn/dxSbF1+bBr+4JFddgpjZ
E9lUhBmHL8iIeZX3xWCS3n4IzzFmzel2RMS4ve7zOlrjEb54UlB7tR2i4lSDL9M9
ITNrKVGEft0U/w7yyzn2UEIs9ZjfiDKDoHgU+qMan4TzqgtkQrJvDqFPEpZlW/oy
tczv+UvA8O/ZWn+zf4UALp7IZR6d7wONDz140+Qe7Z37FhdyYryg6CceZdd68UJU
reNxImZhAjoRLgQEQ1IRNru+p+XgPaSCnWToeFDA7ohLzaJ+AgdqbCeblKiO3yKL
7goXwV7UkHuv6g4g38a2NQLxRJo017GR9tXJzr/Y7yFsF6Y3crW37p4EaC5j/Vwn
AC5zxdQDItQoaNczy0JAmkeK7cEkJqzO87ecDNDP+jjNW5RCDYpx2iqq7t8zwmYA
8izjJ/7Ga5S4eyu0qLlGLghFH3tYKxbxYBlMfPo4iuPUvlO6j5ljiz6pfUNg4I9n
9EIsycbZXXWRyoVKTAz5JdZrDjui8cyQu8ibgBItIT+SdRsW5zlEu61THYHo6zxA
z0f84lFgakhD5Y193phj45WzD3wk4pHXc/l4lmeji87KEN3hdm05ngvlc+wWKnY4
ca0UtMhSiJWWw2143fgPIgL8xWau62nr7ZxUUeR+BR+BIvmqlxKPEg4M+XD/FL/n
CWKN2c7L6tLoW3sr617bo4XTXFB1GNkVmL31E7wSu9NHWLkLRu9xUvrTxAEw2+x7
`protect END_PROTECTED