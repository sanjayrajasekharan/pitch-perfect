-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
bZKa3IX7wqetzPIubueXlCsJRTlj60SU8FoONIDcxcoSQtzgkEQkHrfVEtGMe43j
1GrahmsclfECoPFDhcYN1mzFgv2ht7K6uNlJIw4KDFHRX/6iY7qOvwHQxf2ZrC2v
28LyDKAipXcVpUFp5+gPunE4VLfm+2oc6fCEK7CiUSM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 16528)
`protect data_block
xna8OBA8FqEN8/w4iIe9Aa3OL2qPe0Z8H3O/hxr7kr9gRM+QxHQ4asbCxABf1wTz
ZI9I1CH1c/8EXX8KQ06KKfQEDkbgoh0KyB2VPDRZlW1j86BpQ76FTxSfsem37v+H
7QwGTq+XqR0AjcntYtWc9Nv5JU77o7RBXHQmu7jmDMMTGUApdvSUTNuxJP3dtgGk
+nUBGR2BCrvtnWBoSMLfnXRZFdJOfUaX8hZPsFLBSAZy8O0thsuyyMQEc2eGYIK6
bgL+hmle6QvksTtBtsjoxLPHrYCMaOir/8pi3ibRq42jKp16ppG6E29c/aPp8Q8f
qTSUUZPJKcE5ubKczwSsq7RRqWR5tv/Is5+z4wksXmi15tnE0PESoXH5Dh57uBe9
oHXgdBaNy5kOqKGwqujiZXy9h8G8MImpTU5Wv2XJ8ajOEXhSw5kUL9f3Qc7b6Wso
BWM5/hR6hvVZ3yEI50s+ejqVjY05YseK+oo5QtY2nIxfH8o9Y6/YmqJxSQUftU/h
D9dvWJq6pBfDvFwLzEKdTE9qfSuvdMk/O+wjUMLdgd8lZtl3nxJFLUOhRQVH0U/p
8wK+3/+97U0wQ5v03/r/dHc43CxDSeIv73dtqzAqA7uGgIb6dD9HGpAK4wnJn27O
nfTdoEoHEIrm5hE4kxqEtMc7j2M+JoQPR9KxD5aoz2k0gB56i1NhMUCkPvqJD9pk
OtHP5donJzi1tiUBOzLbGdvNKK5p+C0ErnLd+/SH5Y7fiCPxHhQSIHhFbgWMvXde
SWn9G5A5Y+2GOzmLPPZthmsz8nfGUlsasYCxdE3Im1gwplGv7bZLM1dt1Op4iiQP
V3IKj9NZjvnRku+v0wCjvKQflRWALZkIHjF4Nzg8qy1EMf2XkvV/OEDSFcNIJPQH
DZ0r+yuVqaPr/LQUeMzYoRZ021THXxTNN7eGFV9UN6mJK0duB1qtyb+nTQM+Xiw4
DlW5qejWy+oAbOBbldg19m6Sb84uTcT/Feto+jaiXvw1T2p0YNSw05HROhWYJm2f
Q/JbOc8XAOqyJ8pdeT0n80SemVlxBMildimjQRnjgNUDrXoa3ernPkZ9BG2sM1hu
1p6fM3FNJbOFObCfVlXZp3qwOuUX/HR5GcLYczoJ4UYJwu7DNpcB7U3Lpl0jDrQH
vDIvzqlxjT713Vpw/5b7SV8PZ0RRnsmraGPOwVvSqB9lrNIta17fI7B63t5u/Va/
dSzNLU5dOhla1fHIrNmIzjA7xaK/dRoN4Np7ZrB3f4/SbAWPMGh4IOZiz4eA04ro
lJZauQV5rgcAQYRcJMCQc5i+fMunPNn3pnnj1EwRrd9GxnunTDqCTZFqWwI726yY
HJjpVOyg3XtcBgI8ImWpKRE2gmxJgG/5DTVZNf1GoL/DTGX6IJrOCp6cSqIszhUe
XiqUF79CyoaeeP1HxAdGmWsJ2d1cwGXKa7tXq0c0XSSdMlx84WMQ0puxNdKZD6lc
mMd0lB7Fyg6u9A8CWfyYVgp413TSya3qDVh7TuUTNul6kFBSEOqKh/lpB748rGuj
z2KeqBxs6M1qL7SFzvAMoTpkLXyfv0X3auX53eEX4IdSVMpXhT/+8Z81nqdqIIFU
FbSEnsrQwuZ7035NcMqXk29vpLjsqN4ZAlmgBWALNp3cYp6TxBL7UkIEjJw6dvzV
Lf6dKtqdAchof1AejAOSxmFZwxzLp/gsSreK6DByrbWhdKJiNce0/Fr+V/sYXfKQ
k7644hbbUWXHmCDaxj2vTY3qx4ozh2kfEsBvHKX9QPNEcsBlSGIiickKgABh5xSb
oA6v8ijwD8hgsM2Gj1hcg7q2xG3Czk1ZS8JOq/yWsZNFir6dijM/yvygHxmIxlMy
K+p6LvUQqg1DV1Da8BzCDhZkUf5ms44yYdC056UDIUNAjgNdaOKEzKpe1F8+1tZs
6kwUeFzm64pxLWkjPnzLEeCt1zDpdce0FJ4SfljqYGZuTimju/9FXVC+WGYj79nx
EEvfKtFMR2nzYqkiQI76SYfoXg4wWPZBkDuQofVxsUW6uxjIc3278U1lOUdnw/2o
jVaHJ0F8KklOzKi33hZ+l27NG2lON3B3sfVHo1KPNuqaLz2Z+yl0f1WXIGNzwPlW
ZnvBpxxBwjw0rAJda9uSI0RwgMjxsKeimMeOb3h/7GJ9gxnHWo4uEunGH4fnfXjQ
3T5QEzzzxEu+e4jElkA/GDikByj1LaWWVnI3MosGEueUdNf0kXd2y9sXImoQMV+a
uCdTX+lvU0FO9MfbJbn9NjBwgZXUayvWx7s7U/k3HsJgeFfAM5A2mYqeFF7644B5
p10iOR7/KtHQ903X6QDScWr5EnuYoXEtoHgC04vfR1COGLIXEaEaszUS1McOVFs/
ck7moigCMsKbIezUnK/q2T23xy8rxvMP6B1iLylNCJGws5H6CU/sjYVvcNqgQyMi
9UmwaM8ePSQt8fewIi4v4nhZe52grCf7YBHpmuyTIAUv7Fo2OHj6X2eL/VX9lN67
vj0B35GavZm9xBXHd0/i+o20nZS0BN1XW3AxZcj7OHYWjO6Jd5SUT8Lu+TLH2I60
nJlGxjlInDlQQJ/xRW19Ci9x+VdBabaR9LtqZP2GJHVB3Fy4UmU4eh2JmnvOnaJT
EQLjTX6yH/sgfXtEnmc1LWFTL/FMlL2EWxiB+VYhEWCKAZeRktNq/CVaJXi4UVau
2NV7uB9EGJM+dCHYPJdtaJWHynFNeM47BOn6b4w06Ssew++aN3ZNaeaLqOAAL24i
m7y4PQu9MKxLbS2ck5ACBkHhViwgYkelq3eWcaE2DFJoI/i4tFX3lva/xa5Vkp94
qM7KdDETB7QYccNMPKfy/skA6zg1fdLs8t0Mlu6Fpu58rtJ6N2rhJTkCDC4X487K
MqqwlcQLcSebhgaSfdk7hkE7h4q/Kc0vSfhr33Xa+1OEsUxXlb1ciS1yPWuQ3q+u
ZAsiPPVIsDoLcUHCWEmKmi55Xucp3A+HoRTA8fILS2fAKGfon1G02dat1xqrnHQs
naJ244fa2thU4LZvhRLkBBQZ98RaRQWkdhqLqx+8ZrKgTLj30lFWqijc+M/GmZjL
E8tPJy2mARFTUadzH2c5hf2l/V2zyNEf/gBB80qGfBy/3/QzdrfeycVDFs33TNpy
eJihHZtnahGRhdkVbK+tz0R/gC/qn4RRAu4vmQNIFUaVTy1Kv6zAe1DXGzjzJtDy
GkFYAlFFOvhLPk7PXXXxyiCfEWArgk59WCiWVtPp7DljzLli0b2Waqsxf6OKvaLI
Si11Sq1Yqsdn+lxpymILHE9ttU21Z7ozKymVm9Mf067X92Aq5CsNCQyFYMQQ4xrI
CdXVcJlTRktKa8iG82lBiJgtN8KNzCs8JHPr5msq/MM+KAj8y3FyMf2lY0py+lG4
zWvu2xhqdVdNeNiQd4EATLgKtAk2vLxZ/gKrSYw62hv79PT9bNRI8po6FrJ5pE2X
tOZF1sv9EWl6tgi6ZIpJFslkGW6qdyv3i5iG9/vNiLWfx6wDy0UkMElIeUH8z8G2
F9EkTdZ3Si8X9CTLrAYiJfTs8DiSwMtbuOzLqsbtjHnp3Cs5yplVto3dqhxsdjot
//UsnutWSonpuihhnooohIpsDjhADlSm94qoDpO6nUC6nfZK8yWKbBsNzI+oOZs+
KH4+KwdbYTQhPU5zUQoFqvSJvNQhlrJQoTS4mtYCI3GYobUV11qUyyRk71d99Af0
L0+pd94uS+XQI0pGpb6UhA9twVc0ltaLh4ENT03pcDCCA1Mx8lhKUg44liUclD/a
SNPPSrRkKRRqsIZQJ9TFBQPtiz9hJuRk9SiyE+6LtiwDmX7VGITmozIei5drYiB8
8P0iKFAEON5Sz3VtbvMmhSTBMl0ERki1XUVt++UB/4uKxJ/Y59Tudp5wkcNEhyw+
0/ZyGM9S9WOIWj2ydYTEC9ElBGgiE6uIvtJVZSINm7gAvp42L/koKJocGkDkBK3B
SdT3H5UMV2M2b45534xfOmXDhwfUIrzk4Y50U2PijT0ALJGhb2y2EOCOqI+qKq5K
/SOGXTZeRnyScv42GZWrM/k/cACZSDO4JXTTqprFrkdjyWkae+lXanHWyzKtM07R
TLGrFpd+MDHuLhoGCQCimQj+ifMv4rNCGuutxPBExJaqbXWiPIzgrPe4wyPtw5FE
6EUU3bpe6t37V+fuhQ2oyiqgOGHXL+Lgteh4KwIfldZP2ld/GN88pe4Rtt1G/+Ym
T9mF9M7OdBrnQxao3yh9QsqONWwwxQ7t9T85H0mHmNuqt4LNtTB2y0b6atyoVpuS
R0fuKz0TEijMsy3WOlOF8dA/JSsuxennLX4q/470GGLRYqn+SSLtDPBnFrK2MHE+
lIM3jaEd5MPG6MDtYBEuG/FQG1/RUNonWuEDHcSOcoqK1o/FAlb9IJ0sADBc7xvd
FaTBqlNB2h1LshxKQQL9ZRmwEXLfyi+JgDFIKxBTakNo2KlgGEOEdk/RcWkTSS2B
SNfn2quA4Vi/t1Z1br2gAjZRZKqq+8C3YP7tw4GizJw46uu51fAOzq+PAg4JX20J
lZXAo/bNj04IpEG8u65hz4T2VzNXhm8PJ+ubFVmRn/KpVE7wV31+Exrgvbv6kRmK
aRiug3pLfsZ8SzLc+4/yEPtvGABuKZPhGOPmc9UY51vAr6Z4e7cTb+MFaI2nmIAa
FRSEyj27QfIc93xVgWj4TYf/eFjpJLhCqI/UbZFTn3u7Rt0jVuLDzeAho325TxbW
lxa/P5E5MrQx45od2CzWRl2rVoeDoOmXNpEZfD8SlU+LsCKTLgyKwSFKy57koy9h
JZ5Z/mkLqFoO/cT2oqX9uaCssZHDjqT9CrVoPxpunOBmbPhjYu00t3MnUr5hqGpB
mAqoM/f0l/n/D6QUdz8CX/rSP5nVg2cHGqFS9wQzbdhhdKDB3ZnPJ13KScz5+d2G
VLOnOp3WuzDinktawsavJUBuRo1VvyIaTPhEPJ6EHrg/EhnsL52kv92e5n1LBbBp
RRu49w06YV1UizXlDIP9b25kj+HYF3Z6S3x9hSxcoWsZ6Bdu8Z4R/lLR8XBDX7PA
K0uoWesUAjNmKqnh4FptqL4T7g9pVkQDTO/bAkZqzwuCUIU7hdz9w9v8o5jewVt7
ldI3+4A//TW9Azkrfm5b6K1Bw31jeQZR7QUEbklUcJgRpvlSjCn1Hp/acR8HfMPa
mAzpKkIK7ozdt9YPDCQfGC4tKdYF45gWOeeymI8Og2f4oehECdLMPjTsTRvi5nGs
g6WkZCYlCHWc9nl7+Ys1LKwbiXJ/iLOddBRmS0yjhIhfr4RWZtl7sMmweMNGIT+I
s4sQXzagqaEKLlkZBHTYbIrzlPqy3a7FlKX/T1WUz9Thz01uR+mqCEOwzLebvhjx
0ovA6ACE2mlTcz4VGu3V5xyB7rwHH1xPLxo9+7jDMPGDu+QbFFKwnQ+Jx8dazhtz
frWT7E2FWswh2xc3I1HI3HfjCZgUX1UncBOfwAaAQJ8c6QFL/g7Yrz6GyBBC15ZK
Y0Im8D/IcS0zrnWVSKJggx7DMIgwcAB4flV/vYbHW1qSWNt8ABCvg2cYNNKiO6pT
9J/esSj+lgDs0Rk7Bq+pQ1rkF3LQIeFG2UzIDqi7STyGq7blSGxExQnXTOSyhm8a
fKvUZv3VhNtGLwTEhD+AP20UDWcnJU53FYvIvSc6o9XZNxhma7WZRiQEVIRD355o
HcXzKuh+DfsQrhgGck4w3Zmt6RTJsEtupy/IK6yAFtl6mQYrP8nHklpemWjGztTf
ju6RYilj1YN2XwQdb1LPhFsOyvtd8hy6At3Cdg9K5pikCWzLVInMedKFO4/pmbF4
LtohGYlgaXB209Pc98qCnmGwULp2x07G/lUGI7OKG1OYW7PxEyLRdUDM73huAaLW
dmufqM6XKwBtJ0poeSXd5/epRrB2rJHN27yZjIM4sWXxnqX0wEOhFJA7/K0RGhuS
CKXPge+e1cWfZvAjzFBUewDXMCTP8vSrDxfDqlEW1szjWJvUYMTS2hX2+f9MsOHg
Br0uuc8XVO3/ELcAiyLYjVVtSvPYtGcJlom4RdsQIn2kptf1gq1UDrBhW61f0lJK
k57rBZixS71Pj0lII86wcUpyXNMM551XmC0GZgs2r3ei/iZBJLcyMKDEDhEEItQA
LBmCrxmiTrFD75X5akkP75DGCWBnEtMWlKnIz2W3G4Kc4uFRkjStduRsCt2ZFjN0
2RgOev/YD/NzGjOp/qs5SdnNP55HMjBq+UsFc+F/cwX8BONWxO/WZRpeN4Q27OKH
s6+ukZOhkumpxyr9IGTGoJ1/HFZjwtYpMRgNcyISkc/dSvNjvOPIYEPtzFe0fSmS
UPKaS+1m/GkDrhNijYkL0xh0Yq6+NWuTgPkNfPzZsHKz6YyBE91qgtjYyH9ucuEl
em55qe7VYx9irdA6Lu6gza73+7tQ0mMVC0KG4VrKvb4xplenNC4jaSXQMGuILVdb
92gtsGYZvNlUwJuS4dzhj2NThxN88ilF1Pzfpa1YvtOM9l/WKUXXlyDkKkvNeO5P
TvbsnhtDY0ePkL35rfSogAUENOoc2LbSTick9i4EnRmR8D7KgHqK7wMJiZNL6njo
hlomETkYoOREY4GtOvNtBiq8+QHcj4LUotf9oc203+NNTaNzkw/uRh6w+mIdtFnM
jtcrzuwjRJE4W8hyx9v1rJ0Ebgmumq+qhw/ozgovXVmTq+UvScs6VHMtlfGZML8S
Vob5/budKRRlQsBqDV/BPmrSVw+kwiHJGE7Ju2WJNJs6ff5m9EsbzTa1ouj+n8cB
QHhs10kY0UqEUMWnLDLTTS/wE2zVOrRaVXrqwBpiK9YFbGCkgD38ASduWux7463L
6cg/8z3mRgPJGfdPWe+jSkl9QoJIGcccs1buxP+2EiVDlFJ3YK7y/jBVwljCLOLO
ToBcpZMcAhD9DU23+ignrx+7frk0nTQoB7YxrLrap0YD/Zkv5yU1OF8r8VbLUDfu
hZc1WcFCu/4DT9PZQLSVwSwvy6Rzgbyr0P6A+s6nCvClpNuLxqVjK6L1V20yeaI1
hongoUrSke7KyT5kbIsMYZp5J4Y/AvuWtzQT5uGvq+asl4k8f+cY+rp8H9LQgiLA
YWTz6YqqL73OX99//JuJrgJ9q46dF2mLcCpcabWURAzdMG9rLnQg+ZL+25FLbRvs
Nk73my7ndMo3xKbZI9QIvsKRoVnNiLYSEN3DHSX64GITopcgNTmQe4xOT5+hyBca
ejGNwwqMeLjUleHoi7eb9t9uTMFaE7C9A2myVIQg3yWI8NwSJDD8++TjxSfPmH4x
9MLUEO+uU/jgrrM/8gM898hLxKHL9skyeETxnGzpv9zczE1rQCLrrGbAbzxZIXIJ
DMwoGIVROEbMKHVhJGRe/hNXHFTh+iclJH6kGMZAXDBe0Hd/G5LYlsHoGRtkMG2T
EGvmjiUAbBvOmRuRqTUFNHNCrrDBP6PkDZi0vBx42ZW9C+FuFVC3iavNVKXfZsNx
uMWZ/N3L+8WJcj9Ev5uUZyS1zqYWkDyMxRDong1m9POEM7OK064n0EULRBLOB3SG
OlT8z6J3S+o/rjDc68ExExfJmQLiqrJinDPDSfvCbi8RfJW//dWH3bZON54pYwFW
7frGObUXvs91490x6iWniQ27LMFUgujouUcj6c4TR0NZXj8dnUkDxY3VXsQYL3Gi
yVJb+oYGnUDU13R/ugI0MILdcg3uvCf2aCjPlIytJqIkFAGPeA0OEk2XWVBKSFaL
60M/oU8DTsamig6JMlO08PQpznYTC/osD7/unTXtQ7AUr6L3muah4s2N5iy+Hz4R
i8aYbEYgD/oxVWtlE+l6cb+RqqRxtrmfKt1WVkNetlzCbSutdyEAFmxa9/Jzu6wI
K4PeW0sEnJSQvBxHJompizT5XGjaJ7MsS2/EkIyOWaychRm3kqjy/XlPvJrEmDkp
fg1n/SbFGIqiGv71O08W5B0KZJliofsbZh/UuNV3u+baMpk5uWOG3orHEnijpDdu
RM0vEThIKQcuJt0yjNIUt4Yiv+m4JTNirEoXf7BfjuAcVxqxRrRM0yuy+7YwlwvJ
6LQhHpbtRMUDrpaBc3n6ToIkcdTuAJiFGJYGyYJl3lZ4N++MzS/3/1aEufleL570
NbNhcw4m/4kegoYlTW01VdAOmpmGWwn/NO28o5hSeCSwLIBREq3Qr5X3TlQp3DnH
9tjXxVhG928FHxlyyDG0mAsErNi2yYFfEoyFAVDev+ORSpi/qe0TF1+KQxLPdl0N
e/lWJA4NmIyQoGKr6qWxNwhf/K9jurOkdcDKCH9QOKRnSYpotvO+UdFs8KiPKqwq
cG0HVKONselKBoxXZkfy9ROp6YWoKofKSNmTwHLxtA44rfmdgQp3ECeOtGx6WQjU
8DkLN+qfCk+6KhLBTGpzVlX4k2khr5tMWHUyaF7XaUPQqqp9RtnLxDQhvcTKwvLQ
/TAUBrCwTo92N69tHvJ3HxfW7LKWP55ABxB6hw/4IPp5ew5UmNdwCFbjNUPVOCG2
I453BNWBZ/Ei3a3vv8KQPlgMS5VtFuMdRktk1lLe+bYvgj7Ysg5UyXJC9DKM9yoK
V30DTstuVnzZ1RLLHNC25DKQW2cWXlBgBEcEfojJakJ4411MDP+pIgno61ke2VZC
xDM9hzi06/70WRKDF2ikSiNo8QMJytPXiu5EQc7Dz/CSXZhC1+jaoApc3NbMIS6Y
2/boQucYxKjkjHnxwn68sytCyVFOTqieF5XbxAdItL1qEDOJPD0Zm3KvoIMDUui8
1+CLRhWT7etfM2GNtdzEKqhlUyWSY9YhCBD4FZUgtdGdL5c9QR7Oe0UPVK2TxczY
yzQYcVN6gC2xsiSzpz1TdC6NOoPi+rmnr40zLbjHQ2KItGRPy7q/PS1EgeJdcw8S
gD7RGoXPyDuXnRlV2DrXrOprUtbsMdhY5mSBskt1V3Z7R8JLc89qabm+0dLwso6X
SItu4hbKie5u/xKPPxLNwu8/xCrEc5Dl4pi4n4t1kGbeB8L3CGrYJmNd5hgpyrDk
wwyAssFOZsBh9Mw36jWvkG3ePpTKbdlcrQ+NJ8W5hVrqmaWMaaSOZzyEUIfevsRq
zmbYHHXbOzQvyefq9RdhHwlc1tU0MS2UQWA8XlSl9A4f3LHlM1nX1qG1L1sXUi5U
OyL6ZSAArLQUAocbRWnoRW+mfMBamtbifSo0bTklzIfkAIjJzbx3s4yq6IW7VBNK
6OwDYYg5R5jqtSOBj1L7m2rnysk9Wj5W12YGSXESzPOlLFsNpGvdK/5hQlw6vina
mOEd0EefQZvX60cMsuTRTD+Ps47qm4DzdGZyE0bqZey4b35vac4nhqZ8qV6mV04B
6B+k7Do4llhM6tSAN4DMWrBLtSQzT/dD8IdvN3lVH5/J1TYjf4HVsIx3P8rJEhyW
T8COpSuUAUDWEqj9Ld4GuEA2YOvBjYZMdr+qPiyV/gwABsvw0Z60+J9c/8vhzC5L
W4uxKAOyIa+Btz88TwLgu9RYqr4j+X5e4Eu3PYadc4nvxz6OGbov0rKZ86elqq5i
hcKpLQOLhbh0kxZBgdKABSMfzNEmyh3p9VGFZqdMaCnak3nQUuwJhRgQoAW+JsD3
iZDfvUyFtKvjvcEe8njFepUWtxDrmOhtmi9CDSlngzmDvImVsGN7/bNsYBLs+/uA
jdv0vWrpnoSeRh6GupEhor+Y/8qEdvuArRPBE7zc1yZUaSBYnVPnS85b66L0GeYd
TegrbLsibhMKpJ/dW78IdiDA06hYID6QItVRZp39gh+H0sc30+W14yT96AKl6lV7
LrqYhfzx5XfqRJJm4T4+3iNFiz3DVdQ1CtJQpSIYnFSEm5revuQb3j0Vcnfcn07K
/yT6M/sD/YeyA+kvaY8/vXLbA1BHOuc+/i+6vqft4+h/3q6MxhmkBYl5BZ2Kfvz/
g2A53XG1UIZaNfuvt+0ZKpW6y/2kHKUmKnQyp87+OkBeImfa1fO5MSRt/QDw0F5N
gF3DU+DIYRY9p2Qgd00AAdX9mHMEXw3B3M85owR++c5sQ/vYdDt/XZl83YeEOMJ0
joc2ybp6GoopRmmgIWDu0aE83klnXN5AlzEwvkhtXfxJZMrV3kL8H+9OJlogd9R4
eV5AVGLbwZ0eyS+W0kkvyQVHUU6RVj+Nz3inocPb29dz4o5bOA5r1+gdjKfiqRJQ
hSdzfjiIDIR5YC1FMbqIr2DrY2gqYA4oS8T2hoce2NaI4EiSPloe//QCFRyvBmtS
wOhlRz3gq4flSPIDQereh5BvC6RDn3OhFddNSbddxtXQjKL3Gl+RO+2X3bMN0j+f
5DGhskgJfAyYonA0jIEJ3vMS0MFdbHy/hUbvUF//n144FGwt+WNVqb/nefLn+48+
LvnxFZ/B9Eh5OlJToA0bR1dYTnKQhX/ptdL79XPnP297A0lSW4Liflwoys7/TXM0
2kZHFgNc39oxjSWv4nzlVv4DpGvy5cRxEPemgacPIsBYU7u3c4+XvxLHyR7PGwIU
APEBn0kbw8lSbAcEw3brMWNbOEZ4rYZpC+DOV+R8gNwf5v60ddpH01+Ke6+ie6FH
+FKzHE4MsWGjvTyKeLo8R0IzRu/e19de28toWFbw1iBLZ3O4kECTB7BKOWz+0H8G
EY5PtXpME1tdNHDelut9G++b7DVIJ6YaWWbw4IQkUVVa6bKAp/zErZ/T+rVvvuU7
6cTOjmb3ZcaucUjomEzfpd/+uIOLgohsiaIiVB4NnaXgS+PC1BTYouAED8Ak7suI
ZA4sLyNK55aFhMggUoUtPAoFZjkOhElGeaWVQz981/P9Xgwx/4Ia/QHPvzFzdLHm
rsf+0g/ykib6PJm2Dfg/pUVicpncJEO6Om9guof1G0WpT43CuVFiY4KdFG7o9M7x
GX1fF+UZzK31gsbdaJprwQBQ/tMHkzViNfjz6cQihzFjGKKkBI02wa/+lDCik8t4
K68OOV5RuS+CT4I6KIQYFLt/vSxvYzQu8O8wmHqK7bthp8P5Lh1aN3L8eG3YzTc5
6ciYlEzASrpvDcFYVER3jwZvFB2ftLh1mF00IrGTOEyWFjUiPGS/m8X0N+/JClhi
PP4lh7hiOcwWcM/nVc4CdSZWWvEilRLWYRkU7rn0kJVXQIp/tTwJ0Y9zVnZiSkwq
8SJ+TDz1c0TL2Qp1daPExgPrkeRphq7VzVVQvJl6YzbZDIvK8BO7IiVfwSiaY59r
kTqg4ngOj4yLKmaUZKqC6jLz2iWWY/RIxWoBXNOWaWG4ugYACmstSGVWvkVo2Aut
JULOr6M5XSM4Qfj4RBYp/lkLV8b/AGeS6XMCpF8vO4qebcUReTzMZf6YZ8RfXjl2
X58nFuEYpVhT84fPC6aJR+/nbdIGCRMB47ld3HwUhfGJuwG7WNt7Yr/hDtqV73GF
OPiwwYLn4Lc8b7vK5kDIyZLVnubWamGO1dgNjLKxyddQoOiFmf56xl7pla4Anphg
R0gL+JPEMRh9syuE9djz8CA3Mw6itaS/avHT+mcigWML/Cdf3JLFtbaAplvR8zOX
OokkLxt0ZLajKtrMxSLlkexoA0I5dT1uzM0qoj+GbubZyUfsr8pIOmx6ZtGMqONT
llJBrppF7hwrYAijszkmnrj2/0Cq4O5xAtPJZTkcBsYdonQc80MmqQoOzf5CtlDG
3c0xo4I6Az04LXTc5vXh3h+CzMLSDZlIXQw/xeib7H1CTRZqxzgxSDX94j+4xo4l
nX3EaQkZy1u4z1pXzsKM2rUSjvw45OJmfh2FZEMq4zginGnAR1t7IzROm97dKJTf
lq0Uq24vCL+QJoPqg1ITeGYOsF8rf5lgsHN7GK74BJf4xHN8xdQjBeb0LSeUie/u
7qWKEAxO4x3qXBgqvtHd8e1RPRuxhK2uzpesj4ucXtB+yPdHETUEfWS20udvzFXF
C2oEZ3Eq5egNHunhwNV6gYZcgnabvg8tD63v5Q1eDO0K9prMeY5I31MLpx6IQTs/
qMLoxLnikYxNoDZWnOrtZo7VwWQVJkvip7I6R6a8X7GeWUsIQM3t6vf3kZZA0+O9
wb6cJhjQD0UDmaw/+6EcJ+zV0OlTQu9qAOzetOOQhavdzxM0e289mXe45luQgZfU
F9YRJwfZpRALOGEkEU50wwbfyOLVJo8NZx9OYt8JwCYLaGvW1I68/fNTHgUYX3h5
X/bziLUe2P6nO57jTpjHbYcQwfcacauABj/8B53Ad4ZcXHkEirTU6P9UcXWcD+R3
h4ULILFLULoocOYcJ5fsoIEzSmoA96pZBla3aSwSzhwoiSA1kvvORBS2gJFg4yg7
30dnm3aIHCzTx/lh2ZevnqmSOSMKLwHo0lyBanv5sEDa4zkByxV5MTVOA0GNb+6N
61tNEf8axB5pMoGKyqcBHtBg1Z91iAofO6e3CMzX1+oBNBI/uomiCLZwjJmkCXFM
5pKP6CmsipXftL803g9CwOxwbJb98z9Pey39KLGRg00EpKdwc3BvQYIfhbq3af/T
dcE1BJT2y8KOxAwSqx4QW+QyU7jgS0HXMN99aZfRkGHxYuZ+rQSDIprwCbvM9YBc
cuRo9gvq631O1uG2vu3nUeUjjofnO05CgGcD8fpBu7WsnWsi7njmtFC9Bsuh09/G
rvjGbdY8TdsoW1Y4sKfCR09ERstXI7/j8mLIqzI1aGRiVCalFsP6lBPZh1HeF8x4
h2o+fcGYIAfmCnV4nMMeG+V/vZasfv6eNx7FQQMf94v7bLr2Ag1jAymoyL5LWXYa
oPYx9puQMlOkK/y5YbXIZzcafzNoO1eN39VWTmYuOkJYm23mDTVZOH6fUxECuIC1
fCpqLgKiHsSXeietIJR8xcWyTFIuQwEIh7YkQGgxFVgRqLuOa4Sd1xEBs9dNdupj
fTiJSWfVURax2Mzsq6PIUqIsYAcGlFZZ1HoPVegrK5gdJUW0TkF8v3qo2+NV6bAP
iSDNQK9PoEkbnP8hcadOCTg5+grT2MDuoLJEQqnE59sNSw/hwRxLRe0y0RSbyWkF
dbIREmuSotGx2qcZGy3Tb4XXn9TyRrl6X4WUCKjgOEsFaleVxZM39hRK2YXPln80
GwBQO0QjJRi2GCVh8m8p0vu0QoCbzp6xsmFb0rLwsU36FZOiH/4UBHEE9NADn8Dz
hv9RTzkRUhk+FjAW8bycHy1O4o2jv0HjEZXFwN3rRrzt9PVYIhiZPYpawGp9CR2a
ADO7E7eZ+853fRlbh6U3cNNLMbBxTor/rz+/imu9cpI0j1Ang2gMfKSEapz+d4ug
HFkaeHPuxBnDvwIW7cgacN0W+vNcYzF2sHSGj0ny59bcRizUwfX1ZMxZVF9LC2Vv
u9dI6vTFRcCTOm9lVuMPUnbYYGWu/xiPiFkNgz4aEsFIgLKsXW+XYEpILiIBRkIT
ECxYd4FGNhdfULOw4KfDAD/pwv1UTmZB4w7NDYnPLTvMe93oC8QOghfzqnofM6vg
pnJnC9QqsqPowy9nC9mAb6toM5xpvZW26cCnZvalmgA5knvlOJifdyU1vvpHcWDh
fp+a02ldsWbu2t8ikFae75q+WjVj9BWA41onl+H2u+JycFpQnjUp4DzmGkpt4anG
wFYDoY7Tlrp5wAQgsYdCXiw2j41EzcN9Llkg623OBfINiVKygpBQjAeIUDfo+jXK
FF+hqhqcvN0ApUhJmV6CzKkYAPBZLnyTVe4e15EZr5K6YS+lXCvWof0m4ghriYHU
kTLpeDkQpLYQYaI1CMhpKS0LsODDdrCO5F1/d2hDqOR4W5Bg8qBXni8fLggBAgmj
uSpWytD0wSiUGhxGxCPe7lkuMs2no6XGm6UVFs/K2t5Cowzsfy0qjhVodqQXiy6i
CKp3EE/SUJAuHupU7u62wRA5uryoHu7Z3j7g3OhKU9s3zOK0IGY/4p/VH5k9+67d
NE6McngAOa/qfrzWczXrjHr74g9ItnpbyXfUEFJw4D0fL6VmyLHoCKMebDN+aTUe
XQ/XU3kOl/dJtAE5Hdd+eejn7vnPwCnrP19WPISLGN7pPogJhxLg5rLecmNAlKKF
XdP5J0dAD6j48vqEHm7qklsLqhKqPFyoABE1MTVZYtZmMjKNyIpszuvtvAau8Rci
/+H46ONLvp1loFlEbtKVOE+VgqLqNC5+bcpVYscL+Up4A5o3uCirOiq9ffMXTKJO
GSCLm9JWMYO/JRlmQcmPZ2P27Uh7eD+ClOR+ojYKaCU03tbQDjaMnNZ8X1i94rh9
4kT32kkdzBZ9WeaJ0RIANe091XzSImx7WJk01w1JAbosI8srgKoF302v0v8Grn+l
ZXfuMeGfn11slE4bD9QU1mCv3XK9+bHxM/aYUm00i48UMu1miydqH3ji2JJfkSPX
3DC+SHtdGtUNzd8geQ7D8i57wFUJFRcQ0aURdR7rUAx7J3vUa0FEkTXockmqyYxH
CoWk2D3KkKfx7J0KdSMuWleQbv6ks/7So3BZAsqPh3hM7zaB75lJHVhcMjpYqRmu
i8CNKBTmnJaT0hyDdaEEJa64a/n11KsdNd38IyEk8Rns331V2aIZsXPNTLGTXD9c
9son8mScd64CIe4fY5mqVarv7yuw6vSJHgmkdA+AJ2oEEn+j5mF72HtYflSNrYMw
dmnYj6bHUbrFLXuJSJtcAuAKKHZ9H7yTMxUs2FdJiBMDq+Hq8tdVmunJ42NapbTg
8euIJJ0dhAnoPucTLgHLsRQORVXBtKi8IOPvbt3NfiY3GRaLBDndp+ozY5RNVQfD
n3MmxoPJdJk8fiGhvNANAbOPYDvmIaeyiZTvCAnUcMfJBeW0Rs5pgThSV/+OPygs
Ag/YkSsyaSORMj7tL0e04YmMkqFsckpOIIdABfVPcP00i5/n14nO/lF8NzsfNQd8
gRPCB15vQpOY5UPjiQqApLAvTTgzQ3pGrIYJXyfecAZnaXNvrMHHDBDwpPDxJZRd
TI3itjtUaKAQn9wjOCT2hAOesuHpx246FleT1ZAVNu+JqsBDPPulaFyT/3azouUC
XOdehVE9tq3Cl4Ko0H01SC0RPxqYOqHBnews3PGwlHfuyihMmbAwvbRyM6jqFxbQ
WrSq2yemPii+CV1mJeC0DFgyfY/V+jb2idPBghlhOz/HJiMbqzUQyW5TRAvUNmcp
kg07pMgIOlNlF1IJTYGPbsT8uYJlEAfLGY1zT+ZLVZ6pLkSKF86EX7An2V48tsO2
40+7VswjyFBPqj+6ZB4PXuN1TiKcsjXPgU5PGE+Ko/VLN3QQCmPArsbuR0uB4d9c
s32eFWxxNgJ17rAJ7lCrZr21oJwhAQiFE8+Z7quo4+bntFd/lMxRQDBnbLdC9Xos
+YBDnCIkxbULKi4HCUqskeg6shnah8jS/I6aC6juFiTRelDhAUAEkd9qSmdJLDZh
ewDesm02BxUnKs9/+/JTnyr7PFw3Pyb09B96dNSMf/h9wmM6T2qC/vU8vPVoUQpk
uSOp2rrcSjkIoQahP6byGI2hzShgOx/677XvdXq8i+ZOe3VKN4ZntVAgOIzZEPV+
TSXp8LZyWav5jYmiNj0G/gMcG8kL1H4ELHq7Y6WKSVqQ2tEPSE5TYi8BY8UnrDD8
zdUgYIgVLTlCMguirfOqoze+t/euFOe/qnZaCHAYkuOUz4Yzz3/3qadS0itNhCY1
CKxniIoIrMSSoCwxKvldEkGQnPRjTsL2vnQDpw7Blr7rTze9gPOTCesP7mSuT7Cm
PmVbdPyg6DqY6gUTKB3KSn/QdmpQDFxEEqJKMe6W3trMZO5zuqHqfmLEljxuIWhA
X53oqzDPWvjqEhEqf19iPfS18iFiFbfJClRBFnZXxdGrixh4si6s16VgfJzDUxq9
de5gy0fUDLmkVQhlLDQxZ6hNmdrx+Udp78yMBvvaAjiWAxlqtngzjsc46XCKMGua
lOCYnM+Zx4kti2uxhs2lxM1fvxKDyTwdB6BsYUVL61Fk2qkikOuc4bOSWDTK20U8
jQ27z+gQVsH7x1O2Z//Z78bxu/8Y1/3a9cjwfzkVy5ZBxle0YTBdor6iHICvE9NO
PiHUW1Hvv4+VQCs4krQyByZKtLpQ0JBSfTNThoh8G6v+I4cutIaqMM2ZqwCAkSJN
9v8yr5+lFRvckuZqzgTanT893H/u9nR+iiGb9w6j9fK17K+Qy+xjQXfg1X5hlqNM
nlm2W2O3xmMNNFz+BYP3Ii+MgiQnszVrZPXKP0QtwEtP/0In9P8NXhkTcVyspMOl
jmTf9L77aQ696tinqAoXzKmxO5Ux97CRz0iAFjuVjYQ9K6lu+Gva5MW0hyK2lQIY
DThWCC1JbOXcpS+C72KY3TDSMDxJ+mlfe8VApp6WwiPpo6oDyulvQj56o1Atm3Jz
6lNj04K4L6oRO1qmgI42jHVaAJw1KTH5pcZAoe6nuL6UAvjIHg1HYxZg6IfurHu5
r+hKYaIPWCDuGvWxL5moqCN4GrrgpAZEmPMqqerDkbuRMWGTO9oVyLSRtOx6cLop
s7OxxJzrHHozCSnr5VZLgp9gh2GF63Tb9eflyEGaTfDFjSJl2VCiNA5nezyaKGAb
ykrfc2pDBwqH9+q3dQF5DMx342upt+PaUQZ3p/gMmYmgaJ3sYCGGCGpovC8Fjvxe
ZTLfL9F9PSh+pm23MDXYzKgBE5TWeIni8QCT1y6YrxILGQaD6PMcm7/fSJF9vzoE
N9OMXNRjL0Qz2dAyN5fDoTEjnvQvCjtyu4ge0SWJh9T22OfJYrQqsVnXyLw3L8si
Fa9B0mWA8FwbHXR3H73KnHpjS2dvd93s6b10QuG9adx4R4RbU/ojXmNSvf9aDTmh
hIDpR8BfXdNrksdasHrmGxq2G+obwlsoGL3ee2Zo2MAyN1JRCFNvHXWzgVLJzVBO
7dtpuJJDSik5zUkqIW4BRdCWxLb2KWOMFKsOpkoD/1GonT6GIHF3ZSvNAOzkUJRW
3te18k4zzqGVJVguwuyhyfk/4+p17YTYMX1o107OiZUms/jNF4qLehjkwnAJEfS5
EHiOJcCSM69T6TXz4YEVUpivZaSnzCzesirXVSzGg2+sJYzH8/9p3J9ZaYQnfEMk
wHwTB5m4fWSR9YIqhco8xU03jfOyNa2tRHq5o897TpQWvmlce2up4AMBpd9uAiEa
mhLoA0IBhZF3yCuwiyGSlAv7Yqe++5ObBgQAJs4gI1/JFZZGQ9/vMhonGghAhUi9
Ylrv3gTY2RQzUTIBIoi7isM7W/hX47Ua5vtWkbukMn56lwWCdlN/hQ9ShGHHwjlm
fjjEnxv+C+H7dneVjWvCQAjN/E2fbiuLHdSA/4cp1jpV1q2TH3XeEO7SRSdOUy29
9M4cjbZl2lLNZz8PyO6a9/QqU9ZDwBZXHKebMevNNr0Y3HDLTGr+kHcIwElXA5mX
OKZU+Uz1ImY0JO2l5QtYvTS1PlhF6A84F9iR0z6gig+iiTWo1nTyQGyRUxAhHE7/
IWw8jIG0Xa23mFbNULWFcSsamF3197c1dzXLFJI5BhoH0okHzmZYRTErLFEsWkeS
jpAaRux+Gt4FsVYLHLpkTyPz/F2ExPJEcQ12zZPVNjpBfigEnZBr8U4RqWsGD6gx
ZqReAey3lQJRjWZbVMBheAD3UQwg7MA3n4s5I4sGAzlm6VLkVInCs90EavnS6wQw
uksvFH/qPaKmDRBXYi1kXNSVY/h2GTynM+SOpLZc52WdVtt9X/dHN8u1IwZv9UpY
GoqlzbVdM4OWpT/7kAmuPzDb9UgpQpduwcL1Jplef8BFDIMT6Gsh/Aop61QcvY3G
xQ2MtsmIUropPd/fJdW62+cGUKxBVEbUJM9nARicc4wnz1Mz7uH+fSuFeObHpKnb
nqGdKqXXiLi6eLaOcOb3kIBpmt95JbrOqPfwZ3q4kw7/ydLFGCcfMNXNRQMgVHyu
XLSLPJa7WMTd5k77OSQ37YqbAgotJgIxaT2iP5nyT7bYCFQzHAclR+QdtiwAfTJr
IHt23Cx6RV2YbawHR2brPXC9qImblJaybqEnx3rTTlDa9JVQPeehL0+liqwByrXb
ex2KmAtKLqIlXzdFnwTBr15w2HYVOZfe9caro0c+PDRFJNOIIBPJUnA2qKd8yoDJ
9t2xJXSdglqw6IY/hd/HgggT+ISH5GAYidHgFGsf6Nhg50fg6V7n2C0bvZy+01gf
SLZTmgBq4c0ve5s4fw3QItDVBj1OaamIyqkD/FGhZmEu45mkLk95PFSXOopSrmgE
tAhOf9H3GplQg2Jl0wHi1mxI2ADo3yDA9rdVUfPR3lKpx4NSlsRo1GpB6o0JVVNS
rTBfTlT1BFfNdfZPUjDWj2Ea1JqC+hX0qoN/TGuPtnArKNW8IALyA30j/Xok46jZ
rs7B31/WjyuH+4CUO2sVCN6oVn9sBQS2/SsYF2vBYsn+8QczsNYTOonkXcBXQA2q
sBYYSF03e/i/fGQER5M8FTH/EoWlkwGm73jEFcV8yJ4MxyaxslmasudY7ZquCg3J
weQsQleX8W0uOpcnjmsXasXGwk1eYY6E/Y+7rFu4ayegJp2Rd7d91W31NplJRELz
zpyoF6eGOFQRks88V8hGM2fYHtJeYjoOj0dV54KbysqZNwmseJx5yKzANMGdSB6z
tmqJbrUVrUjjwr08+iaDOeXb6fJaEWoNd4j4s6TqRVrhjrnvTyQAehPr0DK7qeB0
AoyfQ/EVoxomLG8ZNvmAA6QpH41J26a/UV9wiyfak6RweAsIwHFP3hNPiT4ElxfU
byD/E5yTegD4FRFzZ/PUETSl4o/lnjKvRHuZpgNkaCpypmXmiPHjUGGCqlHuXB2G
fbN10jwOSKTTC4+QtW9mzUIPlb6GSw1Dr+8eANpZmU1wUjDQ8Nrh04+ZdcpmgQF1
uDw+upfPn9R8mrI6W80R2l6aUJZJd/l8Ii1udW5JANpGrBXPE55IXdTXh6d9WYQb
g22i5e+wf5BGdyC7wkLHTk3e0VVXUkvSe4lXfOTjIq+9mvjJ8VVUrssnb1V+yr/w
0oTzMBe4xahbf2LtOlQDKY3u/lx23ntfEgeLFefJX4OxCJvhzUNOeuLCRx/uvLWf
3AIxZA1fHujnzN9+106cY5AjqnVU07v0LqxoIjmB2I3ef5MaxIyFXMpkiLvJ0/fJ
27682Vd/pAZXI/zSuSjktG7A2ZvcM9VGZ4m+ND5QmVt4wymD7H5nenKLJgKGu07b
FaTKCYjbuvN2KxX9a2fRagBNa2Q2fN+pr08gRD4r5Y1VC1Wj+53whvPEpG7z51pb
oHFUt5h0RiKKUXCOTEEwMHDLPGh1PwLklYQWfdgKHpcHSH7gl4SIiYbyGvpghIeG
7Q9AG7HmxyQ3WCY0qmfmGbKuSb21K4o5vEvsnUVBcCXDQxgE/feBZFSYuWyy7RUa
+Q67KxVC5L9RGdXhoQON4d2Vquq/CKNlO5P/B33uUjcCcUq10j1qXXs2QRYkBjee
L8BMVLleJ1iRaC112/0clrhCNCrfUcN6Y7scQgENGco8F6AlBmSGWqF1k/RYMnbz
T9R41DtlvuciQkRGr95+sqbDrrfF72PF0vTs8XmTUftxwe2JoKUvl0pBMz/cKUoM
hzJqebSC5M/hTfJgScXtVl7uFueXA3pxccmdFjxq7X3LuYX7abFIVmHeZ1jcbS5c
FJoy3YzKhSzYtC9msoAXeaLJHDC1MZlloJHvm3tfBib0/NTYQSLctb+0o3z09H/n
62m3pMuNUsgvolbcW4ertNCErzy4E/XKrPlJoubIHLEH4ZzXq+NTTHk7H2DeIsvx
Bn8pr4uoR5RrUtMU2fTyMK6853Qe5nKqDXqriaCUFMlElWcSHT0miR9JHZ/TU8V7
fvv7whKAG8KLbBmGJ3hoIycSG8YxCw0gvuX1eJV6cfR7+ocpP4BBYUwc3yB7JnuS
pPWScgWpRmqBVKHbugmB3dE8BG9aIwQbcdYw2n4MzmsGM6rg8WU4sSW8zsnUhs1Q
GCmc4W4fFXTjbtyT7I/CpZrTKGDD3g0sMwY+zQR2PTSuMtW27eauRGPfaWZ0FeWq
w9mDGoyHVxYdQa+F+BtmheRMZHGP2iMCJWWJhmzvKtMJP1cSZYc2/xjxNaElOdmy
HJXBy7JU8QlS3HYTPaygKafbjov5sfCilC0niKLURa2fnNIaCtgOyCNrxLD8Undz
h6rpW+rsxsGfxYvenHnkQDTbTqLVKRtim8V7JufxThYuzQlXaxNeNFcanDTOO+gB
wezzRDNdYYU9uTYgY2tjzwdLLaqDN9zLHjHf82aPHGF/7UkDeAUrYCTNnExc2sCe
3V7q4bLTZeyPIio9klajMBJ8ZmqvK49olH3j4iWaGswSyfq6+2my7LvsMA85mC0q
BJ12jWRIMJAGyl619Vn4/ZxGYiXbFPy3JeI9pm+fPKqt57ivfHfK4LCrrCwBKU+j
SR9vFUkmQyQB5cIgxFp9mBMXn/dWW5iIySphW+T1D44TQip7k68NqE+cSBB1PkEL
NKfbS75peL1JX6YUb/UR1eacVIW+u9mT9nJELHkxEb/QCDH8c3EazWMME2NkUy9F
mjBST8792Bm4xL4k1S1YS9lW0N3pglF0c6RntDqXdNHR1Coc5h48KMF1TjrLhJNo
kjfK110ysC+vPRuw1XH75iqSwGTp6mV8zm3/Eo3EGjBfhnpcx5Jxr4ngGFKEqvUE
5TNXSqXpGIB4cHmpNYXIX9ZZNB8mPa013AXYXqhFjOAh2UsK2ApIeIu4Pmzehsun
oRyd5cA4eNU41oB27aZDtKI3jBXUlzUJPCmF0jI85Nz7pXZYHY0WKg6diWoF7Mnd
qh2NPeCR+sqWA1ls6Oa0gazVcDxjoEVKEeEoQ1p0TGnpbnmzAMTl/dWtfa1TMedb
Ofvh5LZCUkJmX3OVJHweg5Qj22I/1ndeO6DIx9wpHy52vGiL5R55lHzRCICOmm6i
1eK6mw5IaPZwu5NgUeDb9tX+aGhb9FCwaoRxDvd35qQFmyTsrjZ1W7h270XmHxGe
EOgC0pPL9GJRZabuvK3jlsEa8sxBIRl+V5Y357G+MOEh63lBOgEbJgXOlybabO7k
EQKvT/mEVY8CylofEjxBtQb13014Nv1o90/+eS2NsHMdADz2qm+Pgz1MUBAa8x7O
Oc1T6WTVx5xoxeH/AZgyyqmMPOf6THIDpjuDOWbRwhp4DUPaSKa9GkUV2y6jSlXK
x606Zqi7sgzPcT/LoPej/bGp65mJRHVr0HJNmKiL1NKOy5UrBY58/kI+JLDgXlaG
8he299JIPZqmUq/tCC7BLBFc8sAAEFPMIrR42JUvemrVycQkFdpdFyVZj3y4SfR5
sQL6TFALGUIwyCdq4RmBxG6Ph5EuGlmBb+jbWBWqwi46gImmT+6iy+oM/E0OjsfP
1WvLdc4waIdx49dXoioflNeDGzv5hW0+DYC8cVjU6xY9+vEPZIUNURUZJpMDzmZP
gz8FXNtMWls5ALmGMVA/P7qZr4M+pCZHlBHeSf+iPBEmo4X3FFmo8kgGcGNsJtSw
QOj1v/sy6UIN6difkqx45YgR4fBVGDre2yH7wES6CVT4VkFfs5wAWs0gJcetU6D6
N+etnUhMje0jhYgU5N5KOkFpbLdv+wlrl/RjR3uxF60hfmThuheOvSeOmPefxFkO
0+TIxqB2tQmJcN38mJgDqaVf04rye7MInKnmaxYRbI8Mc8mx4kHY8ZaoNrDgo4nI
KL1PRjDYGfLb1ByI8rIkOWA5xMY+uJhg1G8Zbv5qt1MLh7WXKlu7VUT4xC5jiV6c
KUljuo+51/HvApbLA22pcXPhDKzoUy28y5EoLSjLukDmNeSdUlQf2Eggwy6Ep6xH
muWvhpmXDiCRMaRco+GAAan+o/UfY9uMHbaDnC90Pfn4AwndYoP6gZbaCkZTbFmq
GIZ6W8dytp6mOGathYYfoedzXo7eG8UD3vee9NvHbCRVB4XMX4acslkgpUla3G34
7Ym3foqilfFTns+fJt0crcgiPyTgxLMYfxJxKBw3RU1iDA5B3QOLDSi50SOoqSLE
5Yqzyvvw3YApX383y+vXV4Tf614T1xkHKEcd0N2JLNsyF8RRnCMDr9b508Urr63N
nsJpKboMejix8M2/4lssNQ==
`protect end_protected
