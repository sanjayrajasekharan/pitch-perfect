-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KYBvcEPD+Xgy+jUHnkVuZC0w0UhhyMJDEgzBOu0xPwL1ak0AeEzTZH+lxJN3cBdP5fTXMieuBRrd
dILWOivzGCDKe/ZFYgrffmTLGqYeP/u9cjwcXRtITRJI5bq8KAlyvhbDCqN3XDYgVZ+9SXCwMZC0
3sJRyyZhIT6yvKEz516mpWiq56FL5PaLEZgTqAZVOihuYz6lQlN9Y2ByQV7ZecoBnyPYJyU+cEAQ
8uoE8GvrlcL4dQVR62bFSTxHj8Spt+W1PwTJRl43zQSNbiBUgHC35ucBeQ37ZagI02xQQfnvFcfr
Ttn1rcVD95ajnNVN1CrM0l7zD+LFBnr6k2m+FA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
OsEfpIxyBp00+74+JeJOqczqITH/ktvaT/Kp6L9uIf9sZ3bRSaF5JtPN5Ls6I2z8pIl1atY6clRM
S80w9XRPBrHD+s7O8hiBHdbmmYkYw4+ELru654Pe2FyNYxliDZdmjv27X1BOUfAG5z74A6kA+gNb
0Pvsuv2MJSlKhKhphg+SYIY9XbDwvo0odawPdDPeVnhbQedPC9qF2/lHDsoZ4rmodLxX+Q62OY4J
qtgdORMCWdxeyY7wg//O3Av8EPIDofHRwNv+IjNGFdAQLiW2iQ1PJuJdtJuqKiRGkShVUpxRK8Mp
CvNzSps6TjTPeGxfZ08yLx/f+tcJ1T9EbUMlgwCsUggaBBL++EYG2amUcIJYMSccdeGNUrtegbfg
cdXJaE4KuRB+UWEj9sT5JheitqpyZeymFT48FL78eJB0RXYHv8qGqB3uK5aWsMPG1FkoKLT1ubpI
V1sKPpmbnDdTCJNGB9rEIvmaLmiphIMY+yByCYJcsgbX0GyM8mGlHBqDH8/NZkts4MDIMXx/VkEj
JGGUWS/MmoawudfPG+ZKcUDtGVqdGXjdctJ545k0NiFnySWpVDe4mmVqzNf2vDikDRoIhYq9MYoT
DiL+V0XIAAHCUCDC6MupzSswYal9Pb29NAyTNfookzhf15iGURQi4+W7T1DNcTlDBcCJ/oAy0j3+
fE3bpg8AAllbPoUI4sosqaT8N8s6WEzJxpF9SkJCWayEw7keECLSCYg3XqZiDw8J43QYF+QEKOdf
0SP1ghVgqY/rGqY7AfMOLlLUk7NA78pA+LZioEFy+xfs5z4vATN0funOA0huS5oxotm0teD5xSPZ
FH3/iqSmmxQDrPN92tEnX1NjMgVoVzBhkDydO/5S7bWzGWBWiZXCV67V9l3uWQGICHK9TWH3OVPS
zoe2SAf212s5ZVbl6oW2zMbAkorOp0L5q0VdvFd3IBwTvlJmZqm50Zh28/Xm61v0rew9mHqmepxq
6MMA8+oYYs2B4Es02bmsvVZ8HKiNC3xK6iA9qyWgq2o7h6bPw+vdaYiirRSq8wC3P0YU7Yqa3fss
+e58ItA+lJl5sPi9+9xH4dcfHjYaPlPVVc7mfn62oSh/NoljkOHYf9Z9+hDoWFq1we8ATKE+fHoy
vp7KV6M855u4Poku7pZr547Qkc2hC2TG/fjf6BmymAnxTlCM5Lpwyq88pBxd/vPuMxLKsoMJbXOL
yS5gHfsCwOHnRcF8sBXfmo8pSe0LCnuj7ve8YO0yCk2EjaaJZn9V8kN5aLy9/R/BXvfsHJTsTe7Q
oFWvOEXSmATunpzGJ0+GqKQ0OjnYjhSF693u/hw9PNcaYL/QEVGLLu0291JYdAzJGiTgHSrphAQT
eiPghXYS9FKALNIO8G5qXKAZtAD+EzS+o2vL7H//yJOvg3ZRXQffPzrAhl3MhVYKzc9U/CFSghlR
hVRwxNmCJf+KhXg+4vhvRWxvvHr8YaaPK5Ea5WWVHyhWdSG9tnPAbbqtAfOgo7C5XuWEt+lKs+0C
CRFK/guU9dpxgSVbzVr9B+3IIvCgME46MEWMxeMlesQ3mkmmUQ0PoXHp+VRBk0LpAOCgxw/iUhjk
WdeBxM7/0Yo6XBR+a0PFNZj5kxp7rlR+WlmLGpuqD2BlVphs/c/PJxK3IUcvVWB2bV/EH7/1kf1R
iTjSGOiPVvSpAOO6FT1+tiWUYsHhYSvT4ZHzOJpsxVT/cSoDpZhH/7MW8lBGziRDDyKSZRPDk4rz
UpLYt+nPxuVeaD3KDGS13LtWEB3K0OboAIpeVhD/Ntg8y1QzHOteT9xBTHf7A7d6tluQ2bBtGjGJ
5B2WoMM0Yy5NQ3L0ZhohVk5FL/tg3s7H2/I8Bv+NhpVEmlegzuKTNgS5kEQOmY4W6s6ITivSABM/
Gslf7EmfJwG5QsNx5WZCtF8BtsDzRtb3koQ3ZttDtbE6b4FHB0W14Qt2XwTRMTzZMR9X4oxRfczq
wANBti+QjQ4Dpd0U0i/ehWtl5dIhvaG1gL6rZBPpNGqIojzAbEgdhl4xr8aSGVcbjXuoGSp3LetM
JtWr3JrXk7mIS4MzKq0h5LAH/hpdngTAd0S5PuVUAlPohuce3wGo2VSEFcfnRtnyLi6nFUfXm6Gs
TVjYAl0O+/AZR6xxWwyxWuwrKEV3je8y89dWVWDODTn2viXB+G1poSEpU6ftP9Gfa7avt0YHo9AC
zXmHv3GaiIzIl2V6JJJM2cnPPCxmA883s2bmGN9WtMptzsBmNfhceKQBQQlgdguuIfBfvW0hSpNh
KgzgzPSQwDI4pPgkXA4JCX4DqKyS1r3IZ+2Jm2t51FgbS8jPUqVMVnxtTxljyK0plhLEzYkHQsrL
Zxxrb/wnDaRNUgYVXWLAo9k3ZdbU+CQ9vYzrSCnynoFuSqRW9k9b9ZRDSEjsss0EHkRe9yPLtD/Z
Bo3DJ9hyzCswEgTWkZASNyEu+rIAOjfQtw2mTesdF+yYig7rgMZ4I4ITaH/Xn+3Dyk0OliNo7Zhd
89QvZbr8acIgdtP7LKHSlj8bGV1hjCerSNTN/MxXE5WiSs64dCN3Mq0zjtI2v1CSoLlei95X5+Ey
QB/aNVav8Hh0Xko16vDYi63pPOM+ckrJRaCvYFwXQ0UwDzq8OJpO1yv+jbrpEQTNxqOX1C4eLZbZ
kzWRy+zhIzy2sqClYtgwLziwblyoyMv3v66IFO7bMmLXfkdzursBxFQKe2rulkEVIhwVrXns4Z9/
pMFYfTDMLA3WlyBwRQW7wD7HKkqhYyZ4E3R2PjwFaKDUfdH0hq7qspGLx0Bs1ksE3x4aRKsE3Clm
tfaidhzJf1lLM4hJ8nkvVCq8oTmfPcFGrGzDPB7W4RByBK8dbAlVzs/1d6Yn9THPYn6BPIpE2wmD
aJdy/DWNxI+SEcPHl/2yKFhigzz7Al1bMVjssdssUhvEd21SwnXJ8RQf50G6pMeEqg3TXPVxbafF
LKzyEa9eK6hfX+4wonwqqU/Xthpu1eZA0BhwInnWUS/4LLmASHGD11McYFqz911UfPLxZoPaNnka
NEhIK7U9CcVC79mUsO/GVKUrw6yFegCi6PX/KI2sP5+hrtWmX1yEf6h70KdTLhCIOA5ETDTX79rl
P7oRTiqMuJxa5CwB05SdJlMA8EpKp9L7p9YLF/j0ozAB5xBZjUtzSSde2Rnt6/e2DDemmEHNlcwi
AqOXlaW7ckZfxTkbB47IgzCQ4dqKQ2gPVI3LuKj4bcXGmeyK4bgcTjChIfDke4Lw7uU0sJMgOsMS
6TDpl13rBWqGQSzx2EGGLooHsNFg9WbFW+tJ6+2TGH8UNjpFSNI2/Zk2bot92dm6dQe4dwStgLvh
1ham2VCFBMOVOsLAT0X+J61Bv8h9H+LXeGxUGRb0zoawGpDyFtAtf5KDyN+cQmD1slittninO4Xd
JwtrNjEve20VMTllb6Rqtxn3BZogLDa5sJgX0LDAOgOl3Heu1IQV/j4e2HooHBjrDOxxYwlvmoHj
NiSTbB5oM0/N9kLcwGNSJGObCA2D6d60iLnEFedt3IdwBbKmAMa4Xa4ItZJH/+jchEG1XIEzDHbI
n6ciB8sj9xfZnYdq7qvQuBogP9iRjnZ1yoBXv/PyTBBdq+n6UtXFc6Ick1yJTUFycg9cdoILBzgv
Mdb3rrLWTc+n2BW3lUZDUv3E60QXh+Egx6HDqcp+CJxBjVYzXmyGs350jNLS6j2R69/m7ryDV/2G
oBgpE+q3jGwyhZQiM4ulqRa5KgACidRiVceLTv4lz4CvEF6dfHMQBOCWXk6Z6zhdLGO2xX4w8lu2
EhLndHYeKVhW0DXDkjtRAB1fG7+o/8nVSrS9CDDapJvLWRiMzG17okiwQ0no1OJUKVnl9nOC3TNc
N/N5D9NZoVwSSPVqQkt13tl/GYkp9mBbkNKn+uQN4UYBUTm3cs4ImZP72+mnxtLR6l+n/pHZhh6j
pS3xGLpJOrEAErtJtR7EYHE+QJeDfHKGGnhSzX9MxqcW9o+gfefXYcDpxTZsPfcV9BsYCAvBijnW
rFyF/joNZRnzwFbZzHyA/9qnowbTTO3QNP4o7MiErfKy353xJyeKAyxl2IHGdLGBZmSmO14drZoE
y5WVfSfWFTF/Vush5MV5OvpAwyjXJzGrwnQzUhffA9+EGS0EpWcXDIpFwX9crGO+IMdEDZhE7tWN
0CDXRAi2PK2bVC4GMRDK31iJhdj2oi62+twLuVxVzpZXz+8BoLGVtcLiJVBtD1kTy8VY0z/G0t7K
BjqG4b4N2tZB8Ze8d7LqGALJX5pyGfLxJpMHdR3zjjxEJ5zK0dixLMoW90cv2W02e4MZwjUrJxVE
AntCYwoCQdl3LEQXY06/XIS6LuoHxPlZZeEg9s7y4rZHxY/qOWuWQ+VLKvExJ3Mrt90GUumd/fLm
VkUkhN6HjGzeuu1wMYjrcm0iioIkq4k047AtLq8FK8HBl1lo2axaBTDkOOfDWkaKXHS3O15s7nMM
HhCpkhY2NsLE2qtk9suoaQkPPN04MfmmWJgCVrBWN+GnH5XNnzdAKI9rT6BC+7pRRF9RWjh+/qE+
rpOjtf15tm7C6OB4L6mp2gqDcdOhbNPeE+y/lnxkihTfFIq9f1AtOUkvIuXJmYztikJAxayfj3pt
qTv4JzIQKSInhEMNMoHcdty34tc2UUMZd7LlpBVq74PxqsngpmhUQRkD2FUUFS13Jni32FMbYB5l
DHSKqOIVXTtYt6TbzffBinH/ZUD4tKfh5lmQSj08ePPTBmFvRTzCaRKti2UTZ8qae5S733Mkdbdp
3M5rb+3/loC3Ws5iydNyQgcdq4A/kQwi6VnPx0GVobsL8/xdc6Mm45NyjEcPeV2XmRowJtpzoea5
pfMKH7a3lJ6MIr7skNVzcMHObV4A4oTLPGd12hxm/w3HA0yKj5QQUX2DRFkgTdrWVoBdoeHRpGYH
/b4fPrgP37xrbKb2hFm4XPxIEeE7d1PdzEv8t+CwgDl5ijMo/NxwhHO2BNrUcXvGrg6062LI4w/B
sz2tQKfWXv7DeoqLv33t/5NU6su2evRbTfOSo1GklgXmGjl/l4wHGL2Li7uYwLLaT67D07VZTPic
QQqCRmh9EDDroNLYWlPpD80xtIjvT55S2Mb0hfSA2iynFDCtd6Ewsnj2iVrHlQQhEJvwET9ztHHq
4W9Lt097Xj3wwejQK8BfPyefmvPmua0hzHX0cAkE46o6ZbXHlIAD3Vf0MyjpREvflajQbK0KZsc1
oYAUSsgWZOw489ZSYo/ivf+x+UxpJSqe6HiHyasXXp0G94AorrBCLiM3siv+J33eX5xmuBay60Yx
Z+rZA9BUqfI+gPWgdf/VhVW20c54CFi2bOKESoYb2lfukb7FQlsw+A/wZks4XwG1rjxxb8Qo82hM
iGqFT5PKarE5+GlYnK5WVT2cDMdDMUJpabO6w8P6GNSG5cS2uajRjc//D3VUq63sbUec6YXc3jk9
fP9vog2l2U32POPqKbyCBOE0q/RwGR7IxLzNgijapzenZ0CguHcCEC5R9ypoCBRKf15Ij0oH/BuP
MVVUHRqIQqDOiMsIeJxJOx4Vke1dSZlRhk/Pfw73ZfWzwXyGsWUfJixu5Mswk+1lWcdgbs9NEijD
FU7Mexq1esPelw1jkQEpQFf4pHgSasAJUXjZ8zOC+saaRu/uEIX/V9gH0mrXwFo9bIXj7oFwZVf/
4HGodSAhNbVjrD/Xazq2c3wQ5/H3hdc8f/gW0S8CPjzZEl7UAgbvWYPMPkwxv8E2wVaCUp+PBIy+
5V41q/zHZWNOZJYlWVp3Xw4VOTiCttpxJaU+9Pa4MkarxsEk/IIFtskoXqGtCMliJdXR1T0ix76q
gOTmatTzWzdSad0z17ILqvrDSKNiEJl+noFcLuAZ3QynQlZZF4NOapCRv8i92v4rBEPuCrfkaPPq
2Mlx4/+kNlVtmjD6A6cQzI5wdB7IbVsGlok0PzdFqLG9eh0pedSrnOy2w4lbKOB2mGeR49hJbnKy
J3x4c1nYznGqusO8lJZKax9g4x9Vksg8PeC3DHWeo50IXM5qLtjXpLyp/1EBdW0Yc+/+w8Kms++u
WfHwLW6EGfpblzkxR7+ZQdbC4ucu8KCr/WTDktHGHFbT+anSup3gGl2kcrsUw81YA9qU9lNudhAl
3+aKZW9jNBdybzUmuCER3xD9UIAFjBc7+3e3zexSlsFLanR7JDHXLlxHxvfuzj1zYsgG6Txr0w==
`protect end_protected
