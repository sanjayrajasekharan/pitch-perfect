-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
h3Rwz3CjBbtuDlMUKfUs7zUF98S8VmtNU1MR9HKTmnjyDbq4v9sNysAYIJfI9cAG3T34GnSMHyol
N+rkZILZ4x/tbMrKcgXp7rNNpv902f+bsrYXa1uqz9HdJq90/nVjSZPBciFwleVZSuSMaS9+kLNN
V9zXp+ez7Vb4tBbcEfNBw04iendG4zW0yDc5s4ilzTZuhD+j2YVTy6jQDZQuJC8UuLoOIG3QEZsP
oxPNAKlmY+GXpTV96/TfUoGuiaAVnbV785PQk/kPNR7ztO3usHFU+Z/Q+d2MEUSKOVOrh1y+ImKM
RLeEgbg+XvMIxRG5HQ3JvgWZOXkgibG+4EEaRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23392)
`protect data_block
Rl7Z7muXBQN2PkpHcdnwyeCqySSADSs7JvoVm7/T6/AkNCBGroarkSfwRW5jzdDrHLlPmhYBJFXu
e7Pcr4UVuCsp4/vQ2hp/vPCrNRF092AdgrMZlw2AJS7WGmYWRnT6motXNzyJgAyy10gnVHJdQtTA
+U0ai8EH5VwamCIuua1sKqj5mP4jFF5EqBKwyVj7Gz+2WRBXwZsYaZzlpMuWIOOsHT6lzuoWlIzw
zW0JleveGaiWP4INJDLTY/rMRzNRXRBcPN5sEEJszS4/Z9oiXtpfk/fMW5L/+QcjqzozqER6S9bi
pofMaqbFcGhQ4rgY2d+3W4kFguini6IZj4JOa/eRJoXfWq4Cd1DTcEOTAUNultNoJ40fQNlPRESM
pVCJpw0g+5JkpXIMn1WTDGv/ocYchg7l0shNAh7WySWzDZJI6nE5TE1rUanjH+bcFTR4/O3LLjHa
Q+Oa54y/EVMxwDMSyYx1JFXtDaVDM6LbrqIJItsr/HwPj+LebJGdvh7xZ+r5sDM01C42hfv9k1aI
+QoflcDtdSTIzjYHGZ0MNVT2fkBI4hSS4YTqyaqN8EEzlYTAakxqTd1weqJTMHJO/qk3ZgZ2+KMm
HLYZNQa0v5W7xHgevgWyICMWWRSRl/rq+C0BNsHFzYjlA28HPAnpohwbgwK9WMSTAu0OHaxrfFIU
Ae/PFR/dG0tk81htK2fE40Pr6rhIOuMeHxdUGA+u2gYsZEa7ti6JrUVGqUX1IpmDaQ80K4m7LzRm
KLCuiNMigNSAf5WNicTq+s1JtZ/ey5PHpuHyc0dENZ7eeq5BQAZryw1scp9DiqTTuT+3uyg+ScPF
1RFRIMWfocfIIas3T5yU/46pJbsOpBNu38kRhZz7cxLmk7QL0lwou086RUf+i2y8IazPlHLbwaIr
VdHx/G4nhsW9+jXK28eUDevmR6yn/3Tb3U0X0xaYqstfhKkK4mPZ+XbtS7OxQRCwAXDEYrixs3jJ
CkKPPs6DVyilKeOOKGJG0C25SbRBWLBoRJpmJmh5igGPamczqV52BNsXWavSxRjWhULMYL1FOn3L
yk+sVKD2mBhuT2tsllg0snT1Gyhz7WOjtbh9333ZuOlYQvyxPZI2kOIb7otGtxM5INo5mJI9ATDy
n1rg4AJYmDeeAwJsYsfPEi2dUy6EczgLRYq8ZklLwdelWxe9NUcQyXOUHThahNQ+4FdovNQnA3v8
RWzDdQmu7JXYTgv3derOFeCtD1BFrebKkeM9KUpqJDQR9JkqhryVuTkDsTnH0zc4SWo6A/wioMgt
q70768Ruau+k6EftywHbHJLW7/oCy+YZnMJ9Cpz7I1xQYqkAVQmg5D1aVwSdcf3mPYSrURqSzxkN
Tc/yFaEQeG5fA9BXEj8Kd6dM1g1uN78tClycmXYR+YDqczuAFztNLq51SPHKQqqhHx1LpsehgcHq
uOKT0aV8HN+JubgfyNkykmfn6uE49b6hTYMv67ufq9F2bjGtxYvEnvANYtSY0BNNQP/331gTNwgB
2a9gmRst6xKrsCBXgIghNRAxdAu/K+WS2MFY9IJbQZGePBXOCmms0LCpXoHzxOGv4VebvWflW0wy
EE7UAimKqru75hycwLqffWJ8gER6sXQ0luOL+jECL2f84uaI0UfKmSxyGknV/i8fF5+fwxMuLiBA
axSiVmohZlKko5jVeWfDilm1DZHLTvrOLZ1nlAyAFQ7dH6KHRHAxwRDo/oyx7bwe55Xen4gm3GGm
zEZEb9uvYKFIebpMMk+Z2arHMkdb2Jisr4hblQbtKJGy2cRI6Kz//1XNHcsKpWYpLUrssuslV+MP
2MovzBqHn/9KcAntDEQJXkHXiDTw/AZvgHzA3M6+4XfLr1Q2gzOfyZsSah2sKLqRizoJJNOT95Ak
epa9WkUxXa4XC5JELzp+9yHI8D74r9+xR0jM62QDVfF424P84n1pprB5A8LrW1t/fVPzMi/oVE/0
wPCWHjYm/HU6TPOFasYSOdB//ijNDNHXLI8fQt+MqUjCpt5RAktOUS5M0fVUJWBkhgD3wW0X/kEs
olUE3MCBcRADjwyIFeQZohnbuwVGFVrmqNcPctyLDbGpscDurT2yijOm75ujZTRzNfLH0tBj4QMU
cL2nWANaiTrWgclMc7Xe/2JNgZq0RPe1uuGumI6EJ12su2UUaLzhS1IamQrareM9r21T6woxoqgK
0dPcaSHbbAMjkbytANDr2yBceWrquwyQHa7Nt9rP8bVviyWICUvUdsz1cl3csLd0rpfaXmRfu6eo
c3uMjZoxJJaWGLs1MakAJyXJnOiFFZGP5lpm3oXuTq4xWzxuveYD0CYGpauX0oeqwY3T1sawb1Ic
PGHHUS1B/Z+Mbap899y+7Px9htC88uqbizzdvLuJdfV2sIVM2JTJX+T7H+kQJLrXRJH9BcMFWNtD
TSomhE8Pohed8LLkZqWpqZsSQODA4xTDeubiZCq/UJi1abFfZr+nu+F9YIi0/bRSSoFA3yUMgTfz
bp2coUFQ4ylTYluDORjDkRB+fMXcScuFgB3anOf5krheiF0nU0P4lLQ3H/xT8yQLs8o9/1l8f03e
pElkj/pJsvd2xPrhr4PfEkWdwv0Y4uw5oZumV4BfMMLnScEpAP0/2ILTh0Igm8DYOb3IiZXISUxp
uD14AozLPop0S2UElVCueTHtOD0ovFwTNL7rBBeSzYHvmC01AemSPyVbxZHfVXbsxeFVbv+52rOE
CWkiXJSyMl/OqLhAu9IW0+c8zlzr9/mx3jwUEZA5m+io3zzeQw+wt3b5fIV6zJBJ4B6nrysSzDny
QTuOorm3SeSRaC6nls6agnXgzkfk8M14wb73P3boLrxPQYvKHe6XR4LgThrp9GJBjXp+rofmweoS
rxZgpmcn/8nxAO8MUoxAZFErjidVPVJxazmRKfuvQ1YCXYoTuBFDIj9aluex0SFbjJ2Ocbn6CyH9
37yfaoPhwLns0cXIrx+U3mG7OvoiIVxhVMftGE9w4UqOxDBA1bYwv6bZsyA65PI4vgRkeMkn+Tm+
ENu05RsSvGISiK48Bs7qFgxaqOr0x+rwHusVTN59u1GzcaKO/mFNjAJPjEmS2kJX0t5mevfDjuw+
4N6ZWKVUt/0dDChDea34CCrXGK7YT1vRFweaF9z1Yo46r952iFGVOXTJKsBWD40ut4ehSE/Itnsk
xmwFgCHcEfu9Ay9Yl7sDtAzk8AaMj8Hr1Y9vWOUxaK/KogW/MtluBf9m5OXwdgQ39PqeMc/rKY8o
cT8oIdHfIK2+7xPYpH1ppfq+MWKJptUJFuDY2I4xsV/S+rA54jDPCiA7FCgSOeot/Ph8nFMzfdM1
Pv7bQnrWW/RTf3T4aMFQELgSBNaTqYuuzytwby3BgPtGXosx1pruliTpTGuvk8CHodzkmQQYE4th
sKZAZhOyTsnCYZG91iIqkNlX/+n/2Ki8B3Vn+pXlh0fv1KREoW2exGOwzk/Ub5Yemqw8r+JQl1fu
CmkZJP7ODGC2BvNbrDJSj9Vk7eCzYIu6ST/96rLxsc3o87IcGNa4890UJpIw2sH+sfSeeRmfzf8o
hnF20VE58DQccSgviy5BTsHl6dNv6OL34wp9IaqWxrP6a2aaKCB+pX2MF7aH9d6FOUfTqHv3x6if
l/J5hjdQ7AWAGun7gNBaZuiozpC4Zhpiv0GRYdeGZ1eo5LHUI9Wq+wT4HK92FwIBXNHy09AQ7wpL
iCHZ2/0JOCnsTktWpdRicS5rs9XxNXfNk0LZooGdkt/GX4i9z7CO8davOO1ja3Tl30VvcT8AC0C9
E4pd5t2E97oQk07maw5vU/veeBAM6FeZ6RYsyi6xPPiGFyvexaCBc+27Y9fWnSgflJn020RC5bTY
szBuI8vADNdbLc/8aQvBEg0TELui8qKkqFO9QQEXtEFpSsjJmjKK6mKnsf0RBsrIznWL7zqgsLwQ
TqZrRYcBQmkartBBQBL1r1u0uo0OamGXTLpdh/kS+QBvblq2VxlpowR5vWstG20MCUuHYvF2j0y9
SiOehZaaWbUudEQVTeqTFidE+h82sqP9k1kPfZsHY7yG4kR0FceDnwLbDIEKcunOBwTrjrrKaruy
VHeR5c+cHe7m54O3646duZ9mnrny0N9/DN+ggcavsTGXTZSVdlOAcUmM2ruIlAfyvtGlhpKQqvex
7UrPTxc0U00h0IpsyQ6LwzF6P85lv5V1iUApIUEIkIKUO55J4xRy3tsIOqcXMSQTspt0hpuVs3nM
IDHaRxbsS8dMZArwz/VGmi5BSJppoCIs2D6zZqjuWnCTBgO0MejXjXY/crykTJ0Nw1v8ZX69in8O
xjea06LW8B0so+E4WPokxwAxSimGvPV4OTG7mFdTQdQhpWdEwdML1MI05tlTi8UwKIExIcRe/nrn
WQ4OIS+zS+QHx+CgXlgI6Nh4bkpkT8aUq+0WLKdygg4WIQP2B5AQEvCJfue3t7KzsSgbxlDUK0LE
EYMU7FnN1XkoFHB05pT/tT0OAzr14NRwOXSnvY/3Kix9EwnAakUOLqB1PnPADglgsHdK9pA3lJOQ
5YI2QOerV+5DPhNYaOZaAezPhgrJCFJR7lxRAJcB45KqdQi2989LCIPKalLo6+u+kpLP49+xtDA8
mSNbwDnKVRDqrDVarLVhMj43u2Jx22havJ6j9cercDXwCZH0ekHpr9ne5vfcUwkKh/d8oKt/WfMu
qeibnQVDph9dVM6l5iykOBpFhc7tFS6I3v63oRSLc1QDy9HjJ0XPkIMoh1KfCaFCmVp7R2yFdTLY
2J4O2tJc16Pe3xKA2QtOkcD4YrW3ZQ4Cnpe2C7Buue9jo5MXmfv2kJ7fzxNn+Iey7XZ/kA+U0B1t
ar6U9uF+sC3HpgPK6BTBZylVg8uQoI3jHEHYz4xX2PLRzpBpcxpnoEsJqHPehZ3MQZiuxx0Uc6+m
tpDfmisVWWd+5WV0P4sXsiZcMSrxwiHJE2r4FaZa+1ZjzCVxhJyDJywLYSUlI26D7sWGLFIkjFWt
TS+EtD4Y7oEHpsZ/1/JXhhO9UhzqmS9Uif0C/gIWqoj1YNvih9Gs+FLD3S16ule9k/RvnMuvMfuH
cYhbkAbhMuKx1D7rYZjMZxLEAsXKZO9WD6BplbViX2Bv+G6wsqEXvNr/7D9HSYfRn3S2Q9WfYIqK
WelPO4KjPya5E55whkFCNJ9Wr1ZyoV01Dh2l9NhPyNSz3rGGKV3EfpBpAamM/HGiXLjvp5UdonZA
Wyl9uUYoJPKci6LQjD5xhUGwjAr4O/lmMRSac6GM24ZmdJM/KLHBTTry5BQSRWx3b53dPG3etmcu
qE54THYeTMbSoWsQsuSfzVHPPh3/ZG3sdSVi2O8AbRX2WNEmRGOfEJzKP5XbjmZYzgDngFBsyEzY
rTAWcRPNrKWXbLlhjrdQ0sNlOpNZntYsYiEmKldhkrrfIdW6CMusRGqXXaOb/rHm4klFJqAmA9F+
k7AwZ0hBs2qxtRXy2ldDsTJ1Jm7evD1AFtbqWjHYu/kQL2OznbVUBgvPiJQ+ICtmjfStbJAhrWoY
jMcackr2qf0AbMVsrHDOqzjtjlZ7BQa06c907c++vojKMhjbuCzkBF4FoA3Nwzz/dDI8Ac+8Tpqt
L679J4CpXfyyAMsIMWdKPSB++7PU1QZtvLyyZyim4aAYqOFny+OeZKdUFozL46q099IGwBaTDkTZ
tvbmtnk7KJi7MWxbsmEREHNAPvwtcCvYFeglRzZnnNUd0A667lz4HoPmfHdavUa2IVrXnd0XgeV5
A2Yl0un6owfzCSyf5RxfNR64yUgLlIcETkQn0Mqlg0nbK8hvR63tH7iafKFsgBizXmGZ4kv9K6i5
KwLxVIQv0HauZ6D1lt94MBoVOaO5M5QP9XGUXtu2UZJspgJApJskpPFgSIC1fvCYUsj88vUsdAB2
Un7rtZ6RwVyOZ2YKryb15TGM2KxR52RA8pAXr81jQIpVaH7bKh7dJOxTs4fHFddIvFReh+s7rst8
eV1lyHAvKJCa0D91C2Ed8deBoKqJiqnJYRzoSQUo5FXeS+YEWtF0dtn9Sfk2abS2tFJuP3qr+CEc
c0jhAys2onS7gQg8pjfyKrgO8/zw+xSR2ELSNYVRw9FfE+IXoUQsoTV7BpP+9VVmKBMsM9ZBFsrt
61BIRYnFgqSa8C7iJGjZkJXT7EYSod/2SiSo/uaqG2ZCgpI2yAfGIyUxvyNv0cvPLy7001uEhPAO
JO8adJhAXs1qKIGeFefAAxJZF9YiRsvb14VK94mG0wjLRQcEo7GHeMs1ohix1mpuMxBYGoPZRDTu
TkTGwq/yVkI3xexFSMyTyht6uf3IJ89ZRVo/ijWHXCSluuVr6UOW9gMasCprb3pSXXbJvRLPWkfQ
C/ok95fVQy8JKgPBg6AWHDcGGFs6WXUMCbGXkQBO5ASVhBf+ZsUkI1E6WhukaZ/6cFVhnEonBHML
XqAaul3ngdUrtRxv1iaa1zH6e+yR+zT/hoiApVKUZ994EeSYeybSkmNMmFLfJ4sjJ1PcDnhxeoIa
GYu+037tD8FP82MMhQDzu6LZiqzD7gPiBQVYbxKNQ/YaGOfoaqcrQO+O4urozbFJ7UBpgZSE//1A
/kkA/XmZQUmN8mD0Pp/DlXyqrWoyXnU4mq1/YDMxoxDmsKQTam8mldYPoxkpt/D1J4digC8p+FBI
I0BtGFlrCMJeq0bvPorQjeZJV4EQyn0dCg8AMrv23KTHjMGJDoDsz/Wc9vZN9/A9hVgwyouIy07K
3VEF67RHh9thrgSraXjJWI84nbHZ/YMN+d3ttEc5jFJ2QTXccpG6S5Ck+rD+tDyozEnk4/9kLi5n
N40eghWt5U+NkwMD6jk9DVpjFOWbvbYHt3oivWA3U+K30XfHXzMOcvy2Z3asW+A0BBPvaTsPIYc8
AHPHwYz+87NqN5w1fV1XtF/wFQ3q8UNKvC0jD87Q5PYcY6YEPaRQzXnU4zJJTU38WNULvdKmxycc
UoWG0qtPco2T1WlCzxuNaqmlZwwNn9kh7ZbeDpM4YrOmK5I50oqXE/D8hxEHyX9HpEQv9FaooSR+
GC9OTzmMI331+MRpO7lf5mwdEKa4W7/0VcRiQcJbYC8gaScVSICA/eBGfG14Yr/dOrwgdxPYvdTj
D2HseUlctYWMTUrCgQgpSd8SMEqXxrPqPvuRPG43m1OBZ9//oEdaAcI4wyDPw90/FMS1D8de3RDb
V2rCJvOZIsieAZZIRLaJb6HnQovREPcZDSzVUczzfurhWACZ31ScVsslvXSyiCTHms47Gpqpl+Ma
ZcMb6tRKy8scTjsAQqyYIgyUvGLwcNnxqbCjpCenQJxSCY9pAZGXEBWSyps/q1U27AwuImxGHA0d
kwueOab6Mn+/xLT6j3vjQxjTq38XaKEk3uREQDqz4Yf47ZTjRdi5BBMKFpvtAZE+BP+LDgVe+LFE
FfMbs1BSYHizmjzco24ZhdTAkZa1K9ovIa3YssoXtym3sQOZHRMhXw5/VqXnicBcjUhnsGtO3/2r
Iz21jcE4y5+q8oMa3erEncqUUemLWarT8cX5EHC7c3my+u0AAuCackkL940E4vQOl4Hiz5aO3a91
76vUnwrBaFntuyLY3mNyfzNWMc8vCf6Kmz+KdydGnfm2mAhu8xMDYNXO0w01KqQwEzpgvijzoExS
hCDz3EoEbUw68BWJDhyehHH2ogjgXcef9BDjnrS6AsjS5wihL1Zp5H2qgE/VOd3bsBI8JFK6/wQn
yeX9jes8Hw4/bYfGB9KOloLbXaPw/nHy1d99k9kBV9CCkVVvX0L0LtzRzTEAJbWrxsA+SibsFnLZ
vYeQ+P2+dgH2UQo/OA9DrVAGDCHcnYOTqRbri5QmQ8mqiZm8Tji4DYuFuHG1Tue+xTH0RWpkpbAs
AdxxLXaYfBHunuc+UrWdpvS0rKWWVgf+0jVAN6yieBKeplH7z5H2DyLZH7QMwREZIZeslzqU0ilo
mPF2/tffndReT3iOPSoWG379bxkmaJuyLQH7ThJwcexUOB1GKseEZbMZ/xnGS3tPPlBnhWujt+r4
vqDhmIDdjRR+kRjJO9ohxuVvXoSlvOpEUUR35kRaIKfh9NORcuP00BAlT8e4QaJPA8itQhyvLOeS
xcQAgp6ykOMOzqupgdaLhfEQHQZgz+CtnIicwkzLOakMO5uOLlPBfsFCLCN6GcGvTK01ZKCFudDm
56e0T0gn29BCvaHZuruBduB9MIA/PfgJCm01Na+uZuwVLii9hys7TlyfkXoO/4KlvCJoOtgmif2F
Ndg0VTAH5rMgOu2sN4MHkGdm7vGvuCzwhDMLGJ32MV7a+VH66BY2Yf4IQcmTeCKw92pDy/AzcxGX
7Vmma2Yv7k3+7cuYdHjgWJ7gXUJsiDtWWt4arHrD3rF09lzZkGRrZ1A93swhIcVHiG9TAUhspzxL
vnuv8CR5mc7FFOdA/WfEBzCXh2YgNrKShXEJiXaj2mt96r+73BfR0mDLqNgHcpeUrkj0Brcw/Wfw
FwHo2DsmtkT9nNHB0QzMkI6Wo8fSlb94lL1c0umW3Zabm544iFqhiubstdqtvwwmYBx/H8j+DAlb
Su1ur0DvxF1lqkiP6gjdKGL01O0KKGuBl7Ys6olz04njS7XTaBWruNpEqQcy8ygQ0ob2cTaJhTpx
XZVIOHBDWJIwDr29fk6z07AGB0dc8XDBiV/mg74oYoa0jrrJESbZecfP499yuZ+BLUh2CPlP8cuF
St0il9hhaMh7LLkKTJrLUG1GqVC+bUWLOlyMveB4m/nD84tifKLkIfizfeOKM+fLw3oFRggqfqGE
LeQhwpmvCnQnsOhxOiEsAbPO1CuRTp9CoeGA2cQYGDjHCUSlHgP9JwP3hzuiQnhrOx2VUCl6ws/y
v95JEDn3S7ilITWEarfK6AwGKZhldRMFYqePMsZDqV6J9/fIkgMsE8FMbdIBh6SHQ3OctMp2DceD
rHrsFkzxegcUwJsY8J4/kJzr8js50P/tsumN/w696PuGCJSUUsuJ1B5zqBMgF8rNZlZLWSFUvra5
hUUN+BySPyWI6qFUApt0sz4PGOFGjsNT3DD9Zl1kWudoTXr8F464gZH1oXqPljnZXSJqjfV6bzcc
k7dBJlRzevsQYGtumjHNe2vt0ps1WhpF+v4fCK7YuuOGy5KROP9uXLXRb4jUXxtTlTpp2OYVZAWz
VulsnGKeHwOvWQ9ncdfGF2AttMD0F+6R+hoaWpyvKMmz4AxAFT2wVgl6G8wuHwq6Slm9e5zEARg7
LCDVrdePDPzWYBm728EvNsKl6+JtSGYksIOPIbflvtazLPIrKI/N2RSpgdibNl+HihEDjPlnXTKt
d3YWZ1RwM1xb2M4JvB3LRpsEXgXxGQhASUkrNELqXPxv8xBQOHoGCN1oCxWa94vd7qDJ7J5NHc66
NVnxEcVehqDHHvZW+LaXKPViGQZAo5pZM/jYXuV8JySJNU8GZ6B4aIXV+Ra3JGxaCXM1rka4Dt4a
740mUs2r6dhp9D9ylXpHCn3eH3IRJ2oNWBKjr4t7LQVjVlRqDFrX166zBZbmtSTQN0aiPcnRe0hs
ehaiifpgiGtkn91F3hyrlnUuPxJgfoSvawWPMotL4JMOFLC0PYTWJr1sgUvftgxmtt6sm8ldI7fd
BuVCMFyVYNtqOdk/TPt3t7Ps64Qzaf0OfBtzSrAvLHzE67ChAlus/Wc2Wq8aPyYy/aoePFwr0AVg
wVWq4lJsdTIBcCXX6/XHeBIYM9yf7fH8+2yAZQbk7Uwed94cbilTmNuBaWB4spb5+CCfUnp7qCiH
MgOuJ2GQ6HFB1EYBGKHlLZ6EeMKpLaIZk0xbzv0mw5Cl0iaYxRVNPLVLOD0DxphxyMJ7vF+jaYsF
8GWlmP6CDQxZOeLC2tBkUpQGeGQB6qRFjgGf5B8GERnwj2JJZa19Ittv23Y//Quz3w2085LbFkJC
EupqfpsUHq+z1MH0We0BodwdwDqQzcTFygtFBk+EbzGrK8zeAWpfzgyM1+0N143A9FFoy85+jEG5
txgsZsgM8XQEHhyczZmcCGHwouPtIkgodh59Nk3L4hVe/U0X8rQcJMTSuhKCnjGRjPtSKjo0g0zC
vPZR1l20OALXJN42J5V4cYfjGVG7vuNoB5Zc4boEc7taSS5E+SC1xsXBSLlK1cUb2gv83MAmH+g/
fmiqSG6wooLIoeewdAZ9QFx2PO7sIwwRcwjJ1Cr25QUztP4DOMK+HnP0fjIZGFSYlqS7CT/g+F0a
EF/IV0gKT0M2zapX9aNeG6ZHUfCjsaL148j6cQeWv3CrxLg4imUGYMQQGpfcUovh0FU/feDsko/H
7m6nc4dZVjYMR2bMfwCcWRGJuZOOuV+K8V4c+rDUcWwzyg/cgMY0BTVXU/h51SGct2hwL3OKV4iO
Wd8J8Co5rzh7rylGtoEhTwNlJ/1vM7ev7VQwnY7AapM/vVYLgi4OuKmGOSQ4kcdMZgKLlqgZQjG4
jWHjr84JTmcb9jK7VLNeo3ATxOyiyFoZgEOsr4GzDH/EmqOaSAO1f+6lbP2K9PrLfUof6OVrCH45
aBvtHpFF+ZP7Il5l9X0zlRjGuxQiwtjEx62DmsZ+0Q5aAW7srPMHuTVwJuEKdfGx0r23tEI+5mfs
EdmLm9pO0eXxd2/IdWZyW7Wlon6cmC2bWM7XnSzb2icLFdXQwGtCtbPipjbK3DkbvPiY/g1s7Dsq
PihwlTyzuvJrTUp4Im7vpvWp4W/cjOOLaxVQBAcJs3UWy9vtXoViYxmbdUfWlimnrMlpW1BEUhCY
NnqZlQ21LQsz265SE0NVaYk/wO+pQ7eKPE4ceGk/77eJZXGEuFxud8BCXYcJcuYFePuhZmusu0p1
G/8VGDI7T/wIKnKWhwe6zwmB8flEO8D1V8OIZkyrDjobJ4DTh/eyvHp47zZAfjrI4/4glodkOK+2
4od5ynRj8ckXdv+e4aVgalOxE7MlXaatH9ad8fs78Zr367rMNv26d0UcEH50GpjQ6hqYnJu754tF
j1JOz+A8FLdGr0YeR/x8KqPsyss4pBNNk/2/TGr0mcSRcfAHx1POXDfLxC+RO6Cr88/HMpN8Yytg
wXh5DFnviMYkQ6uC8kinuBzRHfpOYowa4oi9bOacdcqiDZfBP6eC5mjq8/UANYTVX5iWGib6NJlW
4meC/6PIu0Sro8PxjbnKuINprY0KT7D67SG5fUR/QFqKgX9hmlmgexJSryDmk1e1FzG8RwJQtTqA
L7R6VgwbF2DUDCAiIHkM9ACvWnLWqoMyT1OzBwRP1oLoLtMjK80RoGQS/JHAEzV3CaGmDsmA0QbX
TQ6CqYWxWmcKsAPF2PrOBj/1SmHxCji+6Oo/ohub8v9yWxyraO6dguHROOqjgJHy+AjVlzsPczC5
S+2OuzmnbCjPm93VvP9vKgwxNuxz4UUnWxL3h+bSfhbHHgQTC8RGAyoOXHSYBY7eMCsoCrbTzXcu
jv+y+TuuYr9CzjYfaVDS5eXbhowA5xb4UPKZ+mxIUcglyqdfsDPYEbLDELirYvmuigaoUnCyBeJv
Dwqrm4eiFhTQeyR3/lzG0KD/OHlNgeI8EpadwNIbyoXw5FmfP89W9OGuNNj7MGj4yhrw4dW36Bpo
5rwzYkvCorhCtjqOOxXnZ5KkJgdKoZU3pIAWZv5FcFo/rdLFu+6OiLdSZNLkbPAKMIWMlntAwH1o
oSXnZJMMsiJ1l2OhKsWUeTZquaSkDgs8fU8jScNwZVKg3eyuaVZon08ZnAZUVMrnJPNG9RfOait8
oOfsIs97SqXFS/EtNo8PcTi9ZX4Fi+VgrPDGrmGpos13nMkOcmlzA7k8y1SMJpsATTZjZxpVKa+8
0dQF0qgQ+oqEU/N1ztde3WaRJY8yljqtX1dcQGsGzAbY6bMJRQd1EKfnKTFtvZX8hgfW5w+GzNB6
eRTjEyhQmO057xljqYLxtXwuDp+E9I3rQZe18KKJx7f/gzGpDrMoAjVGsmVwugSKe52YHD/J7ZO5
ZqIw2KU6hxqfPavvEnh8hXeBeMpMxjSriwGgE/ELAv2Hy7F5KLhklXopRjQ2aS9TVpo3qybjJChy
weoLI7bgi4Ow7bz52FOiocleHigvO71Ygxlvr6uRgR9YIwYLtQdKjt8heyQTdGEwFj856D4ILguL
yAA07hNBJ2CD7xja5ETRWzIdZAoTZWUe33n/DTyh/CIeDew2GN/2TwqgWvYYdGr72M2eF7vU631n
JSSDr0FNNaETx6uZyrsK348W+y29dDqnQuhl1nnEhouUvfV0aTXl/rYnBrrRArkXKAwVCrQ1mUGn
yrxWky9vuum87HV7M4WlCTzLFSW77I0c6wsLoCwNv4VmuuNjfPY1JD2cHSsYJbwshUBrqU7BpQGB
9jnuBpA0oRe2ycHQxCJ7M0oniXrbiiOQySeongeyc914GCVniqPU1SYEiGYj16DCaneB4FlVw4ZX
MO7ned3WcxKEjhozy8D0T8FKJcCeCSyA+IW+i7rxhLYo+ObRyUgAvWfjM1WvhcvzZx7sMSwM7vFC
se01C6iOe+2XSHtmNDlAxvK8Q1uUgzkcoSbeKAizrolasz+2nu2/OH3nEfK+cXJae6V15PAdVIva
4rBQa29i2TbxHjcMuTVi4y8LCHZEVkO+Mz3XlFkVby/iXDiO/D3zSglhjQkIGNEKTlKsVXMNSbeb
Q7D1aVbFmBZmZoU0qbHFottoMD3HIR88WkmaFVR7Ttn1gQbXmgjYngXf46eaIKwXYZkM9KQAYWg1
odoTBChIkS1eBXm8f5hgM78UPemOO+opr3QsK5zDMr2/KOwe94lib70lKt1aNIgSid4MGnf1+DDS
5Ji5YwoaF9lg63YyWW1LwXy5q3eVplXj4c0fdYY1ri27ibxvfI4zJvbrFByWKM75GnQnWtbyFbEk
5AzCRnffUUS/YAQyDLbMljqhznXwYJtamOWMEWSzslarQABJAyhlsLyuZZhrsGzsZxgJxVICUHix
NFa+5Fha4vQxAmPMoQALhN74yIkf4v6IwAW/V+ULGsMvVZClQzDqqt/FK+7R/nbRPtUWIhIfcr/R
39VSia3JOFyELLPhxCFJZuWcjplb/jQvxVbwGrOqQKYFNt2T0Iso0p9Dd0q6VSmxU6/vOm0kidSc
aXpMcdOo+e6jtL0y//Jwm78YJI4MWPCKUjpZp+3+5xLKg2UEuWan3PpJ9IDm0V7Txeo7zc9uy3gd
zqcu4+2TqIj6MgrDgb4xOgg/TRhiN1mjNX//yzgNNhNicN9B2pARTqov12l3XnCP5ko3exXcqLHg
IYGSdG3PmI5YCaXQK6RZkHh5qDhho3Ulbl52OrrKykvM9DNkh+F4QBohKVy4ylNhyy1r44ovR2vZ
sd5xEWEWg254fTbPkeyk4jJL/RKSyHw230XiviatNkOrY7wZTQle06ZxyMaRe9jrorivOy2Emkr7
5OwX/G8W1X1+Kcv+FLkUo47Eb1SFNlklVOYAQ0mYLNAXq6+/MoR0EEac0CtFqP2T8frirsfHFRN+
Clc56Iatnuanv8zdgJhOH5x8CiEaLW4TdB0QH0kaX2Ikm6iKY55buWEfZfsFZzsBQFWXGcARs3tb
CEtRLZjvz1q/oG8ohFR5bwzeQB/afD+1Q/epk0nhRgV2PWo2jSYF9kQHAfXVrsn0RyjIFa794afs
a4rMNgY/VavHsu9YXj3rRi+dlP+JZ/OTZTx6XHBtf9mDVK9ekTqcOmyl6l18ugfxUh70EolkcyEZ
sMTBDm4ljr663BCUkpWa0q0boPQCDyfBC1gbDxaBawZcpb4BD9p4MUH6fbFNliJLwLngxXonBj6+
vpO1AZGpr3oFIv1YjGAeCgoD83Ch/qqVChqzwUih4t/AAacC7CeEjCkNCLMHFW5L7Kb4Vaf1llQu
MKdBrWhBjws4G42uD/HdbZEUspRxpdICwURvb3K1uyhcDltd1j9MiVDewr3DRIQa+OG4AOLjdC0W
pZV7r9+v0tu2yA9r/IepMlk7/OQGKUprzzz8tzsdovMcLjuUAEw1R3abajShncRj1uOEaLOJLtRI
0s/VVK/ngJExHTkB2s6QeOjyLgD8sezparNvwPDNLVSP3K06khsr3VDj0BV5SNEd+3tzCGN4VbMD
8WHS5TecH4eElw2QLJQbWqMuXKtRWXG+KaNYv3JlFYXyzhPdugIw9AGIIu4lCJiInguplq+O8ZUo
Ybdio0yXo/qtTGk5vap+lRLidGqfwWxgIWqTVI0+4WXcdnxAzWrJk0NYgU1ZYb7q+KZFMSsq+o7y
uORL6aPUJ2LPo/tMGlOCONS/47O1Ci4/9msSenGiQJrBDZFXamTGUjP7hgFMA5f/JKTvRTZnmo1N
exgSlhw20SQUFg/WGFp85KOOX6qvD+pELxCgfPucZH6p0BV9MDbpZQmjAZrG4EwNOzRRe/P/eh0F
PAuNwJPYinzXr18hMcj33zpUc4Vqx0EQIJrOI/SL2PGR7lVkSf9ulEK6evWmbqftTr5zxhm+fYxj
RDIkNd0vTJre6jE9KoOl93L0oeoz5wnYVXKztz/bJN3Mo8TliYZ8znZ009cKniEaFBxAt8JZvyHm
AXPCAc8gum0BTIrU7ok6ypVg61qSUKu2WoD3zYbG+p72wrIBxe7bGW0QaE3blhihla7q/N2CU8qd
sr4fa003cjdq+cONfwrHe50cz+OcApuxy+NBZ6KBIgYMbPM0cVQvzvc8bWYb1ac0IPlXxuiiBaM3
uIQ/iKJyNXiW6cAMo+/Xy02rR+WYsafQSDiKZ4ZALT9FcAl0Me0rwu5rq+OIMbZ38IYgQmypTG/4
uhiSmJY0s/ivbKz9HMg6IcqOIq39K/iDMjtLlsMZuemmQWOc0Hu06sF7frM02F09PC0ZPoS+ysXj
vKi0yC2Q2uzY+u1EqJFa34uLxQ08UvPmiMCo3GNPuRHQ/vOWJIuY6TNyLPtpZ2EkFZTb96D+mZ5S
8xcc6v2tJ7z+uBoA6gUr6yMlCJCk2lFk0NzuEZ1v8pqMOy58jkja0+oXBbAV5JWKeOeAGuv6y13M
xld2lNjfe8LFF0etQ2cMuyoBENyiXibVSL+sXA6V+xT3LStYCewXuS3KniODrCYs3fRfR7ug8T3N
931vizcXJYQ/ocnX5Kt3wYS4N9Uu+cifHUikw2G9acE9NsiD+M1nqT8/lrV6D7QBa9GmFMPa3t1/
wRPHNnATuF4Og8uRK8AUZ+jPa0YMkF/+mm05Jw70uEQwXQHUnVP/FN58pWWgNtdHy+wj4JfsVU8i
Hr89uaW9KB4I/d0bEUjvuqNgzU2N7WmL2W3BcEfDSUOOpIlEHYJd6IMyctss/X5kFbawb+ZyZlCC
fOSi8keDm75k4kMS4i3p1OR2klSNoZO6vt/UMCUje+Fh6/ahx5ou79PueP8y435jQ89++s+F3MIO
U3D9GU4/SamL5Ix61EuMLSb7Z/rXlj+Dn5sqLV3CF1haxJadxKqq/0HTB+IgVIV40fRQFympr+le
KuyAmgtRBzSWWMrblp2puNqIUFk4AwPicDK097+gXK7QqG8GaFZRUWhAn+b2bTKdWmNIPpFupKge
bU1okTZonz2hbT7SDhiYsfaZxp8ffMr5bIBloyMeh9Z6NA2zhMvkjTSgtCRGs/DC7B08JX5m86re
Peo6gViWeIuI5fRy07+n656m1nZDZsk9jYJmjlPj9zOSGARM5w50PXG11QWbHHsY2tIKiNx9Dio+
0TkswlRW9eGgEsphGU2EI9vqq2fG4PmJZlM+6WAaocanOqUVFw/+0aE9wht0hiKBM/2nKM+B5Ycb
rluNaUMH3Z3GCR2gKs7Y3uh33iqw17f0owxVjagswv7EZYg7hNL/rVSQDUvgAwKl1NwHS5z81VcE
dNYM+7BqMhikmBW9Le5udFqtMzJtvI4AWg1+mWpigNePxJ8KCrvQjMBMatLja2hcBlokuoMmNDWb
kQojhhZdygKho1eZQstDAqciQqAXeXkQR++pWslodFy8VcQnB2aCgzW7bnOzxPyAJ/PGP7VfECQ2
Y5B7/9HoBzIOsyh/AqGa6IPdqIxR1KxFJW0N/WO1DmlAZzzIM2cEsmweP5yCiy6adNH0DhS1RDef
dtU2/FMCa9l05dD6Djyh+plFT79ViNT9CpE/MW+gTF//Rhvrta+EvndTrHYbgI+ihWZtITDMQy01
x7VbUNWBdEcxZW3X3pTWTCgXcecALW2STdA7CZEXIUgf1XsIEPYRTHpRmu/NszyQDeqUphueuSeM
+XbDPUueC3a1NCC7SFNaR2L+v2HsPd8L/5LwrQn33KR86p/CjtjODe/W+xRfC6xeee/raTIdb5HC
8HWDuB2R7X72PSsd46lIr7oJjc4qCEDbGCjm9BlOBalUE9gyF6jxEsSyjr2jjn4siMhJXbYcRFlP
rH3bEyq27Wvk+PL1Fyr+AERKVDpy8PRH4e7F/gwdpyTJyt6qMoM7uEQ/2ZqbWmXUouzD/dU4on9G
31Nje7JQNLK9Ae3hPJAn8g37jyVRktzWHuTM4BHgYCdMMmpqmrYwS6BiWKgtTaRxOlKZxMqF5L3n
QEReBO/R8RtCNcKV2Gph1ZilsMFSAZB4b4cbOPc6Kx0+mSuSnfDD6pnKyv4RSXgnCsf1c9XzSuoQ
4tWkz65cOAmKBZ4kAAZ8Sgu3tcqwAQ6zLidgWnFyYUVkNdJmLPVx4Skk3u19ZnapjarM+Kjjk6qK
fJ7NQc3vXasSDLIYKB14CteYMf7/S7TGr3xbgZoNpFPUE7YAfJvjCGOIfBeA1BBb4AciAL9NmYAb
6UIs8FGLwg3fxVk6iIsAjzW4gKkDmLVSc229Cr64hMZCGo/qx4ocT+ZvbW3cq0IQePjN6sZWFGWJ
VTMkJ7ewmoeBBFM7R8037byvzjoEtmAhfoaCLtcksUV0qm52W9wKSxNuAP7M57m9+iOIfThtMAui
sXkhZhTZO8iCN03IRnMMNDCe6gTo2V+R4DyHFLQTLEJdpOUf9pyhdzx1ZKl8IOSw7hGUPcopNbrb
epKyX+XAhZZsWm2BgnBw+R8b2n+jWyuW3nNuia33YLsn3oILR4lw0uNLXzSiqUITML9h4kYqA5D5
ZRCsckbUdY7JTLwAgfvrUFWZGz4x2f/k/AZuwhCoBuaz7ZH6OnfvfH8j2MYXtt2BUfiLBZ7T293i
xBOssivdfN16RFp8q4AWmfcN9x8r9LiRVjt+m2karSKAhyQDQ+pzWUnJbdxhVnDudpeKjFEVGJ/s
dYtfMVkw5O3yxYaE2lE8WilMmaFyPAoyyi7lN+hPj+AC+78dAIBywsFE7sypbTBLd4Rp/WTaO+OT
CWpGfXmgpnlXx3exrYSC6qg+e8HUZPF8ANXv6mJK2moqLpHKb23NaID2lAP2zhVzsV6faQ7N3Eez
i4nfABy/KxsrjYZj3K34HcdsjUNrHusP6dK7rU0SCb/V+WHAUw/XZQK6hh//ZhowgnuCpjjDGa/E
BtouazIom1RqNISqur851qt/c+MtL9z4rm2t5a3rE+H3thz36FLSJRARZpuB7jXfkxHHBOPik8cG
/LaVwHwudlMRQRSkI0UXHHT0tX5YH2utQl14zTSc0EseVPUG/AQDP8Jq5YJemp0Qr7BlulKHMkj2
7IOTWvXmyBas36di6GSxCZHdZkDt+2l6kzrZUyLIVer0VtA6vyq4p8IHH6gGRnP1bKJTBVkRyil8
qf7rZ3rCW6TtEg9iuPNFUMlA2B0YIG2HyNrUP+anrMuauM2xZGBY9RJeLtgYC9/Yc3605H9DElun
GAu6xBBffA+RYx63xhCBHyRPqNbpgKzZb07925tM9j6JmHfIL8ZlseByPFq2RyVvG0FIMOOWzpwW
02VHu2muxhv5BmKiw7pJWnR49407amOkCp9PUMZt76bOJe590igJ9FNnbdTEzSj/DBa/bBfUwQ5n
MrO+Azorb/8LLq74ZxdeG9T7GJ4QdmmxsmGto89VUwhGXdTtW/TA5MovtrP/7iaEf9epxAeSXAXD
7EbnMibHW5rawVVJww3Vem6u1noDI1GdHPIn775TaTH2rx2G2giyrIwYZVALggRWFXt5c0/yAbXE
hNNJ4SXexGk3/fi4OmvLJ0KaMAhtH4JkDQkSOGsk/VN5PLhWwmvwSLmndlXDkrpUlyI4WvpJk9bo
Fw6tymrCJbZKohFf4sDokUzXTiOOyzTNhWApsasc3Lznyy3QNUpOT6gq5GbnwXlgmQmPulqYs6K5
jPokqPuH0PYo6JbDKq0GAbLF4c/OWkc9uykA2z0DE0I2LplHEzGB/CFQ1b4d9lxEEESxL0Gd5nj+
w8x15PE3njXwTKg/de6/1YzFE0wb4dP8Ui6caET9gRQxtTrBIJoD+fyK+ScArnVyxneOTSCi6fNt
oR9ToikFY1ZATmnwmgV2LINheVnLMBBY3yrVhlPYy4t9I9YIuUL4JQtSjrtFps2JqkVKxwfrfxKU
ioWbMnw2e9mPyV/Aa5XaSEVeqK1XugZuU5nC8OKTEWVUg73u/ZQj4DuCiQ67nlhD4cV6Dq6nV7lg
skA4O5PgCddpVpfg46yX2g3g6aA9cBlzzpd8bi2bH1YvCFG4RjIk5Mhgp/k6je5NpeUCwHy2cpXO
uf0f2EyLsd/zmiaRU5t6vJsgsYz0tth0foX3JhzAv//P4qEiSI21jijkDM88jaTr5LmVDlxRYCXo
2k6rGEu4A3gwXDJ882Nmxs+TSSVCpgVSr3uDJolBDgnGm4+dWy76mbkwoWjR29JLjiD+civYtI4y
vShnCGtwfMfL53NeHjaKa/uAAhcmNexnoa6wSr66PftswCC3rGoE2OvYfxN+UKebRRvuF76HRvTT
5eEGKemZagD8ah4GbPw12DMmLSe1zir+YJ9aiqHQo1LriL89T0cuEFrqTj4HavO39zqpIeawqAMS
+FaVhmT9eVHLnjhWRAryt+fHWjGAF8e6+oNkHucWRXBdhG35VDh95Cj+7PTe9MOeYRbWa/MyG7Gw
T5WjYc9RQ2HD0sChK40ETclmBVajOD+8dRS9FRtWoRJnn2OmF9E3YwUyiAtn7GrF5nlKELAdEO4+
5yUjn/d4uXtzzhuMzwkXkw1FvXDy2AiWRg769KKM97Yh38/O52panfgpKr1epLOl1L+5y27d9jo9
CAFO3B4EMeLcRAp2htscs0/kVH08Q6WFM7aYacmjY2y6ojeoI3IyGlrZdaCJXatezmp77HJBTFxh
RxlVNVDBICh3S/3cJgpnLpOhdKXifhuXdNBifUpXjfnyn+3mCuWsBujJs8FTjkjczHSd7kDkJM9V
TcNYqHYB74azleokHC+CdLzz/0Vtl4J8XDAhsfZJwaf+0vgPRObkTvlNO59EHwfZTN1MoPhc7Fe/
SwzHT6tMeXQeI5GU6gJcWzyxnQ5PMGHUdxaJfT2A2yKns/qiWnGQQnUrBNp//U8dRcaPXVh4lt+n
uTXSdl0ZZ40oDrHWuDxgtz7vQTDiO/oW2C6P9XFKtrU1RjrjM24kF4qN+Z2TCAK7oF0lXXOmj6hC
TDFG408FC8fmI6upgu6Lte8mja6eYsw6t6DQAJct8TkKjok4ICH89mmzjSjL3kZ5NbU/N/MYvdUJ
SZoXwUitwaD5WVID5vCv3fywSg2gP/qFW6UVMuNxWYFRFzHDB3HTMo1mABOj4k4FgIFzH+4veuKn
c/DS+RtgPnnMOg5GAyGS73dYwZI1qbX3nS1IvpXO5gxb+/KgKmJZQ6XHONpYRrmsCHFiAJ7VlpAg
yYy4jaOb0Ybl4899zX4nZlFFklkTx2iF3YjmW1Zt9L3PhRyaRO2kpKfvOn2ek4laLavjUm9r3oiz
Xh8wPj7291LEw2lVEaOoRiXHln/SkCGctgNb+1gL+OUjEpOnjESickBg8mPfRZJ4IzCmOe7fY6Iv
yXqmLAWydobItEEC3mrEspzFqyAZq0JswKQetBnino+FNdCzrvc/ARFgevRfwiGgpn6UOvfihahr
UYm8B0ooYtVxQtcS7s7C1uqp9HhJ3Zl9P4/R88lKV9JV0LfSHfLkSmAmWSayq4UeT0EvzPIqYMrW
ef2VKPP76X7jytNxrtt1MUCWtnDnkiRZvAeht83RYjTtQUsgM4qkYpTt0056BiNJKeFfMID0hAeo
1KadEDE5AZ1xI66lUFZqcQfNXvugO0MprJKv1FfRW9BWKSCQHHOd5tAWVgJcTj6Wuq+ohvYXXdc4
q1rdghl5Gwc7jbVLC8UDlQsUxYGMmSJvypUxf4gGWKXUn/V0ftufqjjGsoLV1WTQ/4SdprWyJcTY
2kTXhmXo1D9xPPPGgVFRLFy+aEMcoHhTaDZOWaPydfSUclScyykrUMQyWw8UYPjATu8XYZvg/fHg
LBWd0hQDMQG24rGDm84KeIoomaeCQU3MClz/a0Lfic7lozhH4DW78m+dgdaSPsjrJxaVnCLJQu+H
05utJh6HN+u+CyRCVy+69eq8cuu9jaeZOiNMk1M19h40pWzMQLhgFW5HkVR8uPIOs4/FhtKSVQdO
6zTMJd2zj3kaxx4g3RW8pAvE/U07RiYUJ1iciKHiBAfIOGUVW62DczUZTx0qsEDsp/n17cpRSaDs
LRJPcFhx/9KB8/5Uk9xCcP2wBN6J28pBrCiyvjlZotm7k72jJv25DZNBEsh28kZiG8gUZMNh3+Gv
Y2WmgRTCoNxE/bRc8Go7Pju30j+gJcz+61tugpzz+OlBJ2wjeoF9ONxzo4jFo71ApCWHx5RwTFau
4xdzAY/Ed88x8Exwba+G1Oe5k6zJxjTFSrVhPvnrsyyyLOO6Y6vjleloslvVv7OU21bg6GsEqRGC
h6HC7+BgkcoiyNszzYo4/t0YQAQjUZlQLGcqVctCqcNKz22UAVyjoPg+dNEOiPw5x9MPQFZzpAZC
01/2dQ718dgjoDqXohiB1Hoj13HI2NEJD+6FfZEE4Yn8iibQ09olecr0d+b6Fzen2dwNqOG8Qz1C
UJfNAAV318d37WZFmWshMYefYRJ7KAigJ7gcdk7FJ1nMule06n2aOoTW56s08vT0T78Lf1Ur9GPM
qrSOQea9N2+1PlNTenqfgio+9/IS5NRTi2tzZEIhOFX+YGE6DShcycPHz8Leyen6yhG38GP0PO9B
OV7DqdScrfsDSC8JPCIwh+uQLOhBC9hA3yCqC8sH9OmUhZyXSLbuzjbpPvY5jjUpjgBet9qo3cLC
1S5ENzvBMiE8qSedYHi6c7YliTKOilf/BEvkP2bzLSipibphtyXhX1p2196mIvueJ5g7nZLMx+5Y
Pm/rlaLiFzgv8AnwV44bEfBBu4p1o52B6csUIKT5DMldvWb5gAlUdqZPebWmG3VxXSzN+mYCZA+J
o5QKky8AYZRpmeE6qlVehWuK/EP8HapYou5Z/GyPZDmNcB1UYGpuPZ5/YftHjUivbtXkLFQ9T1v8
0U5FI3OjQSM2/Z40bdKJDJ3WPYsZ1c235l+Ud/rwkNFnpDq7oS8R4Czc3gRRVL1gaIV8PbRoFk2w
oq1NXvqCSAoT2osKfy2afpTZwOrpy4oVaqM0H04UY4mgT/6mpzLwwuVd/NzhSjKC1Fr5hm/GbCnu
SRegLuUrU2+U6pU/sqeBdbUX02xoHq2l2lHckSsbeVphw2hpOBEAsQSl0Gucyhr3slWSa8AxlyO/
qnNARISrpfR2imFQ+zo2dDn3cKvxfGCeeHtmejF0P8tqcCU/ASh8SNVEdvXzxOyrFsqj9Cl4lDsz
x5CshtOPt7QJZrJjQHVcVolTXrGy73d5BdSWWvO6sVgrnWw/vEd6WNLEL3YHEJtHId+BQjTydn+D
HdsjLSePTcNlCJv86UiSDk5THlTFVhGFbG5WkwCDQpQXIPiIUc/gbLgtawzRFlFq8k6ZdSBTEAzW
ORn1q7uprmtSnkETrN+YSGxgaWVW87tyPFfd89OXPIEhq+k7wVqzEyLkxIoZ9tBsS5U5MCT9cP60
R/IhJmYDMyIQMIsRpoNbhlS+KKauWWqvzlAlXPgF/GWh0hQ/kZwRGee7DbA6+lcSQKVun8EU3QMC
PkLMPZfGyd6DbA7nH/beOElY15/Hxk61w3r9VjrJHzexgA2+RpkSj3uJqX5u8Vq3ykheGm/Wics9
USClTMcVwY/3KkfiCiWdi8khy7eL4QwkHOsfnDkT1EB5/eAxWe6sExfGeSx8w/4h4hoU0k5opIFG
mLRbDcvOC8t9Xu7wvGN794bsohYhpCkzetN5a9YaJfAVCpGPwerUi575A7dIXHRVmBaahXOoKjis
xSIw3n2PEPgcGU+nD1qHtbGsusIaN1Mv8KhE4kKrXNelZlV5v9L5gW3s3Guygkra8Ob+kDrSgZD9
FHVUenmSGVZ5arrjj2WOjB/OYltpdK9YBc/xNRLLt4IoaQbVDVihgy2t56Kt48raMtHi37DLEHqc
9r9U8gVfEFcwUNAGRTrV0i8hzzGDJqlYE+PATuUtEoM2E5YJpC8rTDg5WdjKbQqRYgb36FbPJImp
5y/MHbGCf0XtQzcZtb16sEJofsXCRLSA1j8wu5s5XpaknRMlZDpG9aHh7YYE51jmtj8ZdQFl/cH/
c70tAAIjgzwhkiH5spg6Q4gXEU1INfDJYFWxAEZDTdEgys6mAflf6+6xXrhyjsu6ZbXM776eBMg4
xxEodFuwCNso1j7AX4cXqeTZaPouG39zTk1UOHZM0qUzngBoGYAlaExrU2A4DPjrBt6/LW3JWJ6W
3MV5OoPCJSU9zb8uTgTYuACELMUVfFHKqJGjhk7miIJpJgVIrK3WeRXtBgquJbYF5cNG+1WICmfX
9acIUyRSD3tQqxauGWLbNovP8z2+2do4QOyNL0M14itDOiz/uobVdpRx/PcenLUoPsfLs+Av59FN
mC5CZR3P0ChUsbyj/uyG62INYbV3xnmlPGyo+cGynzJAfLFc8bmRN6GCSZFaqKL4fqGAwM9baK2l
VG6emsunrB8WzGQH0ktRzdvXI7zcfIkP9ELV/s1DRaNnGUrGeesTplhMdbhyhpYYLZC8mEh/PyJ8
C8VbxavidJxVnMO0Dktz/Zl5zMdhLzwyBG2cpRRO/wswrjo2x+gYxSOVspn5H1Pk2+w3/rAKwNvG
ktJnMRN++2nX6d+3N95SAYkV+fBzVH51iC99+6U4Z3GLsmaB1z3kuxIxDuY4KhE55I/SK9QQylRI
Qr0VIjhdBsXBDnGmkyggoXR6cSsxhmzFpEyPWh7tKrcCH36NZ/Al+MyvwVNZTEVy3S6IWZiGZXW8
vih9YhoXxoiRycPDK4fwGzy6P4vrxCYjZDcmzcK5hh42/J0wl+XSpX6u7CFFM9yPBlBbFXnVvltP
ClHnpH0UUob3NKMFvxoY/NUPOCnpAxwhw2uQfznUD93yMu6JUrz8RsdjFTVXv0Nm9j9DLwyhU+5c
AyxvT9NFr9U58cdMtIBl1tp/JxYMDSblSfWkHhv64+33syVmkU8zzL4jvHt7xmZM8kNAM+w7Uj59
gNy0vbO0jrAK6wQFfA99ZMTgQz2Uz2c6omVT3PerourVqFKe5hP9fFImaQddsi9YJmBnQ2XHt4s1
MVSjciOoJd1sALSFpgb8OCIUPXdDH6q6kyPVemx6fQzOyE8QpSKkuXsKfmgvHT9RDe7r2oZGZpkT
C5jfbMrv2EWRro6Tk8BO7CTowLsgOBmnQot6WvPjB9qBVk84Q1E2dUFGM02fLU51QicTuZvzXNuL
yWRmGsW0DyrPYwfxNxw474dLqkMISggMhf/901i4iBqVHbiubpP+ZxZDGW+yNnU4j671cbYRo78J
LbN8F4Qjy0sci7hO8uuUdcchvnBPRpD0Rgryq+z9qognDP48IKrEnFWjpfOUJdoICN7C8vB0SNc9
fphPn9aHVCSJpXtQxiyEON4BS8Umqxi97xlb0ZNPOFQT2/s9YEWvfPtEHZN+sV+sOp64V6tAkkFG
C65wR5Acj64iu/zbHbzIa6GQzi47yp2xvn/YTk1mvOUNKLGI/fjQFj0fTo+72KjXaZbo3UZU1z7/
1QWCJ8anRPieYu9IB9zydANIvoRENjE8Ze712qMJ/3go5u4QPQCvQeBUqaaT9GAxSULYgpKo+Xf6
Rj7YzR17BWL2nMi5jBAohPrlXc7EdzVgdot8qzr7BHJtaWNmIB8K/5HUOD1uIvQZqig//4WgmcZS
CSn+KvfqX4lTWkiHYUGMnEOo5iMvs/NIREO74dni/0CM72P7TItQZ54ZZ3aIytYLbTApAjg5al0D
mY7NyBjSyDX/o+ExvHreUZnfvWDAwbInmHaflLo9Hy/IlFNd3mqyKMu1szlwID6d2vKsG0OxLKw7
h/Izy08S3CiwPQfhXzBRLMY3wmlnX9s8TOxAb2R+bteNW7dmK2wfH9hc2esHGI5zehCZEMHdve2t
upNRnLuDbQ9srOBZzDbkkXkL5daFM2BFgxuXwXIWSLs8PMr4iPbQ8dXMwBEcY7XPOcJP7heTdPq+
5zEXpqOMz0FxR/Q6NTOpPOcduoEU8tQii277oWuv6mw80+1xUsYte82b7dBDEXo02y2mFFv7FRSa
UGW0VJZKrBmKhlnTb9G5ESIp3lRrmrOWnr0vGLUeLVNTinuSHch7T0zWnSGou36YQV/RLd5deXlp
gOQMMFlDenpyMEdL/NefBArgM6Itb5l79CztipOCY1Vj3eYSArbdRrTAKCYLKminvUvfHMlf6aAD
LI2IcdUGjXF4nPI3U4J+v1nKOEPzV1kePQ9wQ2YN1/onpuLL/ykJ4vpfRj/tRByoZGn/DFES9WPd
8B5hFsB5Og19dgMm4kiIpifcIwl44CI6C3+dMWTrLf0V8nh8eKqYxT5oeiqg1i6Cyr+6ZZ0D2tnp
0yYi+ljoLXvCw8upVFLpOTIxFdY/Bhn4kqxikpkdL0g5Z36reEVRkfaoJpPTxqjozd1vyvtn8Fby
X1lvLkG76tZWC0Z4jakBPlMb7L4mST37S5/g6HwTNCgGK7hZr7sYmwFaiIAsX4qPQrcPDVBjbMEZ
IUp37mDcX0MTf9dK0MZKFUMcEhML3vSaK5Jy0Fy/xgHoUMIB+bSH152qKwr8k35aU7+VFdigxj9d
BqwzCDlFAGNDf1mFLKeTGi9Jah/wZ8zpcp/5tDERrGkO9v1Pi7SqW0UlwcrdJuIW1Ym2Xf2bIr5s
39acQe8cmJBun6je3TT7mHLzNqHiFl0xdqpCn4KBSlD9uH3Lhpy4xFq0fIH2zulGXxi8zedYgAzu
1yZPD/kZd7kB1hJozVlYaOs6rlunM9uKLpNXxP1gZCYcDAFZRKzt+CKZfotm2NODLJ/znLk6Aplu
+N8SrYe7rkSeNGMipQd2YKYqzS86GAM52kaZn6Vf9RmHfHAHZ2hbv5lo1ysqHK1BMB9QLulXMmoR
+SjfajDDl3O/qETGyrGrvJMTlx0alKIeEsNT9DTctoZSq0xjNkWUMHNz+daIGw4AD8jmtmDrfliM
e1mvoW2ATQCWqp2UL1VnJkz8/VkhKogbm16kOSEmOecFnZsAK/Etbup4H5N76vnFVcsIcPJRXF5p
2ImmarM41H93CDk183q9Qa5ULKirQqfmyzgUefK94Hq0UYayRkpL0W5C0WLMOxD7nvF7BHvPNTwF
zRKEtu9Vj6n2UEQBm10NivbXEWk/g4N+sW7AwmMUS3MRCrOudc6TiTsZ8JMuOf17JB+9AKKyED3/
301rAlJQxhxEZLc+UFmSlUuD0zv42qBnBhveVZARKa+AUNjqtiy4d48rJrlwcVBdyGvfmMXq+N1b
sE3P0ptDTgFypeiDllURdMlkb8KmVjSUH2R++994PDIZnXAcKNVxWgWfyrDP5lzOY8qKNOgBZjZg
IB2sTJXR8xVmmuG6y3iYy8gCVVmMCw2+ucgu5PVQaS09LhdJS63+2cvZnsSrujsDBETvxlshAta0
qChe23I+xkIIF55hAS+1FNSZcJUpm+m0gt0lHZYhHmQFqYYagEnrSuWw4DRXPhay3yt2iswOAF/r
D+CzBdydIXIglxxp3JLizmU/5YMTa0uuHnefRS0uaeNh8BBAStK4IYKJ+Lr1lD+dYjdTK+jwCFHm
bpHAuqgqkHwTQnaQg2QbgZyFptPgxvj+42YkWU37jNb/tfN0ocWPxg/nLrHEkr5t/y5XFPZ6FFUk
zD80r4KEHJkbf303CGvTsYza8IwaVf7sit7KhzCZ7Fj/jewnVJwwF4pWAFxFd7cXhrTSGHqgpd/N
HtQqxhoG+ZenjadXhduvXP5V0BoFjmRHPErH4MGeMona7x5nc7GzEq9Swoq+stjarXt/RtKOOA95
fW3y2lu/cmViMnxyj9W5Y2CnpUNhwYoSIvzorvMgGBQ9N9osyRWdYJ+CdQgficAKWU16GQXEyaVW
8J1lcPXLLFei+0CzjqEkAgAjdlnEsJyKblGoQJ+xlkYUlzCZVJARdYCiISnQQuz7St5DMgThMgbv
uFZea/Tkh7NO7XYsZ+igSNE+nUZf94+TDyTJE/9bh9Z+Jr7ZYgkAmEchYumvD2hTMzSb2E78ux3w
lsHClphsu9N9xzN+845xk5wR9hdns12D0hjPXrnh4JVASBo1KRUe3fZdTh9y+E+5irsuhTmpl3io
jjajq66f8m5jahXxxYwWrOIQH0O3ZH7z6hMkT0OxioyQup85+dYoL2KKxJeYQSD+bzie+YkeNC/V
xGarVYCN82+T5H1KMSi6jhPH/6X0bt+J1YH6ZIG0IeZr3K5+4sTpQrF57ma/6f7Ft34wHWcWEkQx
Yoi647yhrUVibSBZaorPz6JAkoqZ52GNRUvOUI9sp+D44LlxJYHrLVhe4HIyVtMG63E+bQ3yNU4x
ayNcC+kB1g04dGRyHCKpTyiyYJnS3Jo0C2c77IG+qUdYt3jRklQQ1tuZD24DnxhR3lt0xdbDBtIJ
17iTjaeCBNIugtBhZPXhG8jqv22enP0L48ibFc0OBE6s/YYbefbec1526aZIUGfz2ls99hR8nXmW
RShvPC6siHrSzyMTSti5ppLvf/0nPxDUQTdTqivKempYtP35mNuOBToQdpyLnSpRwY7WMLdB/vNa
/By9VI7K1OhVf/u/TIJYBotM3aV74U5pv8DJxA8aPt//Ll64GH3A20SrMHyJN3zSTku9V9co+YoE
ANyWyjfTmu4eXstoA4Lphb6N5Elts94JcO3FJTo1q5Krcv4uBDNbyEyqYhtsODxtoV4XQCMwPH95
/WVpKAAXH5E4ttEs6+VVUv8wD1Af9BdMmQjAosW/7VUJXCoATJiEgfB7urSVxrvNwrQ9C5UKZa0i
zf9Nhi9ykF4oZ36HmwDmpFYcYkrCFZlgLxqwj5m5eEjiNi5682XyuAGMFPeeuyhDzBR2mDJBkyvO
TyngNWsmKHM6HnJKkeonUkR8j+2yIiva4bxZRP3E0SDL32+sDHxmru7KtuPpXj7Ezm88cOGysooE
1acZ7eusJTRH0Zc7wCEkdsKuKVWmDpZNH2AlrRVFbNrkOuyQbeClSFNpSBNxCbWYQKms+BS23Arc
hDA5tHWubXAASygzmWroUgF8smp25pZXmvcnrXymOjtCJ+4/LXHcinRPyIbVDiM24L/V5q3wEuyy
rMF6O4Q+2DxuuX+jBfkTZ4BHWh2TUhlGFPYNiPXjhLov6+s76RkRZNOh15Y2n7ircVGTQQXDBHTR
jkWEJNiXPnqLVUZ/6NWAM0uttovLT2PgMdwdqIBZn8vWIyuOWtP9kmiPeq7sSd9wlORZlapNyH/1
xSP2S/85GVs7MNVyYvVSKg2eYGWNsECgNAl+WGjKJEHwke4q8blN/ONgdvxfXDcXky9j+xhnBpXS
TmgzkkRHt22ga9AMSLg7ZuxonGsEgmuK1dUIMztKReUXbxDmCpHFVTFpKYCti+DGA65dFPylrSxZ
/nBZ0HYdv3YSJIPREhIeOE4uURZHLzBUrEzgg+1yvQvGh3/aAPp83tFL1nPAbIbOc9NtV5S/m7tH
wh4nhimwnCRgA//ONVXuj+9fhoBF/Lcch4sa0sp/jmIGCaZ1oDc9JhQjz6UNmyD5QcCs6XM+38vv
94MQdRKYsyaw+hQNtHg1pT/35vEbvmOaFh1RvYFwtt0VnGIhcdVszmbP1fB4thHKCFj7F7Ndw2MB
0MemwopZnqSwsae8Fs6Khe0cvXAb+nJvUQCV+Q8mLqmMGw/1TCWynKWUFlxwxkhGqUu7OfsmeSV9
cDKKsJ+L77T9AMc/u+9WDoZz+maSnYLAHexip7d+r9qMjJeWS4iR86y3Y/gosPb9v/BhCppIE7vx
4DB9ud23vYhY8/AbunAV9mM52NcFwRr4Oa7htxgI7A46lcRfYD684WWGjwx3hjGfvUEI6WNJHMt5
jEpRpIKArWOwwIjj1VZL03BztvOeTLM9wF6+JQwN9+ZfI3oWstd1PfwXuetMX413dWHZimw9xEgl
ywRr5azaU5GmkWPWm8JO601L09OOP/s9dVkjsHGwcuELcUvVN2R0ROWje+uBk030R09DbN7cndv7
8ChJNpbNzkMs44kQUqPN/jIiW1RBtf6aXDc3GQqkrY5DjiJ3iToXVQQA5iSSLIe4ufnv0bopf1lR
wQQhsIm2nf8dygZ5XBN/s1pMSHQjN50Ic4YZeF6pIVySTXG9oAtQgUjtTI9H/+uOp+vCYI9PInBm
6421pTsv/jSyrP8Lu+JLgbBN99pgT0P7czix3lnOAfsmbuuzH5HEkPFOXXxCIfinafiT1lxirNj0
hlzVFo1+qLtlNNagooRHRmgeL+fmyHxpffJC6kRCRd5aRGuiJtK3z9eVB65y32AJObvLb630qI10
tcTiOSwOzIGe1P4LWu+hTH996ZP+k3El1xas+WELk6tfVzVyfta7bA+4ybIwrhPwcuT106h5b3N5
4ir2DwTrWHHbBlDI63RZWwyQPAS0iWtYbNU6j8LrywAvPzlHDuEDYKM0GSN3cJ9ShRTgn/rbmfT4
yG5Xd1ZTav+s0vqOtdEyCjkSbl++1L9++rwHiFAvxoASx7q9Osz4tuxDr7SMidqksiT3JwlLKVV8
OcoAUMxBv/DXhpPrFyds9iJ9/38p05Ba/Ws31L1MLvQfxYtlqPXEKWjUo6jde3UwsnkkLTcDJK7l
C9B5+PfJr5JRAgKMcyr/lq6FNqwEru5Vs/sZe+bvuAkqEBKAMvOIFuLR8sFUiSlMI0SNJL1kCKDz
1CDygGnMGbORAlgyXCtihFdIRAtw1Pu0IQUWpUsdt04pSlrW1fN/BWPQ8kDXYJHEYGXrhm+YDuT1
K74hzr+FugvylqedWGvc3ne5awuIsdqpo8gHrwXmEpVEUIuCaM91oZdjrhQ00C2KEtSmDUaBJN0b
nRl76k8yHjnntqjO/z1G5ZedTELG3eYSWsZ7RiOk0d23TIyWRR9C4rVK8hhuKhm3ehWGO64yKWSB
H0ujVWAPrW4OEow+ffKvaczckKQzUL7eZb3yR9womV5c78UmIr97+BlJSzoQ7pNubEBUS16/cPLr
WrzXVU85yETXhSqCu2V52IxOp5VpNcHcxfiYhyGpZApF5xp85g5r9dor8S9Z31OyaDXur1zjZU5C
qTLga8KPhXnzsLSPYztRpxv/hPcRuNFd8w4gHOOFJwcAOFqThBqhs/OcIAxbFLMF5UEyK2IcXb3J
HEyoXkXMGuPLjUHknj7RcqwK0846+qU41PTCdDjwygyM9kOsJ/IMR9EetTyA8IC36o6cvE2rG436
wHInarEuOW553KVFazhqXl+ws6pgstDeUPosltj7qRuv65zPxwFmb3COcT5pbrALCdzy7AfTslEP
ZH9mdqu15fhpHB1OcB+rqHnX3sB/FF8ukoN/nka6Zy1NHNtYIpY/BMvDjVZiuVHvU6/ato83f13D
D85llQqKcQ95wBM12ihkdt5jaDH6xyBjA29KAxnbdqaZ2zZ4uSblm6tzPzxOJcuXYI2X+A/KF1Q1
/tPhwfOoWRM3jKbhdEqH6osMYbNQMP0OIc89f7QpLeg+uqUJwCom2F6kaa0raPlPIYUC+AZcm7YD
XW/7npWahGkBnDiKr+TWp3LB2IjZP88riRPpODB0ua7OvPjKDti41pb1HbpPobSJlcdv9HRALf9i
coQvt/kV9160QBj3MJAGRdPEvDKB93SJEG3KQXFTutJeg8MJ0aLij9tnB5Km2WZD65qDN0wh+rPf
caQoIm0SwJMJUuroRppw4P9Aw8FXWrgEb6EGvopq8rp6aWpFqu6fjiOIZzolh5D0XAX0bjaik/nr
idkIxh5n4hG7DeaE0u11ZXOyFgV+zzH5j3bcURJRjcPZxz/yW7ecrSQFmJLDiXGwARzOZ2seMFnC
pEF63u4U1hsb22aCTt8wRDIStRHrO34VqGz0/zxCd5cfrOlbvPLtGT28t+Uy6PfciRB49TcpCyuE
9S6y9fX+59t3pSK64xUVlbzO0lEiULO7/7hyBbqcQNiCnaOehX2TF6xX1KkKBBhMfHLPqxtktryO
ysg8//6+HntuQd9iUyRxfT+TIUn3tRxb0Fr2vH0yPg/uiYEFXjPX8RS1lGKQAiWt5nACEezMUPq9
c1N0ttdOGhxOaFq438AZ5gEw/nuZYcFO7NUXUUCT8n2n6daHuCTloV/oehkzozuQnNXjqG+qMAG5
iyBTOAnFHAVIQazS2/Da5uDC7I0IT/BsiQjmwZ5HJTOEIXRN7J5GrPho/9g0sL+KuooBXL6b56zB
UmfORJ/eOdnbPHPcBBPKyJ4WE2/0kjzJCSJ9zWkPozJOO5QqpvnPXeGYzb++jeYeQ9oVVgiOd4MP
FlkIr+3nsr83zNPvATdVhAB/QM+9HXuRgvF+uz9oNY4rQ4VN81ZEySIEUtViKeu0bPSz72Rxxxc8
Xh+fy85CLWXggj29M9pQ0msVrNwpFtDACRLsJ9nLgEeABsnuZ+/23d+n1kM/nOEa9wrmSQZzjU2U
EihSDF1ejjyToNP1hkldWsl+thAA6qmrxEI48WqTmBs3WBBUm5LyE4cMmLO3Kz/6PeLlxeKE7+YL
LgNGEWX2ssihOg5zQNkikmc3aSJe/94MZMmsk2XOX8Lzzu9zG86b5HXw/+/6gffU5dowVC7jyV9Z
nV9MQf+YPkbOuNMPTRTz3hsNSG5sGXeWHerLWACP9k9wqpqkGw59uZyYLHbYGhhbdyGBD8I6ZSZI
990+2vUIqpZt4sMil06stxJMg8Ftkg==
`protect end_protected
