��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�������B���8���"���FE�Ҧ�@�Q\_������C]���5��1)2���� hڻu1ǯ�C�ƾ���kT��_W�p.=�@�0�l!�\�F��'����e�4�Cd�����Q����ǒܝv�D�w�l�!��V��<�1�U��Տ!E��!D�6�4O}=E�t�ՙY���#c��$TS��.�4`1f�ZG%�?T�k�u�c������rj�>�J��h�+���܄�k��cFա�T�/��^:$H����zSA��.+�~~oav�r�6ڌl�ɱ�e�y���12tc\ ��P�,��Ѫ�jM�Gw(��f�`	�f"���0��Sÿi��s�?��!B	��g��	��r�I��y`00��RՈ�Ԩ,�@]D��R��7;������=5j��Ptz�"Ӽ�oR���x�:�&U�[���7�QF�4�uT�v)�q���ܩݦP���f�u*=�]\������sk{�������-����0L0��R��5C��]T��唟�/(�Xl�42F�PM`~�98����*~��2 g�ʀ�qh�M���+!��ʘ������^s�WM�C���VH�#���ۃ��Kxk�@��~q��e��_�����l���*2��@И�'�|:�!2�j�FجA4t��4�� g���(�@����+b���Ɠ��[��xtO�?�_����d���N�D����8��@�N�}��'!��敏������W]�.���lgw�!�_ ʤ
#aĐH'��Z�(��/�X�[��~r�R�߷5�ϓGh'�vH��I�f�aJb��%2X�KZ�Ɉ��&�p�)_��#S��k��$N׀�7����+]�w��4-�Jǲ��{�p�U%�B��@�R���,�!����76� �#��"Ų�:Lr*�{�U�g2�y}��Gy`���D�����MD�F�^��8 �-ש�"��:8���v�F'dh�w�� �zÎnpk������)�6B�����by���Ye7i��3�����z�����'?���X�ϔ3b�?���9��d�.��틐�/|�u��q���L����]��A%���}r�~tN ��l��ü\tZmNsd9�I�,
�)�Dvڲ�3cjd��Q���<��������f/-ԋo�D�������<�M��]� ���}��=[�"�G��"�[à[��_�j����/�d]hì��-g��Dwؤ�g�>N����u��.����8��� >p-+�se��+@Ԏ�u����8h��m� '���v��MWϺ���d:�D�i"U�d9��44�8�ol��^�"�r�fޓC}�茉�^�u�B-�	�[lԻG�4�Ǵ�i>dGbQ�bM��zL�,���nY��� �h_�hM�õ/¸��$�ϥ��i��,ӒT)A+���r����lnd"4��=6c�$@{琱@���4�G��w�x2BЧ��Dw��؂X�%��t�J�z�$���IeKf*��v�:�_�g]������u'�Z�3�K���r�؍$&������ʺI�.@A0Z��}� (���b�M�2���yG���?y��*5��O`ݷ4@՞I�i4t����c.Д�s�Xӿ����D���AR�U�S���V	9����HZ�re8G�������-$`�-'fo�l��� 1�X����։�qG~7�^+����t��(�4g�n�^,�-�>����TU	_/4�
�)S7���oX�������A@M��V@6�Ϋ}�4�=��2��Ruo�N�bʔ ����FGr"���>S�i�L�LS��xUёrw� �h6&��oΨ�Z�߭_X�3�]�^4� �˓OS3jO}7��
�3�;�_ħ����ЄxLN	���@w,T6x"�[��'|畾�ȳ1�E�C֟rذg,o[e7�䢫O?�k�7N�r���ޔO')�F�'H���Ӥ�ܣ���ػ�-j�Ҷ	xr_��j���7n-�hdɒ�4�L���}Z�)v:�Ϝ{�|Bo<��������F�I������J�?���2����9�?��dvSי�����P�kօ�oj����"��p�`E�
sXa;����F-<��L�ւ����n�����G�#e#j��{/�< �`��q�6cm~ �v���k�5�R��ǂ'���6��m�J�c�K;�0��r����t��jE;h� L�"� �j_c��b� ��5bX�F�l�s��/���
��-]n��h���bj�
IS�N'w!�Ӯ	��vp�;bM�q��`N���=.k���
~OV�F����5�!B'��8sd��,��2C��6lgf�}�ős�Y��GI��h�zЯn��Q� }s�l1��.���/��g��B�N�<��#sf֟\j�J!R��|q�<9@��~��P&-��y1>љ7�?���l�g2ߊ%��e���=YJ���\lζ�7�����v���v("���Y�e��J4�Ov\Ȼ����P�8_
�Q���c�`��|�^�W�.�"�۔�W�N�|-cbOk��2�+���+W[��!���.�ýw��.��r�b$�<l�T��i��,χ��З)���y��X�v�Y�L�^�L�^J3G���sF�=b��x{%��n�~���Ob<u��n9���U�<�eDs�=�:��Or��T'��`
��W��_��7�?�����'smA;݇f�n�q��J��=0���F$~��f�8���]�-��5lc�=��5�~�"���Z'X�6�����Q�`�[Z2ġ&u/]f70�ؽ���A͐�q����j:,��P�|t�pR]�S�gy�	]�-�y�mE�76���W�ʷ(�X�[��m�lZV�ձ��ܓ��*��^~�7'����*\�P_�ޮ�K8���~�+����Q��8�l܊s�֯ϥ~h$�k����cX�Qx�)�$a�[L#��6��W�s"c��DQ�T��;�ͭ�LFi��\>����� ��}�P�"���f�e�UyX���5�І�>��"A�̪+��d�����F����h��p)�;���Ͱ<�,��K�$I ]ee�c�$6��3hp"����\l�ه( K�4D����a�$����QR"�/��=�4�Ad��<Y�b�6�@���טF��Q@J��W���I_o¾�i���K�
1 mFu��ZF�#-h{؅*�����=u�HUB���,���D҇x�=�C�r��1¥�"P7Z5�U���8����K8
z����=s:�fdPy�ag�&
�{#]����Z��n�>����t��su���H�!���5��`c�uZg�!�����(����t�^�dh��F����Im6ޱ�
�1�0!1u66�)oʅ���K��z�`Ih��MH����|^�s���V<f
�ݖ顤h��B��F>�G��ܤ4��,���vd//q¯?0����w���[þ�³�:�
�S��E��|���V����o�
��',}Ј������Y������ "]N�hy�U����XT��#ˊ�+�_�Z����!�Բe�a�P�#� �j�q��Y4r<�|3�Z��e�k))�rI�|e>��s�S˖q�Z%�!��,��=s�J&'x�BV�\�5eR��#b� ܦo��*�.[������>����a�&���Y(��� v�d]�4	�L�4C�m� M!o�0���r��jm7
�����#��9��װ�{-�TJ���	l8�����-i��
/�F��5�߫_?�/JK-����A�:�{��UP�ְ�U�YQ���M�r�Cf�$��n�e��8OT��~.򔍫�9Hy�X��?K��I��mT�g��gG�|*zG��0����=�>?Ē*Ae�U�5����\[_t�c
f'���05���;nf,��|�S��9RuI�%�"�3i�C�S�����N��,X��/����ZɶQث4�$�u�}�#�s}�F�W;am�����O�|cp1�q5]ĥ,��7V�R!ѭ�C
t��:����
7d|��L!	��/2�l�T����$�Z.��Y;�h~U�'{��^�3�}��!T[`8z�ˬ��~n� MuН}�g�/�ס��{�1!�� ��%U�l��_�W����;����U<g}�oRP�<r��A�z����W�FՌ7>�xby)���y�C�����Qbj��슇���{�4~��!"-��y
n���9�B��c<<�p[=�AxswIX.T@�ɆR�8XT�D����V�Wo�ҡ*���\k��ad?��`���:a�K����I$��a�E�R����j��>�xd=�
)i\fVI%Ig��O�\�ǉ9����q ����a�w�����x.v�u��c�$���G��۟�
�^�;�MGm���$�.�t*���b@,��z�n$��q��7#��r����k��P��Ile:,��|�Wб��L3��e��_4��>����8n%$�uVTYO���ge�)����*6�B��ҞI���U�^*��}k�Hn��ν�q�ǎؤ����!�P5�L%�l�����y������0�*s�x=~S�s��+<��e�Vc�u8�%����*s򊱱�
�o8�p��9�іL~����/^��/,,�%a�b����Ջ��s���A��K�$W]���Yt�����i�+ꀸ��Z%D�� :r���Îm�d#�B�U�x+��"{�q����o�M�ƚە��ZU��H�Ќ��9��u�,ܾLz+�bD*���g�k�A}�9"�E��~��ݡXrEq\p��7���)�E��¸�3ưw�Z:�j@<��?-��@���F�Ȱ��ӱ�1���J�A�Z����}L��r`��)����=��D݌W����Ĕ���L�T��%ʉ��&�]e��'�� l�k����{�I���!���3u���0��Xg�յ�({�ћ�~����>�KÊ��od��C51T$B�lZ���R)�7LY�)8��1ё�]P���� /k����`��GC�kv�~���XhT��k�����k=^�ʙ%�<���@�.��.Y�;L}����6_�A`��� 	�1Q�8l���l���#�cI�KLA�jY�
}|�7�9[�w�����i�����C	F�t��;'9;k����q�oH�e��g�e����tڊ�P� T7��2'h;��:�I4���6W"?,��xU��%�d�g]�'!b_���}������4�0���j�Nր���4
i��,�$��R�P4U�����)Ğ#L��������[:�$9��3�
�w\�a
���5��'w^$�#EYۆ�s9�7��lV��V��x��A�Q6hz���O�P�〶���Y6��O�&o��'"N�S���hѮ՘����%&�;Y:�&��!j�ڽ��I���� 
��5)�]�ٵI�$V�gv�N=탛u�pDiNB�$?�U�~yG�0`I����-���Q���s��yB�_lm���Ԑ��^d�����<�fC�T�����P �b"ns]n��c�@p����96�p��wbZ,9�v�Ч���[I}U@�q�F8#��K#�Q�|�KUs��h��Ž�#���%�Z����JŁ���ޔI�FIp��!�|��(�/��I�g|`s�]�? M�$�W�ʳ\|�����N�E$���lW����cpOɌ-6��^��$��>�l�fXE����c+�g�����ً`VD�a�(�xS�P��!,#�%?Wm��C���_��SI�U���q�Vu��Ho	�]V^`��Q���F?����9����8�m~.u�Gȷ�=����ƅɲ�=+�<@ϸ}#�n�^������]�p���v<��--}�5�hJ�_T�X=��D��?���5���E���{���7�@�@�9���d�2�#���d �|̬��h�E�C^;R]��n��פ�k�8�M��:�X�s���2�\�٭+��ԗ���f��1���N��Yr��~��\q��߮���9�.��\O�t���oA�$~;��O1���s�TS�;��P�@q��C~�ao��:�`d�fC��>`�����ܵ�a�t�_�X<�1kh�<��q<RԳ�E�a��EM��
�,���sB����_��zѥsy��hʓ#��y��J_���U��*�4ĹA�Y�L��W`�Z�"(�x�5�"?�5��oj�|'k�;V���3��T�� ���lW�vv��v��rM[�:6�~�e��]*�z��IY�j~�u���M�Ç/'H������~F�O�r��(��`���lB��]�j]+yZr�6�n��M7�^/���
�r� O����R	�C5z������7'pĭ�?�_��M�]T�Gm�@P-G�a��m�{29��d�>�t��.$.u�F"'us��Z��� ��
yB��LJ�{hEa������%çN�s�ȣP �Qh��,_|M����Ӑ5���mw �S���"1$���Ϟz��;j0�d������Rs����h}�ì�́��%��b&�p�����#798�l~\������γ@}��@{^�ޑd��$�����wF@jb��c��H��_R�|΄����="�l��diISW��y�d���k6��[u����R|4�҅��Dj�J��ҽ��i�h�%��GZ���:�����Xz.���h��#q�T���)���