-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
MkuRnrIxq8FAfQwz1OyQOOMqnlxgsGTCvOgkrELP33Zd39nMq9DSc9aYhGHDZnCA
NhxaG/kJwTUfI29WRaUWny08qny+CHzpx1lyKum5GAmWZj3E9q+wqZnNpkD8j2tb
40QNcpdbxt/5JsS2Gj1BTmo91R/j39+D2sUQSbrXF00=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8032)
`protect data_block
5Uyzle3dV4F+IOI2QrNST2k3Gs1gynj9ZoWCV9y7tRiagJs6u/rU2+w52cLSmLWm
cJ9Ih0N9ULQNactjJ8RbKfwcRaEhjhb7lcCGeSifrF48Q2rY6RoaIMHzl/V+dnxt
CR603wncK+k/821q86iBFYDpGMIWYJXq9couOSvBxeRlyxRBhxCTdjpCjZ5XA5pA
2Qa8bjYUC5C7dPhfhCy5JPVuwjtO58V4bAUDCRpVpOuHrMkMxuWHLitXKJftR5GV
io5LXbknJoA8GsVxrClf05RZpG+7feCPWyOHioiGSx7i8AiWD1kQLvfr/dXB71Ex
4PxuktwCbwyAMlVyzGpOzWp6qF/FeqHni+kklHhR8lZHJ/1fLtrZwMjDekMuIljU
Hl3hqtcUk1J4YEpofMEsj39rhZOyOpeTHXBrPQykFGzCr3GVLNwKHPHY0zVbHCAu
eKWr+YsP0WgP/qMQse6smiR2W06iu5uisjDwuo1yTry13WgQ78UMs4Uc21taKVzR
le+Yy/lfsfZuEUPkg9ldTphHCqs2+wgXrc4kyJgYMkYCcdicrZBPzuZmV3nJf2fY
h+Y3z70Ua1NsJeWWprLDQhfAMwnIzpJPXZnTPwsGkNewHJOExFPoh7AqVdLQbb/W
K1T7O/STd6OB58sUUcFL3fN6OShJeDynlZLayzHWqgyM+tyxIvKRzerR8Zb/4PLM
j9hxBaugI/u1QW4m3im4lxjg+VcXSPP0CkUoZumkHq4M0/8pfXidh7F6o4ge0n3L
qFEic+iaIpt5I23zri25Z5bjfMU3Z2UGoYQs0cat0XkQcPRYGg5zC+beEtuzuxaI
7Xvf5LgSST5IKFLL1un/TXjfn3eCAMc4k3z2SQHp9uoIqA7C+3gTPQRco3dktJax
HmpLbZOB/6tGai8f0kKPPBY+/OmzeGGAbunnBoJimEojQRtXjyr7k3yXM5Q0zWNJ
3lMd6fgfnmbmlcgA/TT+ajSIiJ0ooN1WUlcFBogTnvomnPrwcTIjkwEOs2yncZqW
cuAt84xxTzh+JKKluBwGik4V6GATw/Crvq8uMCba1SxYje1tP5wxA3l/wdIndxWE
8vZ/YtUZK4WMfTB4KVOHsb9b2lju23PNZFSk7wQDdL9BaZXHaK+3dWbmOZNmbPSv
eo1v+rsDpNR5Mr/28OlJUv9C6s0Hdc9uLM7TvZR+slDfd8x++WLABghc8ESrvgBz
3WqDUiD0OGIvYyCgHp5AStcffLcCxcIz8DH7oaINm+F84dMeAyyImRGv1+WuPFw5
IBnSIAQhIags8EBbmxGGkJIUimXtV0KJjOhul9c7P/3pyPjJ0WqZ1bVUmgTSPghf
62nHjksOg5oYeVm5HB0YOpSuMwqDnOc9Fzwz+pINIfZTmLmjig7ibo7AS/xKgF7m
ES2hCp5CdJDLOqIkELP0qN+Kg0/tKFwkdDGDipCinNP2SU9f09p4yKFA+CkuJ9nw
vSp7ODX1GGX3KJSt0sAXFUglGuaPjwt8mdmFz+lwhfZm5ayvKrDdUOEcxZ9W/IX7
krRdDBvzbAQ1Br9XNqqQ3qblXRpQQyjqU/rU7soG+AIDfJY90sGLSkC5ud0UtH+w
jjnhexZtHyxWMS7K69BuC0WmeXS4hJeJlfj9OPre+5s4HPxpIsugxuv6t4VXGx1H
a0uJsjtTFQFNFy612+XsWFzDikajug12Z9hIsEry/MNlyVeE+NgHGmDwGw9XwIki
GUXAlkf0LEWUsHGVhNtik8J276PLN0Tpls1Yz5rbm/AIY0IuWjwVvNt1rWKknSDI
1VNRqjmvsyGiZ6QlNjVMiTnzMutjiekQiIzFHWBNC4d9XrbKvmNpAh5saPwRloJN
wajbgjp2BclFUJ9tt6lQUZvYIsvP9sT2wkEPUh3TtPaDoiAwRrL3W9nHqMPvRB42
wXY7JnPXlCHwrgdJ+CgtugesN6pgPsYmPglVK0DTIJz++RKr059DxkryHF2qxlT9
2bTkQ2/tdHiNHz65RPrE/yZtaaeFpU6v+7axaDEg6dYN1MblKRxV2QTQWBmecSym
nKLlsmnPSPRtl5VkB3AKYn2/KZWUZ3GXONN8097u2RB+WGDmj8mB4vPbhmBPpxCx
cciZu2/8Rm0/ClA3NdtD0FwDde4RUbNd3eDIoobdeK0WgMM2rNnMAGCZHIHBzLXv
85gBNiqk4IsYDoDqbUc5qFDtHI3y+cXO+SzfD00xAkZWn9NRabp+I2toAIdk6BJI
11gqrlm6cop+x0OOGKmAib8ovsRnQITuqb5gxB8f7nO0+PC0dt/4oMJ88UAoq481
eeJB7hdaoMfdt2RCV+8oEhc8CTVuyCzLfOQZc9rVJTrKSw6qWVWw17Qm/UlSBNJv
INsrarcvVUHJ2SmCZpO2ljjdUUjpjp/1h16sHnLW6u5tDFhjQ4wsiQcbxkj4PI4C
enUOPxK3uGd9RlRkRphg7PUTaGqJZkMUZFbdwcV1fIA5Xk0kAsv1/TWKRabBZooj
tOow6UXxDq5gjTOi7L5MToO9+o6itmHyTDspwWViuXrgZbXvzOIHkynRH/sGEl9a
OdheH5AE33WxqBPgoC3VoSuihq0n3qtX+8BO6w8OM1pkiTYy5Udh9x81pptTWlwf
TcMG7mNwyv6kTvtGxugC9HP38uGMyMCrRV7nFMg5sg5YescQi0T8EUyVaKegqp3q
Sr5tCdoXyOgad0y0RIZilIEoxUTdSrP/WSts2FzWgUwT1AbLha5tiqzS8REyv/T+
YnpoN4xIRJPj2q/WcTskGclHWAZnHPx15hoB7DtyrgxVmngwG7lKs2qXAo0/WxUA
2u9rNM2+34Luug6+uOSV3eYyzlL2+d8SignhXD+s+KVSDmhxSNuF/waTmdGJ5JMU
eNiZ5OyXkbPR4jsDYSZhg2mCOGisQUy95c9u6TDWpTZpLZdKsWeX+b0E1hETRu6W
soj/T96r5PYFMRVnxssH9QRqH6O6oGpzIVKoZv/pQ39zr6Wejakna6ECp93ZpNJG
a2JWcWpSpKA01biZO7Im65ZGGIJKY7fsrSdJa3EAifhftIRdsuOqeldC4rj/ty47
ps3V7Mj2taP/70yrF1SOb6SnhK1B9dUcUnPfTKxXknUq86YK+BNqN4C8vo04P/hu
RBgA/q9jHywmEqJR6/xkHB/bZvDHX5baSwbc2oxWPcfx0Nm3euUXki31ECa75Tpp
DGOuzRzcRxIYEOKWMepKj3YYKkmYOSpIMbUwlfXp/jYLwW+QDcIY4wEuWUxOKZiX
/YffmfKGFIjBd8fzloVfY+WMFmHOIVsnry+dUu2teGaVn6Lepu5V8UxeAgK9jeuM
/XKxYfcpdSHxVhr+nPEhYOEmSXXVfnBArcIFg8f25uBkrnp2Wl5GOptt0gEEvUC9
rWL/Mm/OhOzCwfRapkzIq2e5YXIIs6GbqakygcmY43zM2BChO/H3A93lqa9rkwrh
5RU/0YpBuqkytWpg+B+7nLzOrdSaJ1SOfPgY3yhtACODGLOiGtTpeijG/6jE7sX7
rxwo0MxavTlBKBvuhTJRp5JlEM9QKKOwW+OQd4Q+Z6TBuo5GBHitQSelPCbaooRd
KQ1kVqTsT+l2MySXQOuJNhcnwH9ljjnu/Rae9aRcr/noni+rkT9ljsqYXQoWzUq/
9y+lWiDmIEfGGu/QKhdqVRA02gntwOQweNwzgVBXVUMkEily1wlHA60GqZ9TwTcN
EjMhYQ0A+GDwzpqTjpzlkFzvWQ09x6Y5IisLFptEgF3jGQuNM/UHyD5NYsClIgw5
3PIHl6IHgr1hLq2srnfMOs0y6ojAeMJCLtkSDKV5KSABFSDDN1pqxzdIHQElF+t8
X9w+Qgz1Q/pFhGanssgY90GOcRa+Jagdf68wpv6P4C3wOqhb64sjjayOs63SnrcF
D+lAYHeGrYxH/zAlC0q66JdcG0K2BGFbjo5oz3NYbwb3yF/4wD1BBhSWx7mUdXhD
maNJRhjY4uKWth+RBtv2BpJwZwEUHRsbpMJCI7sxaGs6F+GdZEsRgVQPn5h8bzv5
reRcujmk5aS0GMiKY3sOnKvqSOsmH1rLV8A0VBkcS+exmw6knlVGjQB4oiA1QQBZ
jGg2HcdHXLyCeK6YWangKhE/O8/DYnPMLHhWC7WoZ7E5Juu2Qap312cbgITIghev
dQEKdl/kfMC26tX2gm2Ix5N+SC82BUblH9FIvtXBDn4ncErwO5RXgNTavSoxKVhZ
rMjT0TbkEqBxMwVMkv33XvX39ya0ioB/dCqI/ecM/PvuQ4bNDSzDzhtByEC0l3AZ
HgYVM/FoEyFfljyMP8hPifCrgphRv97PB97ifpgBYIZfONpoVajYrofzHYzPu2qL
eddoU61d1ozSRoNxbd304q/j5A/jcHQWqqvllJXfGJYlArNPYWCot/ZiP4mDS76/
fE4JxWIKI0shu7iEfyqUx7eCKY+Q2YFHclxJpMNctlHFt9KOsmOLFmscPA0QhW7A
h3LTXL8rq7Pw9XKPm9TbdjCPUX1EqMcIZXURejVDZHO6rslwFl0WDJfLyh9HnWPh
VmCM9pRlW7Jg07+pF63XpwxPxDEVeJxv5urZ2acwFTuS6iHTRisqlLZqtaWVnlxJ
hDx7jY+NAEyz8DdQgEXRanhKeEVuQ2bi6wwJQi1nxjbIm03fjg6WdWn3M1ArogCg
Sa+C/82vfDmPrSA1xftRy/JqkOCfx8D54BtwcAQy92cNsoyxF/NL9kkBGL1zw/3z
va18Vk7ajh7KfEGqvcCj4Iq2jZAwEW+8xmolPRiV8Aeun1/N2rmryi1tdCostiUL
w2IgaKc+yGipMYTZ04yMLFrBpmhnf98XbQbYblRS/imDHPlYn6Hnm5LdCf3s9PDf
bmJJn35ejoqKbVDGjPev5otZB79gNDn55so3ybMOQW8Thh3pmDQlNzUFpnq5prXv
sJsBBH9Ogqoyg4BnxXwgv/CDiJequ3uSc19l/fc3g3yJT9hfaFvrV4q1LPNbSrmX
qdHS9voqIuiS5lIFxk9PJBk3D/gZ46cHFiH2L5Feu/TivHhK2775qQPbgjoDTQ4I
ELUQoopyRB/uaqbVdFlRSsWqaqt4mqc8P0iGq+TdTuazx+ur6ocF0pDGkUHpyj3b
zh2xYIYb03PnuBWeqEHGtPHGNex9gaxREOVihBo1n9H5/VVJ6ZzT2gEdxgKPdbO2
dgZNDo7R2YRz4b/BMmcDrADNH6ypvcdC+nZaDQlJUWDr2+nXiLn0piUstkWoW8XW
5i5MApCyoSGblvPA/MXq+kCUyXPXrqwt0sh7LsTCqA0Es+yTkvHNQ6UNseSw6m0D
yV7rXTn0EuaqV6b3AcLAHrQFJhkup/M4M5/kEAFOjiWLHz+Vgv5iu36DOBD0u5nD
fGNsF66e5kNy/HiYrorafvnNy8THUumVJrqDIGquxkmnjUbE3EIViYOQxT0uG4Lp
E+7VIzUjggXH0DXR+2+FtVB3yf4NceRT08ekhyfG/HCLR0Yg5kfCVfqWu+VYh9oW
4foQRsN/NtEyytQM4kN3yxtQHwrMIh3qgooP8Htjs01fAHesZKiceJhOWXdteKJt
1mbY7smfANpcAeNdY478nnKaqLAjQscKwEKNcSJfjlLBXsNSExINe355q/X0cxCE
4RKrt3/V4W0lyMyuXY5jhrhb/Loq/KDP1NOTDVpcsMDICTRFJR7Nesb031zlfkux
c6yROa9TU+XW3O6ZXirk7dtmD6+siHHY50y60PrVZGn9s4/9P/pYmg9urLmyhVvI
aB8QzBArPlQflUwwXATELolMrt5PVK4Ebly2QbaMb3EJ/EQt4qjHPTDluguoiwDb
tLW/s7FZMeua97j/lBDlicHY09FBALlYVCq3h9s7JwBoq0dao3rCaRnbrb/RxLzZ
UBfVEAI0zu4ZaVKdIYNyAOXNKK6PFBYsTOIe8tL31PfPWChyjb3DbKNERIkR40KX
wdZJ0KkGgD45WRjOXYzd3Ebp65igg9HrdLV/lxhiL6VFiNn97VXaCU1KDzRj3c59
O43CdJbzkaSEXJaGQeHDqoUWqJSZ51qvsCkjPGFFSpIG9aLca9gpnOCbMZBiEBkz
3eWin28GV3nqV8gHJRAX0V1/tr1HotccoXfD3A64r21nV+A9HtG++X0c6lKcYQZm
b22olwyOHlLAFZQC2YdM8fvKkcqhUT7AwH2ed5RAejdMAwB+MdfY5tK755RlL+aP
WM4fXvdHhdtlmPO00uCusTxh8BDPnzoxM12HqnHWrS36y0ZGqRRh979lxknjyQuF
xcbYVKXXjYCGgLEgYJ6iFyo5CZJBwVbCeVKPJRLZmMxwW2H96F3cnKksbFT6bzUk
vLa1Y5HfXfpcfSAWrvUfugzEkxK1QG5Vj+rm5xRu4ZyAszPuarA1DhBezv6T9133
0Os/a1FFzPt2BQiqcNIpQlQHNhmqY/gtRFtIzpbfw/XZtmQRRyaLPAuWHp7Ow5h9
HICkcPRdcpIWoApm7SoBmOKHQ8Ev6GOFKXDpwjaY1ObrWaf9kJLSnH5t7SvlbbO7
Ex8z6Khp1ji9elD6ZFyc8IzLQ/bjO81amKbPunwI+VnxW1ceh6+bw7C0JESvWVdT
PHOzZVNrxWlat3VJx/OqdKnJLBmU8BBXAa2vRKkOScBf7KP9bnTklCpaw9cNSHxy
xmrqyF9g4auUeEQjdO/iDVY1ruYCwqJtr/Fa7YbktLAHT/wJX8m4Z6QpXEaI0VJq
EcoMPsTJQGOqMMLLTz5k7RL2PfSwOeaJuVvgUl9GvVfNod6NAJtXJer+m8Mw7u0U
5h+Wgqt/aA3LE2R8Be+o8zym7WAYWkDgSj3ySo1Ki8l1pmVWXqojFvn2DeyLitA8
wpvoVzrEzbhPwIubFKZ9HE3gM1xSFFbKPwAGhiv5Kw4GiTB249sqHkr20dX9sYcl
9JYe1UEjeehsNlSwHt+EHchXbats85/eqxHlYXESBpj8XstO3Hu+jF5bkPdQ7wDz
Hw1YdvpYNIzM+KVBCGB8ZWM3F46cI+itFetm1Dl10RLjOg9/DQ0RouHcPuTlLXbU
7LytvU+IL/mZuN2y8CQAuCjLvnbe2uMDLCqY0QhapoyImM+w7PbpK20X45VnGje6
eHcMEjFbXMNvRzwS9BHEAiCz3HdGNd7I4jDOZmXSlO882EJp9a9xzgfiFxVttLn4
7btugXGUj0TlZxp+bb4Qvhj7rInCvH9CJ8nbnuRplc+Us6uHi9CwEf6iDtzN//Rb
GKm0y92v2+r/flg0qqT1BfG5rT1bQjtgSBQVwh+rNCB2j505qiK3A4p5K0MF2qdw
xUDFjtOuPfYpST/qRAIjgOwobTs76HxJ+zZonNCVaLeXX/Do+va7mzwBc3CmttQ1
GvzlQvfItEanXof9VHWbvV6DFecbTTtGVG+omnt9Dpe34JOeclyhdxJkF28IIoig
D+V45XLonwtdlre22EiggGNNy0qtfMZuBdiFlIkwC22akC3XRjxkhbnX8tOpFc9B
Sk4PcXw5Q09X+t7X6fHGV7TfihlREHIEnqyadCqaSl+Yl0MAUhnVVRULFHbLHtAz
bxoSREee9B4MBLFhw+tVSDdm2wzlAcnB5RloTvYgUYcNvOZ9SmhZh9pHxMTkwaoN
JjgCsprvuJoZlHwDx9gP95qL+/Fj6f077+zRbswXTMnlJFNTlDMY1fpMfeMAVoJs
/dF1XS0osrLZh5FUZ5xqLHaEF+LoT3DwE2v4ksPP5+r5n/nMiqcIsrfZ6NXpinzu
tC90EqD65DfiRjltWFodaEf4piCODHQH5QNPxz2W8lAHrGrQVveaJH4g9OSFmM6w
v/9wqm5iczIrxIDdcttu572jNYQLTXnE5JorMTRsk7eJV14yqxHKXtZ6OeCQ7FUu
rJ5qFd87C822+B88x8DD7jnBo8aBL7paKZo+5KFHRCqeV///WAnGO7HgwUGcjSFU
1KORNLhV/kj6RTpRpmexntETK6QjjENsTeYzbad0We7jeNKjutq+7ECsyLyfeeXq
rK03LWUVfCJDwFBLPATbo1mlkeqZkLXx781JmFH0H0wXkR4g41Ub26zk/7B8C/ev
Lz5BgtYo5MrJkUBYRR8oKjFx7htBhK4JTN58MXHI6yCEdsqXo1n5LKbA20CMAgsi
nXIdB3EeYrOIrAiYxJTJDIVkpMMf5Qs3cQI4YYdJ0Br7MVO+hnofGa6qsxFN6cwP
oVR937S/S5f+Qgn4Q5khsu5GI6vH6GmAZEvoWVQprR5Rimktn2Vmfk0sOdF0qrMG
aXjVTgTLuMeZA8Q8RHPd/QbUQCAeku3Z4eC3kW8zA1D/pTguguG5TjXa6W4Bb4Lb
TzV9jlTScFQoj7wGkqJa3X8vvSEBEebtcKR7TtofNm1mnoxrcDOl/E8hlS0MQsaK
UiytwrJIOMo8laLxTOoUSJlGIjh+Q974jcwB5mR2Gz/w6iQPTmonDAkWERHohV7C
yUR7TjhY/6jrcpIZChiMVpQ+6XwrvZLd8DRFKPPjxkTWmlYecvKEb11USA9r+n5b
xxZdNRQGpw3sa6hFfmMVaAZqI4bxKBVmeJCZj94jH2hGjcx99w/m24x1HkWxX/TP
SeJrT4FtOA7xBLx7BlDyM+/A6SET3TCn+E50DvulQirL4WKkcW14VXhDFRyy6Itr
bU89hai0NkuPWonQnXtbRo7RooYqdp0fQ7UFNFA+VfewsBtgL/CnA7s0Vqlb81ZP
AfjH2MMXrGxB5kKNk3NdWJLW9jtfpoWNKkvFyCUip4pa+Lx5/PXqylOYILpTjmXK
W+p330iyqGQX91PMM7iLzTEViKkAu4Ls9wIa2e73k6tPqN2eW32nS83K1tsChFkb
Y9Qennuhgl5nwBQQda9Dzn0UOcvCr/1RFXluVnhoJ797vnuLIwUD0fzlqLpcpFVj
Tghk9QCChH9HtOPcjhBrwmpdO5h80jt3l3BkS6alGzW42C+OeC8k6cBShFcQpuuz
3ibBlGPaaSB0i3CT1ORat0Dr0FKbVvDYCQapYjelf1yeExf0tbfAlJMZDKNABdMW
dAg8CskebrtThG0FS+toFU+uJzmdhOighlis1ZNlRvRhwQ6kj54kFyeOEMrlnFBI
oJ3hLKvhGLeiqmdYr998W6ZXDF02wuQemG5PDtVWM9n0fkCSVEDuedLx6er2XEQC
8GWF26nsw1vv9ZvZSyhsyRC+5LwY+aN1Vcz0kR4u+M8Z0bVSfGy52IrsQQaaw/lR
O+WdDV3Yiwtb1RCHz/AsmLPmAb9NVFi4VxyGsFtpfNKvDaXN++SLXoIjvZlkjdPX
8NKMoVG3WNernM6babd1KxmZqHjzZcuGRGW8LDVev+h+jQkKMaByb2Co2ecBpqtE
+LdRmTQCKwlOegkTYj1w0STm7jKC3tIsYWALZYnMh4MTxC59GIZI/djegBTYWm57
bdX3t7Badem5fP6QELF5shVXu9dEX35dKiAQ2vC5jxQ1HZ/5fs55LfBkohzRrQV6
gE/NfwxM1ckPiL9PClr7b1BFlFVClmdZZ0nvvF8vcwmsfxx928ka9ico7rmcyjKx
GeKLdl6LTpIM5TAED9w/e23wVDP+xOFjpoVrnaObeQS6xFpBrQycRIl02zECsPTe
o2/49ESRphgRFHIhu+XQ9yvC5/2RoY/TlY3nUGGUWtJRDG0zRRO3Dg15sIJo4D8D
IfT2qiwT5JTDXWMGUn1LQPUSad5fp5j2se2aDupwE9VN0T9NWhA8jKxywnIdKX1G
RhQ++8DNg8NaLlc+dXvmyahBTHJROjhjczyPZ/AiRQ8kD0yE1rGspdFcBJL3poW8
7KRhPrFbWmDv/k5NHJS7j4Grvz5c4aTwjdwA4wFr2h70mD9QJgIbaChuv3gaLFEl
f0EIj6ExBl2p7+VJBni384V2wZxV90YMviR7C3kvUKNvHdV5w6bc/O1bx7MVSCjD
q1WsHUVc7VfcWdqjx9IUYJJ3YiZIKXWwWRt1fN005Ic6iAGFrU0wSWDgDvOr2Rsg
mWND+hgu/lW5r2Wcx/WONah8BYxKojMq1MGbK2ROmeYXTEf3u7hzHQwFLzcvJWx6
95tCMfxCTf1rOCTlBlUy64tvr/NhtSsOJXi/U3xiL8gYVPhh87loFZpKY1VTLz/X
4/pjuQcYG/jtA2jMbdYXxESuBevRgcj1cwIPwwT8QKlpp+eC99ojaCwWA2PmO/XX
S2DnqKYnxkw9A1SyaNdUdOdY+szeglzHngkrb6W5EA1EScQgSVkDWhtl8Dk2a2nB
1akxRA01ip1vshABO4rwo5lW557lmC6CKmuwxfZClbDh0ygLpUrY61PB92thHhCn
zo93QJ2TN9vixvS8ezye3sb8bTJxtBHZhGgJrXQG01kL1udlZ596kFhN4btHC2iD
25Map0orOgPB3qFLvDNNxhwkGAozTMKTU0DScZ8hTpRu9SXHMaUSQK8Q9FZVhCeu
kBtfUqxv8FxLyUCCDOmp3Gf2SSlz6ntbcOTlP8jsMe6myxUoHzRJuGQB6uuLy5aq
20eBEndatFyToQ1tdhTGR93wV0kZ/qz5WfnfAYTj9hAH+j0cpw3+W2cdu0SZFE0d
7/6wmd0zgJkeA19I1NF4aS++qPYH1YWTHpOD9nFWPcQlxVJxXt/zL0Vu5xaOJ/dE
uDko+wlGy9fHg7ReUnfbrelJnzov+7czZ9qpizk4qT1x0ajfCxqKf3ILrsX6u98+
G09K+G9CyPBfXrCpexuU6g==
`protect end_protected
