-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
eXwq7y4ljKAkfB7djj79IvQ3nPjXbYSII719dCoDHFIXNiNiZYrr4+/Hbuf91WOc
NoSW7IdWpVMB4LmFCSi8cL8N4QeEOjmv3D7GoYsyq6Ao6J9Eg2A1Q2xPgVd4l7Fq
Jy9GJnEofSKtxXXK6IYdw3H8TY3LfY6l/uMWuubHng8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 11552)
`protect data_block
D8YEHwQG9mwWVthwRjZlGhfM8nu+G3UGeNcpHNp1B3zv0/Hnxhk7WZHNGfvEGRYo
K+u1zorUb7pwEcv/5wuQ8jF6XhfqSDCzEmKNWG+kGgbP+SaATAGwHerAYxMLNIKY
+XSLSRJb242EG2mpOLvqNANetOR+r5fK7W292YlBszaZIPsZumUiDtx6pX3zGg1m
TXTEra+Yu5bmbqgU1411t/erEJhaYGH8ij54FJredSDULGlTpLe88EcCaunxEsAV
jobVvUV41DWdI7CEn9uQt8Dwltf/0dqUJvN3W3ISkvMsEg9ulHQms9XJCxkUIh7K
p69lOchImTiNnhV2JoLp2rYwcxZFw8/l4Ed9FvAiHncMp8q91rOQ1XKDzFnpAu0m
iU+AgjeZJ6g549Gh+RhGCZ6hJgelkWXXlF578oxTovSKFiN3Z4nAcV5vCYlhUXb1
qiiftMU/lIyl0FTQ++eCg35AXwl99RN1dJcD5oK6A4Rd6YMLAsw9wkKh1Df4v2vK
o5Ycu6WU6nkLFOHxEXFV0uxOc+VEcV3tQrr4J0mdJhNCwb+V5esL+Mv6f3iCCuBj
JA6jLQdbkfM6BTWHc+2UVhBMT9uTcFu0eIENLpqy+vOJmrQtHKgkvIAN9/GXvVjB
VEbIjTA8NjNBaY+aCCiQGy8KZx/mE0sWPBpEqK4jRH1iAWYHuuMpHnTrBfZ4qdF3
WBYZPwREoL5t/oHbbfp5ZWUyiyLxX0sLGYJnGsXixEA7TgBk6aM4OQVsZJ1gTpib
39sh77v39o78pijjEgfkg9j0CZRzaEP4p/Pmt81uWBmcxF+nQUAQHayOK9odUVDi
v4ny7o4BgGbq173coRCLkTo1CeTUMSsckpjY6qVP5cEFbgPdbd8uB+/hKmoko0p8
iXU+KRi777SwxIjHP12aee3zo3AnPr/ziQYeYVJfUcYT13x6P/imP+N1htHmXnLy
c8V+dnC/rGR4D9gqcQ0Xo9dRdNNhpDVHaB3Twu2ZTxG9OSFdD264xi/R8j/SoBOG
An1bKYOAGtkDNRjgo/MEDs080FHold6da4tf4dGMygPpYZmcAPxBBV45bk6Vl7X2
C+1LFWEGzNoaubhnDDc5n0YxXdW/DGv+0yGyBcg6nrm7IOEBX4F1JcKHjCzH8Tbd
iaDKj+8NanzOCfFafTqyz/dOasG/Z9g9s+sVk7XZkTErTLGGiBlq/20tZOEkj+ud
gZUQUtW2dTL8tmZExslTzRB4SthJ8shYZONc+IRhPyVNTyVaHGSb8auaF4xahAiv
JsA2VEVtp+z/nOIRKHSNaLYKazKR+5zAS+QIXWCLrz7Uqw5tMPg0+F3KtkZ8qoU/
EVtCcJXxGAqfb1dbtNNoGjjwxbh2VgxzQJdVEE4MEfyzfKx+QgiBeGiyHhYbm5ab
ulgllFpaa3ail8RSSpmYOml2eqPtKz7En0kIIQdFTbOK7EeCJZzYECdBFCeDMAwq
S+ZiQYUphKe4qM5r8Yu8e0OEJUbvVLioWRlcV7Nu8WTpgV5CL+/nDRK7JX13NfFZ
8Nq5V5LKF3I9Wq+MsvhlrRxE2Oz0vQF4ATRgUQJLPxHqUSHajsEM1gG11+o1ppxx
2yy12ncZkEBuKfQb/F+xqYiX+Q6mtP4bZU7h4rtJ3Vyut0oDGU9fdNBfkSL5vGG7
FeivdPrOHaGwyH+gyH5aF9ZZE3KXlMPKdN4dptjnOXm+JBwmHqud4eQyadAOhIQ1
+3AXU9zXqfGucq5TnBICBCSXQJthddpLWHL+aVPhp2Pvp0mlCwxwMaFTeR5EdnHp
qgpqTSd2s3fiZc0AcHgwb5OgrnWm7IrQgjOCtu3gmyx4ZtdIgmo68Mk5cU631e5z
0mmDjXQzQHVdtWkB2qkt6rnANxE49gnhq2D5tdjtzzyON7fdzgNY+Eo2R4gBrohJ
zkHlOwuU0KGnF2EYpeejQCgRsSPDZUQrvPbwc/EDIw/bTds4n3jYEZueTMV2BSxy
FS5V5t+sPzgX4bEGYgpBl03/rpIoemIZvMVzXwr9LNXagrf+XQT9RCPFFSAd5URm
uz+83gcre9kFLye5nIHbt9I6vtHewv7qQdba3Sxiltsl9Zw53brrXvfuC+w0URek
xLo751WdQ5U1GkHn2cGQcuwsC27VJ9/RBvuLa+qQwUyGDCNHMGe+f7X0L9rboWUK
ftfexDFwzM1BPAVT0VEMasPNjJrp53aaqO8WPEStS4OeJVMo/DNyHeHMv1tMzGVL
JUzzOMtw3R4QB+mTmq/uFphYwdxK4NDRSsNplhgv2cTAIjtW747s0JmSlanMUzX+
CFCy1c042qUT2F/pOff8XlnSLbjI1YfmeZutQ+j/6lvE11p2vPYsKRvNn1YlvPl1
LLEAg9XKN+JgOIWynk1a8gRwDvJj0/oX2rwCmwhKzF7JxyVr25eoYl75R4RbzoOE
jdsY6sG3AyU5tzxUt0C2zspdIEz7nSDDsbXOlshJkqkTJVVvzn51e8D9m7wC0r9D
aeMapsDO7Bk9xiPCyYqYDf/aVfNVwpTIINQkOwea8eftHRAXmekSMQN8yxI2PD2j
TfSSYwbZxv4u0uVz7IM1RBe1K3ZwvMfTWUXeMdOHIUqAP3ic9UnyUUUKxmiYGEGD
/7x75nK+PF6s29lviQkl1tlJGg2lp0K0Pnd7kWewadueKRAAtoJxb/PM1wGeA16z
XEPmw8hxvtWjCh16GkYPj85h7obmEFYYCcl1eHMJ8IitQkYlyzNEeEp+9dN1Q0td
NCrVIFDPAORGOSFLK/xNN7RBJCiDstfVKVQdAWsWqzv+vKrQLsZStCdnqbL6GNJD
D6S2TLJ6PEX/x6aa4EOT0iKz/OJxVr5uA2JBNxTBQFFS+CZCeK8/9nZ+cCaFBdgU
1AKSYd9Opk37th1VisdwHrWRcSnBaoWX1P/KVfnt6rX9ydp+/gUqlS/SMauTYLQJ
d2TyfWnDUvpeWZq3xtHHvJk4WkzzPiOQq+gaVceh1A/EdFYRM7SUJvhHv3lkSxBD
lpOsf1dxQJzGMnSG61xjiPkugjTflGH2x4H9TOfXqhs0lTQRmJQYorPRwVHjaNU0
bPpY3mbU0LPZ9v3iH37LNSwOoVoHFw054OzEKBYmuJpCz8Cp61aE5BSmj5X2Hk4I
RWXcA1U8ec5oemKxgGB/sc2FXA8ZvWUFve+nJCJKB4PaRyF92hZyyGtbJnYTCxmL
30mVVzajc74bV/4+scYXuSDUB0D1PtskSKeNIbQB7wM+ypJ2Pb9G4E9+syvmlqwJ
nNPlGNfKhfHeE2O8O/Yp5DOTQ97NFOZAwGrVlBlhwFRvJO4VUSdyFHN342XXtnlp
JLNkwnbi1fblqs2YMH4dQvpCFu2XJhMcghaGh8kDVR8bQgFHhWAlyI7maeTtT8Xz
BChnmEoeieg5k0SyDKF21d50fYpS7t/gvtOG4tdlp7BqE3qkgVswS+iXpS8Jj3ww
p+UCFTnQvokIXq5m2t8M0erK1QA9EA0tiWBSh3TR7B11yCG0DRTbB4rm++fk+7kp
QGzVv/HLCZAEDrZeDv0EhBlQCUyAAdJqnZy3Yy5GJINecsHic+1d4O1uny4EI1Wa
hSjrk0G+fP52AY2vzh/yYMQBKOEtf9eU4sKYhozecxeI4ppv87m/bvPgXVSN9srq
XX7k7nK9r2RI8O7VFNQQg/9y8Y9RWj/j4vNjaQpQT8CBvGkQlNdn/tmBs/D4rL8J
uEe9egHh5Sb6fFfvOL1VpivxhH3RkiosWqfncfAbYumvibzbZqveh0UPV60TN+Qo
kOfEGmrIzKkBwLsIZMMH9prPy8FuN6oyDPrWI2CUNUWwwuAcwFuCiOhf/Vxobi47
e8xbHEuhKYBtbP7qwOMqHEuIuRdqs0FzWmJ4KFC97qVuE/T5XtxU9wlt26sv7Tbp
mb93hf/zwC2gDfjtDW228FO8kGLxDfnZ0ucJmp0ZpTP34Sb3fZGgcpStY//EbFbL
xfqth4we3KMwHlM+9eNmMtCk6xpMu9vWvaggzH+7vRJQIBWZaOTZGu+kU3UMrO4Q
tJ1KBJS+ufswNkxUy36oKbgrNT9Br2PPpAoxRS11HAaYOITsY8cAnH9bHOQnrDF4
2DDEyXyw1Qwl3UqJ6SLJssJeCwwzRa3f1a8oY/HwQwAzRrAUFDzarNBDLO0lN8IU
heA3SlVksekBT+nEwo9rSKhIyP7h6gHhsR3xzswDakmQJrhWYhvskCMnVyXY3n1j
GtFF9wJOx1GKTTlTyh0HOupdmCdu7HwbIm+5NbI1eiHrYPsV4+unIAYqvVGRMnIY
KxZhWsTGj0AzuXxkYziouGe0W7dhmeduvwvFZ6Zrk+H9mVYzjUklfy5ryBWQbEze
3IUbG8ss52PX4zg/twFyV1BTZmHCltbxwQ51QcB+BUfdshBE2IR8DJ1NXXK65GA2
CtykxhmKZ00NyWHod/iS0VmqntdUM8EtANgZ+hMdFJztrVWV+J9je+/8oKdpoAW3
t6NMTmRM5ZCDxcqpz5GQ1yxoo+urEAkhqIB/d/3ZD+myJu3HaP6AwlXWC448kQBY
FsNr8lCHAgFdXcfTfL+A38UAdT0n3SsJe1jeHPSUb27hhdLctDZmiuTUr71yZnmL
JCgDR2fEtgtq3mjGZ1xaFoaCU0IMcmvciSllHlRyrlDEILQKZktYvq368UpMfzKW
RRN46tgkzruxZYvhaGe/jptn64DDrpuUFW84Y3Ai2sKMIRXUoKhdguaci391xbDO
q+mzTHVx6lpsqF2WpA4KuQSzwLsnTrRtEP7sILNQ1TM3LhEugT3SctM2n+vq5MHt
fj7/6Zrw0f8GWllF4BtyvvUtwtrYrj5xCbx9+mpW0ILiNAox7G64mryyu8TCrW2F
ueDdJY8jg0Tubxnd9uio7pGEsUo2kIpNWlqEWK9lstuZIo+yuq+HPDzdkSfBFIV2
E6eYjn77/RxFOEWPzky4z+caDVXRn5j6AL+HsBctmwRzJvh+02cqugGtBeVBnvgZ
cORhm4eyO6ZVdcjze7hhJvZKmAwUyW8jbvwhkjX/09uK77j0bQLVF45wJ3IFxZNP
RCp+DuuD3RPOLyfPhBj0UJ1+R4s1h2i1ESm2il0HMxhg4p8HMxmh7SSfLc6mJobw
UkioIynmk9aSB/d/+dSq0/RvUD3G9+1mLsWTyVk2v8FbDHg+sHNe2I+BvwVb1QLt
WEzrNRpOx/zxy2YlNQkF/weAJ5HALJzHb2JzZlCFzIEtv74zFY9As1AMGblqHQpr
YSmmdPSI+i5bOkCv/pYoOMwaTX2zL66AhIdqmj7oUiPf4ZKOikIXaFnG5fxq4w00
ucqyoVNkCuIIRA2uCf8EkEYEMq7JVfWDqSRaqgb9Untwd0oZm4nc2ntKB20HEgIN
lAPhGjm4hrvVpr6AssWyICdLFJMM7g60YeAungqSoYOJKWbCpKW9OQ6/+/DYfxfk
S7lfMxthQGwN2QwuSzhtwRe1F1IY1oF7MfBKa8dLj5btTb0bRbhEdtHwGrlJ4dMf
NGt6uL+6GF9u29tsAOhzT91DrWdPTKQHPWK/dBWz0T3q131x+rQcW6IKROLPA3sN
dhuTWZcWzJE8NA38aA8aQ59MpVABcKCL8MOicZ6uyOyRPEQV066ise+eXRtCdJyC
pBQD1bqi0DRCeqEdpDLYT3f0ZNxv4AdMZupt/C+6ZM3cOYGBM3pybWs6cl/xEC+m
O+jdJ1CjIUuEpczpT72NtTx+9d3GXlG+akIJc3+Vx5wD2sOTi6BEMTwLcPhSYVqi
eGCKtWDdaBEkMmgf0gHttdrek/0N90bLq7dB9Ho8CiXrZDbpIgxQkjrE7+GKG49G
7nWIKDyzyroVYmsAYUqP3Q5okqGm0+GwAbZkxcoLkBBjokPg+2uWtyfBU0RlxkYP
fv4oCHrPc1w3FLMufExM6T8aD7ouUKUFHECBmjbVCemx+dhfRrkHjn/5h2ExpM9H
Sd5SgybxcepV1Kq6cSfcypGpZLoj4paa1LzO/uL4zungqB7+9rTjMxFStQQAT+zQ
CYwoYWaYwQdxgsYnSJ23gB6qK4y31SgGIuHrXyj3iFkhsB8Zstaqy4+KZ0HlFjrS
3WAheBeRxPWjm5DuHVGH3WU1xJdrCUk+S1uyOmIwMKrnY+dhS3IxcHWa4ZPVtNO+
n1sS8EF/G/YXM5Dvs6k0Q9nmm8oAPupxFe8PohHCwLx8gWalJgbn3QVIkNCQ1Y9Y
ZxY8H4lQ3gGOV15MernbllPBFGGXnQx26g7j4HMFPkB1fTK99YkgNrOGLn5aKl0r
cILNI6kGa6sbS1fqkFbAlQFUfxckJNu2xfuhlwt3wPiV+dyFd2ej9+9K//+uAyAg
Z2trq27CmRJrH6vXrwvWg56+VM6oHaPTwXOE14vQQAm8Kx6D4kTJ5/o2dCqrm7so
fMZQAE1NJO8Yz2TVz2enFvXo4Ls1W97FdEKvPc7ISixkPZ1qyLxDJ9xnU/+hLlx0
/zE/u1Erbw9tW1lqOp4gw5jmTnD7txV+rAzGm7qQHl1PWMX1yGmJmynR2P8GTbiv
AceauwU2qYRam8Yv/3eqc+vvhWnhylKsnoWApU1PHSpBUW46dxQZ4GXkWiwR0V4E
HJC+p00J023vZY1n42gyfTRAH4+1n+LbB6pntELgt1sLRlzjq9EyAH32RtaP7H9R
SAZmnRLDYt/v1CJcGwvXrW2GmSHZwn0EyVJ1Pze32tOGbKQMFhGWza7m10OHWGUV
oZr0KHBFrjxfwWiCjLT0xSwQ3UMKLY/eTTZnYUbM7wIOD7Oiu0PKEhgv15vgVX+W
BhdzmRKkpVwEfpebxSJPfMjAMWtb3EeWljJte7bZ/UfbqsofxYY5Y3ZyMroh3AVB
Pw9SzrfowG9ZbBtIibL3ihiUlaonaNxOzvBQ3zo2f9Zk92Fuz7RSfq7UmNfLb+x9
18/jYz6mE6v3kj5qaLg9yZGHFi9MWN57TicebRiBouemiiSrdi02uwd20CgCpaLt
WbdYGo6UM7u1IK9ScOfA6s+QtaPB8V8lk2vdc4rcOcXarugTFJJ2oEifAuO9iZPf
6yrP8vbw6kjFavmLS9nkXW41r9VGsBT6lL/Z9Zdi83iRyrbqAlrObXvcZkv1uBS3
Eb7hBxSOj/pwp21wNM4Rn44V4En9D5nFF/3FKZriZq9b1h7L6GABaWswe1sAHdQy
Ewyl5gt1MwSJE3b/jBBGKFfmTRuzspTydw3wxJcDQO58xH1rRuxPW4VMtktuprps
KGdNAKGXW6+lgDGSqWoFzjfJtzTsVe6sDhmlvOAZVeTEOPiFvIRaKKWcpBWvXvJz
RKfN6VhMUf2dMeoWjI8XdBtNvqMwfuKtTru5Jisdz1nwt/gfOfVMtC36B4dzKS6x
dtKRegKuJ4Uc00UnWTMV0wxJRIKLHp0QMpz8uzw3dbWOHc+gVZFVmaGtknD+1T0I
iAYFafnv29qRpax2t64hr//A9xic5czjzVCjhDQQfhZAm/W1Ue+TItQmZ8Rn8t/P
ncNc0sxEZYngrw6NaZVWUvkLjNJ2mD0jfAPN8KpVGqsifX6XvkvNTaPF3OWz1Qwf
oVPHUrjJLejnybyW/v33JWKZ+4SrrZtvS10lQkjCgmJvtzJ1j9iYi2w7axdVPSAm
VYMEcUM044iFLgt/E8hM2YmyLLqyRkEusNWh+Dr+EISZgCwXpCaieL4BBVmlRfPp
Szbx6Ojiym4+HgVU7XSkgoJQAJBTjkLKtIyTvHOMvZ8WXR6oZtoq+iMAln4MNFUt
ynJ5bGI+Yo77LGCS8R+bAkWiTwvsZn6RsSjwKBOOEdxwrp4wqmfB5vfDAt+k6COD
hnHFYSOMkFr4fElJ7G57+m8yjayCI4hCytGuqlfZ1moMxjj58P3oY5dcF2SLAskn
UiCz7PoP3dCzaiwtSI7EsfVhNLlclTXfQgb3v4q5lr4g9dVw9B+M8QenUfm+ukOR
do2Cos0x5PwaFiR/JWi0x/guXg/zecMAV/OgkW1DExRkZapdDdIJ4ORYXdH+Ym4q
tQzXJthddndXWLo047xYZSjD8iERItEyi4y641RPkMgItJfWWkuF2YnPN5DbC3aK
yvRMArhi7Xqv2rNE22MW9pzFNjsRJ8P7eo9I2TA154JHYFsdov8i+neAsdko6wqW
QAWxl/bpZmqyz152i2y3gDq5B/IU4cVh2IUttgB8jZSaPCWXCDWJsux7oka52foU
q5TJsac0K1l7/uoUi5pBRu+d2N1suJIhhHbSgNmbi0nhcBam7uh7JhUQ9pT/okp2
j/XwmnFmhe/597/psair8PNxpYVX7NIUbJZSrJK7oJBGHZtE8BQGFLa7/YrZrzLD
R0MLImskGPClqr92ydukg3BK0sJGEZzntgzlQAHpYaHOxfoA4Rs5xK3LcplNWPGC
kiieVVcangoglNRjeEDlshlxyGBKAw7hBkpSWOD70QJxeyEMuqHE3EwoikK+JgY0
hoISYTCoPbEtbbA8iuTWSYylTFbhgKPzQXmf7iO9dLNlDXs7Qt4DQvbWRwpx0N59
JlgU8MiloZxpOXwCeAtwLUXXJI4bRyC/uslAAFtiYcv/RrCObZmdn1LR44uOnm02
+XqVMadYkJHV8pnIhlbIfteUp8i4mbM99YXjR/AlMd3zLq6IybO5sBQig1vSKlkW
R3ZGyaBf5bFk1+IyudwMn2irKqLyaW3l3O+KOXNM5XtG/1WHrDZPuASlmWacNcAY
Hj1ZUhPA0Y78UMa2aH3qfwQwR6F/rgTuH7aeGDMnnEPKtTDF9c9xLKAUqX9t22kM
3XYx9cYccm31GZpNvh5LZe5WC4d6pnB/Xo/hzSH4ppxRnAZQL0AxJe7Bu7ogFeJX
0e4WeT5TJxIepgb6+QYUtg40QVCma4s/IGi9FaVHQWIrHRHZ9h6xaTweTVgcg9RD
Mm4jZ0MGWrNyvb/gpwqMI5s7D32bMa3rAoQqozmOIjPvp/xohXWR1pVz9gHxkFz0
40hS25+7gu/+vXb0APCLddx+yr/gGQO/Tktu/AYzp1uHh0x+li8BlsizfPK7kK60
Qg+ZROJHksSMHEY5ikt5e6FfWJjoaE6iEI8RKYGdWeUavoo+yS4fT6M/HJfOK3Ki
c+Dl4aWsN+RRgu+Zg25uqLSg2aMLh2Sb7IVetbN5N+KpOPPN+XAwNj/OdDkaki2q
AOyC0y3bBcrrGFLRUOjtIm4t55S+tjtVtYLIReCy3nZ6Awtt1TVDJfdnnJZJ03ye
PNLsumwBFpOwHyp7hufZcm/Qgsp2OCyFmMbN5+JUWc/dEcp8mmHC2oZYW12D8Shs
BgpITDfoiUK64A5/PHZivQOZAaMJ5wBnycSBgV6RBbWN++58WmKb7/HVM2e9ZzQo
3pVfvtgnDoST15rZ7y/Qvgr3DFqeYSOmI8lHnM3OgT+uM2ge4laNm2B8qyBnMJye
nP2piUKutZ6NPgYrG1D/GJmEENSk30iSHYLBRy21rDskUFPe31ENplct2jT/xxyt
LUiKMxSjV8ZiU7OLtFcjToWkEB/P+AR5B719hXtE4bhtduqBR/IRJqsHrVfFdKOq
RYeIbWcL0dENuo3mb3NkjG1Et0bcl1nL9KF3yY+1hQhk+3db0NtqViJ+CMYyQLFI
P+t4vF6qKFly2gu+TBF8U9O7P2hN5qJ9Bx59CzOWXvISmQH8of7ppubv1LIYJql6
9EEa9kwBSM/IbZAi5sugFkWeZU8XWpbCY+K3giRz2ralGHweQLRMKagmFSmTCeas
8PM/eYIEvMuzKGezQ4BTVdzAZus26x1qRr24MOhciXfP5/DcT0xpnVPD6rZjBGAt
sdvZgTwhm93p4jvZ5Q8AskroCiuGMwXXqjsZf0usgHt9CbpsX8HFy/Ylo8so+ESd
8bcdpNbGFgVgAsON/Ljmm8kbwV8jdEDSaWHuiFcpja5/ffrS+vbAWjf1fFd3xmEZ
GXq/ABkRp4+DDnJpzWMQRpOHHJClIkhNxBvND/w4Dbo7gqM/Y3tNTmo1WDettx9z
VKsuAWphWVQ570rldbPX34m0kszkWb851MzXmAI/nqbCoP6luU/JqHo00R4BNVUw
OPvYbsOhTJzIoB6r9sn8MFNm202wWP1PtDIXwuLYZ6tbM9g0QIxOx2OyqNYRXMqw
XeZfqStb4s16+BEOmQh71C/y8mzFsGut4h7aTAGVzkAgVxdCVySJ02c7uhZquz2y
Q8BkFnUX06TzQkXt4zcY2yXcSv4awZzl1Wc7gj1RGJBVB5V+lsX7xC6+w2F/kgJr
x74/CvA5Z0J5vAVBDmowP/BdN8fxU0tQamDfd17H/C8KiqK99ObOZ+7ofTdzy1FR
qdRPNdo4ok/9pACPqvVvm9DQQn9Og+hNcFR0EpTIBhZ3fylRtbWpQu7Jkm65dJvX
43q8t2yDBtjYT8zH3mTeO3cSWoMby4w1i2I+yeBdVy0WLr9fHAhC4zLgZqhGYrb3
xZaOQbXTyaKf+9Wfb8rCcZI5kaoB8mrLR9b45buRzYIqkkLVqHodpJ4ihJUti0Or
4Z2L3s+nNbuZ6I8ouE9FViPpLfcPYd0gr/7GvAvt62XWZ4azvkMKCSdJcnvCg52u
j4K8YLYjPdcnrvHZLOBePuqSs3QxcIF87x+V9NzGJN6SAVBvgJIbt3YvbDlZfhP4
UUIyMTxp6M2E6ZNoUW+VVdg7nLvn3XFsSxynJD4LO/XQ1rgoWRoi3zWARPNEokRW
4A8EDYmkw1gTiZC+w/kpNhDl3rP0i3gIeBAH8cEMytWfr6mqpknZA5YdNMcT4BWO
8T31DgIhROWhANPgjy6/GHmcQt8SEIHRVeDI3vF34GHmjfb7qTv+7/y8SDptR9ix
NeUIAnZW7S8NDRlh0dY+eLRdRvL1f6FS5qGSGlKN5rYBfPWHsCXiE6HVREG3cShc
bfOPS7XPJbgII9x1TTZ5cyJQcWewysCkLNi2Wwjku1+7b6SdWxrA8K+WdCp7Ah3V
N81Esu3VPCK5mDiKFyYbLxX7V/LFb2EQCpLuKSFz+9IPKMY5tTf2v++kVUbIsip7
PVQAc4ULlMNWtRf99RW/ow1AfAvQz2XjuBAqHZPpr/F/V5qjP5rXhNkjw1GyPiwH
2mNjKaUEfP5ERpbf2i5Xs4YhZsgitx5lelTlhX+X6Uqb2ZR8BGYKWioeF8ZPcz6u
WkbA7LRU3u4+ezLFAp4+/+M9cr6gU2o94S41ntkzT1X0EwpJEmGNkFuW8PV5g1+7
yit8sdzqLPhE9LDZkDW+4nfHDmwNm8EZ1ucdcyyZg3Fg1VRY2KcM6HKe5MZ7fLr0
WhlDzVPAK4+N9zz2TCvLWuRCFVwmnsyz1AsFqr5/jxG8Mp+92DlqCjco6/eKi+8A
svyr7kxY4oHH+32tsRKKbEsPf/EJcKz69cZGhNoUEt7J3Qzxp9I4ln6cqVzm4fGK
DAJPaH5s9s5p1iSiG2ECJh/hpcK+NagOhngs5Iu7fTiiHZxVO+dDr31JwKOQVJBN
kmmHY9FTEAMWc6GdeSNfUFW736LHV/YR1VfXJxB214Ovuda5kPsTikKgPpEq+QAK
z+6NVM0SF7weJjiYwaRZ1J6+xHG7MLnl7ZP8ZKW8uFimKvf3FfJ43AJt8zvKJCHb
bq2p/DMQ6809NkSucX5jRGsSuOXML36FZlLx0FprEopGo102077daOqQJLvTZV2/
701jfjOala4mZw9Y3Lnpop5tWfVa2FgeFU4/XSJ+5RpF6yLeayk+kA2xP/eZtVWk
iNZO6wP5PD3g93205P+lmUdkwDQlkZTwbth1C+/AFwRWOvPQnzfSKxkPgKaVBcQv
N8ubykxDp0CY2ccrL5TCqlNhJiznm0ue5N8A8F2xJKyse+Jdo2+IQNcVuIItm6+a
VCiQFX33XA95UmVUYPbNp4lU2ziQPrTdDXQa4ovKmoZ8/IKHWsyDwEdrAXiknj3T
jOtGZ/xBtZJeRNnURturH36gksixvbBRQEwlbKXTzecQiolmnT3ofVFfmopAjZHb
B83Dfe+dvsTx72hINeHDAB2kY7piLi8UyE3ZGMcOe70ShoyPUxIg9kXXTV3qOufq
pv1K3N5pAh/pdneUCxUK9liYRYTJO0oYySnr1kPTmfxYV6u1C60XWw1bO7E3DEka
+kI3AuR35aEKLmUSqMWGF3EEDl0XmxzzCvLzGpC8mWKByrhadZ2PMft0bsAn46Pr
1CucVtfOMFcqmy/JFsbT4lFBA/fn4MV3ytS/XcmghEv79CUncCEnTf/YGTBKl554
STkbApkIvUekVr7WQR4VVvgd6TfDxYcwKmVJnyQMi7PRTJZ9yW8Cl91aSS5N5FVm
nWTdjsOsOsJDp30lkQsANXqWwqYPGfybVa2hGh81XhToRrs6vGRPx5ghW6ILOJ1c
FS7+PKmKahL6bqqrCvfyLRanlMdz+zvaSdWOdPuegMgSRnjFQwm47CIUJJzxNkge
oi+Rhunegwg0t2+0vW4siIYVBjrPfBPYQ3EBpvD1HrIbP1bON2bQ7nmhbI9200B4
mc/b0tRBxswsCr/20PqYBtjVlqSxGtejIKi+1Bxc3gf43zlWGESs+UlWge5MdwrW
6vokWdkaC+JKaeVRgvo/EaEEdhNswpKkApn/Dj5ELKgVfxU1ue4sGr/ubm+WgxZf
2ESFQZsqoDnDr6XmDoyJsFc7TctrZHUh/B7rvixf3vMI5t2V8u9cIz+hHuqkazbp
9tInOPjTie7FyR+6hRf8J/tOZx8eTBWnzkLM4l5HMITSPEiXje3r/WRiWmTrtXrN
sSqeHUkHBK7gha9tZcjykqxFrFmunI13E0MlfsHXV5KDC7YaTSPAjLttOBVxW8Lw
aMulRmPRGeSki8APRm4HqcPWxjXYupzJMaOpxTaQmCgf2hbZyeqXZFDkEyimx5xJ
0UWj21wlDIq6H0jy9E66UZqVfl8ycGslpsbKPcj0pLpUlwqLRvBXnKvq796JgElJ
g73XwRH1VFj8P7JU3BRuOWBiWGYAQM+D2bB/ZsbQTPNHMFi9qBFvgXQ6llDwYkyl
5dg6+J2pfCZ03YTZKsNgZIYbk06xG4Nf9j1XhAz80mOBGkm+QDqORG1b7h1cYveR
iM9tlfTSbC9OuQtA47L6AQ8Xtp8lXMKJmXa8TSJErdZU//2TGdsMlkiSlI56f/rz
03D8EGw38ksZPO3bZOL7TulXivRqf/eJtrIlcjr4l75YpIOoAgjsXt5267bYUqVF
DsBZ+MNWs84xKW5K151dMj6mQI4WfEndUh+Lo2vEjy+cRTBahVScX8WvhbCLkN2y
4Sd3lLwcwMh0F10urMzgmFnfK9xyemO5ChjZjVry/Z2nY+tdJI5kRnY38RWrYIyV
wNOQRa7QwCtHDG1S/gcimIIRYmpG6Q0T2SFlYXKYKO17bQKNtj/jyoVjqocnK14B
fHedqdyY/DvpA3gY8Xs9fj1b6ZtLbLnwIKCFaDN7eYBfHT7SeFmEayKchze9JGbM
qL1OAaE5Hw1H/YFXVMqlt2yfKulABXe/iHunGGip4afcc2RkHxT/Scdyr+huVqkg
kZo1bdJQBLH8VhH++3grP5mUuNifkFpOvzyq0vq7CCp36pRQQ85daZ8wEPo6j8pP
wt2eluNLOpnUD/Q7HSC3Wovn857kxJcdRKgwnQvmL/Y3ilOrtgXVGVS0QN/KntkS
qQwGqL56nveZ/d72eYoWFhvQjUkWgLAjuTjxQoHgzga/NZ0JCqbalJ3QTW3f/mLK
8Bbg6vaB8ZEmCe7rpdIbMl++6cGsxelsGRUSe/t95DfaWCBNx3H+JaqMrvohWyIn
Laktj0dnUAbQlGBDqHtaY9M2YCaavytdEIATvlh1gElDHrK4Ovx+OTLloEgZMqOo
qRcUvyGki3KlJv4BBjrp6izw5SJkGgFXz8SSnjWxlOY+ciZ4a245yQl8Apb/n1rU
VWzymTDLGAphgpo/WxxA8ErGMav9RWLVb/R3XyasGCquDPKj/mzl3MvydDar/ySV
1foBxf5t8htZb2H6Rvo7IpdFTqA7+Og3C26luJL12IZMZLrKPCr2hO0TszM5x93S
adFsW/wUQ6WjCPBndBTUenHSO26fXj4YnLlONA4HkzAZ70bbO6EZvMDtaTK2v7Sd
+H2Cl5WB4A5uvFE6M4MskGTZvNwV41PggfW8P0T8n01OpOUONfTywyKGMf3eBFGY
nL8wyw4BIKlzA/fSSHL6R+qV6cPSjabMbqtUt0RO6lSy9tkM/BeR8lk2ga+nkf2Y
exSO5rVktXWKuSmY6J1xoESjhtLMgFt84GN7YfyliA4nhY5eHzqmL5GSHJsWspND
1Ed+FFj72kVGcSn6tuoixLYt6WBSQmWSO3Hqi8i+mnxmHVVyhXapHSxhXsIb4Q9X
a8PPK+8ascrGmXu8CT55Nb9S4cVOr6n0yJvRi7RRpyHyRHEk+9leSoAiROXCDhDl
OwjKPGbCaz0joHLWUipRfkK5Beo4Q7dgH4vi1oDZiof3nqCGC+t+62ENWnncCX9N
wZVp4qwSTzVx6g9CatJzqaXRs+Lw/T6PP0yGucXp7fZH+8Y2nicQX8zysGOXaMF8
m2e4hdCEqpLBhS3U/QBhx9nm65ZtBM5qonjKHWUDGR/rSEc+rn6M4VdkMjdq8sl1
/iFJjrePeSH4xC4miIjRF2LCzEUn1XN1L0mAiwKT+fl9Tvi6+oAR4ERkQfUQwdA5
FPaUyJp2tlknYW1VUj5dbUwHixstWFJEDDjWikly7iP5rOC+gAso/v4HUx4B9n5i
y4WKZRMvimZynphTZ4/j3hhTas75biyHXctB+ZAhgevRfl34sfVCugJtvbdLIrmP
H9iAj88rGTq5BvmRBGg1nqMZu30KbM/llAvbOVE0ho68ewj5J9kOKZkEOtPvyqm0
nuB5ZXHO04dKDn0HVHv9c4C7IEzQ9WuklsFc6DLLMkj/tZc5n1UkB5zX9Qpe/Sik
wBsDOPTgDKinZ6fEEvRiMDS6VirrPxMPreH3M6e4B04Csm4ZTVnikL8UvgvnUnTb
7jvwpzrkXTATcFvMNKjKhb6zFHde2wfdNBbHPN40LvvcfmI9S+vbmMWUXr2UJ3bi
LYkjPmanlo6QRURCy5HMchi6T9i2zfigt6NmOEMKoOoHWp9YHF54LQnJ69WI95rH
jx/o+/xqhf5kgiwwCl0uXDHPZSbeJbPnEs55DMTWVa2NeAXc+yrKpqscqXjEsn1B
7dAQ8nT3gPUCQTkHlD+5VcBdbB1oW9TXtgwZ3ptMf6YizPQ+NsFuy7thLIJcAzwm
PNMgyMIneVSasD4riJIy7PM6h6yKmnoZFpxQ6CXLMYcHnTpR9MkhqvvGjmukSOXw
dBwrjcKpjdd+3H7XoDbqJ3+PYdfpRajHW4vJcejiMDnnUnwuCMegRjo4RYgSyHdr
Op+nUb6k5u9KU+tHqrL8+o8jXTTj52Aq4mxQ2wsS0tc=
`protect end_protected
