��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����S�M�hkF��1~� Ά�``0Hɿ��b��i�<�1�SzFĐ�48��ch�iIQ���H����:4(c��_V����&��}�w9B
��T#�_qx35t���D��<��R*�E����nK�N���������19N3a7K�0~��!�@ըfG#�=V�[��&@0Xy8�U�N�
�y��I�S���j�kU�,���87��u�:]q�Ƒgh��8�i;�f��ܐWq�Re�R^Y�˒�
�1h��{�%z��1(Q�,1:k��S�pv�p�$�듮Z�����C;�y�A֚��Au��*��1�-�_��e�(� $��d8T4���z"�������0����W���j�Eզ�$f\��W�t�(;�g���u��A�j(���g.��=�kz�7݅cִ10m�OɅ��1YW��F�O�`�,�w#{�iR�{���X%>�w�?U4�re�C�E��C&�i��r0��vf�8�ԫ�ft�cY!h�����Ϸ����q�ׇ��/j�"(@��c������mI�kru��)��2��*��0�r4�������i:3a����-�������g=���\6A9l�6ιB������:p��Y�Y�[*i�29��w_�\�&�h+!�)�v<�}�!&��V� !/��y17�&�ţ�*�Ҕ} �2]�H�,�nV���˻u%x��[�n^j^���XԞ:��
v�9Q�����3.O?����Խ��@��5�RlCN=ۛR�J�%���oP�PDq�w�V�e���?|3ʆ�ꊆ��#%�P���ץ�sJ%C����o;�`Ԗi��CM�+�j�ت3I@��fUh3F���v�J@<l�CpK�Am�'ο���q}%4w��gc��O�M-�hоC3�T���32���e��j���5Z���WJ��)R�o��[����͐��P;f>B:�f�uP����n7�q�" �#���A���p3|�KZQ��$�xA�[Ќ�Gґ��:��	�Q���*�����f��F����g�,��u�������Ae�\�ܾɍC��Ǳ�rK\��YM�˺���/��9p�e�-"�>|�%M}ɬ,r/�����ę�H�=�ؗU�elj��	�*���>�zɅ��t뗨��o��p��˳�;����MW4q���i����yG��L��D��!D�x��Οܦcߋ@�O0���%�qYq{�2�ʙƛr	�ȺN�*ĥ6eO0͑����<��D[臮�|�w����v�7bq�Y0�1]/�G�#vsH'b�a�8	����V}0���5���h���k�W1v���%����I����1�~'���}��<��4|�JƋ��7��b��vN��( ��ύ���2g�XR4��S����'���lN�����`S	<���ږyjR�(P�-ˍ'���Ԛ:3Q0�O� =�A|5����a��Ŝ}�I5_���<VW9:̇�0�.%a\Ȁ5���q�[$�����!Gv��sT�����6Ҭ�i'n\j7Q�֓GX��.��l�.gջ�����M1�\��e�>	A/U���L��̵m,�q"GIKt�a�{��:@�
��|�IBE{;p���K ���"1��8�Qw3X�Sgmִ�2��z둚W�p�wVێ=?�;챞W_�fmI��a	��̀Ֆo(LR�+�=��`�����A�)$c�ś`���ǯ!K�Wл��#)[�q=Ú8������¤�y�i��Z:���$��*����`	�,��]�Ǜ~D#l�MQ��O
�@0,B����yT�0b�3dn�Vʘv��5uM���U�yS�q���a�԰-&a�1��mtAZ�x��w�G��/� 5L_U�Hg�����n�.�a0j�S�d��������Kw�(ń+����o/V/��b
������ ~-��� �?�Bˑ��L�x��_��g�jE��ezI��3�u�R�|��fs��y�MLD���m"����z�i���gsr�y��V9)�8�1�0��a+�{�K&�H/-fشɶ}��K��(|4-Z9"6�a�I4g��_��9q��!j����eg�o�F�Z�NM�Hy����>b��?�b��h�)�9"C��uo\�"�oP�s�ۼ(W��9���E�β����Oh_B��69:y� !� ���%�pN�C�7���Sg�� �@�Uv�o�b�
�4�ѯ��9�R"��_B��� ~��O�VV�+.�"�N�
pdX�uِ�(!D[ک�.�1r��Rdsݔ2�V�Ζ�'��U�4�-_�#'5�w�\�g^�.�畵Xm���U ��RV�r��\21�4�|��ň��)Xu��$q�)��{�ڮ��,y�2��`�@j�׬Čo�^��S|�ig�i�ؚ<�,/�7c��7طX9��v�= ���wg���;.��܈Y����z7��TTy-]������ۖ.�s���ҨfFS[L�xnݲO p�m�#UL{.�,�#E-�>)��;�7�=#2�(�_�&\z��/[\�Z��@��^�B�,^�����:ݎ��z t������� ��ʠ�z3���87yny"�
��B_����E��v����iG��lA�W�����\hM��rSC	1H\p��(~��۷X�.�Ś�ݦ#(�x����ȫ.��ba��W��m��2<�e�Q�_6���
��_�/�E��<��?r���R��W�TIJgu����r�]�D���%��D�i�35/rdeᑱ��hQw0���8��R��u�u�e4U���;&G���U��ڟ��z�*�u�����]�T°�� ��\�����\\ST˫��@2�������Qi6?�JÓ��vcӡF�汎@�e���$��U����9S�} �)�׌c-�P�Y�PL�?��F7 6�V�� �Ŗ�I�å_u>=��ٓN[�	��vBSڂ��J)<Q��^�_轢)}!���"�y��Ķ����ץU�f�f��
��ِ��<���ʠ.��-�Y%ς�����ӝ�+�!���L�b.�h,�"�C$�~=�x�C��S�0�{���l+�G06\�"2`����r�G����ZMPV���]�}G��'���� �͊�kWc����A�b'��h��'#8���?u�#��.��Ge=�|_OP�KAs��>�Ko@q*��Vf��Zʙ�a�r&�ì��o*Q3���<����?���u�|ե�FȞ�z�%����-�c�VznS|*2&
������?�>�
������������V@�s.��\ Fe�χ��G�ϙ?#~���h��)�w�;��\����~����n��u��mAF���W��
���O�	�1�\�~˫��>���OC�d.�9�+>����.`��*Y�]+������Fu`�)F��9�2�ʹ�('�W�ψd+�2�p*��<�3I�N+1M��~�v�So�L8�dK�������]�r��|��9-�"T'����;��+�*:�����qY�����pq��ԙ�F�=��^�)��Z/I�f!ně�Z{Sq���Cju�V񉫬}A7�u�6K�`�P��.bGGr��Y��>ʿ5��\�Q�go�����N˟,.*"!�_FƳn�Ϧh��Lt#�gQ4�"D����u�HqPhSf�����X�\埌�8�9
�"���dJ��w~t?2Ouw5x��݈fA�e��q��뮹��wϬ�KB�8 "}��z��xg=W6,~�N�R'��#�տ�����@%�#Bc����^���S�S���R�M��*_@h�k����O&w�
����^r7����qV%!�~2���������~O�q7F��B�@ۋ־�q��O��pG�D_�y��ٓ��#���(�=EQ�>߀m�t�Ѧ^G���&/`�)D���uň��q��$<�Gdj�E]2
�-˓t𷝌<��j����aG���X'l(�FV��@:���f-Y�GY ?�	�X�_L�6@��?9�Ј�몕��F�8[�ݣ�oN

��W��7�-ט��aj����<�=Py�WD7�Ua�*^�]�L+��=����#�%�kS+`wW��J>��z@�	U�tER˽�e��t�c-�5k�aC9��%���h�{FR���4��f,nr�г�A��x�n�g	���[�2�}:)%��j���A�F�1���5��zf�A��``T.�鏯6G�0�����)&!<�ޞ�I�<lQTeC�1$Q@����{贰t7����C�8wI��M�k�+��ᜋ>�qƍ��:�>гD	|�dHmjPREC�l{�������t`3D'�C����+Tp ?�}���{S<�f��&Ϥ���p46�l;7l{k���ע8�D�Y��j�7W��qu5�	�Y�lt]5<�]!y���/8G�,��ho�b�{�:��y�W%�	�PS�4W����X�����R8 ,>�$�X��$���E��{��j������G#/�����8�R�ێ"1O5�#�]{4	�AdM%&�S�G%�2_v²�<�?rB�QI�|�2�K�un���H��b�H�������X@��S�4�@��\���g�%�� �?��?�sjW�ot@�wS��	�v�8������֨�~y}�&+�)�l��@V6�f��6w3GT>$�T^�ao���I���0޺���T�cA6�hR�B<8qi���掄�y�"�&���rh�>�ȟW���.R0Q�|�N����j�a���y.��}����oz�ط��oI(̔,Ks��`6X���x�a��g��<I=َ�$qe��&uI�2�o�ƙ��Ŋ��{�Q������F��:ȏigaZ��H#��JW^̬�5���H�ͺ��O�"��S��+�x-��c[øi_d������BT:[��G|3{��#�>_�s��������D��-�V�ۡ:i�N��=���`�l�)�$O�gɔ�R��L���8s��ǆ!��Z��U]��ӊ���������nn���u�Idz��h��{�@{\(���������9.�7�
�Ku��^-�i�IG}4�($�[��p�Q���XD�����tuw������3wB� �\�HI?�ܷ����6��dLO���t8���!�1/�������+�*X;Z�C0[�u�V��r�r��yWS$Q*9&��Dh��o7/W��_C���m�� �aE5�"�^�ȣp4�@�����X�h���ڍ��1�]����r�lH�h�(�\Y����J���Gqlue��gL@m�99�TzǙs�z��e��������'� g���<3�hd��aĭq�0GuG�Z�)�t�L��~^X.ֶ<0�*�Ԋn���렗ћ�Tf����,4��Ȥ��Xc�'Xb�:v�K�I c42B��9��!�K]�O.t�5�Ď���W��*�h&&�F�cNm,0�a��i"��� B��+�_-���b�͐��b�ƍ�=(Op�|�����]�Q侀nd�#�}Gc�:w��g����A�&�,ѽ7|�#�����99
0�d�������������K�u�p�b)|.����qE�"��I�sS���{���j	-l�G�اP`@���^�����2`��&����]ڷ{R��}~�G�nj�����e9{@�%�*3�l`q�J�qB�q٘�ݝ�;���N��|(g!�wW@�W� ���`.�+�@�.���!Q0��0i�y^����UA��9x��~�6�d���c�lC��r/\6��Ls8�zG	�-g~��p>3F��j�
��^�ق72�|&;��EW�Bl��X�t�H9�כ)��Z�P�v�j�������/�zUkQkX�����T\mMK��j�LZp��g�.�wr���B`S�6����fў!|�c�a2�X���zȓ|�yQ!��?k~�����}�.�L�ý����a?r��c��z�b����[�h��\��A���ߊ������B��4>k��K������y�pf�E<�����W�Q	�qL�d.�0�=v>�qv]���D͙U���V�Nn~�5x���A`)_�gS
���0�X�GIT%r^���O�"�؜��+�����rG�ޒ9ܱ;�]vV{�;�W���X������K����{�H.*�	l����;7t�d5F �[ "�EV��k�e��N���+���'M��s{?�A2K�,�,ll�=�7�%��UA�֔�P�ŭ���ƈ*XԓƷ,��͚LHr�"%�gl"c��&l���;����`w�Iu�s�Sβ섃�c�演B.���w�3BÑ�љ���⦿��꘬'2Mu�C�1�FI���^��NX�\ˍ�g�FE�̢]�ϼ>i����{&ŒǊ5��S�������k��`�vVٜ3I¦|�]1:n���䚨�@��n�[l���*��>�N4W��zh5yCl�c�����dsD�BN��SI����p�>9����=��71n'��W%�]�v�M��RU��`) �{���+; �'��x�f\��!�����¿��yP!���w�r���]p, �w���:�@�5�'R�8�8���y�Q��4^�өV�R&�8M��CeI����d���P6d��vٳ�X*ˢ��M����p��-���v�|�#5����4��h��/ ޢ�KPy�����}�ߪ��I�'{y�u�ޅ�J`hF���H��{]�����z)'	��9'b�cH'4�Q�'���5b/��ڬ����&$5�g���/
��
�m�өB8�.}L�h�u�T��ǈ�Qf�5�m^+��ݢ�0�[Q5Z�e�#+�z�C�k�x��n�.�Z�9�Զ7A}�m�'k9p�Pث^y"ȳ�Wy�fEJW�/)5Ng��ᜎB�w��O�e~@�2q6(�'�,�C�+އ�ѳHAq��R�>M��y�Ɨ�����2�������-nc�6�RŻnF̦r��}&��-S�������_*vI�����q9��JrOa��g0�-���&��w�]
��+鹂��k�s@��s����8;�qz�m�qZ�o��K(x���~�\��5�\'1�%[\Qg:�2��B�r�uʄ�P�.1&���vΏ����fP���,�E\���$o[J�q�)�v��A���+�E,U�T�.�w��S��C�
���,�B5h�/����MX��P�����an3��rg<t�v?v�wrQ΢�nP�6��.���CX�8g
ښ�F��������#��Q�LPz��:�)ٹ*�L�ZW��5��8�蜇q�
;$��� ��~d����H���1SC�Ɔ��k�����J���$
���L}�T��<���EK8pE�hia�h]o<����ǈ�P���,aJ�.�,�����̴���Z(��x�H�Y�D�XAʇ
���;���>�����n�J�9[��.X�q�����;�YC*��7���T��E|��3��q��dO�a���G�Ξ��M��K��k��i"- *m#�=� HWj�qdn�uL��}2�-�zKscw��ߺ��b�Zu9��3fL�e���η��%�N��o��i?7=&�%��j�<�0��W`B�;���_��/Ad��
�[��w�4H��su��q铒5Na�^���5�`s���%����@O��Hw*�PI��Ίv��t��45A��'wn��k���}Y^?�F��Ơ.6��(�r�ѡޯ�>��b	�G���'������l�>U�Z��*bȱ_Wp�2�~
�^��y�7���SG�J� �kPt1��*�
��M?�(݄��v��7�v�̔f=���V�����9 ^���	oM��L�C��t���b�����ϛ���&^-�\���X
���}�c���a!f�!�'�̵Y�)�ؙNtx�~+"ր���V����xEώ\�\S驏�J����[����.s~���&��������t�5�+o4���Ւt?AzgJ�dX���bYv�G��SLU�W �c���^�5ө&�Dh��ہ�Hx��Z��G���1��I0���^j�e��u��ņ(5Y�0't�$v�'��ͯXC_�����, \�n���
�����nϝN*����^~����RꅒM wŰ��������@�Qv�^?�޸#I���L]fsj�b�t�׌�o3T\j ���d��uܩ���{P�i
�@k��Dj�Ɩ�������|5�3��ޭP|�7X�b�h�̷����kV	1���Lg����Q��;��^~�;t	�xghc��G�6@�d'�H��t\�|ֹdw�$�+�2�n�zߠ��כ�~pH9�G�`�*'�y���F]p9�c6���4[&�R�XH��'��^�6�+ڶry��G��M伧��4&�������R�+7��Iq��t1�O�w��Y�	T~cᱦ#.��+�hO�De�Ο�>�0��,4�m��ǰ}*ֲ�@`�{����T2"�������B�� ��nS{O�NV�%�9Ԥ1�FV��$�O�-�>�|�f���4B�ֱ݆5����ּ$��YL�� (3=Od��Mv�'/��Tݲ�o��=�+v��ŕ�;�f[a�A��0������ٳ��j'(�ݿKp{y9��.hǶ��ؓC�=����.x׫���+kgu����m1H��fr-O�]�����4y<�&&I�t�����G4�"$x�l�M$���æw�=��$�e�T�����:Sf�(Z�D���_�j�*ѫ��ː���J�LI
�(1��W^�hъ0���N��{-�P��$������ �������2�F�� �C�6Ƿ���@��k�	����)�fz{>)Ȑ�)�M�_A���ntog���������^���c�"�E?�����C�܂�.n5ɋ,����-_�/8�m#{�Ն���jÿ�����ߡ^�@�ł�I<�Q��ph�pU	��)>�A����4fk�]�����y��h�& MȀ��@�ۀA��D)2S���D�R
,8|����Ć����Y�������LhL��
�S�q m^�*1Ґ~���i��n�W�� ���V��*ί��O�ף������b��B�i����ڷbiV��7U�L���U�����$s�Un�/�G<�Z@����$:��Ax�1l�ta)�?�S��U�5��X�v�UH�E���(�)���p���鮝�6�x�̒��G��]ja���۟߸	jXc�VIJ�+�~�E�O����"e�D�"b��*@O!{��dDє�v�2shh/��1
uFY��n��G �~��^D_IU�;Ím�0��z=)�9܇�˪N�~1�8��%{�����͞�k��><������s5s7�r \����a���X���8'e�U�>�R	.P�i$�O��_|LTp���/E��0>���M�^��-�kI��?�]�d��¬[�na��Z-'� �T���Ym>q��Ibҁ��#_���&1�ݒ��ܚ�tv���S=^s�T����)���[��(sV�'���b1��tD&�-}V����w&��$'�jhzv����%K$�%�
�Ҹ�`7�:YĺA�@u�=���!O!�F��4��m�P`���FX��@��a���9?+����#S�4f=;���� ���F�GC��[�̅l�N�� ��&k��	I�̋�޺᱓�ۗ޿���y<��59���x��|_D<	�z�YQH6���N[IҘu����n]��{V��j���f��-�b����i���{G���5�?j0����SoN�<���h���Wd	l`��c��a� S4���G�@��c��Ѕu�}�-m���9Ƨ�cb�������Wt �$���"���9�^�X'�������Y�u��_��0�@!�t;>�!��� �"�/SȺo�m��IƗ|���,�3gD��F��;��wg�!x�(N_j8���˃HL���9�;����d�l�sIQ���5y�8�HlB�Z������� ���f{�����T̷pӇ�L�N����� >�5=u/�`����}6F!]��O�}��J		jς����s�E�0h�^��G�7b�Z��-�WԘʫ*z[,���������)�"�0Z�}lj>jv�v:׍��{�����"A?�t1�e$M|BQ��gC^ a��T$ޅ�s^�2:t���� }�,f�@��HK��)�>V���Ѝp�Tb����"cJ+�:-)*?����fT��*n�o6�9�?��{0� Cޅb�q�e]p�Z�i��-�� �003�{h�7� s@B�6'�=k{�=ԼYl+O�G���4�3���xQ ��6�Q�r�}R�mΚ�@��x��.K}5\�z�ɠcqm�Q�.�Я���K��!�j TqQK_$��B�_D�:U�.[��d�Wj//�i�r5�j�����dC��������юg�+.��X��ܰ6S��)���H�=�Z�K<�m���heL�İ�j~���C=ĕQ&_L���9W�Ɣ�`��ϴ��<ˬD�	r�1Qx�Vy5��������l%x��p��N켠}y��s�<������I<�.ϢH���Ǥ`�#���ˁ� `�@2e$�ʽ�h�JѦ��%)��tU�c�
]3�q�1�#e��&��]��nPcR�^�f�v ��4�h4^\��9:��n����G/9*`$,8�	�߿7q�u����������ф��QJoM��E=N�f��r���%1�{/<���}�2�Ug�&�Ǫaܥ��Eꁛ C�ځ������I��$�A}1괦"���b����v��x�lF�`��O�N�|�գ\�#���#�1������?��c%hF�=gC\o 6A�D��4pR�aٰx�$�==���Ūms�M_�'U���+E9��8q=×��ɠ�q�ߣ��ﾓg�sg�����`�5=�8ݹW�<DX&����p�v!O;�'�Vs�B�s[}��M��8�J�-�V�qT�<��	��Y2|!�Z����d�%K
|b��8	���·vA�6�:5��@�5�դr.��yE�]���dN���u6��n.k١:�:�������%�?N�}�zA�����ژ��S�+��ډ�?���\j��!�6�a���CA,ԏb��y��򔔢`5��l�zi�JS�o&�sB^�tT�<(��T���!<��P^��}�qkj'�C����=o�������+��	��[$������y����\�/���h�� �5 I:K�)�B�u���9�~�9 ?&\�2�,���q��ZS��)�i�OO�"�[�x�osn��������/�,؂ٷ �Z\��� W"~���n�,��L�~O5^�^WHh�f���(S�e��V�å8,���H�S�h�9����Nv���?yA m�KX�k�k.a����ߥFX�R��̻��JN.ۭ�)�����2��kQL"���}��ϔ�+tE��Z*����|�!��d��,d��C�q��I��C|�+��u�d���O/�~c_'�oe������J�*n1�[8kf�$ew�;����I/����L}��Y@n��O���q):bk�?� m�.�C]Q�=@��eL��Ƈ䆶>�E�W�Vn������
P�*ꢄf�U/�jV�2�/���>7)��Z:ict�(�b̅�UCaQ_�e�_��a� �qE��*�\䭭�̤�_��v�[���f������.�x����2t�W���j�P`h���=JM0��1��нŨ�Z/���l
Luj��-"=�P6��
r�!8�h�h"FW��^�8�*�Z�Q3����(����Mm����$�b��w�d�}^m*���S�8��R��>��~���}�
��B|�=r3���U����(-Z5���lшJ{��"q�mNص��7E��(44�� �jp����[5�����_��o��Jv�M4B�4gr����� �0�V�v���:3�eje�pG���rZ��s�/�t!ʩ�������r@�Q~��53߬_5�\�)W�՘���Y��ITG�v\�D>���yl�[3NL�V��1��/.��M��^��[�b1���J���{M��)������x�b5���>�\����=�f��I&=��.��4L�f1�1�FfهjD��d�U��*��Eՠ��gmʥ�_���q�#"!(j��i�Uw�'�ӝAou�_���*j(	��Tc�{#'�Zw�N@�d�.��V�, �W:������/�K�!�Ǐ{F,[�R�l�9{V�N���s�V5��<���q��.kb.�p�Р�����}����)U�2�.E�a�#m�E[����>ؔ�/�WPX�=�]+�jO��i*��@c�М�P�~�g՗z�.ؙZ�n�Xnо�g����H������5tz�V�h���+�F�e<�պ�Vj|j�-���/�����+�������f�):�u��3 J� �)�R���j������Hm.��;�<xj(�Bm@�W�ˣ6�u����z͎�i�1������Y�u�m]p4jy�,��c�:��T�(\��_����j
�jķ�-p���T��� ���0ϢD�3���%��L�����m$��dN�����E��^�=
��NM�Q���C�.C�AC�ƀb�����K2��%3����?G:��R�XTH*�H6��Jk�>kŒys��Cg��%�%���n���xr�ps�ߣ���m?�d�s?���osĖ9-���H���Q����X�(쌙�x#�d���0��r�������:ݢ��F�����+�US�%E��N|�YjDX'`�2�+t�md������@~��d0��1 �|�C[^U�ɦΉ��
|#�F.&W�4���N.:h�d'4N۟�j���{�(�c������d���çg�bOvV�{ct��?���H��F:�߷E�	:�>��]��3�Gg�׌h�t��J�+�>k�qi��>��@���)W��|���iê &���V�}v���<*Q���V�*�gլ6
�K�H��m1��bk����2$�%lA"��'��7O�����g*lsi�k�c�т��Rk���F1~��Lv�j^���B�L�Jw�)���U���Ϩܬ�m��q"4�k�7�^������CN?;o��d�.O�һ���d@�� ���AG�~�z� _�5��~���i-_�ܕtMG��m�D���<(7�c�B���S���������1���%�!_�Ig��8��A(���ݪl"ɰ�$`#]>t	`��ļ�NI��uM����iRb���ȱ�k@��Tϕ�u�ng��r2z���ycÖ7���b�^�I���p���zq�>�&�T�v�82���ԏ#���~�Q5mȆ���mh�h��a�iftQ�����?�t��R$n���Rt�?��d�`�5�m6��|���R�s4��M��ϫ�4Y�����K�����x$G���G�T�sm�p�1��zo?�~�8�{]�݁��j�vP�D'|3|��鵖c6�Y`��.K�2	�{��p�aA�x����ДEjVF�G����]�B�}��Ӿ���,��jM�T����#�)ϲN��T:�&�}M���mYL����)����؛a��D�'�3�)�_�h���%���L�4l�u�(zN����y1��I�UC-�������@c�i���K9���B���:N	���ٕN���=�[�9�^_懟{�Xz�P�����*��C�R�ULd���Z���Y�� %���>!��i4�?�-񂎘6T�Z����~`��R����-cTJ�d�?��E�Ƈ��4�wSK��K��{b��^e�)���	�T�`ے@�%��8�J�nT5��9���Y���yc=��6�y��R���mRA�����ϕ��]B����e�ѿ`�_y�R9E���F#�>MT�=$,9�2��Nhi�}�B'S2�"�-�{���S��~�V�Km(~t{b��	��;J΅�8�5��}^h�V�A��g3>/k�>E�@�A�Z���Ԭ@�.s1E���=%REn������>�F��8��G뮑kJ#��z[���s��=�̙5Q� �� #;�A5��Ն�A�1.�����J�X3%�ʘ㋮y�W����\[G��]�	�TX0��c<��h��]>�5>@�4�������+���V����*�W<]S��<�6���GS����6?��b�g���ʡ�Rz��)����Vgml�t���������zp�D��3��XJR�����6T&(�+����s�0?yNmȊ>t�Cjb��B�1�.n�4"���}2H#�<���R���@��;��i�a�v��6� P'���孆�W8��Z����b%�4����I����;�{����!�.q����O#��`��)����b 4Iq�e["j�������n4�$Uo�Q@%V]!��r�񙋷FM��N�x�&Gy�#�d��5�o����p���5!C;�(�\�f͚�Ԋ5w%��Y�-�|�ļ	ٓ��Y��E9b�U�Pi��:�!YmL{�iR��fx��w�.�.�#�c�6�&����Ȧy�ȱ�������N;uZH�hE��S��]��f,�b˦yE��,V���dZU�'(�yVM���v�F76���|��:�m F��� ���|��o:�G��:�ڊ�s�6�a��(Sz�X�oI�	 �[�I�B��Z�hB;>�N���
z?�ȟ�	�LѪ�T(o曻���T+$LQ�[��C��h6�kՇo���e9[�v�Hs�"t)k�>���$�����u�9�N<��on'�ƹ�T�;ܹ^�Y��_�D
.�EF.�,�Ԓ�+��Z�Vk��'��F�;��ؼ�`e4򜼡�c;L��t�g4�^���Xؚ�gQwi?%-C
k>
���qa.Î��)8��봇�l92c��H'�p��1���|�Z{�D��{iX�_>*�O��OG�����Ruf;��.���cb��h�f��_`��]^n�Szd�L��(;����L����jH��ri�Pd`���Zfa���Y��fi�L��n�a���]���.��o_������`^n��5�/�O�'�4���=�Ur��1��������fj�uDE���n撙S#װ��s��QkȜ�ĒAe�x��Ox�S�HCA~ų\_�J)��]��%ŀ=���L����6x�C���������2��L�cWMn��0~ԯ�z�1�?�O�EM��e�:|Si�'0fIZ�J�l�4�����Ľ�ZҢ�F�&��`��KP�l�Һ��_��(���Cm,�����7��V!��jXoY�[�0�a���{5�#�Osx}�� ��p`����μ�[Y2qU}���� ��M^�^�m_tcgĴ�5	)Vp�s�a",�[�� �1/?mj)4k�Y;�F�|����e�$�Z��G�@�#����s�q9ڮ�|j�j�Qɂ��0!3��.yEQ���S'���G.���ۣ��R�&ʣu�A�?\R�*�X�M�̴��
��QIM�xF�_`��4�����\��^&��s����#���5J���N}�b��젣M�c�|��$������>��w�O�s����h�53�A绠�g�罭�{YYy��J���&������c�(��f7e.�����9�ȝ��	�F�k�(3�V�/��ՙS��o|�4�O�Y��<�x�8O�qq�9!~%J�R�Bx��s���ݯnS@�R�W�̚`���+��?_>���*{�򘡩۴ZLS�5��<,�f������8��yz�H�s��LP��g���
�G�&��6���scu&�p.�w�~rc�E�iE��ъ���}�(��$IC� 
��B�(�^A�lgiٺ����.�Z��#-4�,n�&�n���Kx�ok�@��,&�Hr^UK�0��56W��h+�׿�����s��L�uJ� �W�[�]��ft`=��.��X0l��4�w�6��%ť�����[�PE3��^��hF�񥛠9��J)���r7DZ�XI�F-3_���Eit���Yѩ�[��� ��3�e?�1ԗ-���I6N��e
`�t�G)U��ڑV����ђ�ڼ�7�s29�	��yIG�V僋��+
|k�����y�86y����-3�/�	��x�wm�d���?r�m���LSw����е���	�}�(�5L����I�\�Z���?�CJ�;�$��ye���o�Qَ�p�XO��:ڦ4�1Q��Q3��wQ[�ܝ�&W;��_M�m,v �����L��T=������=`�d�c�Q�_f��r�p��+�8�9�����#���_k*j�S]JIV �Q�(aq��$m2S�Ŭ��=���?�4��NY(ؾ[gxx �s�Ԏ���{�����.'�9��q�}B�ws�����򄞞Kn���
(
W0AQ��1h�"���@��"+g*A})��1&Fl��>����R�4W_�I�$F�=��jq���ք
t\��Hb���.���w�M�y��!�#�C6|'n0�Ir�0|�yS�2<0�Q�� ��@���M��VR"��vf9Ez�irȬ�U��q����|X�<��cd�i��5b�ձ�QO.��X_�A����9?B�F�7эo���?��g:/�-�Se�y���V��k�ȉ�����8$��SN�+�5�}mK����D����9u�����|"�{90��C�~z^��r�JbͦI$����:���ݷi�Uw�r�F5��t��[���;�wR�5#.غU��Ƅ��f�u���ﹾ�#k4O�H�6������Ǫ�~�Z�*�=�S�G����П�52�G�я��h��t��m��i��c�X<�FIڞ�OK�r�}g:&|x�{5j&-QnLDi㧷k��9�nfd�u�k��l�{X�4l���>�ED:8m�v�=����R["�|t��ӽ|$��c���#���'���b*H0C��W�K*�YvuB�M�O����&�N�Р�q�V<旌�t���J`H={�$��wY:d�i-�̅��
}�F0��5Z�~�ۯTAP��Њ�ku��
����ɢ������S�<��Y��(�<;�(bp�*���$�w���(:��+�v��w�l*�� J8&l��ߢ��v�+�4�#}��f������z'�!�~�49U�]�_�c�nV��J��� �Zp8Lh�"!��ejUDu/h����ɋ����K��A��~�J�0s4��
	�3:cq�z���g�*��Ն�(�z�i]l��W�����r��+]�!h̙ΠGp���:3w����_�\�J!U���;�yt������p���{���:��T�+�d�Z @��؎P�w��7�Cgߢ���S=�Y*ػx_���YK��}����YQ�M�5[Sk�l'����3����N��&�a��̗|ܓ\�ew5�yOq�Z��lh�&	�}�Riu�����ƨs9�ޗ[�@���LE�(��`Sr򩲤,8Ϳ�d�:͘a��[>]�"v<?@�f��b��"���v4�"jD�7��\��bƨtP9F,+�p��(r}�$���2aVK���n%#u�t��Em�ۯ����؎��OF�ݮ��md�H
��/Buެ�
������o��C��T����ɤF��.�����݈�������-Q��u�� m�wD/d�P�^�M�e���1^����o�m�B5��u�J;����9����l#CK��$a��-�	�w��wW���f�q���ת�d�1Uw>�d�惱y���h�th���c���.�� �������
��d<�QKa����S���,r.@M��7����qj��(t��V����|?�����!r�@���	�ԋd?��+*ZZpp]!�Z#��E�1�g��$TǠ*!�@0�q�)�q)妻i�S� \ V��������������\��(��"�Gz��Y�ý*Q�� 0EDkpjFY�g]"A��},�QH�>�����f���?����]�E}F�������S�\�Lz< �\�є$����8�[=)Co�)�����7(����	k#mv��G�\Ͻ��]��H�k�p�,b��_�f[����G����3��A���Au�`'g>i��!z�oV4^����dX4jJ$���e��*���8�pss�[z/ǘ�K\˂�]�˩���.Rob�c8 ���fH�rj�1�hz��wd��Z|���W�cƊ˜ӊ�{
D������Ú�)�D*/-SI��\^��M�\a�\�mcQA��[��Dw�U� ���֨R1n�TȺ3��w�seP\�G�*��l:ϛ��tῡ������X-*	��j�4�@O.�-��F��m8'�w�ʭ/���;��P'�Mϒ�,Bu(H�V�U��*�w|(z�6��D���
)��َ1jvWT�����!�\��Z5�sM���F��#4� ��M��c˯
Zg�M���/����_�P�zhފr�]��}�y�\Xn��I�N��1ǝ0L#���P8L}q��&�w��B���u"�,\J�427�L��!�ŠtH;:&�0�AOQ��* �
޼���J����/M�ޙ�P��CiWe�I	��B㐩��&���/�2��]��:}�h��O��]:g���x�����Z�@!��h<1�r������~����DV����,����_��#ljF~V������v_��)oUW3�����X���g�G��C�SS=�H�2	�U9m���U{.�M���%ʯ>�XT9 ��y���僈b���T2y=ѥ��!��d�c���xy�]X��O�:���:��}E����_�p��"5P?��Ғx$�ǟ�����+.�	�e��ܤ7������޼�<\��	�DE�a�́�ְ�S�R4�1�Q��n����H7���M���3�)�sӽR�Z�~V�-�uE���vFu�'_V���
��w���w`c���I�~�?s����S���@2-ۃ�@ Kia���2���N� ��,ǽ�Ȩ���H���qC`Qv2f�}�ٍ��e'�����O��L��k��D���d�?q����n$�g�[��񓆤2��Z��ܑD��?��%��=�A���L�@8N���ɷ�E��T8N��~�Wsa��Y{z���g��
O��+��p�Ѧ�L3���`< TX#�����7��gAJ���$b1]Z�����]�!�cԤ����y2l�7�����|�d��bU�=2"�h�T�2~�Rt���]8�|leEP���،8�
�饧���P�]��"��:� F@��g8�5�����lkS���4�+2�0D��}?<�k{�@N�8�q��50[>k~օ��"���V ���֧TF��3���G�u��,_;!~�]�����vh���&;� ���E�������rϷ�H�b#��%^���t_��v�ZP��I�+'){���{��Ҭ��GB���9�w�ok�}ޢv[d�~��t�^�X�q��O$z�M��"EE(����b�`\ӛ�q���蛓��0����F��:9(�2���y�����N��$A�z;c?ƞ�#@K+4���y�l�u�p�įVZ�Pp2��GD�
%���n�������"�� ��)�)%�X�$杭`�
f�IUk����;Bk�C��c��Tm3E�ƹ��w����Ԕ�Ʋ��ި�b��٬=��av+У�OQ�3�ZnI);Kx͗��mN��!��JZ��jQh(��1r��3��m4����p°P���[��1�Y��gp��2Y~.\΅Gap���siBoO8̥�1M�'�_>_ሑ�-�kiC����;ƌ�9���I�#z�]���tic_��9�������S,�i���'4陣v��0;sq����/�l�[MeS�ڡ}�hV�,m�S���`�E�md�,�-��V�L��}|_/��d�j��%��
����&yU��`ķ�]>�8�0%|���W֞�ɳ�����?��hox������HH?^;<K�ظmz7�Ԓ�H�}����7����IL�Am�1� ��Td������m�7@������U�u��x7�5�e����L �OV#��ct�ғ7GC��^m���lu|6��/�d��F͎��K�>�6�V\���������R>�d��8�`�"����b����Z���ƮU���t�ʧ@�u@r(.t�ouǗ�_�ބ�G\B��F}E����V���ޙ�ͱ�����
�]������eeS����;W{����۷s�*�7�:�,�U4?0`��쑒�%�5Uu];�����R��I-�8\T
8�k~=S�G�Y���e;��;F+q�V��N����V��#�#�~+�B�$φ�G�Z�d�y�$�2�؅�o6��
���5�G�"��%|�]�R*A��z7�d�"Ӟg�;������.��p�v�?8cċ]M�l�
����z�UX~��_}o��n�T�%K����D b��=r6|G�����q��9�1Ѫu؜�3 }Uba�N)�&����>�$�#�{{��3ZL�p�Պ���U(�O�r�>'i��ߌ
T��(�Q�9�U��(�TL���K��M�����+o8!��#�a���N+�;������y�P�U;���W�NQ0�G��}Aw��(̖�����_�-��Qu��!)`(��I�,�)��T��?�p�<�f�����`�7����c�Gɶ>��%g8_���������o!C>X�}�!w*ϘzH��~�\�c)����8��Ir�==�M�F;��=�D�A�4��C��A?w�|&=�$�@P%k"Z�A>^��b�q�zО�%�4�71U�@�ɌDeGo	i����8�ò��.$e����B�u�i�
��F	@��*|��)\��k!v���㵏��nN��~���!�O�qxE0�� ���m�����H^�qS�I�lZ4at�� pln ��#G]t��0�}N!�p|J�/?W~e
��hl���EW��P4;��Vc����IJK'���:�9��B>��bD�xkJe+�TJ���u��Jrm�N��� �����IGԵj�|Q^c:tQ"cƻ�,F7&jLǌ�(z��OV��C'��[Q7�z~�g�:����)��7{Yk��*I��¬O�>@J�5^%"�ǩ�h���
*|����P���E�'1B	+q��ג�O6_�v�/\T�u��X{=Nw�a�ˬj<����(E9h/{#�1����ƚ��w;��J�~�_G[��A@3;&y�隹簒@�o$4<X���O@P57��Wj���+���1�0��A�l�Z}E�3ͼL}�*��*��0�GcɩX�/H>���<��\$ ������K*��yW��C�1�7�5Kz��u��%�$�-�=j5���@�ݼ)��B�J���|��=�E�KˮJ��*��fQA8Z�����!����x�����q<��uxD=ѹp�P5<p��U��n�� AZQ��$_
����V7�m�{��[��K�+�n,�T%0���z�ǆ0�޷/Ｖ����BǕŕ�`]j��Syq]������|Q��5~竒?2\xҐb?�ʋ
<�L?-����' �@��F���x��su	1�� ���е$�W!�9!�q���q{I ����)��t�nƎ_��I���G�����*���a7ϩ?�}�p��f�籝hM��C}q�9�#h����&���{�\PCt�yl-n0$��ƒ��V��Ӈ�Q-wI�#f'���sH��������F�y��n�-=�q��)cy�lV�醱�HH'��ɤPn���9�/R�
�������l�sY�-�HV��8�;Ct襕j�;�Ւ�{�=%.kq�I��K����׆��T���O�IB3{��p�U���fx;�K%F��L��,�s���H���[@N��N�z�k��V�C
Xn��xG�V�oJ �ZQ��8-���,�0�c��G&j/,�39���@8s�n�����?U�p�������tՋ
�[=i�0u�R$�n[nY�`�����p,̛_nHC��Wj+��?\���d�����HU�m�>���3p��mf�:�m�숀�i<��H�/�?	Y7�KY�Jc��=B�`�]Z-�x ϖ����6�ɖ���#L?�r��iԩ���a���4\rC���CR�?��;�3�|;�0D]L���
�AuP�9a���*1I���7B7����5�#���)A�!�p���OaE�ֶ�͊l/ʾT	�|�#��7'^{J�f\��8LڨC�ڊ���ḫ���?������Q�����u3VДR�%a���r����`(qȥA�2jC0���f�x�2@��W�v�����	,����X��J�F��K�"3�1�<^��cN�Dg�~�S��o�m�:z�P��7ɾ��p'�P����u0Rq�(k�tKz����� MȌ�z��E�s�x�8�a���NWY�[�ň��r�~*��0)��_ j�d8f�V�B�\�������_�ГY�\Q���2��@|�~�!,��jWM�#v�����6��@0
p����n`������1,��+j�ɢ���	W7l%��ɞ�+��hq�V+E>�M��Z��?;�����(�̼y�C`k�7�h� � r��ɯA����P�³��ZÏUiA��.G�`�X�ʔH4E ��p	�i��Xv��oH��(w6���B�r&�g�.gG��-� �X��@�l��1eK�eY���i���}�����W����1͹�풠��ƀP���
>%
�"H�NI�Qڄ�,V��?�8|��p�/��%M�:w�0��ե�!���k���=�6q�=�ʮ���\؇�,�r�L\�u��]��!"�*(I|�"����9a�MK�����[&�A�5(�#�B��ʭy�5{Uk�z�*���l%����^� =N�A+��$�Bt�a���U�:-�[���UAJ�<���/������C��Y�.��}`p��5�lh2��n	S7�Ճ���=9z���(�oR8T�3�
�+߰1~
xG���m�NЫ��B���hI��X5�gG�F;΅M��v�B�8�7@g0����7A<�U�^�k�H& ��G�f��wClV�/�B�yg�h�:h�i����f4 ����=e�!�`t�P�����\�t��߮��CWl�;U'�~c��[L��l��Y~#avOi�����-�3?Ǣ��R"(��HK����K��iO'!w/y�_���̛�b�����-�26��5�/������<H���5���۟~��x��A	�da�D���%���8��+�Q�\>޹w����>4�b=<�F@*�Ma��'��Tm�"���؟��P����
L)�~ww#>��BZ}h&���}Kx��N�TLB;��h�m[1(U��e\�XS7I�������q�������j��|:W^(�Шv�8&Ĕ���Mv6	b޻JKU��G�"a�! �Zq�xo��6��	��m�~�"���Ez~=�W��؝
:*��ȋ~ !	j�y���nk���ژ��V�\���o����� �	��d�(��v��� �����l+�z�Cq�@k����cv���D��u7|�I��[�ۉ$l��B�Bf��(/`�tT�IU�b�	o=��u�5(i/�`r�Uv<"^�3��_��[]�{�a�>o��Ą/���;�A&0�-�w��H��k��\�M}��?a�p[L^MpĎ#'WN�3�*�t��DZ��^V�wv������cx�%g��~V���_d�ݾ�������r

Y5�e]��m㐘��G�c�[��\�Ϳ�E{���=:��Ƽ���R^�9��]2��\�8�9�ڛp����1�R����\ �>�1��qF���o|z'q�{g���>�'�>2-�`*_n��.����8�7�Q6�_'Oh�;X��S)�^`��`����޶�P�9i������s��"�_'����r��g��/%����l�\�P �	@�����F"�9�6�7?7�&�yae���(/���9���j��Z�f�LD���{b;�8�SM�5M�gK�S4'6k7_�m���fO���A,���_j$�,I0�֙h�a�k�R�����PZU�h���}�'H�=���w���U�ZL�r=+Y���(���Tĉ�
�<*@m�E6���`���C(3�L݀�ȶݰ�Ѝ�"�*\�M����d%	8��}arO�=�gg��?���ކ�^O���im�6����|0�HƵ�Q�t ��y+��8�Al��\9�7�[���o��_r��t� X�;�%j{ ��C�#f��Z���.�*w���C.n�Yp�mZ:9?����	v�8	�� ~2D�<K<؜�Thf����*T���e� v!����HɚԌ��9��0�&���m��7D�Z�t�n��Oh��g�1���`ą]5F�hv^կ�� =	�k������7j0��Ĺ�!��Y����6���+�G��Ȓ؊��T��s�X};�v� Цx�D�g��k`c���mfQ5��
�`Gdje�J0��'%�kxJ,/.{}�^ �$<�K���=��?��]~��eՒ�fs���>ȼ�z6xQ{�v:��'Z;���S5m!�G�o�$ή�7K���wm�"/�C�dk�Y)|�֏јs3�1.�,ry[cV���]T�s�!8Oeh�Ol��$|9�ڗ%�'ڶ�����KP��Q@��0�sf�t"í���R2�%�c�lM1���A�TK+�𑝷R�������c1o�m:B�E��à�y:�;/��3�ŽVv�	��Y��a;�%�t�0Tܣ�?DW���fM����⍭��:��"}.����ƪTi)s=��-O�}ߦ:�=��V�@�}?�[a>+����ܑ^+Oo
��O�>�U�K����	���B�R-bp=�F�:(P�M�����*?�_�[�w�7��\���l0y�m�5(�݈���l���,� H��V��6�]o���vD{��n�\�rYȦ_?N� 03FKXƲ5[���0~@��-�m�.���{7f�*�_�_Å�߸(�"堬DT�}.��M��Ȁ�<�8�Ub�H'�t8O���bF��E��������*� Q���E�S�-��¹"Ow*	[����	��A��]���|�'	�n����ʸ��6�������3?�]E��������׉3�>I}�1��sg)k�E*�"�jUHr(ro9Kʨ�Wbk�:�G�N�U�z7|ُ-�]2Bo����.��c��aԒ�����E3I#�zY��3Zr�*`�l�����
�e]a������9��Xڧƹ�>���s|g�����x�a���p��͙��в�9����ӿ)����X��>�#^z%4@��/�k���el�W���>�7x�w=#`�+C6(`�a����8o�9�^Ya��
]3�1�%� D ��c��T��	i�m�� q�t^��r�0���p<R:��nk(�	�U�����䴪�ɳ��DZ���Q�:��! ����k^<���tx��JȦ��x ��<� �P �c-�t87>p�̂��m���"�,���Ӷ(q	{���R����(9�)׀�=Tf�eʙ���
�I"�����$�U��(z�Q���{E\gApy@�u���{D�*CI�'�m�Ƀ�B���ݑ'�2 A��)�bJ>��|�Z�&YT���\�^{n o��	gB�>]��y� �B���?͎B�=#I�v�p��SM���=[���vM����-�����݉}J3cMu���l��*;��\8*�`ήFk �rV��0gE^�OH��<E��	��ıH����
�s���P��~�Z��Z�(��L��e.Du�V`�����vh,7m��h}*a��Lp�J'N%�-
¤�9Q�ɼ����b����׻Hɻ�u8+}Z*R�1PF�T8�濠���Z\�'�m6����r?~Z�p���v��~p֐_Bxa�����č5%鐇�gD��&���d��9��-[L����6Ԍ��4O_T���";܁��ڥ�1�fY�Dfʤ�s�r_Ê
�X
0���)�h�-Z�n���yXj��E��Ʈ��m�c� z>��@��{=Q�o���e�t����>��n�������sˉP=H���#�'m=E����&��E���]�SL���F_�0Q�n���5J���s/�	�)Ǽr%BL���u�H��Q6v��nl����<�_`c����ՋF�ڭ@��c���Σ����S�>�p�([^�杠ɇ�⃠Fm앟%���J�N�h_�����}HE`~LK�������Iڔ�*��/�nT�n��Fչ�e��8��l:{��e�_�R.DBY�,���\�KՂ��f���;l����)�4!�L]����f_�#���\�r�/o�$�ަ��*�P�I֨���Hyp񂸴�a*�7�׃�f�$4�o�!�"��wI��'1�������;�ѐf��7p��ZQ�`��wo����J~^����/X]�V����ŔB�M��b�������k��2u�NԃP��
��ce��:vRu�85L"cS��,�C{ 8����
�]etJx-���%h �SIO� D�r�0���h,�
�}�@iY z��1+���G�sg�8�I�ʥr�Α�z��ӃFNɭ�������	/>o�ɐ��~��%ʽ��	���Ό!0Jj{���1=E���� ��.D�Z�w^�O��w��%�� <�1����L/�k&s;#�vP�C�&:Z[>�y��,eSɽ��؀r1�q�qԹ�t�z��"rk���xDɫ2��ᠷw�PO�cbκv��"η����O'Ҁ�8F.��4H�U�b�9���m]��{@�H�X/g��eZ�k�den[��u�9�j�e��9��g�\��;�!h�4Ի,UFo5ȧ��K�Prv��G̚���I�py�����
s<e-]����Z�xC�����
����j��B٬u|DiG�˕L(���L���l	��X$",�QZ�KC�[�J3*�7���l���~�j{�=�XZw�(K�z���O ��e������c�]I,��V���8��=�]y�LBE��J`�BE�@r���{���>���r���&��) eAw���.Y�7�2X�ۦ��mi�9��~S���>l�<�NZ'f���,c>��ӳ�˕7�^j���a8st��ml��R���;��Ƥ�ٍ���2�bv��w#��5_��p[�{C�w��z��k��_�o��(:����tS��<��<I2����q�aE@�X1Q�p�n^i���	�a9n�qt��.��D�U����?�G����	;�Qɳ�]�C��9�/Vڛ��s�;��A2;����}K�|&�q�i���%��1`Q�2� ��X� �q�F4���.�L)����E��,j�O7�isfv婯D~����Vg�R�6�g�2oح9�R7i=yM6�ܿ`�'"Y��n���-yڳS��d�Z��r�]�wW���(����#!݁7@�M�9�-(���>Zۤ::43�� ��C	�$�N^YF$%��M�s�rV����S}�6�+����8���v� s�Q�ݦ2�@�#j�X�tmA��8)��N6��.�M*��+�!�x����g�}u�V<�`���q���y�A�ՙ�X3-@兣v��TF��W����⫚�P�:���� x�}6AS��${��戮���56���Q�� =Dg����9�=g��G�bii�RU�z\�o�z���Db�}E�p7�������+�hDB�Q��)WnH xr���b 9�Op��^ T���B����i����ۍ��$�x�����G[aſbг�k�5J����J����$��O���t/��k��3���OэsjN�ר<f�odl��Yg��_�֨���:���^(�[�5��h��<c�?C�����T6�V&��DP�|-��ݻO�e g���k�{�0#�S�w�ǳ�+�,���;�#��Q�x��QGz��!�|0
�*�����
�"�1BC���[p
��?�e�i8����_8����W�8�K fs�}} l��b�ӞR�Y�6L! ��{ܔ��ݯHF��������S����/��U���3�>�����χ����z��	P�5��S�|�=,�- ��Ո��9����C�$('|m���W�A�b�;R$7��W�?�a�1ϯ_K#��,�p o�vG
�Mt��^�(��<�|�'Lp�y1^�F2���y�,iS�aO`(F���]�?/�n�^�"���ρ�ޅ�;�2�YSB�-b��ik�&FZ����]<;� �a���RC�fgr[��`@��v\Ѕ|Wݰ�榹�	����l�8�T"h>���=�d�I���j7j�ϟ{�����s�H��a�Bhk�����O@��ɱ�7��:���f���ֺ���I4L�2M�3��H=`�U�ĺ���P7�V�R�b�ֳ�.���yL�R�C��4�K0���ÇD��	=���F���Td \�\���N�`+�|CTζ�i�.}����B��=.#T�ŵ%F�Ң83?E���wܬ�~�c��*��Ԗ3X�����ߌ�~F��훅����,9�Xx����q��a�;��z'j��`��-��Z�X�v$Ò��wk���x8:?��^�\��`�^;/���	���b��d�������!����u-/h�8gV��W	�:��"l�\̅
����p�$A������"B��K�o[-D�q���Z�^Ҥj���7@��E����l!� Fɴ�I�B�M%��mu����@OB��&h"Σ�ݾ(�wiR�� �.O5UJ9����Ԛ&eXS;�Ob}��]�y��v%o$ZV�k��Q�fB��゛��չڿ��;a�<yL���өg:y�%�s>��?�H�͗�\�(}SQmv�WQ�)�A�=j:,��7���"0%+^\jg�ԯ���Ґr �c1;p��N�􆎳���cB��9
�V0��]o*�A�gmhۿ��*���i	��o��n��}�;�.�K��ݘ~��o@�Ǣ��&Ҫ�zh�b�>��X�1ߟ�`���Gf��d ��A.?��\K�����-)�UJ{�\Nݫo�������{�^�h�wfrA"�:!H�.r��3=3.ࡽ+��˘`�.��uS0��� Q�y�8px�V�\KJK��	�|L �(�%��^q�5����Ɂ��ynj���M���p�/��F+�6��jU�X���t}��M�(��ǴT&���@�_��|G��#ݵk�&Wߢ����>(�Z#����k�����"���!���bͧ�P#Ө�m
ah���~U�Ǚ�]K��Ꮰ�>�=:)o��y�!Q]t���۞���9Pݽ5���ͬeD]|o���>T�.0������`3�O�5���D�H���!���ҟ��_�@���?Q���"�m/�VO����9��S�̓�r��	.J�	T�@Q

 =�C��Af�i�v�T�m$��t�Cs��������hիW�V�ېƯ�ʕ��Dgu�H(����m��0x���b�e�<�3X����q�?�z}�������1X<	��'6�ZK�o�
82B����U6��s�3\z�nNV�U�Τ������7�uƑ½y��EL5[�����.z9��)Yn�b�߸l�v����V�ek�d� g=0�(�f%�	�0↪OK"a�a�(�d��:�Ł�1_YA�J�iǪ�n8>�!�E�~��X�f?LetA��dR�0P�IǊ���!&ߢ�>��K� ��'O4����얝��	��Y��rVͬ|z�^���W+I0e��p���v�O[o�����rH��$��ڏ�p����咣:��jfJ����C��x�FpW�������-Y�D �Eғ�p���Er� �-�x�%�ua����5�H g�tQ���	�����=I0p�,���k�� ��O*�x�+����La�/}�zL=��`IQ������BG�xH��O~�֐n���h
�U#'Q�5;$IP�<T˭1���lc��ǣg�|hx���+�-�~���^_c#��A�RF���Q�'o�+�����V��*P�bČQ��sK|Fz��i�ܑ�	G���� �o�~��Y��K�}]��K���Ax���#�;y[f6vEF9�5���*�7@c���N�~���`$��E#4�"T��#���+�7�o8P�0�Y	Y��s]?��u ��s�Z�W��Y/69
��Vy�T�FEi����B8Z�������%��"XD϶�Jx,�Z)����Y"���t�>�i�F�)D<�z�X@��b�y�� (?����4�J�џ��:����np�ޘƃ~��J%�H�a���p5��Va8h���ug���_�]�����c`M���K=�o��e�����rͯ}�v����������`ǿ��*K�M�{�;2�Ǩ��u"-��m��ȣ��$�i/C_Ù�'�_4��]{2�<2��T��]���v���n�����S�G��j�?�
�KtqeՑ��<8�D����r�Dt��'��?\߿D�r)��xɹ�k����)�!CxJ2��5�˜�	E��@���tt�R�p�����3�*���� b����UF�ƿGe�+�H]jD<*�U����!��fW �.�[��F�M�+�l
U�� �3��:1��Q��=���
����>�l6�e�qC/��,�W���&H����j��ܓ��!�ܤ�+�0ьR�Q(�G�i܇���U��NV����[$�f)8	�6���&Q�(ʬ��g�zT�%bc�?m>=��y��t{O�m�?	O��%Ws:{�̏+���t|@u7ś��T��\��P���6��HYn���V7�a����R4�=�Z����m3�,A.d�?�a�:8�%Tbm��E�G�n`���[��J
��� � ��}uY7�lZ�ĂF�`Ɵ�'[R	�h�>�̜��o���EK&_5Ϭ��2R���?�-��d}7J�m�X�5x/}ylW�L��l��u�m�=�f�L8��bt"j5k����
9&�'����h���w��wId��ȝ_>/B��12&H��-u��,��=ԗ�%(}�B��v��j� ��&��z� �Ŭ�W��^���ߨ��1��j��VV	�J[aiIq�s�m&��Zqg�zy$��qJW7��B�+�/��k�Ƚ�������'������%�� ��D>[�&�<�����_j�tj_P�-�V���C`�~>z��.��@�A�Q1V��*��C>��5�<��7�ٻR�m�e��CEe}j�i��q&Sv1��3�ཌ�(Ty��z�ƃ�r�U�z.�I��6�}�ӑ^[����_�u!�VZ��4pM�����������Ӷ.*��甁^篴V��8l��`o11Od�\.c�{��s2)R�� F,��Ho�����oKI���۔I��ĥ(�5w�SjI
�JI��=Wv+l��<�Of�(�)s0o�K+���#���������wZ��5;8u0�]D�Q/v�zs-}?����Ϭ�+Dm���������H�fa�B�x�N���$�-��<����j��D��('\{}�Y��Ow��2��n�uv�C�-L���A���;��>�@���z�'�]R��7W��]?AH�n�I�]Z[x¡ô(*k,�������or��:��}�h��j��iu_}.R����t x�Z�^/1�L��~.l7�Fa��i^���ǭ/�s�Bg�_����j2��ISZ.���_��R{4�j��ʄ��k�U&�ʔ���z`�M�Ap��A�$��I.zV���&g^�A��>����8�~K�?U����=>a�0��r�x��^� ~*�!Pn�ꗤ�A� Ф<.�.����w��j\Bfl�J�LM�̀
�B,���	8u9���4K��zj�ըN\��(wA��߼_룛\WX�}��xY�A��;�B�:'����E)nV����,�m����U��UXB�<B$�2�����^>^B�'w���p���9�-5��&O�٘��sU�c� �a
j�����Pe'����!�H�~.��]	��F�>EP��\�Ԋۜ{��5�����G�-u�=T�'c�-\p{�e�o�h��H �w�1N)���M�=�����R�A�Y����Y/tIR�p�
z����Ң�]-9֍0�i��=g��{ɍ`�`�R,�lY��#c'�/SS�%������A��|�Π����t̚S%��40���mm�3�����ջ>��L����z�ASje4Y(WE��$p{��@	��l��ky����9�O��B��z 4<ޮ�J���;���ÀY���|������z��}������2�����u��zɤ��^T(�m�HJ�ާ��e!�Dj�y��-��X�NA���f͘�3~��ϸ�'2��r�(�7�#� ���Ԣ��d�t۫&���=����/o���Gנ���w����9��x� �|��o���/��������B6ʫI�X �~~�N���]
A:�����~��Y�FXī��k>��Z��,�Xn��!�򐊛��XU�r��7��"���yQ��	�d��bઝ�La��"����W�˘�'Y�����u؝`S���6P|GH���Q��
���B?����{U*��8q ��I�֛�x�}��{K�~�#W$��6q�~"�}T�#�~0���ؾ�ʭ�9����:XԪ�ϯ�<�#���$���z����aN�ڎ��(xG��#B�|�WM���������:sN� �v
ٔ�@�P*�$5`%�| �+�Qo�?�l��^W��$�ɝ����D��*��v٧#�nŘ'l���`�}�0"�v��䅱�#��9���p�������i���4?w���jm"O(�ҫ��{M�~O����.���ht�D����W���p�T>c�d}x��r8�j;��ɑ����oE}��/2�i6Ʒ�