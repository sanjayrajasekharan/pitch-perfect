-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Y2QLoUYHHDR5p2Ql+/3vnEsOjOo79VdKXdg1leL67O+5IH/r+n4uy26h01DU1CX4
LApvDl0g+lYZT/9No3XO9rr36iFig0a1meC7fbITSwZsAv6Rzlr77v1TqM+Trp+e
tDeg5fDKqBQSC+Cr5h5srz5YXv773e7cvgdxgQ9i278=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 22621)

`protect DATA_BLOCK
5eO/CVGjls2aXXRIZ9FLuJOirfb6Ze1mQkBmlszUfRQnn6YTTYmT3rZ+jWtsIxUy
t+piANh4kcPCyuDxdNhpJMdpGrnUxCqLp5vkGlfnss4nTvjC/+wpkCUgHySEmXE7
jFyiKzXCoEF73Cz+JA9aNmtEjWeCwFAonJWTavJKaJNpbR3Re9JTa09eSd+Kert1
a2UjhVMIKT5pZZd1Q9ESyJ+zcs1q8FSn4WbTjYSe7sLixjucDjMVYt0bAado+AI3
7zQ+ptnEGZUr8wTOQS5xYehA0cDQvxID9M/pVrdY4i0q9FekshIt/hZpltHRu3V6
hjuUSe0zLoBg/kR1A0KBCG8f3jaJKthVCXjcZJLitKp+VvbjcjRLv117T5zVX4EY
4H5jIKVjcYe3av38hXYSyNq/Umc6rkdGsZ9TyCeG8meQtLgseLbkDffle+TLw4eO
Wyg9Ua79hKDeIBjeo8bxWmkBcntspyRp7K3RT1895yJ9s124xP7HVykxi7ghIrcv
CND7ov+S83Z8x0vxoF9ztJYp72TKaMzIyB7CQfOUCTXuhFwwlcqE04I4w1wUTH5u
AnjcK29aluWC5ljCMnEcliPP3m6OFw9Hjz1G0U4NBVdhgoQr1VGXKarIqgHzeSXB
MTHDCC5yaLcIPVN0/FnCzahnJHnINBmg2Vd9tEU58W3VZH5KpRN+Hd6YX6TQF/j8
TOYn3w6yi8zrA9iPtUykh6W3ELn2BZd5Lz3ShaJdIdeJ4y6YcGa+8LkuFHFddfiN
+NJMK8tqbb7DNNJl6RwSVCr1nywEN0o+STN/NuQZtw+bTJambECAoPArRvpKLkVX
4SEgRHss/6ZjOopCso/A0I3epOqb5n9ZozPL38wBUfrOdSAviSQDeTzjMS91ukHk
CbKBesP+S8emtexTJmp6PDeTZvmFvA6c88KdmctFfRJ6N1Vdld28PQTOPNgV2w4j
lPL+8QjHYwuEFShJiB/axSBqldpqGlVWK0fKPZEZFRFbKTZWesqUzvDf/buI+Asn
ECMg2dI++0Qd/XdyAoMtIb+6YvrMjOc43PWE1iL66cSLjYUp5v49k5WKSgcghc6q
IlolJBayya3ep+QCpuXsyLol4pP+anpzkSmnfX6DWei1CRHcPR9NBfZp1UkYS3ZF
y1vnMvcpCFNkY/00dHzHxbkCKQr/Wyjq19zDtmohhwxaw/LzD2rf9GoTXi2l4iSf
iLdi2HTlIjo3dzYyUS24j8WBjc3zLUUsy16Trp1IGOne4gSuTrVaQMtmt1mKyJ3y
uZqbvyKuzzvcheeJpN5+QlUaVMCqqIFToWifADNV9i7s/FebqjuGei4zlps0SFfO
Na8FaF+z0M9JnR3NV3qFFs8oW5wRpi+6loWbLt1LsYROyMOODmoJnv6tgtjXZrEE
HYO8dGft8smrhO+uyWBuBzGLzCIauZrw1WEfZiftIqCE9jHQzdXOZzfVWRNDOYzi
4LREsRAoGOCCcbLya7VJRua1q4BjusZOiWjGffCx5VzVrCxwEescvo1O8JH509fb
xIf6S5vTaIIqQrRtN94g+yG8H8L+rOTqCb1w0/p2NUWr0+T2SlV6/m5b+yymto06
TtqH3KflmBMrJYMVVZ1kw1NHBMUbT5gMWa9bzKnC9qlEHQ3xX8CQS0N2UpQ0tqcT
d9E0peybudRewVT52pJXPFXj3j7OpHj46X41zH0ZpgLz7SGl+u+OUYHOT90Epsnh
cXVE8nGfmxjefh1MFGvFKfiovmf2RtcFy8GTV6YG3fuWVXCMgayvZOEXzJkkoiXy
Wxknwg1jj3UBVvFPQN2VF4JkK7wMZ8IQsgIYl55z/yROpWz/1dqZMDqOErFYo2Sj
gEswaiqk/oi0ajABn7PDPS5qpoyDI4J4Der+9plMKW0b3PtkK6ncas0YE9F0JwzH
fC7S6pXvubUh7kYD/dhhxlkqDkPh/AXIO6OKCWv+69AjkiqSGurV6krPdGV12U6k
kqZYxo+0+ST4T0APQVvgnt6JZB8T/zzVvwI9qpKJub0bgE9fs9EbmWQCBIDkAYV8
NmsPOG4ccQ7pYynbUOuKSt4dwxYWSePu4yjjSeXJ1THhpAvjzuD4fygPcOnYyWJv
FVpZ6LcnpLK8EZzEAoJ5AiBOdDMeEqxUIYALLG3pwieEdGW2AMkpewd/aTWSJPno
1PB1/0/5rh4OhowCIz5qOgLNdW0kD71ualsGdhvtyCigx2W29GhiI4aXHq/8oFF2
hGQDTSBC5z1L9kU3QZ07gYOeaX7Z4iAnAaevMot5xvoCl8sy6ot8I3LRVkrRwcCZ
aa+Fqbv11HLWOmsy+ClTl4By/1A1KlzJzQ9SDDR7iC09xd03tbOuIel0eA3EthaO
g7cJK53abu1JtshLWkLnGSE2a1uoIqMp6enHng74KEelXCJRZ8rVTMbtxNngr+4m
pcOGF7lRQlYNXGr9FyY6RPMu/psifBUbL0ZiKpMC7cVe/4WzxWSLRgmA1pgwI6cV
bUjmJwvMBoj4I9+2cufeZCuZ2hrC6ifiGzE0AtK/Brk4rNUYHXmyVe+pL5FqSYqu
g7e4/zDycvRZdX7H2hh9X4CVC4+Jb1c0hzDfT+FpEUJZqtIjLx9iglXZcOo47MQk
1m+BVO84I1Db5sbUoDJHQtI9RhaECW/eWEfHbg2/PZbhqpwn5OlQoJrxiHymDQGf
EazHqOfM1L5nCxhkEasHc4UMRoT4yj9nlwL0dwejzXIC3n3pDfcXfuNZxKU1x3bd
Q/mpTTRdfINCaFBa0fbkJFIkmvKcVJt2pDIc0wAmImB7l6QxIr7fJx393zurLKna
2NQcloQXMdkwjk7bGB0S7ZX8PwfhDZBqAf9YaBvfODNpoVD+S97nxGL+7TfVR/zr
IPTiwDsY2Tr5nxkzd/WcxZnHrGYVArLYWW+pvQfQQjKtCmgOLExOv/wAoKB2QUeX
uGLCY+s6bVUDLtF1+L1lF39zhb4QQxu8aBr9JbHH2b2MAkLjACLwkxCsYysM5Dkx
NNEtV+/tc4SfQPZZJ8tDwToYCunOx3p68oEx6jMLorhHfmUUzbIxgeQIpdT95mIk
nQ00oyVuDB2uPp7LFxmUJYMgAH+DsK3mI6KhyowpaVWUJLEt3+RxqRBNVfntuL10
XLD33i7w68jb7wWWtEI7YUBdBrS00v6uielbGHmX9QN6DY9QuKX5b2c2l3N7RGNh
YEiCThCMLqusSMPfkUuXORTbktedx9Go/1+zJ3aYR4ZUEmHeamDDggAo8aLpubEu
2HlIUMYrJbgXdyUSAolXi70XfHkDo7TPxY2zPxshAK2zxTxfKVS5uSZhiv53x1eG
G9hHBHRYkGds6eXZ5lb9Ty/3zjuR6JICXXinV1HB1mtwS+FBcw6HmS7lbnBbNBDy
ApjpCsM5CODqnc1bNRMRr1IsVef6jHeqcdYgtgetw5K1+bTPnE0kvYiQv+fZkdlT
6EJYtfPwF4EyXu1eNVKZvKAtQ8tASnremP8S/gN9N5e+Q2CC7tNxtBMDV5zEFBjR
XsTAbMXi2rfD9KKGsuG4zOv/BJNPTxEqSgRyHlebtV+UH6xZEipVmUNlKCb2/XDj
V/cKoZ+Pgoa7FTN4w/nu7OwzJQmiSX7tMcwchLlWvuwDEcVs77g6iC74Qi6WmKoT
9U5UDxH+AGbAuUOD2dyR1UxoMQEFU6jFz8vQbZxtTU0djqHqSU+hZD84v/6deL65
S2F0omEUe/uB+7RMuFJGtpvPJmoK+lCBbQjZg+vzHrR8EMXWLRf2EPxSidNPemzC
jJX0uy14misNlYc2R4PB2/2LC6HIA3pD/GeJndkX1rchWJ7JN4d7/54GWc3SgvD9
BYKCMXcn/fiVUJOnzD9ogXEd0a+exWwro0b+OuGNHF/PnGVM0NbTUCbUvQYSrUJS
L81wt2W0yPPfd9y/UtBRXje9OK5+V0W7x/vW7BjJ25hInw7GJsUBp1ihEXHS/Zm7
xD1T7a/PCLNq8g07CbH54EgArAeb+GBeBBXEDb6xRlVAQ3kPD6ebFxIigj9VuGG2
rOYANcC2stsGxYBavDBeNUsb5+TEnhSwyp2FZrWeQEuYaVGm7GlCZ1Skt0SOKM5Y
6ftNa/AH0HlmDTiApyRa6/9SIM5zu7Hi8HkzfRETSBIHY8Ew2wr+qIhVpqzJLV+B
NxdcXNc4/tbxPOfjGSZtnULLANEPwrsJksfFzNl8mkzUzkyOuhPUc4YyXpNC3de4
EYC1k4WUZIvuWNOYf41klrWCj7KafbPmMGAwQWzQHfIk8qp3JedWr5C40LG7zRgE
nXCWd/S8IkJfp3H5H572G6GiQv4qKNZUnx8pLZNDGquT9eUouVfTjwHm2/R2BChy
8Pmzc9W/RpG0uQjZ+F01ZQR8xt3r4oRqrmfR3qkQrEpSWqEH1JllBxFYeNI8WF0C
lGdhzQtGAeKJM1ayfskt06uiXzqBx0iP9vGjcbviFrEuigVGCFvS8+ACwxQROKK8
UHQy5+y6MW7HscIuvUZTp4tdwbBjcMYJ7m1T5RJh98EPy7htFeuuzF8Mhy0kJk3+
qTzqQM2IgRXHGnxpnQk0BGxxhN1mPzvwGhI2vKjKQvDh+3if6ZZzF56H3SrER/yG
S6Eewzrd6IiUqebZhH24tbjPc+GuxPE1h4QkyQSWz2pf5Z0O4dv0g1iFRb9Y9VFC
7W2aINcECXa59vvLhMLpXpGZwSIs17dxerRwkHIJ4ajbO38HfEOchk5v6EzvTHBr
hCM1yH+UIT4REu20C74uXaWdU5oEWbmU4F3MN0VuvaNsiaksm3mJxrlZR4xNUh5b
kmAeG7vcoECnQbGXKWTq9omi5Co5PIIr4fUZqFSsaiV44Iu7tjW/zUeqkI/+d43q
ns5I8uyU4/HZfjK8c5m3OEERtMSlNK9YRtMI3WSyWLUORpcZfjth2QkvnwHLkGxF
neGrU9zBKFu+G2tKas5yqkXzy09+gnke5eCqobhTs/bb4IRkbRbtrKJzozETO8J7
RXnipLXxGUbCy7m6kC3DFnXFNr6iMHhWY6W49O/5m0ZY9Ujp3eDqaDkU62H5XAjL
ruDVT4XJZ268nYt7quvLnEJU/Yg7S4GvqPAIGqCzZakCYZQx6RHXiPXyYOlaoU9S
pOHOPJg3hIaFjTQhPYdjRrb0E9F2A8OCSQHP2nr9Trp7BJE/JT/LrXLgKlMui/nt
wcqjx2JfHdL7w5Uqd9imJcDI8QVq1xKJhaTq+lbPpxIChL4DD2pE9/KveHmNoGa/
7D1BWUgplpMdpZd8NCAN8stYr5MBblB/+2iRkYOtRduDjh56tWnyASyPKI9//Hts
H6GBaiZckM2RhRg47ngKRj43sLOs2gH2xwTBb43cGZqdFufQdsLUBnvuGze0apgA
qv2AKluMZQM0AAPzz+hzHA6HmWHbSlxJ0jsGqll+/nmzrBrLHT+ZCsoS7pxbu6jb
gAETyDRibqcx66fXHK2GaV2Jeyc/qAXPOi4zK82vZm54W8d7xTgZIrQechnQZhIS
3eibDDZz57UoQMiEaLtQETpRRshlcYmC45kEY7ASxemhVUUFac0t9XA9wfGIsPga
z+gIlcQQUZkBUFzvwa90P7/DPza6p1/MFhPrJ32mkOd30EMb4zUl2/bn4ST2olZV
fymoT4OQ2NSGNpV+vCK1BehamjoI29mYs2xGcNTmhusR2s3KTYhFe0O3tMgyrqyB
8Xox4VfzlEmkG3xsQ+lfxybWeGG6RNYikqpSVMCYFWCfQzKAD3nmHI/p/L2TgfVI
tKjbrnsBXpWRih7I44M4lVh84FEYTIE8xShcDTbcTMhjo+46uj9jciMyO0H3LYfe
B9OmbW9I5bNq9asXi5Kpd3hu/dmZ/xB6q9UfCGKB3QNg5+tS4PGOgZh0DBM/TRH1
/Bmgly+2N96ov8FdbimNylR0Y76qUSovzD+4yNl5vBUtfxlZZ/AEgH0/HZYtjrqr
WSzIsZXfv2662WVwo5/+DoIt7U8+95V6LT3lVnRc/50RvA5MDUxnsfD7PZ+anOEY
rstc49oKt4t8LsqYPl3nvgY//fa8ELE2FVW0mtPFy5NDm9tvBzTVx6zkEj3a0lxZ
aNgampc0LrvMBYdIncQNYRYATPiRlK7/tZvShaeJbRJfSJVBxHy45VOGDtgoa/K3
zZ23ETDj/jmeIHBb28IuyenOCPJbCL+yv0Av4Xd9ZRxBxyd+5r4OYnOKm9fZX3GE
2CowkHfAuO8MW86MVeaXiJ2sJOYFF8Hup6FLjziTtsGg69Vv+ATOwXmmfKaetVTy
SQPI6hgaXs2aMDVMB2eD/Ggzk/RFTNM7MskXNFpwnwdwZhYZtmj+m+eJ56WlskJB
w+1EYv83ZOLtXVn8HU52ske7HQwHHtAsYL9tpfxJ7AVmjmiWba9ilpGyCxuiIbSE
L+/E1lnFx/H3ROcUzvw3lDEAHiSFyLJmmHS9uS2qGWd78u1eWa37IC2poG46vUUR
ToFBAbQiGb9X9fUW8PnGnDZXReLp/D8mqA95QyUGHoO8rknC8iVSfpBKa2roZNko
00vHOMxjKDhl3puf94TffsbA5oLIq24elXOkUnulU8wS8raNMnRphYZNTg42yEEg
xLkPg1tV19GkHjyX5Y0jM1xQrBhO6bDLfG7qeTDQwgRXznyL5+udl2+T2F+iiahF
pFEQ9QkDRXlwuutB9cIwNTeAfOj1RXfa2oBcobqM8M3fB7lHzZ88jjTeCkvu9GCo
N5dBd0dprNiJE8SJGA8v9nPe2fIJPRuASDbmRi0a3VbO5CFI8UFDJmSeN3Vv9C9O
rYisoeT6qNsfs0zirzfQpx+D/DSZmQik0QBnRFre6hSrRuI8VCy/RE/+KnNZ3JXV
leP6xz3VDw+TfpC6hWF37FSZUT+0FvrqI9+0S8Kpq029NJ+hZ+eyAlojHx+yZ1qd
7x2PTB1bPiM2tfz5donUW9aN6+Mvsty0dxf1dr75dVAn95gQlWUPFeqxzwuzGJrE
UdQcGZyxuwYYXSm/CtFBwXO8XNhyZbXhDN0/s9R6Kh0sDfGS5Jy0HfoYSvXwCgk5
bNV1GFjs9AiRNoQRZW8MjYuHRHA+vHIg/P2kuhjLgt2/NA0VJ8HGC2e60/lkKE95
vF1B2IZZ50c0xvEfnTun3fSDgTWanT7Vxl0I/ufKfJVqrlseANzD+ETfr+DuhFSa
s0tV9GrVbK/9U+UIaFmgEvxNroEhXmjp4nWTkRb+SnSjYYZnzBdW9pjmeOdJJnya
xE4BS54Fc+RzDbvtpreJ8+GRMtEi0tHvRsBfn1JsL+rurNuk4hMYw+MphRPdRIAk
ZGnrDoPRZTlJrN/aSBcspZbz7VqVGrDZDTG6y4CCtToHAq3Nc4DTfkNO+WLbePnR
SmWozEdrJ35E4xt6Klj1GzE5JA2ScMe+nePT35Pe894nHHjTG79rUPnJtZYCqPbm
hX4L+MW8A+6x4ZkYAjbroAsml09JP/E5M0WQNvlqHCBc/1t2sWx07vK2RJqy1eYJ
Seqempu70PRZLjX7Xf4F2ynvS+kExWhnFkd+U8a902pNAUHDRmNc/Vmvkz+YFOi3
dpujJiPeJrjkOG96zrKy0QTwJvJF2shXqgUrso/Dv/Qo1t+Y81e+Wbi6FVdRSvy+
mFtSYSMxHomEWr2ugDM3lXN4PRsJvjvYpg5sfDFxwPbGoQHcNJjFqxqRVkqkjZyF
eeSGwJzvY0f3ozkkbXLr+2yw8I374cD+wlaCJn2OoRCX+ElKv/FSyP8+3vjREvju
XWZN8CJl/x7vfzr/rVU+1dpOK0IzzY9QlGYGdgPhSNjICJkmvoOubEOMuKo/cBqz
/fXDx7+wUHsm7z99ixiLpjgShU/i/yjKD+J2D/DWwZuAnjej/nTgBCri07nTvurt
tJjsybImPH78YRARHGWRbdvrBF6HxXtMjUkGdD6SD2CqwQe4qubqStTsLosJW5MD
q8OD782NwJifXy9TQz/O6JjWxqZoXSbM0tWuSwbzT9JVJOGdXoWO5n8wKY6OLgCh
CDSMNHbwLS/YF9WubzIesmgZcP8Lm0cBr991Etvs7iHsbKjTgMTp+sQy2oEjbSeg
4QJAoB0TXhfmvEJjXF2nCCMo9FznL/aARA0s1aoBz2fQ3U/Nsv9FHeDNCkK4svm0
ltZxcuaLFl/WZuj+a0nxNdPGMgt1kZnDtlSaZkANwK5ybVPdNf3uCvUyBtLWPFPf
OToe9eoGWUajw/Dnw0OY5L+oTi6VpzQXBuXD0UzeCFfGyKb4gf4+ufH1R8/aEnt0
d1+9geYzJ7C700h+2ETLAzJx+iw6bKpKnS78lBDChW5I1FVeFiZ5nV0L3xJtNZcZ
l9zLgLSLU6VwAY7cDgAiS3Tce3y3DUFjs092P8SIOw8wEvt/srnSZNYB4sYffkQA
hFdCRqFgBgwFLLz7V2pSxyLcJCbPHAcj9vtlcVtACuABjN6F7XEzDnMQEAsKUf6/
CdTT7ow4I7oxOP1Dfz4LfR8ggZ8gLKqtJw+so+iHnxQJgdQFxxXoP2iFPo7lNz0m
oGqKw1m5IDaxKLe1kMh4VNILPn5Sm89nFbgnPsVF2nzHJ/tLGBgJ41O4Xic1W3lO
gcWhtne6UT1JLNUqZ5Ebng3gR/8ymdfS7DlPxDzEzz6IH8Knh4WZTYfSr1jhxHim
uRp/EkwJpp4F6UFm6WPxXjC5rDym7m9tCl4YQnFCfiRlvOWxhZRq3SE4wPOE55fB
YEtReBVu77m4pBuF6HuWzq6mnNqJUKebHw532BU8j/D0BUeoA7PpBPpyCgqSrwjy
y7GHjKnE9ednTj5m7eL2LNNKIrSRA5Xh4O1lc1/pwrSYfEmubjRafdZbyqt3KB9v
S2Kyto8UafDuMdvpFqmZSZ1YTEtqIjKDsNJbSGoMh7lRZOABvTkOr3+Ojytu85Be
aazwYwV/Cko+dhiDcG9jN2t6KXxo1SX6+XC5dpO53cDq7J0rwn9pArtaSmoFrG+T
YwHJzIr0ne8v9AXNEI6wRBSfrnyarMJ9GlsJwxP0GQL5NzposTjnRzf8MP5z7nfO
taTp7sGnNMV6jbKPBDV8tFPewZeI5d0MKlOWOWzMKIyWbREnxs9zUZXqUjG/t3//
gkgI6ACja6/nWcVwyH6Xt4BwIhg6LL7zeAiwRYB8mYV7wSdSsAHPdn+m+NRzQtTK
glBfbZB8MvoP0cnIN99acIWp1DNeWf/EV9a+MdbMkySjZ8m6Luy2+qaeA46+iu7+
ZMZkpEvN4YAprwdVtHZgvIBOyHdG7+Ek1la8F//ql5or3h9TPZvQMEDJ36K/41iI
/SqXvRSMRTA93GXVXssMpK3KOfiKXU2ab5HX8lHwYV++8TtAG55fpJT9Bo05Kggj
1ESB3f1xvqxLbFfQkIMK2RWojKNkSW040DJCdKUODIm5RiPEmDOjCsXBCv9yCkRz
/R+W6QTqBXVLjRfO9ijmTiAOq7NhQOXNNQoznZrsEphwAEETW7T1tkDLcboOENii
QXaSAtlJz7x/DmrHBCB1ofUHqq4nz0T3OIEWnpz0Mee2ewmtQQAyCfrWQRAl6kRa
qRkNClqeRMroH18zc1t08YZIZd9WazlFMdN7sI3Zptz4NcpPnDthxBpyYTWdcbq9
CGYXpth39EPNaOZ8pbmvbM+Dz5tmFs+F4dlLbNUHR1MYz9UQ3taW+xi4f2OAm5rG
bJft1yquHY7wmL9/G9qhclOZhzC1/4ET/TYUuBVZfT1bfwadkTL612xZhthbFiqx
yuqJNzGylXo8pozQWsLiKq1+PMG3LFBvkT8pl7eat02qRXkmCg1f+YMHLMnAgA2i
lib6gsvwFreSuRGrrXAUyuf7KgNs+6wqqShQp38etk0L9d6vNwMwZ9mmHyW98rB7
Y8F6jFOtVKKjGH3jSfWvqRClcWDWgxMXUs5JCvuia6mzGEToQl8P/rgLyGXa9VCA
bveOOe+UuWcjDWWXYLCyM0Z1DR4ZkQ8uPVH6KJ1ZbDzi6xBddqHl//gGZwCfwNfk
8tuNwPUYsWj1E1Tl77YgxaiOSfgFqvyyRLxLXlwekAy4XXvLHovYTUgd69oPBrvy
n95+S/NIigCp7EDh2RfUJu6TdFzyy5pAjG83i6MKGaYpzUu09vMa+ySM9qiKMJZt
BAN+ECRhlSgCyWwxVOxxEESoW9Gbl5k6yUVsDgg9RhQUz3ATb6/icqNctkXr3M04
xRAhXSnuGQsS1CGgAqBtqW7+A6d0OD5eBE0h68sLjqKba11rfUBiC2qXpqB6q2Tb
/SjihogFkAXH9Ri6D4ZG6v39LVz3qzThmpZLUf1plo1DZ+iLPUNVYeIfMXNMC/gl
32M1TxlnYwsuswGNzqsMcgItJbZLGxzX/vyXUTDUFWbHE4Edq285ubXtJ3HksfsW
WXgsZptGU8zPxIhaApEcpd/olN+mT4KfveAIFMHCuyQS43gtsOrg9sMkgXL8c4l9
1ik6uXXROYd6adcXmxRoe85pSEHhW1JfqrwjqeIxqGvfzC9rR/rlsw4HTkGc3Eid
90QPD1qgcRwNr0Oox0c2z0CQ4TLnPLuvm+Bp5I2+mQVM1SabpB7E3nJWjX4ouyXU
R5179CSheyNYdMpB9yqpe4JjT+zYiXDacJe2Cz2a1yKn606hrscGk7FXowFMc8eY
jmllXje/m4VeQMvIpLyNLkEiKnsqFNqoUO5X0mBFPZfAhgrZEoOv8OdprsircM7w
LiTOl/y4SCmErk3/ROQ/Tuq2GX+EVT2l3HqmSB9G7yzNvogVJJGS5yhqa0PoSt7H
e1tvMMRxlMpa//0DEQiMuHe9BDDv33c8bUMaWhG4sJZijAqPz1e1BULijTlFcyjw
6VdTjy6jUaps96GuVFBsGaVeJC2K3LE8TjXbK083dOlqZlBglPYyS3m6FMVG+izg
a/YvhykNLTEfX1G2Np4waEjCY2C45UhVtYm+F6nJqpAWU3GsPnGqPEHMcTgha0yQ
DyYrbjCnzaxMWHwDL7kKejC6F9IU4ppUKkKkLcLYaujBcNMXK8vMFGln8e2/05lH
VyiIpJTTO1vUNOLQW4eIFLT9FWVZaM6iLreXq+ox/005uPP3ilQGbOrgjZNd3DUC
n1B5Gxp0sZ9AwKcUCI5+xS6KahEiyCbD2PSJkrkm6KBksqb89+UWZzLcLv2g5TDp
5t1OWLp37nk9E/c08dPkrfMZP6StUnRp0hXF9XzMzQFz2ONBYXc0JGdw0QThCtdv
/IFTe5fhYQR0pmfILPjtnUiWAMq+hEajX1NfCtTNK9gmory2n1nS4lCk2FPlIjqy
X3SNVVFHCh/qWcmkBv7T5LYMnSuPx0eh2T4DJxTxNGms2TJKiM5nmHrO94yyRJC8
f2CbsuEFZpt60HJT7ckwrEI498Xr5RUIoD3a9wbpjL1Hg0FIJeSsip38563+d/qx
zUlb9JlWNhNGOjg/xE6+7kF2f0EiTcRJ0lVFJ4+yFXX/UJq/tkrWg1pweMst20xT
L0VXothbBmKpLGu8En9mfZzGQeeZUVvEtzm2gD46+gtTGQNdsCuDXlVBlYEunaRw
L5JBPTnsBI+KKWWMS0lXc+LnyjpTuXOsmp9R+I8JWxBxdYy6z4hD5DhZVNPmmEGt
SPF7yVCZVzHTmxhSXl2fj8TC5MPRLeFOQC5eB08AvFXv//vrLDKUP9iYoaaLmvg4
DUsHMCEHVQemezby3VqwWaR1JxhKO9mMoacK+zS1ectxtzVkxCd+pw15FK79YG1s
XA5AZAiVrFKjcPlaB55s9wZ5XAJAkTsUHU+YZNhRZSdjmkhvUSIPPWrfO8x20HE6
DDfOZdgzied506OVgLBcNOw54la7YW93WPk3eopUFQEELjXBwo68s49rDAeKKnNO
gjSP7HyyT3xA++wjQOp6OTbcemz4guHe9MhQ/BR6Wx+z1mWZqbFbeMZdKW40z1wX
zCtJR0nou6wv3Fd8nGkXJ11BlLKP2Epqrud+Vwdj1TCZTsKjpKGn9PzEqPCB3wdv
q3oGlxl/Vh6W//8cPCEK0Cd0Xk0I8piVEaYpzWuHznGleUiOcttYRK27L+LHbbMf
eAc8EAQPODgENc+OR26jeny3Y1RKhyOnI2t41DLid3I2UM/1/aofFpsAUYaUTMtX
NbtyayLcDNkUfvQu/mxxITHj+YGFgDf26oewcbR64VK6JCZT/TTZccey/6r+5k71
ecxkMOSF+hZh5MOgf4XGoIHQnZx82N3RCYrdaSOVajbfk3vicTCZSmn0NYdnN5Tl
KKs/GyLCwT06r7sYMk4B0qo3qqVT/KGhAIBEE4xn31u+lNmRF8WaMx1y0tEiVRnZ
tBj68oV3TQ84pHQmpL4LZCg377m08O2NSu8Xqx+m3011RInwY7X2/dnfzApmgefU
Q3j997UcG18ZK6/lhw7QAkDIutPNw09/XqMZdkOS46o6jhe5J32px9jNiW2N50iK
ZgTMjpHNDZ9rkSQkRBKmWgVs0waoHmbuTmXT1uLowLwU84ZtkY4L2oq1heywC7MJ
yTqivyXS63pEBvvjdDoh7VflB83ekPk6zqKUDFrG7YMV00yCBUVVejTfsv+q5qjR
/4Mxd1/5mq26AH77PH0s9NDp5vP6gwT1LqC3bgJx7C6Nd1C+EFdZSvfakoVRgBC1
w4zWJ3CWG4E8PfXXnbS6aUCR04AtVdu9r69vt9nVW79c+1YfROE8K9G50r18P9nD
DZ/6daxYjsZsgPQ25+zLUXPlhtkN6g+TG07V+6k0rYtfRvHBmKyTXno4RXxwXp6Y
Zln8Q2QyqrgirRkNYLIhmSnxOFRl6NBFz4n11wfGZEhzRUBGlBHUzZEKKxBwt6pu
mURrw8NXraRCiiPZJ5eyxuTCHYMpeotWeW+9SikYWy3Jb7opksJUoDAxlNz7KQXu
CY6LfV+CfziSW8AsAtd4iLTxbElILI4NY9Lrx76fmDFHuKO7krZZ3cW4BFWRpZDb
PfwTKLv8otfEQ5R3y8Si5nVO9k4m95Ynr+8KqfqHC7zB/Q0pVhqzFpDwLSZ8ifvN
vtM4eo8CRwKt58D2Da1D7eg3ySewB3j2osj21U7523uDJ5KejrCvt4tuDGNP0c8W
x+buxRcJySHE44aMv0MPpcwlVzgrzUbSPdaKoq5cSru/uqRoTWXgkoFc4tB4IWRQ
FMyf3ZYkxCI4J9bJvsMJuGbonxaaWmKROYuL1HplRDLi0F9rG+11eIc/3Q1scsQH
ARl8Gh0nI2QkThVUK2e0auWyNm5EEYc3IG1ePTX7+qETh8LOCQjDRJnzqVy1K9f0
0xJr4jjhM6AXjLCZvLJrxpfMwgFUdXk6lsAI10GYvin20+RHVrIYSwOyENRz53D1
nxMfVX4MSon68K49EtNXwZkxn2dB1+xkg6DrSw5C2DwT8eZ0WyX3+1Oe08Fu8wFJ
wOnKCR/TstCmssqZoymJN/hJSkPHwIZsYRn0MItqMpeyiATgzG1RnDydYR8LcIPh
Z8hQ88KfSei1aTBI0mvQGzukVU4r0igngjRIKrNBD+JtxgLSBuBkTEmI0rb5B+Js
zNlgPxrvf1z3LnWRFw1cCUZ2R20R8O8ZU73eidtVhgtQMCbIxnDNDBzMYn//h5l3
C6fvMTKRxxZFQiDvz5ABOi6k5RSqhK21M5w3GdUwghsY+Rf+S0IbH1l1U02hft06
9MKgnPdPUwEnnt8JSTiYmeg6fcEnxSdYeTTcBAufp2cHFupWn3Iv8NA0XdEf/A23
Z5aUWRs2V9zbzPVhGQHg+dKBZRFlkn/x465NbWSRe2vr1qAH4otUa7fm/OeIBD3G
IDuWPOtiSYAdKf7GBDO0mIkkVzrQ4LCxHB2dH7QfBQDWO/+uaKANSIuXqJcy0f9h
kvBlXEiQWOQ2nyMWtg6jUuc24jsYg8w/cUKE/N8aAE9HYLMif3afP+jWaVv/A+PE
IXI4WBiNNtDp4MPdzZEOsuyXn73MKchqIcvqMSLrNs5DY0wXFCHcMd3JvWTLImOW
xDaXEs+7d5PV2k8DIjwJyS0w0akQkV00fygoRFhCQa4V3/eQsjl/6a216bb1P4tV
nPm7TyYrIi6FfQvgyTmMRMFhaPz0vp6aSrD3FXvvR59pyApCj5AQ8yFm55rl1dxL
jZ1Fo8GOYpr+DWLVtR1T2OxllO7Iw2T4xk0PwXoHnS6/KMkBxZcRJdnaRjB9YQWD
c4XSeY0Xfbhjx/C7R3YhVvfsm2Y/pLR5kUBe9Q4ra8iI+pJ/QMPVYNEp/KEuU7Tg
Ccj6XUNnvH4Myt3ThqqhAWdjRTjuL3xYz1bmuMo3MkqYYZRo5XhV5QE4wOdumoYN
HIUYDYzUAx2JawmTL3WhRHbSeGe7mx1pbIV4pPudQ5jqxbS53B1NnuiuhzWFACn+
ZMcq23MhhWU0WndC/kOJrU+80JKd3qWxO/kpgARQfodmIXQMrp5l0S7LpEoQNVbJ
z0o5QSn8C4Tc9ga3/ZOkYLB4vxAM1xHOMP0IHYqiWK8AcC3RK4CasFjhB09nZdgI
fSot71PgX/YWJLiKKCrYZ09Xl3UIzXbcYyC+Ty4NqL8WYtqtYr6Okmu9+j/DRtt9
MQ9xLUECt2Zar1tgNbp+POTxV/jsv3LKhjs4z77OUkJPTSUj6HSmzCdq3RC36aw7
pawsohymFNJHM6aXrQlkbfVJf6F5jLAH1fCoKJUVsRWaCdREA0ilgJiRTw2bWuih
yQDFrR40xFAcyISGG3fXE0a2ohApUMP79NHdOOf170wx72riIO+ePQOZv8xmdyE4
S6mXg2CcDjlm5XRSrBCmiNSP1O6jXx/Fm2r7NuqjO746+f8p4VRuWzZ1TVufU5g3
HgwaR/Dxmotl9LOpCvuhW4LU8RxR8Jag0lc1G1kD3tsM3ntYRQWDfX5jSl4CQiFb
Dc4I9nVMR0m9tFE+sfMFmfzyUB4iSgMbiGaamLUpQe9U7kVkXyk22+5FTydboywT
tZW3EZzcnG/VT3Thd/sa4SdgiKPLmlEqrGj94KkDXZbmldKporKh0BA/TxQEn8LT
rg0ONRNpLrjZAx6nz7R0EZm1B087sC2sd3hQZauGVxRZybz5o9Uzcat16AFsb9/v
XfHr4yamE65R5OZBbpeZ6ZYq/4seiDjzXBUh3KnVQJjcpxbsPGLNTA21P7YHzGAy
qwLuC7XWG1OhW1fW+MLGYkZIaaVcWpeVmC0lDXG6WA9wlXAPbAq0SEhDyYhGz26a
FgPrhZedr1IaDVKsbXtvhCCiOiz9qaTQfKnkKOAGuYU07DZqLWzZPcr7Q726PVzi
3jkCq3PDWaZtk3r5l+DHhtjowJy/Xltz/0Ui93d226iY4nn2TW0wsQ9KHPUl48g2
X2z2nzvXOrbDIWlqw6GUWn32h1VUQB3x2sxmzrhDQ+70NGj2UtCQx7FJRp6jLZly
0o1WoXm6Aet5jqwDDgIxi6FjVruyjomIV2Xd6f5CIUs8lTsoaH/j1CUSs+54fR6u
YprhxPERe8J5ZTrbrRHq6vFsdPxGp5OrQLdOXQRXxiU19nbo+4xf0RSIAPyt8MLs
QrllHmz/2thCgi8SopG9kg6pgmU91UoIn9ID+zJz/TAavPRlG6dFBuFW68G9Nscx
tQtTlXjzGjMUQbluUoLzLhxqBa8ftv6mhMrp2Q4tJF0JVOUg6v7RlcQcrWHZ7B84
xXYDd4oBMJ/qt9X8zfp7bAgXMapoxSVpiCnFSW/uB9FlBHu3hecUJNEw9zlqpLY9
CMoUSV3I/nZKxI5mdmKx46YP5XyMvgNtUXCqgDpJIWbRtJldAUl7W/H+qabxqqyG
0tdfGxJHGdd/5OauZBiwh6x6yuh2JqQrzmXjVyQbkGunI1mNujEnjIIUTJIfqq9Z
52NdoXypdkqnFKhXsPtrAjgf7D044Fock/U+0Bxz9NQnNmD1UEggHjITQKe6CLah
LamjQwD6GqBxT3C3dSLjVsJmt9Pb3RGbMpXa8GKIz/E9SzsChPb2t5IOM2l2aONQ
IUraQM9VAnFfxzc8fO4NQRSe+mRO7nXNMQ1dNKZL8C3X8XKztmhKl9C/1cV3H7ZA
DotBD6kyxiXvAaouGS5/y8SAjWoTNPQryIkx5SEZoVZSrSPpvwpLG7zRUTUXs7j5
+OgpUwWP9uc01A1c5PxV2w9E5gqSsLWQPu01nRv6d++1pxURPQOfDIWw27QL7hi8
zNch3X5LRiNF3J1Qe7hXO3Yt2Aq54e1hYzh2LTfsFSo/zpO7RifPOzz3qAfPkzDH
3qHljtSmoAe5m7lkFy9VvtYkfELqZ/9c+CkqYrzXGl44OQuw1KybKuga206Ki2eL
jTAfRDwXm5wJ4cT1MNPx6wRO7+nNp9YSf3aVDF3WFJZ6Jvl6w8UtLr/kl9C50dKw
0OCLuIfx50W/DxTSdN8Y0kpBbNoQY7KxP8VwcE/JVfGDATDomDCMSA8Sv1eZZsnl
Yynldr4rBEacSX0mmw6ohemGAjR2DAVT6hsLBxIvQqakG0H1VrzYD2XAwvYRDyv2
1R7NC810kgCT9iLg9sK0ZJ6jZEfgUO3bsveiz9SvaNYvwmMLXH8KeAzttXft0M1G
Imcx+2xCn59E5zevPAgbx7mPvc6ZQfbDDHvIpYcj4S9UzWUq4qZAkhlUVIrdJHV+
R9iUODLe3v6hZ11EkOVVjD5VO8Bj7xyLsBo8U75SoFO0NF0dYCrS8EqfuzuhOWAL
Sip1JyLesio14qNCtw20ooczX37S1CCjeLfwoH2gTUhJU+d5lxD6usMlATrYWJE9
mpZGQ0u619O/Nc25AFmX15Vj3GteoCddB1l0lZSMbN4N+3RV9RNoudBw+3w/qhC1
Mbe+slBR2oQXRpX3mzDYsxllQIe5MN7o6Q94U6VrVA9vrA3+vfbT//V3Vw5Qwgno
cw56yvK/BfigbaUPoPbI6WMwpWxdV2q/GT2cUD7IRt5vQR00heG5qbLEfrrZRZQI
QbnqybUqc0aJ4sRHF1gC8bVGLBnFKWFWknhHe5AHqg2Gq9I7AYnRVl4ELpeQ6fny
fbeDPaCF+gIKmkXWJA6C4b7TcoyaiH36AJrXRA5ZMMigHyI8DPfBGRddDNpbcCx0
YPz+qBEu2Pchpr3jpi8KcsuRoRC6ie6l9Fezev7l6pxfEO2k9sKuMd21pf12BAyC
gfoQwDfi3k5PW9Y7i78UQOzzxY3CkFGwJiIDcdIvw2Zfbg/TWGS9TW9S6qm1nh+b
XEIw7bdCnOTfwsSNKQFUnxsXc/ad/d7Hpcod8pU2BnhHkASs3n7VwiWDwQZsZ0PI
H6P3SagppS1KJMDG8ViNJ1PIaLHCAxNRYEtJr1QhD8q990g0F5RbLqRCMWJmPwwz
w7AZoEZKHb74swGIugZCncXJFIoEmB1k2VPMmczlgOxOqcguTFgxuFrFoXXTNGKi
KwgfdZ/j9UByxtRSKiJpVcY98n+LoCBRssMut5NqsnAFXYZ3/VUse4j1Y8sysXIN
waGhVDf+BuOG1P+vndduTcHgyXWLjsOVMceakr5LJe68TMwXxc6N+JeOwPWrkVWs
KyCzy/3UzI6SRBrfym2FG1kkYO7bxJFyhLqktRwv/Ta4H9yvhCJWmAduc2wfguLp
OyxA7/GYRiCfAf7fY2hhczDJHisJ2TWyMjTc6RiJEGuW1wTNfLuISJWYvEBSzI4p
8fPnaOru4sZmZkzIo1ERKiNEQ770v4aLLJS+uHyPD4q2vLIKFT7BToIYhb/kIUIO
M11+w5JKVyCAcYuMF3V7ie0A/Mi+VBChH4RRbawz7pMP7+QjzWO/HDf0FqbAcqCV
pc25o+yu47pUpwQCGHQok4dbvxsu0Yj2aPrD2qJaJASsR+hBQqBenqtFeYlHso4S
Un5UfUAok7xETzvfXfhtRFkngy9VjLaGHBNTHI+XWY4tz0vJl1CyXvvEbkHdI8im
qnNNap+h8ntWjSdgrwXLmJ+iQAOdRyhk13G1zY2OsCz8oSplXR4Ng8X2IwVRGQml
wXD5qWkgX8FNarn0GtcwH45Uvc2pVd2Kt6Csu/qf3HxUiNmUg/C35jYDdoHMgzLA
CaUgFgLRomV3TkV5RqQX0MsPHAyZaFr7tzgRwPsxVJPLpdOp+1SB2/smvIuhylR+
5zIhxANjDUY0SoAygTf94+BQ6LoM4SrMauZ45SZP5kdKe0hrYwL7H4vtBUuuJRAp
ljJzsQjztwahRi8fzmowGdIOU1m3RsgyzQzn/PnVeSMTISEqPab+0zNXLMbpntu2
v80DdF9mUsVLMmlr50hDJUYg8yKfizNOsTbs66qlcy2PGF8Da6sAQARasU5Txsix
uTvHMrlN3pzSvXQ5h+Ahv/61kGuOvc0pn2EGO0Ee24Qr1vqKpZxfVb9JrpN2h2vo
ie+6zT/VRhk6QTHzYhxWfQEi1XT6CS9vPWZN7IakbUZHIuR6fa+6KBgcwL9N4a26
eY6wW2GPes7YfPIngr7LXmaOgY9pSRBygw9Ub+G9LZ+iHwyGW1vVy2faBru/e8vd
clzTF5aEM9Iy+Cry+CIsaTKiZeJVy7I3M0Qb2kipmQkfS2Z/fMS0qiNdhvf1MywJ
iCdlmH6e/MeD98WPyim4KM1cBNmaI8ph4EdPIYqLK80/I/zhVbeLNK+dxAYCFhvM
9giPfXKIv1ONE2SkOlThzKr2RoF3V7Ag/YkSArDLpya+gDPZCYkGV2jrEKAz75vg
DjGgOYdzFWBYkzjX/fC3yZr87yWycUEFX1CLOGafnjA6RZv+Tzy1D3ZMYgpHeiER
Rjr46g+kSnTVFVu/Pky3Ojl2WykjvbadgxxWlsy+fa1bJxrgncV2/tpo8jg2jxOr
ifMO0MDFF52i3bvfv9BheZhYopFNJjHPYldhtK6hPsY53XtiTSfGYFtjVYIR2Utq
/WCLZa/iOZNoaI4AkP9WL11EDURWZKSTQSMeS6ODbnZx0SDcZ2h0E021HiXPWR+I
o8SoNPKa0mP+U2eWGXezBMFEGnxhWGjVpE9G/Dk7sNT8nK2fNmS12y6j7iAkCDYP
AbW670UNWluQGhUPPEwaIhiLB+EosmOxG7eVJ7XzfL5gv9oUDEijFrmHWHMLJBLi
A5/qjXobWrGWPKZrGFjOD7D/ezGgSPm109an0MZ7P7ibSnifvdo8PXjXaPnD9g4e
Oy9YYPfhwgEBT+tVHfyE9Vx5N6V45vNloRPQwNkZKOxiyt/zpPePhiM5UTPksA2k
wBBmOXRwqIThX1aOKGHUOFDyYFOeXjcd03nTbl4mPasKYmgHbUImzMPlTTceZF+S
LDkUfWzTuUB8Rrm4m8QiEv+hu7pZaW/f1zzNnisxe5pmA7DDeAxq/JFVZvxxuWm8
pKCNU9UzTKcBHmipZjHpTPRZeQhpIXhvcfWsIzxvUjlPMMISC5nFNCfyUcpeqvLV
p3Xv/BXPKtpBXQ4imVIbtv9h9DKBPreYZZaaArMzDKkhHf4wPdnMb5pFP0oNOg9Z
HJN7CgSUw3+51bVjKmceA9Kr52RqF5VWW/kQJR3seYf88eVw5T9kB3qrolHABm5F
IQcO1qigqOPTwYBE7QUiyogny/RW1yPRVIQypARmTDeLv2xVtD6Fq/C7X+v/TWr3
tndUIbt0wZhNYGUNGtptAA6n/OH80zzPCwFLh4IPXRMVuBKyuFNyrFVPVYGPghN0
XZf4r64AHoOtw5hYJJll2C9VkEqsrkizMIJN5M1sx39tQcDskvQQBMGnnvRo29O3
+8N2pAwKgPpdHLxCOwGXd8vDkjF9hpoklr6bNVZPAtotMsMNDRClhGj8pn2uKyTl
aHYNzxzb3wspvrWPe7gj9AU7xDDIMHEZ8C4tTE/3hzMkzUK+ZrqTq/K/4bYnMMZT
BihDTgB2tQ9wryl5NOxPBiuCXZ00dDdjhkfvFCvaqjGuAPngKLW8Q8AugXrQgrT8
pSOD/PCD3bcNE6jmgqMsm3Cy56cg4AXZbyLRvrseh1ifvxi27B1A7LLlsXCx4/Zw
cz4GL8htwKBYYoE412/YQivxzfbgfzbHOCuGZYd2K2ObUGRRm+bvg8OhknRplorv
8zDTf7n2yVMziDoFUe6Fm/ETvCxB2xBJS98sq/J48p+wFp8SNJ30cO59tYlmQ7Wh
INnE46umzL0yXXl7nkqS6exQdKJc0ns2hidZMRI0XBe5BoUb0A9TCxIWhd0bT78F
Uf9qDP7Z/9ISrRm/KoytpZZ+YlLpHKSxzXDfR/hv6x6FiImadwmAwNpKwH969uvD
bWNVYWhd133YZzeA1YyFFjKgEh6eEiUfdsYBUtsOlGIUYjQTfqH6Iu+zDC49ARkz
0FW+pL55kYpAwXypZ6HRBu7qkj9CYxym+0McJq24XxUtBxkHm0i3OrbApfsZW7hV
WIs1YdllCo0QaEGeqHzwpQk+sZ7Mk/vxxshr/XBG7zGcwNHXScC9HrJjsYoi/c5D
IYiqJT9mO6tgVQrOdfp9DkMF1IL4WLCPRPJQboy3YvvqB98gMr+Z4dV0koxvDupM
Gjp2fUSVnBT0RdJ+DMmL/JxliPaJ5Un8jBkKsxfsJ35IRzKHcgw9R1tCYvCz1MGG
6siYw6XePED7HVoVXXb7FY5SzUZUoa1hJmKgT2a5WwKtTfeyaFQL73ENE7zhJQ+K
i9WLx2SFQhWmM4BVmeVpCFTmMjMsepJ2f4oUWqkQ+BQjF3qaqpKsUVJ8Mg36Ixp8
/b2yc5hgmmsGKYAhPg7Ve0gYeAiobsqVo1BtHw+xg9id4R6KOUSYgcMOLz7FD//X
7szevjP5NJKBCx553paOj4sCAzRngCnEIf+zXSda4SEqIiSIBeoIMlvOKmexXewW
nkoI4+DuqcmofnZTl+0MIShiWVkFQ62K5m+elhf7YLLz4M9BLtlAse9KsONTaue8
2XneBUX51NCiR/xBNx/sHjt22ck6v34M98wCxyUVeOSFSg2S8SCqKm38+xqAT+Dl
dPe1ZVYGhEk8aSdfkWHP64y9ns3Wz2eliycuOKK0yxLaq/TVk2KfhBdCPG8tzrCi
SPBJi+pm37iixStoVDyf7cXo6+a32jIdJtkHWWa2gz9lyj4DQ5RM+4XiiClYo8u+
lgrsjXjNOThzAhmUawVItFSy8AMwzHukBLxGWmFWWr0sK2Xfxnj2ZwzUP9ny55mX
12LUUaiMDH6BdHElguOoM54tpvbTxZsKFdfd5WnZ8Ogr7EDkPHhdKse6ydkrOKoI
t0NR/uIZ5T3+WtRL81GqOHEMRV4CD4fD/qSPW9dwe+uQR1bnD9T7jmvuUDopSjJZ
SC0uqW1akc5Dg/5IjDh1dFGyazVf5tX4cM3A1btSGabbcgYobf/PB563HNyH4cXL
VOgPF9XXuBjqVgICqZKwoTbIHTux8C9rSFMQGw2139RIPalubwnndGjL15TJFnA2
jl77wf/pvWog/e08sqrowg14SyzQPqyy0cGaqdilXdvMunOBMIWBj9e2m1iZbxT4
OUiH+pGR525cbUtcMOvjviMsK0dLrjrmOxj0Qb6HDIPIGZs3xELP2tCvAkHEbk8a
skvPFrS/yiXJS6FqqVcAzcL+wr6mPUNlw4mQvsRT6Ll0qNAkHEJujGPhRd3mLkT1
61NJJfVpnQqqAJmClGd760/qn1cgbh1PE8zj9QdunFK5ETyE0y0i//bBp0XCVMD1
GheT1irEGJZNCYFaJ9ugk8VFyO91ia5m0rAV9j09gDekFg/9uClZTBEt2zSvgg/T
8pLFcpDD5GfNwrCkupu2X44sn3wUKNyVGMG4dE/rXlbHM4yUUu/FKr+uHb+A2am/
W6XH8fn3HswQdgi9LJrHuEhGHUIFNhMbszxQCYTMXglUFiZqG8CofFFF63K+ztUs
GKAN/qDMfEQgiN7g+00NWZm7KeIcmn0RMMuVfrCIMtgETkQqTQj1gS3u9wWGPfgp
1CUwAbegDnLU5mRAYwpMlyoSxJpKtXSTrB5Kjotl+d/y10W9PV7OXEUu9YooSgl3
kiph7x5Qi8RqV0IwKbtcecArLRRgk/jD3gB93V6j43ZqJbOtCRW0RsEFEjrGZeDp
8sKOayzQ3PHGvhYNM+LibWe9yOnDkdgUZawZfkapzz5nCcYSwzp5tTlslmAXN1tf
vtimpiOPHgKJ7efudWGL3pJw+l/e9xntPXa8XthqRk6W9SZGzycI2C86/goOzkmW
1zAUYmpiArd+okQrH38PwNpnZrMXzOzIpbrm4xZPLZAiXni3aXQqQzNwJTS3B2VH
QFkzPKEHWvXULHtdKqs4mdCV/KjbHxIccK4NGG+thmXYhyhLP9RhX7BmwQP2g3h/
eDSpAlu8qFxYoYZ72SYW+jZWix8uq/021vJbzp7UHZWSh4Kfwdh6rHhd1YZPxDqK
teDTmngNaSwnm7xGi4esfPwCxF5sOLfujHWT2WckCYlYvtJzuU4MicfK7JEUF8UT
aYec5GIRDNSDImwQU3oH5LSgBqlYjrfuemsWg3LPtN8YOPOIzOAz6R0gQ7cNYDsU
w6unSRHZ7UT3DRIKIT1cMyZ6fwM6kTXw3vwoef82viVRlvd72p/t+YXCQGNBFcyO
UPOUvykqkax6MiD36k9kz4Do4coS1KVG3oP9EnWS0NfA6zg/1W20Clrh7Y1BbDNZ
9/FmnnzFsn9maS7jQlyPiWcxrJlxK0sifgvQrwDKNor3YoqVQsg84qaZcKdnheu1
XhH8iwkbtpABD8wC9yDkefZp/C1+npoiA3mNucNhXNwwfHBwETllLsCuLvPecgE+
hBcL8LRX6e4VTgh7kuqocd/5Vgci5jgq2fiZhWwP+76Qjm8Ns0/aXTpLJE+dvEBW
twZiiEn2F2rLl0HYCXYojHklSyHWwh5Dps69T/MTNsfM60qjEKDOhzQ+2Ga5K+ie
62Zgay1D9Qed0oTnEDD1O/eCMFLhEvwNAL9tpzF+xXl2+fh/ehCppsScPz7anyya
ASIAPmpTcZ/EXLVP4W7rSbO368YOgM94kQ4JVwb+BSeizcMNuzkn9RUDN+KUTTcB
BsHHQTNMl53v29QXuFKFhw8fGtqGvckXEtR+sORJxMlrKdB5WwhJ++i/tfkAZY8Z
p/0auKbWR7DGujD+ltIEvFMplR0ywBvywQ9W7YMnHgYxxl8bQh1r0Q6iUqRpeBH1
AyT6NIdO6uvpxwr9FMJ1mioL93OoWnHSbytaSyXrGglQBNo4iN3weL5vYZ+mHqYg
XfC5rRXc0jB1N7BhdsCI5HVUqMAlpj5xKgTsK+MFAIJoIMPIneEG7VfsR9/Lr2FU
PXXt2jfV1CD3awXUg8pgR0WMQ3/VhKyqurQ1sGVFkff/4LfYD/1sY6SawsMVoEdU
YUd+0gfIw3XEHQFvb5vY/i2vZYcepIwCOa63jgPm2O5FlRuahPQ7kAyEQrCiMUzZ
iiZn1hZtmfCTdePHmlVDfqcLpJgWarDX/DLoQ6lRSppXIGngjozUrwzSEF1IPi3k
CgNhwEamrHbd8nVD82LliaoYi66gvoqCUesloQy6//JaEMWWpwWrGy67g915J9JV
FqIUBCHQjoF4e1xSUjPfDxyz9sTeeDR6cRdtyCqSmWjl43I2NHDj9jIo/+7dgZFj
9+BRjdUfnzbPjcsHfVACWC9C4LLy3VZlEoqd2sW+sCYMC9L1X+TYOENeRMkUrHEd
uc2ISAEcMMbeOQ46dGSool2BIiaecQVjdGA23szN8d753u6uMwr2l7TiORJAthx6
pd3K3gWyEuXKHmLdnA9F90f8Bp+gUJ4KIS2Kkp7d4+aDoYoYqnAfzzu8q4HuB6ar
xGuf+tFac30KDgrUAAiPqtD5uP0NYvoVN2wA8fm+cCstTWLYzU20RhnR/Q3BNZZy
aXaPEpXi+/M0mVpcbL4uw1znH+N3exHAxt61u7Ab2Gz5j9YU4tre9bWKeqtVCa3V
HA+EW6EN3cUicSJpU9t5bWlMXFh5nIz+KOm2C/pW916xtILSLBg0ASQ9aPkEs1eQ
bidjHSU1hGwbWJHbnLntabdmZ9rbxsEJhR94DX/2bgA65Uo4OglX2XNDAWu5f9JR
62/z2w0dLdADCZpEKaaI5F1HfAe1mAXEnUa7E55v7Z+829aMIM4eopf2GorhW5Gt
MbIs/ap+o02pUaS3c8t0oXfqA4IkK1ZzKljq5UWj+UMi4QWuUDIGj1sM722MewyB
Jav2tDuYDCMBs3VVQDX3y/tWS+TTGT132pxZQ/dqMOddI9N1bcxhJD2WdTbrE0QE
Mlb8I8x8kE3Bofa3dOGKfHUcc0F/pjFDlCTiQCDRgiKjz3A97cwG6JiaIyGi/wmU
GRFKgOmUbW7525B7H5pm/+mXHY6Aj4mO1ByWRSxaYeAJFirQbgyDIxCZnxYPY6wK
48IcnUnDso+99JYXX/Eec4x2IMCKk7isvoJVdIqkcPN0txULKV4I3Hqq3yOf4tnE
wn+bxKuiOzDYFTTfQx3maR5vJXZjcHDnvrHTZkLFKyuDJ4e0weAHkpWQwap2HIoH
ouV1wqA5onL9VqhPsOx1vX9MYLpC1eKRC8LlouEZpbLQ4WU7VP7gqo184X3Uhkcy
Hy6V1kzin5YrdicRF1U4hDEPJCwQ3W/qq6UvTx2b9Cmo/HKtneVZKjTK1+5Yc47n
QtMIhKu7BML8uFfYwh29D1+dCmV+G1b201osygjF8xxlEnsU3Z1H4YtcTHB2O1b6
PNKJFF+7kL8WVG4/NKX11DXEC/YiIZ2wDP4vgwX1Fgu4ZSSBeIMOkZZFGVhRS0wS
ki56ujstQxbiy+jRGZR6waEgFK0Nk88IDXpx9o3CikusLW+djd+Up/YNtvJcShig
q+4mxzY9/c0woP6UpuGteCgBkM2/AG/vwfG8vMhUUr9PuG5P9+kNKc+saww6hgqu
L3swtFU8x9sRabcz/OmgzWBG9GTSCR3EDIpo5b8dHtD8E6Dn+QfuHsh1U36YPUSm
tBlh3Hy405s2MhapKdbuddEXiIWvzh2wR9+M3VNxjgA7WumTCrNXHKPX6Gg1c1dW
SpPmaTJ6B1KOkybZXK9upQM2k/CIotPIlLA+XTMXwmYuzd7fSV2gvcx6nIkrMM1w
bzqQIOC0EYomB734Jq6I9bu6uDJ9CDPImsqKmg/A81GKDhOLk9j5FbGYpfZqhPkP
l8dRQmGq7rwtDlRY5660c9VbY9p6qkeL1WHUh1BnmMx5hPfZNMEGAS1uF0PLCcLA
4rWZpkDFthNljoyXJ7w7kpvmci2pnWGNbgXVPn3GMHh+xblHUPzjF0XHNQbmc9Ve
BVQk044xZzR+HAjzNK1BHVinktcaFQy/koo3whM/qaguuvlnTeZXrGs7zo434ow4
ouezIJO0IvlvDRgkKEIOrAWQhAK22mo0Iq4f8dZ1aB7m3bUgj/OnVAZSDWblkFGo
IkJwkUTB1DD+GLEZIp+gp7EGPi1sjd/39joqjThsleE0bIa6+LU71tlJ3uEpZ0iz
17mPg6gdTHW4p4lM+M4Ao5SIx8Df1X3OZV+Y25XcvjZhhpZu4YfVciHuar4mHyNZ
C7IHqrfc0X6VyUEw2okU7ggCu3FO60qyb7EQthnGoZpRoX/rGkAPZa3MYhj6Abod
2OnzGc2OSjfr4Zb8CdOQUEPu+Kp6iIDm7DSE7qm5wNz+jMbO74qzUG9Jew3skeYo
nkH+y+F1m3uRtJKBXT79zUwd4r2W2RoBNIY+49zZyEQ51ci0LnZo/F3zwA7kD8ao
VV9Zk4RJV86J1MDrh/M2yxE6pBOgSOHSeqExBDXukpAC1+pn4wi/XL75Ko90ypB9
7OsDDI6sul3ac0rncEi6sPOmcKOfYjv1/ccIYtYprxHaZirZW2zMRyCd/6FovOhj
n9x+18OeigcMC0IM/MG9K4YFKuF41+HLNK48n5ZVddExv/VotrWhSESabQEvG1aH
fyqgJrbJ1TmdxiTFNM2OvWpkmG9pv2ZsqwQwJ10pRhC+3B9D3MB74usbIGsaoKug
DJtn/JlHhqTl6kcTdId+f1Ryf0uvQK7wLBrXLWsSDGdJFzDiKE8iALP1eEoI+L14
honcS2G9zeDbqSv/0Ogdo6ExSPFhQ/nG9phk5Qh00cbxsPV4JWdMBgJ03JnErto9
WL+EnsPpPT9YgAvcejumgsrcuF53wmVznLNZBZSBVpjMEDwFsBE5SDYuXXd+AJU8
74ADk2pj+m9JeBTMjgIwGWc0ECifUJac7Rdjg1Sm5YTpqbq6pqi0dNpQyd9MUtFA
r0xal6oirulqSgQv+AWXADk/ElRct8i5H4r4WIf5Eqo9CoBnxacz7fDDrQ0BCtmz
n8GLqPhQ/2eIteWSY8MmZYkrMIiZzPWFBwk8wn/5QEgyTX61+SXkpJdGdJYzi+ld
aJwcFVovVpdftxHVJS5A7Rs3TIWp9Z38z2GcQbZY19slOlN/8iboDwQHW/qDZ5TY
yEvhRkgmCJ6t7QpBi2bVhUJVVfL8wLjfglCuLL7U+jgilpO3orWgde3Dg5SB8F3M
R3L0OPV+norrRNk3RONyvpUztvA9P03CceWfWpiGITlLGkgkbc0h5fILInCzHUEH
SH1tQ7Ia1RxgV9i6XLhRQHZJQaEfGWOgY6PgRnvBxMb+D+4pWmZ6Zv/IIRtBjQqm
b3/m+NapBOMXayYTyV1LyJtQeMhfd5U9f4i0kXXRh5M2RDOytePZgPp5blSiAauG
FYkb7AsQG+w9EWAG9djKUhFRtiz8fHWliEWKzcgkM5PoElTha/ak1j+Y/JQuD2UC
jjwqexUxvbsDgXLOlFoGEnf/XupwJMzkuz+xzwROB0FE1o6RcMqyBjT9pNEaSh0w
XMe51xDVWR9Pyfo7jSz2jQi80jnF/wOY1UehwZioys9RxLt9OBmpxOYsxfR4p5h7
tY8I9d0a5PZSU4fjESRNsoxkGKy5am/SzZrX7Qdz3/DfhkkUNECWAjfjKBIvTT0Z
qWtKfetQup9eQkOQ/sx/5j6L1hL0FF1WF0RZj8o69ID/jK+ceI/9cu3MiqNTcHd8
8AxhHiW4B0j0LW7ZfSfPWHtD3duBjBxFHRmD0SjpQMMffZ6mUu18+C+hAYL4OpPm
HGqH8WXHnwrjDgLKqkpLfwQz78kgGGdJTTbaRwo9C+bW0/P5KK3k8Shs6sqVXA5t
E/FNkt0fXblG2TxTaDhxyIDFNhiPnRsUYvNAfpNgswK/D9Qdz27UrHZJMP8PWOZp
iGMPatT3SDCL66TJV+Zn0C9VWIzIYW+z557TaP10O54nNbviI7KcjbYe+go0eqiE
v9VZoJpX9F53AO/H4ERv8WUHDM975CEapeg7RZ65Na502Pd1bRBIV+KnbfIueAf8
QQeb00HbES7gZ0Y5HX3E2D35flakYtxC6awaZ6MZq8N6Ex/LV5Cpb09o2Op3OW8M
oXCZTe5MuNv6JDVAq/iTx1gcEe8Iv6jh3M4wgDaBRnkXjdgr/d/Feu2LwS/Z2bBI
+3CYjATCvr1C8B5h5xfiUPUdl3qFixB3MuHxkqEC81fnpWszMgt+2dE6rHl7bqgb
aIG8ksTaPXOIA2jdzI8akDxowNQvCgiG3ahuQ4ppSDaDOD4VSj84giWgV9HQCXB2
yFhyjd3dpCC7TS2ph3ZyUIxziENimzqQy8whvn0gY8lgxIrSxSrJRQKKJBlkRbIZ
Wmdv1WHoPAmHkX8ceGs6qvL7NKTZNryvO0NlketYFvsmxx6MNeqlfF37tzIHGceT
ZcnFSOgtNrQtE1Rx0le7P/Ddc3We+VhM8qyaqvgGfIgFeUtgFgrxCNEWIkT+HUbj
EVOWJfn34MJLGN3iJPWab5UmP1HKZ4WjIXo81TFHga3EU09JqngxUuCtAr3tsVpl
hR2h1mVYagVOp2G2TmBL9fYZqUAc8Qhj/gc1YwqG1DUUNpr4x3/mL9RnaKjQTmlG
UFpNBSM+Nv4B/ACe8YzqYHjecShdIXGutjqKqdLnRmY+XP3rpy/ar5lt1J2xTVC/
bn/SZLwK7TAMtzJ162yxzT3HjaaBR8+txvvrIl4ctIo+hZsL3LKLLuW51XFugNaL
v2D7dnVA2Uc+wNnb2N4j+zD9li1DBH1YAwEmUVWs7b8qRhTZpiX+ohif/tPgGMdq
SM+PDsnljTVNKB0pAgFRg4fyEyopMNtyp2f17ny1efYSp3ZoJ4OxUt69PyvRLvh8
8rNp3f4CGDsWT/v2VOkPpMURsfjXU/KROyDmFjAIjP1FBRWiMkGOLHiOkMmSVNVl
l6VPJ4eTUH5kYvu30G5rBKOSa829M25RN81WJ0yK3zKtLGHwU9un6Nq7yYYWGEL4
d6gTVMB2Bk6oaVcZahhEI3s5OXmZ759QUUYWrwKkKr3gsNEiICtlw+grfaZjXPZg
kYLXQRvu0SQ60mZrJACeUJ6Im0JUyFs6jvrEvOyud2SJfNUI50pXa6Fixz7YrFtF
teub9ehSLm2665X4PQEpb851/QHcNmlp2x65JEi9osQ+HPlmryo18y+Vxj8C5IuZ
3Ee0PQOCinUuZEUOCcZgujsBANKvvPMxYZyP9b84pPTseBxP/N7GS4oh9+Ua/dOI
zJgsR2YB3BYla/v3St43s+WKYCK4eSepRbdwdTAnUwVBpbjbcjiloxtS4jNJURuj
KMQYxK+S2kIP7EVgYK8gxsWlfppRwR6CNI/Cksax0XjQw7PTxDqugRYuSKJ8Krdt
3VxOkhGnh+LtoM1DqXJvNUUboQPBV9iiPP8B3DPCIhvMScFYXZj1lXxgKk3zMCbB
FtfT7jW2P83O2UVQidO14l2qUKRILrf0XLEK1rX1i07vXIRQyR+cQlDd/CU3kyCZ
99VdQLsGz/+2gJERiJ4REy+Ymv8jzPVX1Sr3PLtLapys9qTeqdTzKg6jS1/fD/qQ
y1KelQAYWFZKI9ryRJpMEm6tMI9rHXeS4WSOPTFMTr/2LER+9+eGHSFnzQxeaRGL
BHCuTzU25jUPyPximHhhBsNcRF5fCDRN+wmEDoxiUVIHBjI3kh0RZxsKcn3Ee5m/
iLPkCWj+kPyPz4QArY7J9ecueaNdsZja7UA71p3x45zCbqqd8QE+yrE5kZz7BmUb
u2GgB6aHbhnkGaMLCw7RV9teRqHetH1bDgnAFR86v/6O1KwEaqjvOrPBGtP3jBrJ
ZxG6BoK4dvg6pX8rq3OnuOt7ERMq1OPFxoEMHkYiblYKK0S5/d4L95FZVKl0twyI
SQThJ7W+9GzyGclHs/QooKnZHksDGBoNeuuSUWQRXf4n6cYdOe0UrjPKEsP4sxIX
0jp4cy/F46HBvvws5soahB/dquQZZz3LO6B2Dro+qs5uDj9cP2Y2y835tDmdXg1Y
sGs4IPR/lgJz4HTA7wF2As2gcM93pRqg9+GOR6ym/gzn9e8wwgk317+jmymlhA8X
jO2pDR3Igeh/pyrTi4hvSc2xiJ9LrLXeK7cLYkDGL/CcRqWexiRlcLbiO7B531/s
TJpf9J2hor79cgXFaeI1Pwxjv4Gi7sIIM+TlS0pFtLUBbPLtbmGGoCTNvMh+hy0d
RfrVHBXfnPXQFHOSlfDA+v4vdLc2yKwTV3C0ZDQ+kCeLoEwhvwIEyKPQZBLGdw+u
Cz/nLhleZFs2jgktC0cpDsjhi6Mu6hduTEeJpTGyRPLO1J09R1+2B0T5L/gMsdMG
Vz6uzHBewL4mQ5vuogisgXDRn6WdPBzkTaZjtnciyFJRM7iBaKp9SWPj0NXLjbNx
p2SuMwFW/ALljUDXSYBrOPX3LYJ9MTRE5GP0V2ailSh8j+/sAH4jZJkdDbmDLH5r
GZvriqVfPIwqBaJ40gTH7xLXmAb2f68/LQnclDv2NSTS3/9cPtuTo8A7CcKFeMzT
QbyTRyWMV5oZ1TAMJgryWJKlgKyoFaiGXcQkBcaoa7gt83x94A8SNuGaD6VJpOTa
Lsbl7elsEoi3+9OOUrD/u37pM/MEfdHjfu4nPYJTrg0Ur87AG664sj1Jajlnk6p6
EYgye4kQQ+CV8dnyTUZc6PXpwrsa6cT0/BDUCmYsMsNgHliFo5C3JrsBX/mv1wb5
fOIRQi99q0M0QnhSSkEa6U9ihl9H+Aou5TedQ/XCr1x/iDNoUyu/peyhKCXwck1i
eD/qwlF5rFinkGmJQ3AZbf4deV/QKkcclDPNOPr35Te58qEw+d31zB7H9om9HjUH
B5eARN3i3DvmbV3laAHVYQqZLBt8Mcp6bamjVr2f0FWEE6c63Fg3NPNg0tlDw7BE
Qz6i7lla4czw8BmdPA8BG2qYId1SvFXWq5by62s38zDk6SVyk5Gps+ZDYXCq4Kcl
rdKj1uCxxS4cEACBtLoVm/b3ZlO/eZg7ySDSgjzcm88=
`protect END_PROTECTED