��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q���u��������=]�kN�YO�q}b��9:Mi�h浘	Ü�`�lZ���-��m#:�����sQf{���-����K���B��?����\�pס����V����y�FW����s��(ƾ���g�c��N�ƿ�a`Eo<25ڤ���%u��0i>Y���GZV��eᄉ�׊/ �˝�&>ˊ8O�u` 1=����U������Jn:�3A��9�>b/n�Xl��?)lu��jܐ�y�d��([	 �[|�g��;����Z`���pL����*�vK�gG�[��2?ʿ�i�7~l$��)
�tj}U�r���f�@�S�7)R����o�LX�=��Gx�r&J5��r���/�A4[�d����s���Q�~_���|�Z���OkI��O_��e_�HP�~��ʮ�_�ch-$ׅ�X���B!�E�f�%Ŷ.G���6$��6��;dŅ�~�6'8�,�[��#����'�)���z[N�m���U�f+�����i��'�,@�Q�w.����q܉�.�!�Ó�$���ϰ������^���n���m�UKd�)�a��t���bi��3a\(�G�<m)/b�!���Kl6�2�� ׫Px
�4�F�JL����^"�cMn�Z�C؇?���F�Ioȓ��7�[��h�`aҨF�ʤ�U
�C<�:�'h���������ޖ��+��º[�)�ْ�Ϻ֔<��#@@��-��H�ig�v������P8w,�z���}3�C��1K���N�D.��.#oWJ:�*�ʡա|�n��Ou�4�Y}zbNM�K�Pfy�Pp�����~+��ؐ:����e>U�e�b��LI��Ȑ�d��*u=u��1�c�W����\�(�pz����`�� J�z�B��ps&��A�Թ��p;'�qm/n�V�]����L]�ZM6���T������Տ���=IK��$�7*��3F�|�:@ ��si�3#�e�������;vbZ$�3Һ_��&Ie�Օi
R(�������n��"��iH�+��X��5(��J�O	Nm"���OvA�v
uXG��K�{�	��ؔ�M���N/�#�)㰝����N��}(+VnL�i�����w2�#��|jg��1� �� �~n�v��U��ȸ���Ak��^�\�5��V��E%�@�FU���;aڦҶ��� ڑ���qf/���Vy���������18n*ʯ�yV��j�-���Mr0r�8�k��Y_p����0�wxI���̜W��aR_@��w���X�#ᵡ0~8�A�̉2�������g��`�/,p�dxX�~�8�4$$w%$��n� �v�� 2|ҥ����*��=�I�oL2��K�s�s���SC;�JQɶ�b䐞&K�d�
t�وR�j�V��v4_&ׇ���v2�	���c=��8Y��.^��F��z�~����;U*1�XIZ|S��;}�)έg�+�ł��ׂ_:��N��-��c��@���f{fV(A��M5�\��]��ac�c���
���<b8�`��f(֥��eP�J�eGB���Ãj˺���1� ���d���|���S2S+�|`�en�ڸ�
Ȯ�u��5C��\�#��?q3��z�>Ӂ����u��Na�jK"�#aE�U��1S�X�;��|c�{A��;7@EL�O?h4�	��c􆗇��Ec{�������AʹQM�^V2gS96�E�L���{��LP�v݉V�j5�	�O@=(��z.P�))',����FV��R����(9p'V��.~iF�Ȓ�ư.��M"/I�71���w�������G�IA�A�C�!��2ǥ�J�T�?��%����Z�y~�͙DH�6�s�����3^��e�[�I�0��O l�c�� sSD�e����N�'*�� ����[����I��$Ǫ2快ٲ񏩿��q¯?d �2ꥊ�ڍ�Uܸ��UY�K��v���x]���rq#TL�d���+.���J���{jY�.��o-@��C�-�/�/��2\SP��Ab��oe���O��P5�2�_�fH�O�bWXsxn�M���T�,�w��<?vB��s���u���'�×�ȤO��aY �t��J�v�?v0��J��As{2_v����F�.� _�z�u��_�R���0�m�r�x�OO��si�Q"�u�h\0�s�Ϻ����k-hm/Ԣ�ai:vw�;]7v��I�0̪���/����v��-qσŃ8m|���)��?��qIz�M}9��	}���$Y�Ɛ-,�3ϻ0�,p�����D"��Wl��V��y��!�z���|�:ك��-�����?�#�wHF;�T�y�/�u�dC�����v�G���{?U�����C���ӌ:����64��3��)F
m�!�dH��<:`�,�K#�rS�r��{�i��K�A)�������=���v�F��;SI�9V��,J�'���3q��x.�r1Mk8�4��H8���6Lxr��x�)��Zr ݂0�vP�����G��7BCo�O��5/��^������#��!�t\��/Z S1�-*}����q������}����=�����/���6gP�x�t;��]N��p���\f[��rY�銨>x]a	/F]�k�䀱�s�����;-�He���p�$��@�� b����RU��=`{7���r��}3�?k��eD����>���[� ~�Y���_D����?ͮ(�u&C�v�K���g�M-6_"��(����C@�6ݣ�Z�mn���)��n_��Q\!����xp;��3?�e�	6���yĳ�c���l>a$����f�ᇰ���`�x?M9������2��z�����XD�[VC�+��Vڠ�^6ꊰ��b�� b�֘s��4}�kr���CK�'���xQ���R��H>y@�J���ŭz�U�C���(�8	��ͨ�a�)&���6^nk0f�+GP�h4`c �!����b�ӱS���> ��������[*��k~�����ԙ�v�-3 Q
��$�����ܴ��*9����n��!()��d �$����Mn���.H N����e�[��[����P�$�IE��%�p�&?�?��+D�8�):+����%1~]�s��\����m�u�n�ӂ3%�Xa j�Q���� �⚫�IS�:��:�N���n�=���S�F�<\�w� �4'*�sRPӲ�����lYjx/���`�N�i�[�Ҹf�6v�%)M
CI�����5�G��k�ŬDa�E���	�xuŰ�