��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q���u��������=]�kN�YO�q}b��9:Mi�h浘	Ü�`�lZ���-��m#:�����sQf{���-����K���B��?����\�pס����V����y�FW����s��(ƾ���g�c��N�ƿ�a`Eo<25ڤ���%u��0i>Y���GZV��eᄉ�C�M� ���}���B�ź�Ld����E�sX�����	��l@lR8!�ՋA�>����W0):�e���tw�OKM�2�0���׆������6=�G�.ݫW.[9�Ѓ[Sa2��'n�������҅�J�]�%�{'���]�I����p�N��(�{*s�²w_�&7� 5�}����/����v��#�Mz��v��{b�=�$6�
OQ� �Ș���8�&��y�թ8�,�vy�w��}���H�z� w쬡8u�;&��sVo�.k/��dG�H�n���j���nC�t���:g�ִ��������k.�ZPI�N�H>Ĺ�22_}vn���k�
7�a�-«\���Bs��YF�ior��D� �*�FP�XsRNn��wn�O�#���z#/#��@�R��l�(�2%/};�s3��ܚ�³k��6��h�Z���W�Ɖ`��Ǚ�%��{��yo�h-}�qq����g~��y9ZI�U�Z�n�k�XÄ�@��W�w�x}�{�2�r������q�q���L��ZɆӡ�?(��[�Qytu�����Hfut��&	�L���1 JMu=Ie�nj���5_ 5���|ı�wᅆ�<e�-�޵��gTH��N@>�=��Yت�z(�JB��8}i���TQB�d���J�/�e���q-~P�����������n_}���W����Vs���EB�D���������~��VH�a\�4 g�3������Jb�����Hă�*fTu�ǭ�Ec<�~;to��r{u��	l�T�F�#�����V>��Ҟ�ݐ�,Gk�s� գ�w��)�Z[���%���&��[��k�ܻ=����Q�q.�q����	�(��1��\�� ����-�k+P����x�;�+��T8H�S�ܸ�������,]�(�+�CGDǋ�ݼ���,k�wy!���VTs��K ��_Z��b%�Сq]��.��A������	v�OT5�_Kn?٣��a��c��y�wo��fM�<~�
HFvo���[>�`*����g9�
Ƙ^%�SzC!a8k	��ā�	Y��h��z�x����,��rN����m!��8�-J9��.���U�c."W���	N=9�~���1~�1$2P��r��.�Q �6�+%��'듷sD��MUX�kn��H����q����{�p+@O>˟���7u�0�V]�C��Н�`sv%��R�������&���w;���6�א�����Wİ�9*�"�-z�K`I��h���p<���N����c���(��W'l(��Ѓ,���ɰ��g�Ga�����!g0�u�o(&�4A�&�;aJ�S�LE&�e�T�$��p�������} ѣ�����)�4�k�yH}���G��+�=��3��y�kJ��X|NKE��rro�/C��5?)�`��J"��x�X`On�`Q��˂6�D	K�����1j֤>�X;;V��1K��y=���T�X����jj�@E 7�_�f6L �3���ǽ�,���ؙ3|�-k�0�$��H�9��՘Ec{S�5�۬d����T���P7�32�*Დ�'��7İ�����n��Z91�Y���
�g@5�R6�D�3��i�<:�|AGH���`f�]GQЗ���i����qi�e�%�T�V�fu�~��
�~z�u�L{�ol��T�yJ��z��Y��)��7<1V]-��[���X�{��A�Α��<����Ĵ��ߑ�&l��c��v�*�u�T�V^�j�� Ҍw�R�^K�R�IH9�+��=��;��uK.^(���Yss��7����>/�0���g6m"�.�= �U(Ь�̪5[؃�B��X�G�6��<8�	HOA� WmNbA��v�3f��~X�ʴyLX�,�]���:�#KX�2�?�8ø�����d������w~�45Sp�f-�O�lX��3X@��g�V�{�����������Y�{������}������\l�����CS
׽��n^i-�y�l`�!U�� 6Y��Ζ��X�K������B����]M��33$� Y5���dxrx���d�"���c,�y&#|�����V�l�H�:$��R#��߶�ۊYy0O�@�'�d5��n�Y1*��XK$a3`��LI�����
F�e��������4\l��9��3O_�p3N�ǳ
�6r�]�*���(��Tٿ��b�O�8}��494龜���?6���8��;�k�}�nx��Ȧ�S0[ߧ���m��5���3���6�5�4 kf	B��l�+�HW�� w��g�
J}�[�pS!�R�X��5v��m�y���yVf	�5�C
}��t-�{�X��V���/�����,dU#��-��Z�y�v��Q�N���ab魍���`~7��̝�`�:���'���+��)޽�?�V���6�ý
��Ѓ�Q�Eޛ`�5�a�+؅+�����Q~�hR<�x-�Z�P@C�������1�E�@�1���#V�nw���FQf�ŵ�������f(�0��vd��BΙ�K+=y�ed�?&E=/���DhD	���>$Le"�A�s^Q�p��B���e-bj�X���}=c(�Y6Ju�P����K�e�)B�8���[6ꖤp�ܧ�*���>'�xcL��t��O�cѪ�w�M��In\ ��эi9	����%ɸ���-���-$�"�D�����w��m��<�?��M�5y�����p^R�
3z������:f޽�s�~}t�Y�!K0r�5>��ҋ8�#U�،A�w�`���1I�Q4�WDt(ʗ�mm���t'�#��"����P��C�, {ԛ#��zj@�O50I�'�.����6�C �W���GŁ�
�hl���z�y��]�, ǇvF��QV�+�lĎ#����UW<)؄
�ղx�t��D>>�l[��k2ܮ�z�k��1�+������m�Q��g�ox8E���tP��7�!�E�SR�NUZY?�+������|��e�Ațu�q���;�4��J��n%�iȊg~|���T��A��z�'"�v��b�	M�q�d���H��T�kc������|��X6�82��l������B�4��?��(��e�@����ų�j��m���(�j�Z7��$��=��ui��l�H�1�'ֿ�Y�
����K�{�G���JT|z�I6�u����4la�=m�!ah�U��\�� �r�kX^1	W��T-�м.T�0�LR�C-�>cl��m����gdx�`�������+��6�y����N��HV�[̓�|�gq
�yq�ĭ�d�7��+a����i��E�h>�_&%9+ fƒ�/��\%���/����d�uϰ����|U�}�\��	h"�7 ��)J.a.����r):��N�bKw$�fR��|;�{�-{Z�jst��ї��/�A��X��_a[���z�f>����59�|)G뭊w�H,�h�5H��_}O]q)%�9�=�]�]r���*���jAz���ta��Q@�o��uQ�~5���/�T�v�u�cu��
<{K�A6��a���&4��o���C�݌��2�y�Y�ݚ�<V�՞YϦ�d�����k,Aw�)�	��!_1���v8�t���]v��fc��&1�X)^U5��Äȸ�����g��<�:Vi3���>�\���#C�Ls��6�^�.�(�^	����b��@���4�R-�\�d��>���}Щ�Ig�B�~��;�} A 4���)z},߽���� �S��b�9���qI���>%ב�s	��7��N6̡v0�����NW|��W}�fͩ�GCT�4м�\}e����jkY��g����R��X��v/�د��➟oߦ��Z��*�2Jl�z�>��|�
}�bؘ.����P?���W�u���)����f�xd��!֪ޡ<���?�3Y������J���l�<�a�� �;�m�Y�P���vJ��$���
c����~<յ�O�_�s��4ߏ�F�~\�z-�~�1l����M��M�T�"C5���sЖ�@$b�_���<@m\�1?Q&�e��KOg��\�Ėy�~�ot��\N�c)r'[��_�<U������~�bY�u��VNX�c,�<�K����$/�;'ͷ;��t�oO��ҩ����p�2x`��6�n�4<�+�7���I�J�t�7�7�������d��<^��u`,�2{k<�T�m[�5�kT���l@�u�mL�8�Q[�i�t��|'Z&��{�3O�"���n��|]��M�)9+T|�2HPX�p|+�V�1�D��XCRm�:��Ҋft�K��a��[.u&�t�}e��3�*>/������Th�W�}�Sq���[?=���8��0�U�%x���7m�e藬E0թh��r/)�Q�j֧�2c2������ �nê�O�~���&��a	�?�����ȶT�#�馯�}[�9��:{��f����Fv�ė�1��O��|�ؼ�b�Q������D���D�	���З��R��	x^г'�ڿR˛����mL���9ƘR���1��k�������7���=�2x��ب6j�7��𺈄M��6{~:��
��l��1v�_+�ZK�H��b�ީk�x�|'9�+��+���ƚ�E���}M��&�U�X�בּ˻'#$Z�l��Mf�s\�}~a�g��֣���@��=�ߚ�?tu�(�~$���2��v@5!A<�����DEv^A�)�l���&�&�����G�\��wg�Y��Ԩ�2\u�̞�_��X���B����C����H2*�����Өb {� �$�b��7������ڵ�-�K��ѫ�ƀ�i`~*+�ƣ���$��/�Q���y�aq��65���%:3��O3�����WsP�.-ͼ�A%NAkW� �F��p��Oᓽ�([��h1���f�
C�Y�/�]8#��
�W�5�j�r0��s�X