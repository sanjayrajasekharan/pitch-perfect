��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����S�M�hkF��1~� Ά�``0Hɿ��b��i�<�1�SzFĐ�48��ch�iIQ���H����:4(c��_V����&��}�w9B
��T#�_qx35t���D��<��R*�E����nK�N���������19N3a7K�0~��!�@ըfG#�=V�[��&@0Xy8�U�N�
�y��I�S���j�kU�,���87��u�:]q�Ƒgh��8�i;�f��ܐWq�Re�R^Y�˒�
�1h��{�%z��1(Q�,1:k��S�pv�p�$�듮Z�����C;�y�A֚��Au��*��1�-�_��e�(� $��d8T4���z"�������0����W���j�Eզ�$f\��W�t�(;�g���u��A�j(���g.��=�kz�7݅cִ10m�OɅ��1YW��F�O�`�,�w#{�iR�{���X%>�w�?U4�re�C�E��C&�i��r0��vf�8�ԫ�ft�cY!h�����Ϸ����q�ׇ��/j�"(@��c������mI�kru��)��2��*��0�r4�������i:3a����-�������g=���\6A9l�6ιB������:p��Y�Y�[*i�29��w_�\�&�h+!�)�v<�}�!&��V� !/��y17�&�ţ�*�Ҕ} �2]�H�,�nV���˻u%x��[�n^j^���XԞ:��
v�9Q�����3.O?����Խ��@��5�RlCN=ۛR�J�%���oP��p�^;�m���`CF�zw����'*n��dVj���:�3L�@���w�������UP�{m��"ql�2x�<��~.�0�幺�_B�5B�J��m���c-�BaaU@��@|fܗn҈�q�u^�6�aW����/v�=�i-���B+�'$�f��S15�`���Q�C9l�yr�����(�wJ�t�n]���&��dE�TZ~�T�gӞS{\t�lmх:�ѐ�J��o_]�S��4�U�3Tx�{L5� �[w[OI��Mև�7�*+y�I�eY+#��Ӣt>�e��`����L]
5��ÖF_�wYg4�冓�m�����W'�!�����Q��ٮ��ll*��d�PfS1|��)ɱ�|��/Q|BM�0Ἰ�D�+oa��wJ�4۱���b����F꠰o�Pk�Rf��)��"�]����j*��F��Ey� �]Jp������n�K  嫾�:����px��cqT"���� ��jZ��˦8,���� ����f��c�Q�`_�|#�%F˒��mw^�`4�7w��B�Q^Jb�@��,� Ү��M�1�ZB�|R��d���L���| � wsL%l��6`�ն{���U�{r�R�d�d� q�,�߄�]x��<�@?�������yPW�e� �w��s��3�v��o�eI��?D�������1�}��.q�0�)�1�P�4�6>��7Jټ2�q1"������3GD��ۖ8�fzns������(n�?�>�P�뜍��;��-s0��-XƊ����Y
������AG+�(n�ZC����<Zpd��tO�^@;��*��ܯdXU�+O;B��� ����X��"��Uq�m�|��(h�M(�s��4�T�-��M�6޶��9O/ ����T��'�g�-b�;�Iɷz��@x�r��-A=� ]R��1j�L�[�����cb�a����-��&���0���x9wX�^А(-��͠�g\׏>�20�c�_�}A��:��g��0��v��O+G��������L���}/�Aq�);̸�X�/������F������@T;j����X5�ہ�U0ME�w��Y�JL=��Y,ޤ]a9���;�KK [���?�[&��@���U5� { �(�� ;q��#� ���J �#w'I�����n�V�E�(|}�`m���1\H�V�qF�i�*"ۻ����4}�G_��I	x-�js����T�Y��_�\���smX��$oh��a�S몋ebv@����;��_��W�V��s7wq7_���/)�ʷ�4L[$a,S��d��
TվrA��~� ¶���^�:e>&���Z����5\w�D<��#�P	�µ1dYB�d����X�Hz�����4����:�F�a�ݩLV��yܗd��/A_`��#�Li�RnW��w���� R�V��]�X�)t�8��rg0Լ�}"�d�*Xɔy�V;�G�?���AI��P�x'
� ��P��.��U<_bv�i N�Hԋ����zLV_5����ɏj_.]a�}�� ����C��+�����CVC�ۑx"a$�يY��(����ʼS9��o"��J����6��HM�Kࠡ��3�O�f��5��hp��	��}�Ҽ�CH���7	YE�)O-v��h�$���PC(�2��e��W�`��'~�nEZV�	����~+
ƥ�C� �>� �.9=.%\Uh޵�Ƴ>]��'�_s���jjc�YC6 ~�d�Z�u�x��\��->}���[�:V��@� ��/�?^�W�E`���Gy�BK�c#%L}%f6�Ǳmϻ����[���3����wA��H,���":5l�H	���5�����B�A�E��̾�,�x�=��¨}�8�?ɣ)t�a�Ev?�=��ǜ�mw�')i	d[~7P
�vB�^�h�n|���~'8�*ӳ�˃�-�t������������2�Ǳ�N�Na���7^�
z��+���Hs��S�O�Z]X��5��5(m�w9JPf�EzkN�3�q�v�x&`c	�����������a�Y���B�K��	�
VF`tKu���3$Ձ�.)ℱ��%��P�v�ʕG/������>�?9"֢��U�mhf2~�5wv��1�5���Zv涟��n��4M_G%�_0	'�	��ةL�l���Pl2a��j坂��f�a�s�f�x^g�T]�<�yK�9b6�d]�G�b��X�P��pw�xd�:��Q�WqN���$8#T�����s�h�8��\�;�7��L�i��t%I�@:�%Cw']
*E^�[A?�rw�,]0�%�4�t����Ʃ�v��s�Fz5�[\e��O��ɧa����3)��j�Ⱥ���J2��/7_f���Ɛ�X\Ѝ�D[����T�9t�{q�/�W�}�TyA�����y��A�A,wk^W{6��w��_��Q���R����Կ��/?FF��w��/h�x-43MG7��V��sU�F~� �a9���*Y�`ao��4�J'X=�MCG�F�U�~X�-(�6!t1�Ci��i9�U���t𙑅��lj(2�^.�o��U������-�7�02�Ú�H�}(�/�ٜ�/[�=��_����r�x�8�q���,�/���	��s�U���|��vw�_��Ю[���n����|"�������(Ԁ��F�5i[�mg9(�$���'�h:�������q0&�0
��T8a
�ѕm�%ʹ��s�ͦ 9v�ר�[#߫�h�ܽ	�m�����K��,B�~Ԕ �������:@'w9}hmOӦ_{oK�����ԉ"U��13�K��NWY�%%3��SH8�}֥�}�4a��nR/�����@��ˀ�I��U��,����3N=MNx#Vo�w�̉\U�\ď"�,|��- =�ْ��vB�����-�&e��!�#����~ QH� qax3�˺�j��y5Mo�l��Eq�lͪ�r��/\���P<���d�[���M�����'�ũb�_V��v/M��:±�)�ܪ�4���f��[jx�:���������#��W{�._� ��~����x� nN����4��� �����	j��׃�M�N�����O��5�xj���ʫ��!>�Pź����Y��E��ʸ��A#�[;($e���eS��!�~�1�a����v�zYw���W�x}���d
��XqK��JK�� b{�Xr"E]v�hti��_S0��RSn��;#��u���#�X��p}]J���EZ+�0�=�Q��*�̪�Mwh��`?���5+��jyX��`Fy]8��w�<b@��0)j
�gf��߾(�@�N��i'��U�����m���.����7?���*#6H��H;�ꟊx.��X���huwuP>��Q-�w5I��q[����T�����L��<�$bϦ ��L?���n�洆AK���Χ`��e�,��𒇁�<���o�0Kѡ�v���Ʀ����,�F�~d�V#���R�����om-�wQ����d����J�Y�(�һ��H�\�8�J��Ř=�*��x����/�����V�?�()�d���l��,M�0nzŌ@�5P<v���ǃ��I?�z��p<kD���Y�Cu�1l��4w�,4�o*T�l�R��K�����І���(�M��b��jv�cm��wL�8$�叔`6���V�:ITLd}��D��/ʸ> �H)&��Զ*�G�h�����le�J}����|�Q&�VA�y�>�y_� ur"p]��?�(t����a��}-�T�%�cO�WN��7�:�~y�W�� ��Y���Ѹ����<�Ӕ�yd1���.��J���A�:l�n�*�b��zh��'���7����dhM���+XH�Ң��5��C"zV41u�& 	.IE����K3l���]��F2c�!sk9{��%��tcZ	[��S��F[��q���Q������Bz�@�i���U{�;�Nj�("��S�$�S�_`�&tm�T��,'������_Y7",׊gZo���g쬸-�8��{�m�k�����)&8ɉ|�R��r���E��R�M�2��+��'�a�\�i�7d�r��Aq�g��َ|�V�Z����H�O��z�9��hu��7��HR�O�c��*�2�=L橚+ry�����E��~��9jt��U��e�z�>�Uς>`n���FH6m[�Q���e�Q8�J3�����7��__h\\Y�D ����j�{�`�*X�_q�y,�Y'�>�]	}�s�ڹ�K�L<�Z[+mu�x�M�"=K,D��|�],=L���q[�g�^$��.�������n��Q�L�9�.g0q9bR��P�y"�uO�β�Z���R`&�F�
lD�&�e��Ԡ�y��/ݶX�q>�\+��T,Mj�*�u�l�-�`gBe\�'�N����HN���*�����B/d�DU���>n΂~������r��XU]�k����� ����$�<�K�m��!ړ4��x �ڛ~�C���Q�Юu�S\s���v0���\��R�`R��V��5+F�]S�9 ���=�ի~s��8lX��U���jk��Y�?����u7"ɣ���[pE�_��˹�#h&�hl�ً�7�k)w���s3JS
 Y/i�)�k5�db��yb��ng2��Y!P#ތ�����X��:�bC@�@2�	c--M�bz�Sn���@ƑP��i�PZ���a��
��%~�hqӅ�z��?�ȹE���23O񝷠��J�ި\p4���"W�>WNP���O�w�],Y��U��Aaх���i�_�|2�g�Z��_T<	
��U'�k�y4�Kz�������� ����!h&��௭>��30|Stj=�*��������ѝG�N������l7�n�|[B�Tw��S�~ �Vd6��De�MK�"��&0"$�����N{q��V�3(�jv�����qz�l�@����ܳn5�!n	�u�l���BP��^3?&�E�%��W��~S&1Ȱ:sY#����jj�"ĻW;K��M��;��v����@0��U iCU�/�MR�~���׵ḽoV�Z4S�������#J`�H�|
����m;K�F��cI��P�4)��)���u�:�< ���Y����7ؖ�.���<85*����UD�i�[Ou��Wʑ�:�z~�5R^�'+{$�Pۤ�w��+ۯh�L��,R����HN�Y�\���+���{An���iej,Ì��-IIߏ�8�δy}��6�'G^lB�l���0f J_*�5;aߕ���77!�Bl�u$�"�)P^Df%Wq{�ˁ	��d��	0�����n��,N$F�>1���\n���!��9XH��w�lW����H`4�4֕�="_�-����;�
�'���k(1e����M2�p.�����}E�ۖ&P5~�!�\|�L�7F��㌽\V���X���ȏprcV�ս=��ݒ��c>5��d��N_�4����p�8�kM���]~�݁��u�E5"H�`��ū��ΨY\|ᇑ^Yc��ޚD{b8�BJ�!6����>6�i���㋹:P��2�'��bο��DN&�3�|c<7k��>��W�ď��/k��'@��~�p.5� �t���T�s���d�C�i�9�e!�Sv���1�\� ��=P�.Zu�G9N���&�1W�/��w���
ڥ�����E�̈́�b��T� X::zQv�ͨ�y���mCy�{4oŮ��_M*�
ή�OyC�+�,W�O�2���F9E��ڢz0��ҩ��ȟ�k���P
���l&OOhrO��C�[&F�a#䀡��ѣo�����~S$�t�`��;b�kά�d}���69�V�=���HWl,!�1b�^�������q�-��)�E���u��I�&�-۽)>����"^H�ڈ���ۚWh�9���M"���z;�ġ�֢i��uIA��I�~�HuY<}}oxgЕA�����qO����q� n��z4v������i/I�V�bv^'��,�����v[	���a�S��܃ տ���o�=�G�
�,�a�Y�(i�!0�6�n�����'v S��R����Y,2��|�|�U�}��;�"�U+�@۩��T���a9�����a�M. ����
��b�t���Gߗ��L�
]�G��Y�_�,�;����՜�>mÃԸ�{L��~�N6�,���ɶf��><�c�7`�51�Û��te�ѸV��n[�r�����kޮ��C�+.����v*�y�2zF�MN�E����� z�6|:�����fZ-��#��&$R���a�9�p�M����L���P1�-���g�C#|��JdȠ��)m~^V��!��5Ü/����>?�nT??�6V������)�+~E��z�ȸ ��D�w1q�V�.�����R�T�YP���M;U��5�g�&;��+����zw���mfx)�8�*��z4�Acg�#�
��y�ۙ�3�V��'���Յg���G|$�"�ڨq|`�ڔ�R�f4o*V���+�w�U:��[>Vٝ(����д߭Dduώ�(�\yG�JϳRCv�Z�8t�7���;P�p��J�QV2� C�3u�=�6Z��k�d	N	n���N݌hC������R1p��H+s����W�O�JM���ٓ�j#��$X��wZ|�K�W�q
���`�����p�����>���ᔚuO���r1v	��-��o��K�Hu��?re�#�8e[张BsYep{���0�W�L~�(�[e#P��-�l�uif��a�Nה�B}c�;�UA���FF�*8���?
.�Ӛn�4����(� �4*'������u�����l��qU]W�7�>E_`�v4�6��mY]R��y�X/��+M��0������V�C��\o"�g8 ~_�k�6�|'��f�rζ`�},��]���(�u[Ε�譪b�A����S��1�5�2�4zg�h5�%�d���� ���y�~�z	Y=��]/��ݍ4қVX�� �1.0Ԋy�:����̂�.D�p�=�ڮ�:`�Lubj%�$���?`�V@F�O'S��(����BC,}�ۜ�?0[���\c@�پ�+���6f��.�NڡM�<(t(���x�����s��d���S(!��F\���v��a?�{�z����*������ɆŢ��_>kqz�]s�H��^�����p8��Y���*z��Kx�0&��c����VPE#�����L��#ebb5� �d\��$x+7�T�	ǯ����/[�p0F��؁/:,x�r6Ky\���F{C��^Y@Є@ ��Ճ�L�V�gk�nb�ƽ�L����'�%K��^�T5�V,��/\�w��z1���]��������&���)k����XޑNe�ƅrݸ�P�Ann�^�>L䒔5�S�p��:��'`[pS@o�ʊw����*B�D����_�ͯ����+ۋ-,�-O��'W�b�f��#�D� "?�}Z�@.8"N{�����gpsk<���Á�QQ�٢]u�z�8{�,RZ#u�j+VM�����:c�U��z���=��Y��	��4xV�@-E�b�e[�( ��dr�(��>E�<�:T�u�8�9����.$x����E=J��]��G<�#JY�{!K��"'-b�ܳ���o�'@~�-(���{�-
�ú��ķ���21���HG���u|�8���ej���P�59c!���uL�I�C�T��=����3��0�q�p����Or�љ�\��l�E�O�kWl�^*Ip1<��p���v_b����	����E�j���<����W`�u��@S�@��Ij�R$�L"�˞��1�B9��2��$f��ك�8yS���L�l�1_^St!4���+�w)�=˹le����f3|76\�hژ�{.~g�,	V9R�у�,�L?P��$^��X����8��D�>���f�3��+]
!��_%r��5&��y��S��ͨa�����plm�yq6�&8`��WHƸ�����td��6��e��Qp�p�����r|~c���F%)�*R(ɜ��Ù������ɰ�3���Be���閹�Co9ci�SY@s�Pw��	�J�m�]}�J��c��~9|{��������VvB���( j,G.���jSH9#1� D$V%�