-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
d0pd/ABGe7HUNRavZzCrXfV+I9JLOQ9h2D7K9Wj6LG1OumGK4pSaimlSf6VrNUwC
Ge5k0B94NRptj10bkjBqKXjPsuFQTxJols60/91Bwhyt9wHOWOH7ravgBQ7cZDZH
XWmqPLeVA65CTwLPetqNCB8dJa/93XA67FwX1NRbmM9Gon0hOj91mw==
--pragma protect end_key_block
--pragma protect digest_block
E+FCYDPDu/5TGTRKFeWWoRWbmmk=
--pragma protect end_digest_block
--pragma protect data_block
TrUES+NqIVjnDJtBLvM/RvJYoc+TYsRNlQK6/+v20oLgAMZAObTQYDU+/0cZcqZs
4LsfJnvac/wM1o1QLYBTygOEbmMbSiyiDDCA/CALArx5nJ3cj4jIUl3geUHusGyG
bLDLCeTuowfon8F19m0rOlwCRODeAFp1KulmGrSaf3u0kgMwTOLwAbyG0TxRiIZJ
XUy+u8YF+5jQrnFMfQEUNGXS//uizVEANy0mdtMwIhFUxrGb9jK4NaQj5DISpK2I
TPRXcO5k8CosHWmN2Vp5EdI4kvdg1Z1nrIkXxyLx/aLw8wFVi3FN1K+h/UbqFknd
LN071exqMPQn8VI15dZF9sQIY1sdPx4ybc5OPbtPUvFDTQKRDXuyaJGoSvTVXtoN
SyDKLnjfpHejaUuc3PHn7dAwjVpSqEQJT/0eRuRI1+BP2j99xudLFlKydu4eFvOn
QkM9x+qK8mKl/PsXFmdAZrTFDiIum5YMc/jKk5SyE0EsAqJFI07s9xKSfTnxxDH8
kKdo4tOIs/08N0Arx0opWj7jVMl2kOn76fxqkydSGifPGkVA1McQGWRzrRiwDKFx
HRMZKpywaPVW6LTapcu1E7EUarQZxZtRFirOC9LA2kqjnmj8wQFoz1B/CpYeGSkP
6wJKTInTQ4+heYh3f2nwOdgdw2He+ntSq2Fa9BgLDbJDoHug00TXBAKQv0seKp8I
s5MsE/mCzhi+RbwgwuYhfyP5FkPM9mPIIJo8V+FUXi7fe19UPR4YovlFZ7XB+YMf
I+NyEL7M5jxZ4duf5bDC9Xh3tpBnUh5QNsvebHbSiewDRGR01fwdyR7wzGIt/aao
PBFaxZdMHGyOItCu2HCiqyx8kZt4Py2JPUvz7MdfzbQ84t2zjtbffeJOpZiQLWWK
QvsvsGTy9vQ/X1zLO7Tv5Tj3kgVzM0dafT2XcdmU0fSBHAFk+WMskSqmHnzgiUpj
KLrARbGzLvoT3w5Qu7NlU0EQcI6evj1Clb1VUzB1zToairLi2myZVU8oipZoylR4
GvLcyeGmOOUId1S9OVMoE43AA7DAsllZdWHBM0KVmF21t+Nr2/FN9xwKACOKjTjS
8XLfIZ0IDYWPbEkINDE7GytcKISiZhwcFyN1aI9OPNaNhpMOPFZk5Y5tm0lMo6xg
79BGQdz6CkvpfLFNf6dnM9K4aMiO2YwFEZ9ujByGA2Xu8nRQoeKgjwRGapS+tXiG
ejK49Af5L1J5ZIAaykF1pIp3XEIOcYIwGC31n1BB6cxZ8vz6JewRxIaJ0NP0r72V
vYtCnxFgrqede6vIlc6YpA9AHPTXkgevXV0aMYE61Up/OJj2dAZiFr86RMn5CuVK
Jm2F6JhVis6iZxelOft+xc2ofOO/0AsaC7nshUw8MTb25RRk6CltmwUws2DycWT2
IL/VFaM4Ph2gBc4mgxmqDEXJUCnMpWSiE9jGFXQhqccEtl4j/ELEiY5Jl/4bhJDp
VSZ0nN/F+l2APQwQ34HRcImaMjivsyxeSoym1+AYZvIVQAWCn9C5qaxqsy2f+2wO
xSBCOGI4T+imItFyn7ooEUKLrZUk+dUfxWEK/XwZxPQQi0zCGYrA9zlKakBJINMK
VY9yF+NsLA14veTIX6JFtZWn1KhJrlBUBcpVQK5ont89IxyWzHH960Ib4V6+2vHA
u5qiY3DM2qdlijz0ScaWdA5CyVh3o8I+FsRIeAqe00Yq0SzbDtwuZ08CnleyD6ur
Jo9gqd642xogMiCs5JhOeUOajnqXjD7gzLLpjrH3gINnnvqpKynEL3tr9s+jqjca
llvSwlVWY6acFTUad0wywO5JrSCH3IrKALbXmUr0yjZkyXR9x2l2h/dHpSjcRRPJ
FFjNiLtZ0wgeG90uCd8gqIQVi818GmL1FS62kMq92PayLCtu3TNPBMKw4Bdgm0/P
5NIYHN42IZUO+pLSfNtixoKzz33neUrjFId0qne3vtUwyIegZTx94ssv3B5eMuxr
oz/lxA1mxblQMBg4yS7ptWLIMrUzcqWl6LfRgRGyaypBrMkkAJ0q6oXuvcaGLS9w
wGM27IkCLhN8vCRtDLa51hEv+9G8zM67ZCyqipmsCKKx0FCdnNMhM7mym/e56Uxq
rUogWDx4srJmLZFOPvvj6JGHxGFpix2HwdRz5e+sHmXqZvbEJxm6FF2PZLH/3ozq
SGJ9d9NTDdr5YdAfv8rgqet6XDx+ptcc9ovGJJEzStl5v1UceYZzbRCbwwU3Dhjz
ggFY5IXDBT72EbrbOCWtLTvVKkfmAHyf6O24bldlUxeoTMiSCEMJGTGMaJswl680
MeL/72XsESZUdPhXi89D62XFP86OVabz4VfjGd8qUj43hM5cqBPq8A/GybgaVYGf
/QUMHxPHf5cZXRenpzW5TUhTtrlHeUK6G5WKfkn12II3FJPgcb5RY9WsM3mKjJ1+
yyQ+jdU5mTv8X15SIQWGJIhrRKSfR4OChALNGO/0Wh1lhLCzFHRM0UlaAoOQLvuj
I9OT3cD22NoNDP9HYXsZJ0hlj+Lo7OGX2rbOBZ2+ydRLclAsfiHa3mVtKpnynzS8
yGrtBRmRtyeAiSJtsQFPks/hoMsNlLLFmcIataf6V8koMsh73qEeTAm9Wqd1EIFk
rwLQiiIB+rDEJ+Xnx+i3iRuxXHkF0o9g6jm5SW7+MAMn7cml8QrzXxVYYuN6Yuh4
JXPbvjSAWKLu9x/bymRmU9comk7DVWu/p/Qo+mTGkQqacuc6LIMak8r9yCRDDNvo
UTe1Ij0Jf6m8ZRAZYuDhjzZFyeJjLwDZft8PA5TtxwHHlMzwWrUpy2vsBHz2gll7
3cVgbZFSqMtIRhimcJxQhb2lWx+GyeYA+Je6r+IVBoqrPzbfPRdhvQWwwJ0bJ0A1
y1VbdlpoFJi3ujmRs9/nqEQ11Ws6Z3VubEd7+SOLc8UPPEdN7OWSv7akVfQI4dZY
QtnRqqVR5Vasj9fXgl/Ldms9K8Js6YmMu+v/tneLNFDAeKLuXzc3RziuMuB1IZPY
ISoX4UH3jwDSVYJMWfohkbdf3j6q5+OKJagqY8PSFmm7H/CKI8+ThCRyd5wgjAHC
G18ZmRb4T7+LGde1tBxA4zCzTkIyTOIys2Bp9ovqI39I8ZRhWndpJ6geCw1npYQX
syxWHC7KcFCYQaPiuxNMDa/2Ex7kpR8q3NU+FhhkFSS+E8MVH30rFrst6WRMA98P
7Vmza+O/cglq0tucrU+gq7CSrZ1V9vwpPc9nMjOAnSZ3IEzusGwarwVzCLbDzfZ2
ap2MrPppR5hL8oFjp+BQXh9MQ+qaomYegh0N7kjbWwr4Yr0R8EtWWgKh+6c5NGYC
b3CqipZaZgmAEA/qUJ/YvSpAJGz9X80rWADWtLL34pZP8D770zp00x/hJ48NGENr
xLqCa7w49H0yLICbyF+4Uc/rEDk9XSYHpW7pmz49fltN0siZEHQms2NU7tL46Huw
HKsqByu5etWuhPUZXZy7Wx5yYO7BsRu/6/lI4zvlfeR6L3I2TKeAYILbbqMGmrk4
IHfZnfMPcM2CmeEqyTqF48hC14zqsZGCbIMgikvnc1jdnuVVtuVgqj2FAenStLlF
WpY8QjZJm2BRMLCBV1Fysm7usfEihPIhtoCs7ay9j8OdxlxlDOxqdMIZDA09y4hj
01VCpcGtgORqhRgNb9Bw9KIbg8y82709PZ4XVCXXpi6L9pl+ALElc2lpfrVuEG20
vsLNl98owWpOBDHioBQkDsqDxNC3TiuV9Aisbt/OsYyfM8T9cROP+31eqcIfPk4u
3TdNvoqtHQxC8V3zWFabH0h/3vR58kJ1aFCyMFjFv2u0+KzzcPFcOIUsh8hCd0Xz
VQWmjXBgJiOI7BceXdVNRO2jKrzgK5FPAqnVkICbtdPjtBOf2EmNJZp/kauMAKjh
6QKw5ZllBvpIHuZLPT1n+G17GQmPw/QEMLOEwYOMoa9CBmhtJuljF3SOyeof0atG
ozVrHmy1oi7rFAT8vfx/ZUllNgpUScRZqJFix9g89prIZ1pa+mrjZMLgZL8Wm+mz
9+RboS6ouuha438V5bWnuoAtVnqJQCWTfOh80A/uuP9N8+Jh4RVuv0al2b67Dl7c
46hexo5srfg7vMPL3zhRVRW0Ib2+OiJexhVxbUHMa28odiAl04RbBomb13Zpf+YH
u0TJbUgf/wwKiF+XkmL0kHom+a8WFGTenoJ/GKT++Xkms0kAYE6jbinCOdDJYwGO
SiyhDuoUt5sLN+tHdjmOM/Gg9j4X8FyRThnStK3A9pL6Lj0+TTpU4BzZsT7PF2IW
/mOI+o1tDBKJi7Yd930O6+g1dD02Zedod+U1kzqnWdE+5K25tlrr6RzBotQ8EdYI
wga6kA5vUDbACbuOq0tW+hp5s9Qf++PPWSmnj0N+hy/cEzkdKA7J3G7soKEdcnbG
DgbMml8EnrDIvLhxOL7y7uReSSkUaVwr49HTulIXYkRdyKS54fH0uoiE3BVpxGC7
M6cuItkuSjnyw2eiFUhdcfN1H5GrUg7ug3EwmYcBDCZwNt4wwPeCfLfsRVV1kBzZ
U3utLOD9RX01DNW4OmeAJegxRgttKeQn2qCfisQcuGRgyu4mrAHuoDrQJPweYI5s
bVBz2Nh4RdBwd5ryZx00HydvBgA+TZPd914jrIshazHWhh8Rt32Be2yH2ljL5oug
hmvq6Fi8AKTI0TmneSqQOEojvzCq+SBtdhn3VcXb2v+WPK6MYSoqL8lfAMcjGMpm
knbff1qumgmO/PHk6+6sXkU/mYcnjSFf2jV89jkKPW7HzbyziJ7I+9E0uTrXkNpZ
3XqAlNifwAi72Rf7tfczo+Kn2gxbLP2k0LjzE4gbw6yEmk8Mr3L5eEi/tFPvU36J
rLGuvjAhCeb6FawoW9tstddJY5zNABTRDmzBzuoQCMBWOci2uz++Fz4DtLerXmIU
llr91oTWp2xLLJ0K8xr9XhdtbLFmDf2gvqVZER1nasGGbs9rVlUZC+QEljaymM/g
CZoWorfUd6DtY+ezmN1dEPqgivzyx7PHtFbOMCr79gBLUo32jXjo5Gclb968qNZU
qUzZ5zu0by8pos7v0jW9IdvfRO+wv3mlk73Cveq89vp2nzyqjPeP9edKikNNozAw
WWODBpr1FLOycnIKE/IOsjxZUcvv3BSiJholsnNyHZyDtSlQ6rYdCSdcJIRoYKRA
IzM1CbSqsi9Kgxvc5vy8o2SSLwrvqF5+xia01pyrB0axMjAoZ9s5K50i+J71ZDo+
WwHlRA7ew6PUfcl+Ohsn2JTYES4QEdk5kVJIW0F2vg0ATUR4KvZYM6nymeiMgSMd
xBD07esgn2+nUOtozTFBm8TXAPbATcqcYs91/KXsHNwtX1+XbjCHwzVN1+ZM2W7M
2u1f4yQ0b42Gx3oASZhLaIEKbjXa6mpk7//udJKq23jRsO3XwSI2e6HBzJntTf9A
5dwGHlGWkByNFnNECLYqlFfeaFe5X10jsysJ0GhDXNN/LTJpvdAJeW/8+R40NM5b
+TX39lGhb+4q+ZV0USZIPkD/vfbBqMk/rn/u2vUAv1F3PqDgXg8D/WryOMcexIeE
HXLScaAyzjgMVke4EX41OwQ3ALrU3z0QtavlczNiK51dc6amKSIJvsCArfNLvzpy
k9avN+5mrVquTYflN+AFnO1eLeumk6adXCTMEwpJ78dBC8rALLyEZ93tLjcUNYtu
ep9/jm2y65bYwBSGh89hUxef3Dx13WH+CsbxESdaA5WwS9e/0CxWtW1w1aMoRgNw
R6LOBf8hX9yzugnWFn9qXixACk1ZjsVhhxfv7VTBHnuE5oAcZxlD56XdHbdN+ap9
q+gvJCNmSHne0fcrx88Zr/bxYTde6AEKLxUQnYNcMaMyUIt9DkaXNWWtSbY62Z2J
9/anM35p5K8MXFvnmKDn+AhKJqfS4K/HfyXvK6vSx2VbFymOt4XQie6FBCPqSgK3
mpLo7lRj/AuJFMIX3LRLCbHjQSatoKS9SJ1bx3viJXxLlN2Qnanb1nD8hCFEeUMB
/bi/ytHZIAasXF/g2nszdltKOzSFDi20/WiPvBrN/Zswkrp5h6BcI6zKtYE3Ig9k
LHJKdLbdZZnNIqoidGjlzTlRrLu1TKHcEsZdNhzH4ZPJ8sKzl9x/u7cZQ4mNH4lN
c/lrEh1+L6qSiBS1kf2ZwXpSPRDDquJBPhj+VIbZ8220OqLWki9BU6hzXivHTyrR
QN6y4DGmC3Q5YQvf1TjsCShM9iE4PDBBV7/IPxcre5yta+ChiwBLaBCX8LOTjSiM
hZnzm1BP0MN71IjXSKjIb/+TNtTJD/xHCWR5ckOxAaC4/W7Nx+lFRKL7CrBIK7QJ
frwP5ksk/Sr33c8R/v0OBhCTUKOSn1mq6oKih72G5joETqTApamc6K0+/TK+wt1D
6ii3ndhMhC3i6OuOnFBcA/jad+qZr17/Hvwn19zB8kH+zUox2ck7VYPEdqv1LNWD
V+SbCl1k+DpvN4mMXBDi+U4qNunYKlZvFa8PMNzcBSM5ks133V3hKXN/WgoE0s9R
bC8bW8UCfS7gGp+2n60JRRHhLgW9XvHNbthV2EbnJ3DixP+e9deRi1ikmp9YKLW7
fZFhoSJ2qKIo33wAviUr4qz/wqdA0nkw5OxOzBlXtnWiBKnu2OkmHIWpCtHpkTZH
NqMRf/8rNLBBW47Fj7Vdtnfi3gbYMjcKqpHlgL/EAJ0MNPVKIWoiWhK25awysGzG
eZBR0mcOitHRz7So88LjCwxT4bbQ1VI5KeAuGHfmtShCJnOG+XRArWJv0DH0rN9Y
A9ECietrnsTVyGSs9frYBy3SSzkDVOvN6+/oZKSec/Mga2iuhtdEHp2Te63xXm2A
fIGvwRNzxV19jJUdXQDkw0ngjZPsrimV74cjEcZir8Rfp/7s9FxtiONJ+2KQ0X5n
Es6CnJjpXGCwHSLmGpZC7Ss0jnSbej9udMC4+aVUrV0SxFSK8qmoWBu3hO3yz6Bn
b4bBa5qUnFFmKx0Dca5Jy149vHq0tsGHQmaCyEEa7uicI3snB94iLRxWHfn47lfh
fPrTTeqsweuoxnWw7dBfr5sEsEXWNYTnkz1T9K+K717gtD4zO7vRMWcR2w68THin
3P5gx76YQ/Y/SjkSp2fk+GblN21h2IrFuEXNf1io1t9m7mbUZNoSOVoYMvecA32c
O0wpdhnG17m5QdSWjdmIYNGhD5A7Bz7VgkQW4KUM9FtykyaI+p23r8vkDZ3uKU4s
6xzL3XCRbE9oLUyJgPc3oi3zZcAHgPPBO33nr1ecgaS+kx08VjMKF5jXFFcYA2e5
aR06V1lxz9b4DiceVMWosTYGlzcaAYTV1XNabUQtC+MAn5jDQWL+Wzm+hR+L/k5I
Aiq+X6a1/Rg6DcL2TS6piVf3GB8kuSu+mOvg9G9ZJGnzKFS6/cv49YtqzmmPwUIr
uXny+mDh+TMdor87zM27dyk2gN1JE976ez/nnK0Bq1Pn1m0azk7erKDvHybcDLSu
6NZ3LPWRuTic/jFdm0p17FBa/53QWJ2L0K9v0zP/2jG6rxWgcX+Ow4UtZcYOGjeq
7VPmjMl1vD1EDrPXWGbkL/3vBdKjziLnXR71zhDj5QhbkdPmG/uIqpFtjrLSI0sW
kngmwTdTFrMimxKgdbbp1b7SjBIDhMLHakIHP/e7BnB4XHnCdenehF3wFgj/Z/hP
9Gt1O7+cOTdP9vRb5isO7BnLm5Q0z1J4zgWfnRPLg2p3zb63KkM1IYYhC9StB3iP
ygM13YtqSvkqypd+ZBin2b7pWjv8YtyZgXltWXWsMqrJElFEY+GyvwH2LGUhTlz5
K52nahcpwzs2UTWWn1xdEsqdugOvJtf80q+1zyDYcKFYZJiG66PAhM/oVvLbrEam
r+of2q/wNpAcDNvBIHdd20OnWb/q7145qLPlGV0D+zGqy+Pcclw895/pLy8dT0ED
4fmCjhHkKcgZ0rR5tnss9n7JVj6t0qFnB7hcnyZ/86B5xyWOimqj8b5UbsFprXF2
kAMrj6vFRhCigAdJFR+M8WWAAM90AZahokQxtUUzGUlSeOkQWTst+PahihWZvobh
7yS1AW9lt6t604kQhz4puTOCjoSVkKYfkdOCstQGwZok3unwkeSiUPdmqpV+kiTZ
oBduaMmA6lMQWNjK5LTbTo8/GXbXUH1/PRmubyKP5y34l+e7oOeX36bSzcOjOYWv
U7yObIc3+WQrpo03O6kyev6p9N9qeuA8YWc3FFZbBAW7/eCUJBX+Z9Y3JExQgf85
feYi2mdt8WPdM3S3uxhmaw05Hsb42kL2ICiA0JTqNz6r+otPRl4haNxmJH3L7aOM
YZLnEhAjX6Xf4U1YLyJUL/DmYSyZXPwYPjWTupYksseJztvqaPUEemq6RORYRGCj
BWs/+3QD1xylcrabC7mhCZNmGUV3IVSA3HQOeL3LncHB0dpr50y2xXKNLvM84ZUG
zvJ8uj880FtYOp/Einypz91oO6lteyTllFoKbjk7/r+IjGKwVx5v9Gbwm7QGesCN
mLtsXXcuVcHwPR/fgiTRjVuzHC0ael7ONJmPrMhe0ZL8yCRFkpuY4wWdNP2jTYcq
3i4gDCooNPrKVVEdva+3nGncba2OAsVa36Cgpd8r0DuOGtFsOaLj5zBrgrgCDRlr
yQVOHGR7nbV0SyCF088kveWX2xTrTjKyL/5u5jXfk8GFcFcGR8ssDiHYQFTQPTJn
JBlf6/IO4l+nVhm6E2rIKrRDJbNcX2dwKoOOvOHRco7SPHMPev0WTtVYNPYDxnLV
4Qwt2WpwC3zK9YVxbwajmVFC1bSpC4ZsWyTmt3Gm6AYDlemTH7inh0s4jmqepOEu
bVVm4asfmS+v8qCf9FVWZ7bYIc8R2KtqVXfUnUrahN3qDdBDXuSnoPRsgSgQe1ef
bKf8GH8waonacEdxSksGx9Dqi/hOYTqKYLH/fT+3QMxk893PHr2BveD2hMNVaRZB
05Rtr+hPpiZi3GtJACW3/tNTBq1Bb/S1/GkKjG7uGHRjGsXZlmjEW0NwoEDt+Y2L
u/k0XefxhruzaINKB3PzSn1TyQWRcJuT0RSFObvT1JImBP5YlMNEdfLVAtUwhfme
Z+58OZjR6urTeziTf/t3lenDr6huZnXccVRakFq3ubrqvFpn0Ps0ZXIBPAFQUf1b
gEDDoMqyFUL7SoFaqaKx1ZRrNnFUafx2pUZpraRlfCu6aZ7yKeXH5xvJFdzBqiwv
AaK5M4gxL9E+yFZqg/YnkS8NkKCTZUcLM9AkCfqLZ/rVnjsyosdrl/JNBAqsFWOs
Mu9z9AsQxNJdpeyyltFpSETINh9HXLIrl3dIRCj0orExrFzKRulCHfE/xvgyAcxv
C5ETEuEy8sK7lk2E5EBoLJhJsezScQAyES/RdfulmQTBjjZccJQJ5X9egRHuC5Cf
goymp44cqcwUTN2mW9oSwbi1ZqmkX9D8g+kAbCD12vd8D2kOumFPFjR4nHZ+XaDd
tswb1er+dWuwfr2edYxRyvS91scnLB7yDiNkpW+eArc7Tvar6WKxrcMMk9RRJpY3
pvDjRkAWn5hmX87JI9nYfN9+r7DSln6XVVcxJB8xW8Ab1UiGr8yR2Q6jHesQrdEE
TMriOZmsSjtQTi9lXL5gFRPF2keNUblLd0a9G6Jhy07htI1vPA5dbr6XOgCsPeeL
92SxVb9mWUv8CnwrZXyGLQ+r+S/wOMcRenTO5gzk+KPB1MM8FRQ7xTuLx5yEhUST
t4oW28/uDGejo8Fip4G1A1ZJa7xUOLHUYMIlhe4JCEPiA4LYK4YgBXzwPQMiWoUd
LYOQE9lxHyxGjCApEzYg0uEukWAy9WlmVwGn7jFY3eeHFLm0Jgyfo6XGVoZWSBqh
COk586AnPVWJrMv8HQpLNHIbQO8KkM6H4HJgVQtrfi49UfYgbj0ZZYn96cv2k5gc
rIR0EXCjIirAMBaSMlA4saAW8p11HKC8JlpUst1J7nMxoX7Fmb2onbyZERksGIl7
Z/0U9yVg3jbRfEJxzy4zKgo26wa1ADn1VZhwcExqUJSNd3GyJ/V7F18//vSMZxQM
fFadGX8xuJhQjskdUvX7n0t52+18H7tWwVAz+aY8XPkoYfOwmGEkA0PWvbw1fw6j
uI6phHH+rEXWQhuvkyz3b8IdCrrgOngYJrbdM65b96/aqNLTGUQoC6RBhdUvmdmV
CdU1eWQhDlnAyZkETtK2v5MCz+v59seHeDqHisijmwvQXUXYdvmbvqNXk3dZSRza
ezcvN3Divr3UiOG7tC/wfSW75ukVTp4KoSDHMtmOxRSm8aa7lLlLS6rafwCdjvC2
eVAWLt6swLGnw3L0CM6kmcwZrUdk2ASRUuqT5KrhRVd6bWI3PjSJUnmEA7ElQrJi
DL/lNWZeBgSLH6U3nuOjiaVAQEacHNyQiQH/3jEzClw9diF7Mmn/DfqZVyVdyi9l
1iD2SJCqRlaoh0jGNXJh5Cm75c6jPakE0AeFmr5GI34b9jAlk2QW0JG2uH39AzZn
UAxfXAJowZ9cE1GC40GY/WII405XszJUFwE5VxoVhlpn5a0kXqbFYRrjqxl9Ni6X
9yLOSjwmKBoFB3iW+JFYz0ioQMcHdKe1wmJi1ac18W59r+YODXIQcLpm+Z7lIS3E
7UBa3JmXQUUb8FqcnHHFp67kJy79CuXikRhaAT1RXjZwWMC5p5sKTXWh3/76eGx1
SQz9+DUPIZBTdGpHmafEAft/GeeZKOylowJwpAxg/3X823hddVe+w3g5X8OpjsAS
1GzD1UKZ13boLz7t/4IDurL26cyxVZ7cA7RaprsSYn1vlRuvPUOtNrsz2aHMc9lr
Ir+MpLPkqDKmsk4Xooy+qqNgDu2OzAY2+ChlQVVM3RQaHiTS5TzxZzzTQ/sI1fwl
Z6WtXWACjsvDoQWSg50AvjT5BItrcgBxsz6vV2FuRyYDB/BJWVgSl6DXev22qNyg
bSvRmO/JrEynjtK8zEEBwyog2yg2N7PebD4I7UJXoW9Z9b5qA2gpFWYUbmW95Qpg
3M1aawCuW0/qn6/JUfPU6s9Wo5igWNdt6rCR1Ix2oqANzDRGgqaKSkrj38Bjl2Hq
l64cLI2Rv/pse2W+rUEu9K+L1dIvTXO1RGPx9WZ1RCmI7hiujO0PamSWl723SjSY
19229IcySTiu+7bH9opuFJNFcCOqCGcpHRYjsQvbyM5Wu9Mkmlnn2NqtUhvbcJ1w
CFHm92VH/kG07XsQ/aiIPghChSSLCHDk2wXLhn8jTlJGeFKSIPhHVvWHPZ7q0Uvv
oiDEp4GtCgC+37Cw8yBam8YtAmblXbp7odWmRhbySNbQ5u363biAbq0RngtpgDNN
WUWiT34Fn9QlCwcDMKwc/GN1pgrIa6jMBWMGbyjX8xnBM668pgCQH0Wk7tq6xIOx
LI2FHVvuKXbCguCHOTt3YvycU9FgMHzBxk5Q0mF9ISluHfxaPO2oOhJOgU2Cv9uf
Nb3MlklJkY8A66tGTyiGajctIHLOOeXKm8hiU5mmCxL7lvhb//+xhweO4sEZH2uW
5WOIXGkvGV0xBycXcUowBPhlVa5vYSGwtItAh/coq4QYS4iEBlMPUGp5KlQSV4fA
o1piaP2o5wtBaXqSpZGj5sJUPw5N8b7Qh0/n7/mZ2+miuNg144f1XvvM317Qqsfs
OVo9EGc/vAnppy7iLyeX0CR8oyATsDFqPjx71PVAcfsUpT0o71n06ohbMNwtfFbR
yMDjR93DDJ/+zZHJwLSn186Dd3y8BkJohf90RNu98yfYCOjlbtpP64LTymQDbHWw
mEeRLPIPNr0s3VnixyOhHE076NOI9jqr5V/eNPMkBKK0lx/nGX1nAe+WcXh6v1rD
tEqKAD00kLYLShKddM6ZHMZpdgLLWhMIl0x0X6NaET/K5iod3hhuZlfjX6yslh77
wzBhHs90Hx9cL+KoQbnkikv8KxxRGnJaRe5dhkL2t2Cvh/3lJnoj2mXEDFpw57Ct
GxJO7uJ1WbrGvPfdZjTDvUOynTyqug6159kpJZzSH12l14vd+lRQ7GucTN9jUCzB
tes0WJOHDR105NSgTJ//dIZx1WNXUmnfFL5c8Erro9frbhY7HfztbjKJjJTTDp1d
0aWl8Mhd2044SPOpWIWhvEvexnGAeE4NHNEYowBfmzcOqZlE/wCOV4031sFdb5Ne
xQNwZmjv1mrArIoVILirMcVjBjC5mF94N02FZXnwTgkMAFDyhaE0zjIqNEL8Q21d
7P+h4BvYSUTw8CoTq5MS8ZRkK2aOPkIfSwbwIh21GnxU8Qo0IE6rotYF2DHbZuWC
rmVZroertd6j/c79A5CBQSfws3tToqc1gtBPHNEG03V/9xKCVifPEUGlFRNIPu4+
LWk6jUwXRgkr6VW231O4xAcw7mE2KkxDXmyhJpwaMt02TjBVe4MDv65kfG/Gf9+k
WcIjb1vNXZa+XDWr0lopjsMJA1oQq8nKXlHoloLIhEx2UfyZfkqvnHBI8A56Mm0x
NXMitEsf5HQdfCUBl9ynNLuHFmFHuAxuN2/27mr+n0q3Cgn2ko/KOYn0lTn6FGF5
UXlFyVeUed0AhI9ewZlbG81Yv/OMVF9X2nTlBx0ZGFx0nHMRz+4wF8SzZitJBW9B
n3TBmY/Xwwo1e+4P7p+lRs5tyETIB/lLftCf7vmumX7BYhWUyevVJWIFLpwYUOoc
UkEmSk6Asxy9AUBxCsXYl7ViXXsKdxtTtoiOyETqMTa8hG+Y46YrwA+ufPnPdPe+
dzfBlF6DOEz3cbVfmDBnUGPT/3rLd02mgAhJajS0/kbQsnke+gwwi2QwZKo0m5Kz
ZWo1mE07nAES//ijuN+Ij0Q92d6bNkegEhITkqxaGzthxj4stYJjy6jTAVSVW90d
Iog1I6/3t++swhnhM/SQKGdatQmuNguyaTa+BRb+HwRu+KJd0Sx+/mphtbuolmoA
Kb7vatIzmhwglEK/rkFWDF2aiLb2mcbVJyj7D7+ZG7vjwnI8f4woLX4+OT76+Tip
/XlRTjuOYf+OqbuSbrEh3KMRm9uYfGsUSUpnWig6ECy33bWFP/B5+RS8UTjU/28v
GVE0OXnhaL4Km69PXyDq18zTgsDrpxGYyTPFpaIruBu8C8kDRWnUXcEJA3aPgyH7
ZbQG4RdueU4JMODfPpV0ccomfwqrd6AAgu8Qe0NpCrLjLT14hXbfl2xHpQIB/t2l
ERYuXCpxIVeLk8MCxGToDZ1pAq/mSzdkWAOSKYkCGtwCSXZYN2KXDIUvJmc45atS
zcp/LaR/nIwgeeeAGT2aKQhn2h1XCcnO6CWuRlTlLBBSLy6gB6DZ+26NJkSw5ZPk
O7PHdm5mFNStm+XcRgMmgvVqdiLwTdC4WXq1EXCiLmIP0Iu89WBkF8j1NM7kZakQ
hhe16JLttihRUW89J8XNJiVNU82ZVuZN2AckyaTqZYgCw9aczEDVyHcX7mgWegwL
SlE8nNUbRkDaFNx7zM36elF+q41/JT7ijFUgio9Ib2WQWp7ZiokiZGgQoigwIesq
l8gXN7L3AUrrVwALJOcry3/RGa9cQ7BTqVogKo5jF+mV/jT7YTYY8vCqSR2c6MVm
1f6CUSnPE2SJM4qNgrqtJff6SC95lbqULNzEtt0Xr42XvZ6nhw21KjIeyjx0e+6L
p5KA5rQ2a46O5UeDWRlgEmrFh6G1050Z26zLJ+zalh3ZuNo8IQ5wffRodFdkUIpr
GSl5XU6jcVGqW+1S+LHZTU5A9j3lyTofG8aGXyZ8jYSxrx3RpHYcwlESI+V0PYuo
lGDPqRUh8q3FENqx9tKDLikPTJ0HplFCqOp3FCwKamF3gpkVHtmcRSPWCP5mspGM
BYrLDa8xtSWPtH8yMBOFGshTpMdjSMOirP1oGxGPyEQiGZmWmhQeA3Tf8gvjaxSE
RhkdBmmgUODYIzmZU9cb2m2LcLWIxdv+wA6XtcRCn60JSxASRHAibPyJSnGoLQAE
J1R2tTEx/3ifDUK9pf+JHZSoAz27cMZuvQkupBCtFACPBOTuUeX1jkdN7k28W4o9
lyN9yxGOBc7FA3nVgqLGkLKso/g7N944FYT0pj4rRpolMI/HOSyejEa5HI87gM1j
EkAepclDbv58MkqwdSS7XhO1k/C0a5PaG7ZvchtK+LvxATlaBlYnDeVQm/ua0I33
TBP3hz3tEZrh6kU1mMJ8RzTZUOkOsk4LqCWe4z+XqloCseEHtc0MpkDd1MJk6fZZ
gwJCJMr8zetOX0rRN8bDyuoMF/eslhgO1M12o3wF5YifK0bcmp5BmOQGjGSHgcr2
zNb6cOLaNw1NFhmZD92/l9utu7jWZDJ6MdZFXCJIUaAypWXyEpNlQPIumOlUslhY
prdvwn6sw7VY6MwlVnynZ/p5tj3rhlhpzBFhSZkOQHzND/j228USBv1uOOCVLhYw
0ZvAS6XzPdaoZL32N7Xs0USQZ0AbftWgCHbw00xBtF01zKl8SRNUr+ldjxV3SDJ5
VAkjQWfD2AxWHyQ3fFP6xtZXfDXLJJhlEexnzCfcXotToDdp0bYcxKxotGmZKEi2
/RO+UBQwalK6vsxZeu80RQqX1duoW5eTO/MauQZHTVvXfMOr00vXQ1nMUci1xmu9
IBoIcncK9PTF8UxTJn5sA42qemIsu/3NaYnAihSRyXpKeAGtieG+AEKW3PKdmjUb
2aYu1U+kWwA4vt+EdmdtGoWDmMGKpsP0ga846JyJLkGbsZ5ZGcfmPKHkc4RUMQIu
sU8LmDt4zRzLi+W+MQnk+TVBnIwtU3OMI02+XdWkeKGWfCPKdYqPzZ/Dw+Wrt1SO
pQIO3T4UTq+yOoOU0FUn9uo9pyAq5bp2rErhxj+ua8Tfr1vKw5AXjmeLXK1QXanF
XcshfznkENPjd9NQ5qz6BY+XYWNSTshs+NStwy8N8OC9zVcZnE73gzvXgTS08vLT
BEr1kk4Xqk8vmrdv8ZsT8jvpAo3G9xosPs0Ye9tH+c/86gPnPdnnCT+u24bz3Ymi
wuwzHXYSsgnVeRfLbWUNL0gU0AkhC1lNmt/xH6d6cEEvQBZ+8x8cybjjbuwK49jI
Jxag/x+Q7sZCknprgKx8M6CJEqa/M8sA3cdnwuTma1y4TJ3hut7+xJAo6YAH2DJH
ek8pzh10u9RarArQcomEGp66Q6UHjpzZW/SGgTQSYBfQK42mCX/fPIF+TEshTxmx
jKwI0YlGBAPQPOYZPR2DB6GNqFTKZq0BWyIFGOkVzTTswV1AnOuZs9Ltn3waDqqJ
U+MadQQG7nJfeAn00B0CceMwQ7DFx20bYlk6g4RAJPhw+uE9DtcI7BuAjMxlPQ6U
aIVElbxnrxudZRd6RQiR2TMGBtn6Fb0SQgMNM6tslPmPmoPnrPVdFQXPIPsnvxDr
CKE+MsMmQR43srhRQbN/qXRRzRhdU3rbl/uRJ8C/Cj4bKpWr6VLvkxuQX7qJ80rc
iVuGkBSBWpMO7YSUw/r62nQNx9cI2KWbjx3MFeLjgQ4TT5IKF2ZNKYIDmkwwDjkl
yf4qEDvE2XD6W0kXZO8HxFyDrJSndSg+7it2AiKW5NYCP/dgtluHujFMlRwOScyG
Olh9yzpFkr0yzx8pqpedGzS6lqEgFfo3c3/6apqslYNfO//4ljvPoK0yRmcPLYYN
Qt1UeEWfpOoaqAcmcChciyFpzFkTrsE+9mb695YkHDyJTlyXlIWUgxqtbSLBK/y+
P4C+qbzeCoxleA9IaStUqZBTV9YPoCMpx/kN+Lcgh6YvvC5VuZ0CDIlb98qpGo5F
NOR5VjrWoiRLhVqpA9sv+nkGEXeCYSMIhoZfLFyIW1d/3fgjgar+AwzeA/fAHhC7
kVj0t6XwUb4Ni57353fuY0AcPn52J1SXBx6qZikbj3g9f59zK43ogBifojlRzOYX
kAd4Mib6IXdUq76bIOr8VeAvMKvfzw7v/ld9Fkq/tpDyV7pcBO1js0/7/92+yeH2
DSmiuRBUZig5j7JjZB+VrzOlugYB+oYUVHqG8vNzWLU0zZAKQKlhkgr/zR5EZ05n
ctJXtZQo3guYaeV1YIL4N1vXJNt4MA0v0qjVSmM75M/9fSNldlCf1/GORDPAPLxe
yjwzYRaQ6RPs2HVLJVxgtsfoxGasxrhbmSlO/LF4gE1I2Y4kfqTgAsbRe8rhWFmI
toOoets5fO2XIMvcmigjN1CLVrkSWB1aqyFCE45wnyhJx60f8SjIS/GVxuOYfcnb
4Uj0NhrvKO1FuOD+RWVhzEJoJ6VYoc4rCHm8TDcUmPUahpEkuB5RhEWxBoStCej6
0Yx7iTuTijrqPpxX7kGRzynmwKYVj0BDZ8BOyMwUPPPkt9MOBB0j91A/VJCOUfhS
1QrDi3ydVFrEZ5wCBsWbMKEFEVhPfR4QvOFjOxneOOWQgDgA87gX0wVKd615FAjG
WNDsj1HY6ByB0pJ0EghyplHY+jTqo1zOWd0kHqcxX2oM6qG1EERiFo8EN8/UeMBo
9+P2RTV46BPtEVQpIIxRO40aoickd0CJPcO8EjegLQlTCuJep6QT944la0eUpImV
zNE8GcY+1Ym9MJFxrGWmZFyzaP1df2Oclwk8hznn6MHrI5QbJpyafSPPWYRbX8J9
njf4KI9hJokLvhjITd5OeEsuEdpWJYS52PByXp0s5GHJFZg1c5ViooCVawc3rct0
xE7DMVkEzhClF3DgC6jOzuyD/aiUBfQTzR/giwNOAaZgcKGmLljFaEVFWcszuIJE
ysLoqzqjSpAU3K8+6QRaysLsKZp9T6dQLON18UrJDSLGNvofqBoD/ZKIPLgO5M4N
RhGg78VOX/Ep6FlzY31OaknNlaBwKEYDfzD3AYJQQTp0VXaENoQsJTUXBoxUYAm4
58AS/rTpvjG27YnxFqZ1JbpMEmXuuo3FRh+hwY2Vh6JqLZ2+1wxZ+WH6TxdVzdNQ
Q8J9ImfNwA/b7vc0rvLefZWaaGJ33u0xRwDyP/WNCZtLpXzNgEb6FTiK1emoYgDl
R9a8F1cYlIEyq9qaJa2S9s4noy/iL7+tsFoQ/Fhyfn7t99ceQkVaDAtdldkhIzw9
mcpAHdk5SXcTjOO7uKXiTAE5VeID/rN4nCfbJxSCDd5P8P1RWGvztxu6/MQOxwBL
yCCcQZAVbSbWAoDvVkRbQIRmc3PKf3apQorLV2Hj8p+HPlNWJkc8LPBy5hLmeNSG
vFE+FYk3LiEyXWYIqFOiQ3C/0xnP6+fe8Qsy8cL75QLBtOpsz8WHbazFdFttBGDC
lC0LcNSD/NrIW/TPg4fYCmfjpI2K1qv3hQqwlGLcEnKn8vcLte+Pdlzg8UrCD8ew
PvfXL5BPucwMRUyKbGL1R1eL1iKOU3ogXot0DqA+7cfO4lQVc2jIC9NO1EowANZf
R/f6MBroJG7u605VFj0l3nlP2OG3OwJUigwUkB7IyIUfdCdJtExYXLcwOYg3IGPc
Zq1NaGyD974Fmw7yRa8LbZNz8r5Speu3DpZzfxrxcXETsBNW+ZW47l79BrlFlnHf
PLRc+HAHxuHzzgld1Yd58XZEmtDR974jSWrMaawqRQCCJTGHLhyavScwm5Xm6RN2
so3cUV3yCMUN1neg6pTzAVi+AaOqODGM8JuGM9nvchzgRGVU1K9aWv3Kyy+fr+b5
TIa5EFuN8ZDfufWpT0uFXLyQ1lsU+P2q/JGKgaOoYVSqVpGnnh0BFUjKT2+bnMG8
quLRG/Lwki9JiCMdFkUS8AwcdFj4qvEcdSnA/FkoXF2g0V3KXxH++FdMtTKWNuGs
8sfBCKnSTowag22nuJaLGbaykavsYsLqz5MQQk2yD+TcOK/Dmbdad7jPgAxUfbKo
1Rr+3xbLQiObLwCiaZt4JEGDsRniYAb9vj/vigiq1PBcCXwJD8e6+a4QjT5BxAiE
3i4OE9lF+9Qp66BetZF7qQSah2yqBc+R1koRMb8AObhXIf+u83UcQn06nTPwvNFk
v7Ak5aYPfpPIQ9NrzTjDxRDqvqJjiT4y4WjNGm5r3YuGsyAVm40qfRqERtUloul9
P0lHnQrdptJrAHYmIV/qq8g+crRrISKB64Q299Emv5oaxnOaq8cNHlZrHLnit0ZU
R8E6xx6QDqPMCxroNlGoPQ50ezXR223JYr/YM2ZB5ncvuqwyPBQCghdSpbB+m5pl
4+vwHJrXAB9B5Ar746FHcviEOHQ1OOUmVWa7ogIRW5mvqiA7qwl3M4MjgZ5inXMX
BJ50EgOBUw+Jx2NkvZ1P9v0FMnmP2mJYTegvoG1cUHqDexB3A0eM3OWMYnMf8F0h
TmxunGCnoPwWKplvR1mp1tnLszEnePYB/s8Olo+L6a2fAKzMNALQKahVDS+RpGZg
DRKz+kwyCey/r4jk0UIEKVA1bSSU98OyutaY01NVNetIidPB/ChYx1QB4b934/OL
BA7UIZ+dVTFmOHKKer/How+zqraRqxiRunb9Kmj54OC+hrTa97I3bS8woUN5G7Kn
z6GYN1HVdOtPS5xDESihvP20C/yty3hrO3mGNQYH9D3eQUrOZCgWHr9mM2wEwszd
nQo7t18Qkq6d6ASq6F92lLLyQtmVwTlKqzC9zSOIO7k9DLYZTNSCjmGRVoZKO9wT
xsSeZhRntS/cGa8teda5RmPtYWUmQ7qGcF5rh0aVvQMykofUw0MMgkcgHr7n8IPZ
qljgFb9JXWmTrwZqbQ5eIUd+gpAMZ0xJwjP5AN919HKsGUCoGmwRJJjFyb9cb66i
4xy+R2vKT52OqrRsWoVs0UbIxTh3OBP1bMcAQ0Qz4ICjY+qxoT/bqKJxl8Ho9GXZ
AGvNQdmWmDvm5VkVS5VtZDfxrpfyh5U3Uaa0gJrrSiJ7tFfTJalEq9LarPX746k8
i80YLqE7Gkd6NP+pu4fo8qGGIu1OFnC8NlT9QpVxKSLS22W+x8IS/QA4VT/RPN7+
IYo2Q8zUr5Q9nO0UtI66iXUiiPTuP3lJsI7lBPxs9xU3ebgeq5qt+CIfbVmVH7v/
ImE8JxJ4UtsJ0YZzyNC0/7Ae3dIem/XAkUQ5PGVoI/zSFFc6UQhi6q7SGOwIlFXc
KyZwa/ScwUcx+OMb+eT5SxWE1ooAmVELKy9jDuVgR67aDLYI0DT6fR8dxK+tveo4
UCo02G0f+xEFx4tLg5RcHNFdsp0VWEgS41YOFLO0rfSjfU1NXvOzD/m1DRf4SGqR
yR8P/4/F0NTnnPntkn6Rt5R+ikGp9rXDWYO0a+WPPHXytDv9d2ucj8Y7Gdj2yQ6y
pu5ntgTQG90f0HpdsTw4dw+4gOfNbpQYtB8Fkcp7GCOi76+SudkPMX6n3ZNy7keY
mukW3SAA/7OgmYkSKsmYDhMbhZY3EWIj9xrrkYawE6w8y77rPbOYABp0QPICNmDe
evy9Xgh4QO1OeSU1Zcl58bSfEFTyrTa0kpJ21/heGjkLeInW67xz4AZh9Nw3yUGI
LO9lmYCRmhJmhru6V3VjjRXCwor4rNJio1/x5ItcXhe7Ikz/xvRfn3/cdX78rniW
MCc0M1f8H/HNjxhnFTF6hs3RC4wJCaZP/wZIWXOWbYyAjSDrjvQyrWawyc0Ww2tc
+9XhkkGYFl0KZXbxd0r4h/DDvsyeEvSoO7HHdbjhN3WbKBI6T4wPW6AJO1OiWqQF
kQWXvDKY35RNErw4dYnXU8Z/NajPoq21d3tWIbzeRqG7C8scEtq6Qz/8cQDowX6U
nj5JOf0AwW1lqxBXpN4Z2/4D1+Bn4Ybye4bKFI2EhHZ2LzPszZF2jtoFIkdh/Nqi
Hu2iIPqhsEeD48JYsnuhnNBf3NNupulk2T0vmrXV+5/kv0g47I3cMdN57rIU6yDZ
KYLHlQDpzbsT7cOttHpS8NZaHBEsZNPRVIgYJYN68rQEe7JKUyvKexd8LlKP1j6E
SY8ytFJic6wnHgKS6rC83zT2leQKpIbBr1e0cWn4SF0hgfeZ5EnKn8X6iXSefqJx
jQTcdjD4Y2N0tGOex2lliefh+ROgpC/MmVcUi3/+2myp5TtEYxJxDjVjJ75upDjx
m8qb6byfVOyvtQqop5eHWD6bWXlPZo9uCyJXqf63q/kV3PB4u9CuRWlIdclVDegb
OOZsXn49gB0743HxNJq/SqxuBwCvVQJazR/QySoCB+9TODtwzc3ddC0ja7ujmZzS
8ojMRhv2DRGqdPIFSwbrJQ9MNSD3VUAvhEsbJ2NrU/jH6k/7khlFYeGzS102tvU9
3+H3qM8TTW40HhCKxK1t+XHpCtZvyW2fEcyX8GtR9/bgCK+2ofsNxR8VRLzjeskJ
q2D4cynugTXJwogcv0CDORc+R00bMYbafP+JKEPfr1bSI894+iYnZk1z5icVioWe
I4k0HHJ7GQ6k/fdr4QBnmvcRM/mFJ7bAb8w4OHtTN1qpuMYmuMlOS7u0NtWhhI0s
TeJroKDVpv/9xabirsnWT2qyogkllePCf35USSGH7YAnq6RxrGkbQspgiEfU/At2
00KxABLAzcXYZvI0twg392XuiiEz1j+SLORrYnhOhapORGb9QQflyPP28NhbkNRE
+X/eIu9w8qawzFIF+vRjxztYED/M7ol+083XllFZwWdXGZttSxpIVwg1TWLKbfK2
tvuJx0+a0DN8Nlg8ByIrJtmeox0HIb8RTfWDHP7VOvus9yHFy5+Wq28h/ZYjEScH
UZgvq1ds3BT9I8ThWMJUh72U5JfPJAliBvNQblY0lpl/jDUNqHioxccEINxCUVaX
f6QZcupISbxKpHYGb+Yk7I7/SSlZcZWXyA1jo3P4uUAhmtBGDMf7kYv/7AJAv4c7
rVnRSvaPxTlSO7f8xKsI9NMT9zQJQrRLZLD+pFvOEVjwDEIgphX4BuuJteIdyCmL
M3XKBKMVpiF04HL0GEdFATU1wUcv/m3Sr+bdTCv11V8CWNKrS9YT7inI5lqHe8zA
Qy6S082JaX4YusK0Af1OO0KqFKy5U3pwYV2j4vG2fjOhjJqmQJzS3ebrDA3QfEZU
5Rdfp9dPi0/OhA2PBzSsnrvTmEVMrZJbeTpRZYhxuDCH/7t1B83UEKdtHjuj/uHU
+GQyh1DoA4fNBd1iy4CuhF3vKFMO5Sd1BS1U8JtJhnWUkia/FKzKQIiQR9vs11ny
GZYJ246CnUu7/0rj5GirU1B/Gf0G3y2BcJhZFoxSpiPQQx/L//s0TSGcvGMNBjBE
AG3pW/hqNN95Lo6+UiLJA1l06+M+1aHEwVv7eiM/hki0dEp27ochdUpbaRrV6BHe
sGR2K3470bhNaB423wQoiIzlT4bJH5T9tw8ZE/fjGXL1j6FjZ4sHdLEwWbkFni3Z
6hPhuSn3TQG481zONQFB+XqVwAeMtMiF4dkPy1WIllrlo/ssp+8g0+uMod8WYDCo
2I7emMqJR3eMmEZgjDmtf01u2riTIsBVZXoOhBoyPiFaQVC6pL7z2+XTlVkVhXHj
QH9wTEud+pbmI5T43uJvIiEOthKCUpqQYufmzmmxaTQBcGJ7JIyEUl3iKtS0Gq2K
4uMKKoiMP3LH+eFURrsZ06dxvAYJY2DgoqJzXiHFU1MdWPAC1VeSeAZP87fss90W
ganJRh37cDxAm8c31ZnXm/2GRqACsj2UHiduSApMRwBZRaS6P//0JTU6jYK1UOa4
xI2WwK0Ol4aMKnDvSytFOOmXJ7h6aguf5L64bw/RKUDjFfwMPFC4DU/yyj8kDtmQ
h1E1sIwdI+7L0Go3ysbBV1zUT72O1OvJ9sKMdSGj23dDN9aY3u1CGJZ+gYbTVSSW
eKVVLHMkkDWl8q20SNBuz4MMoNt9mWcnLXv/28akqV6g/4LOkEw7+UYiifIAdkMH
uBfQbakm96KFI+GNTf/yPcvD8oOe5qhz7wazZ2X74nZA/M6i7n5HutYQZNvaEzxR
0pobXkY1BPCUpOVKgPKnfrbctWAIMounFkdTmWpz65fTGV/BOugE70fhbVQTgGy6
7EapgI0W4drdFYClh5OUMX18FO/qCmAcq12o+woa5eY3j3lMep5sk1R/GhXP7BXM
HrEECGkoQotUv9dTMAqGfug/xmLlObyOm6Xp0nBkB+DJmUbx2hbVHOV5ZwPKk0T0
aa9imJckyoeHd0GwuE5TDUxUMWF5TvFDDjfwh7e4dxGLRykj4d6xbvBmAXXCkCFS
EYnCBxEeGzaQ1tFhEyjLnX9B/8bzPrhOEIgvEaS20+RZeaNfWx1RDmlIlqM392o/
jxvHmgL9+hDpR4AmcEEvTuw6iH06/Ue9NDNS0EQeBncL4yUQu5u1BJkGTLbzvtvV
QOxCzKBy9Lt2BQh4q9UVlErEXi5NRvm5sgAd1I1g2+RSeF0ywmttSpTrLLbH1agm
1T81skBln43enxugHNGTgba8fY9q2xyPwTlEhZA6vA7PZaN1lqX/SjKUFSTTZpTF
/bTFf4Q/g0b4ZcfL6usvED769yYtdwUrB6DcbXKz6EfZvLHyaS8U9Ik0yFKNf5da
xtwWRcHq8OrDHwdTA4AS8/kDixcdWI0xIzESem+4Rgu3uJBBnSqT6g0BeUS04hFl
b5tRdCGZbe6sH+SUuFP9iA9OL8odM1MvHVhDnzQpC6SePubHQGSRtBjGZwC/4T8t
gOm4aTS3yKAWGIW4JqZqrfIc0daLB4UFXfk5kGq8W8izUnKGaXj1L3AHoshw9tU/
oliVHkT5K/DpSs9kiBbh5bWPmK77SNAtInY8jXHCCKdnuXjhgUnMvE+hY9wjujW2
32ViQWUAprk8osdDsObSVlZEUEfFBnIGAMXZWoYp/ewe+UaxW9819QSd7FAaY1Fh
m0q7eRIP4fpLoFJWMqEkzuPYfiAw8lbSF7KtBG60C9xkwF3jwgZ9G7f+Kfs3Meus
agUPZXBVjCHYM7fpfFNj3rstfjRzZBt3lQcMGiqgd9PA/OmhnP7T5Bjoa5zY279g
6rTjf5MzZYdHFBEEEIEXxbuaxICwusvZcxFtELbL2iB6TpizBKRkYxjxNNWefry3
iUUj+tN14C0xiEuieLqpCYPPIMvg7nQHXxZWihLDkBPctSO1rsytVykUp/0Ha2du
f9+g3VuZUScsLftuG3qKuV28so2HnRFIRf9UXRB9o0rt79B0rUGJGjve71Mf5bSF
QrjWFFQpp7I46eeq1o2kDK1C1qcFqoc/+Nvcm1D9RMHxEMmAHQhVi/WSGIsjEHjk
HUgLqTn1H7ZNdBesMmwlQdxTL8LAinVWD0vka28xK3Z3LmQe4L6/IChE4+E0Bf8F
wl6d0rzlpHJqa+kOinFOn/zp0IufQMAnmppvY3adQ2IouEV/KX4dow4EYCjtMXY4
YEDYEp6lMcuKc2vzp+nUE7oWFT/LYz6WQt4w/4YvCqUX2/7qaZHEJITVCI7NPyhf
HsGpU4eOnvsrVn3jyWoRgCQD0vsmb4mRtcRQ9AuW7Kf73q/pth3rw6GSgGKk/E0A
lJfmpQ1H63kuHTr3J1ylDTcXi4lG10i515TQQvZDdvb//yBIHJlaJCtrxPuI0Dm9
lqC7/EnjSPb9mrpqxkUlvsHlYJcnPMyNYSm6t9j8oFv4zrmIMa0dzxF8J1bKmAZs
Zeema4Al6qyhECRgesN+EQ4gys9VvhjWCg06g65u/h/7LkJz9S9IBmV7Dx48xawn
XW5aZb7TO/Ublay8lBE/RXaR57WsAi55dnVvAMdY2srZm0t26SrzLTFhPW+NBhlE
YcNZxDLHQ50TsUxvlo55gU/+Bh9/b6IM6rrHpmQrDHTVYtUge2h2t247bALhGQML
xCzC8A13B7PnM7Xfx7Unl8JqXMjsZ7ZNKlavofF7AYOHClwx49p8s09uCMuwzOz2
j5e68F/50EfLgnBs79nPI0Fb7qWZb8afxZtcrHFu6DTBBIOpYuA5AyzJyJm8nDdQ
Ecu0qP3BrNLsqVmQtz2XCu+2SBsBHAIkLIBWWVTm1ZDjMXz73m89KgfSRN4iW5ie
ZAC5r3oOOup4F5J08qGUF5LWegxQRNd4OqundA8IezIPSH8L1Est+CDcn1c0YIOi
UcyWmjkgDdN1oYHDnuk2CBR2v7QdOWRA3LcVjQQgD6sRLQuFrmzpegkk4CZP8gGq
x4JbAZOts4/eWMAMBAqEcOTYFmClNHi/Hadw1+IYbF4+hLFO4tGjGNBv3i+sC8TY
YXmPM+nIZAUF4WpFnB+kxBcxnDoVIK9j1ibfWOHivY9IyzAe/ORBreI40Ma3Xi0D
cbQQqgJvNPPXNWcCapwmATytvDzWLz8ppZ0d58dn+F3ME0Aoupc7q3WCWnSE/6j2
XnLHbUckaQZiNfmZSWoHWa6a1FQ6Paqn+kJcJaLY6URBcP/BqoG5/lXS2LP00UGV
uTaLeZxdKflE2VRHouDLLBQNGXfVbk+ZUI3RrDtqTVTygKIVENrXpmAS3tk1cb99
+mbCDcexekRsJT5wHrnM77HYji0f17yS5eQhejvhu98CUCAznqET8+GyiOA6BHX7
DUsSkqYw85iddIJJYgclOASqWuxL+Y7+3JUn5rEPbXk+mFjaJ0goINsP4ODtbkh3
3wlF7THbDsBUGfTZQ989KEJ5/D2I7DKY+FJF8II2kvC1g5ryFoDiHMWfUkhrWnml
E5s5kAEYuenjuRKv8sL/2/Gqh/+735JUr4ScC97h2X24ItIFvWdakFvlkLiY/9r4
pyugS9FGyZsmishx7VVghGpX6XeJ5J9swE/rPR2PkTHZxo4lPjpqFZec4qA3wnfR
Wc7STtqON53ZcQVdD0WVGDnwK4BovArjNjPIUviwORausWcyxYf1rHD9m45d3wf8
jDcXnSlR/QC6rZovGeGi5kIUG7742Ec13fJpbet6NhqnJ5pMQzeltAZESoI0Afar
HpPinkDyJ78dz/ZLJJBgm99PHjf+rmDy7tf27AEK/avt7fOzui4vTIhWHh978P61
Een41ir5BeeC5+h1fZgwifrQ6wonXMgZZelwHKZmc3qoTNwyq76+ZLg3fNQicyxF
fAn+J6M/H4HxEEhMeKoGtbDcsyilCld1KFwfT5bwshtOxjwM5yBXOxMfnRpToOX7
Uim9qjXauSNc4BDB/Z8oWM+Z9Fp/8pBOaVw+kcPOLYRidnKPBvACgEo3hyRnFXvJ
/pSQQ5eOuZq5Ix7GRUY5RVoL2LARLXM2hY87A/0P3txnFQnZIOQcyeAYn1jC7/D3
VpEaamxAAF8V3QaYqaatbgVEDCq6w4VSjOC72XTcN4qmXXPt4CL3rWDDlHhT9PmC
g1e7lSQAvCrLhUYDideAbAyrNk7ayWcpYczNp7CjKQs08qRT+aGNVtIK8VJHcjgu
U7KbMiEq1vfFSvlmAal530T3VnCHak5Cf8dy7C/U/jc/qvRrr+7bHqYiPQ4eHwK+
NMpKa3zWk4ZPJgYe3LqYfIZEDIOYBxClJqmoOsCS+aJJrfMfWX0NFAexlVd4pTqa
twoKa8Xaa5lzGnxScO2IG9wMHtWKjsw5O07aXs5krCO2FQdiQCcbbhMpFNeqp07O
f44ap47kFrxe5fAlrMjZswPemtaOk3n97/1bBh+OibiXDNsZD2l6Fk1SQiklf1TS
jKw3/tHZryzTc0ANFRPacYWwTc0DueKFsOKzCIhCitS+WMTaw2o7Ts97w3bLMtxx
TuW2PFkDZsmmosdS+yVodv/nALG2sfVfQrtrOK+CsCy2oSbjvZDwLAQc1Ocszc5t
S7iHWgPNRkx/m8nk4Av55meAoZXPjeoD70EuZNVqOkAj6tSvbRNeBgXvUT1pkc+M
K3Tg6jwYMqELBRIuse6ThUZ7DkDTueSVP7qB+DtTlNHy99VvipqrCH2MBrXGTAHP
AvMWGS4ZUT+q4iiDK/jZE9NQRv77eXXkjghX6y0D07e00wxIlXhZf+AfwJFJpWxx
ATNFtgt1Xys0L54qZjqLRasS1bKKDtiidDFL54eOkJfAGtLUo1YsBPSoaATe2iNL
rWBpK4jr/9USJ2K3VooIG/+cLV1zjGvSPRO3h5LllP06ih3LRW9pHI2pXOyY12fF
L/mPihAx5ZcxAWZsMbSE/3HF6fcTI5xawXUtYnt1LblqGzViWwDdmUZOYUO6zzMO
OGcSQ07W1I1EBUpuPoIMdS4gxOA5xhZMzUkd9O7o+NlHPewGPN53ZMVhOc/s4Fl1
vAbPHhMl7oJrNq6ouBYXY4JgkLJ4QapidYzVWXn6Br2OQDdNojzAp2HE9UnfMiAW
qlal/85+s9rdoWPOs30zRXazt9y9CbaQ9tldI73Tm3EjPrW3rxHECSZIglhPOusA
RmsKkY4joAU5aYlK/S9EuNGyio7nYa5bbNNb71Jlg5AOBh3W16RMOvuJZZBryL7Z
p8YpI7kssdKwaw1nVUAMhVV1/X9pd0XwRLsLxacooxJtsZ+BO2LWAKiDzFCEsZsm
aoR/pm131O/Vfcp1jtv6sa8ly6tPzmAUqJpqq576kCNArkBeAvZmL9gmk8Cgyzw1
PLTATBNhxh6UGQ8IMJ/5/659mw1IuWQinUCxur7r6CHnnStAyiJmwOB3fajAgB1G
LNT8RZbqDOsmHHVVXCxGrcuO5N92xYwtt0+Z1KDeTU9NO/ws0HollmmYcaP7eqWx
naJOfNuKLoqYL8d1/o7EZRw08h8pgn7VlNIgmzxbRf7tM7xssoBiIOIXQrMBD7Dz
RQS5JUBZ3Mr/L4bMSuZdNuyXSUAb1hbyScW8WcNrQ94uD55xRY4RBTyrf6DW4H4A
nnhN+8h3/AIYPGmiiHrY1x+QAoJBGZLK4qnzGYDs19tZTjbNY7jhGFxQKq8fmiWh
hVnrhVxPd0n+vAydxy7qnt3FHMHanOaspfu+U9tJmkWGy34D/j0wC6MPbSCmFgSb
Ni1bpUj12LlZ6vyLdVkDnO8wHc8s8t2P3G0kldICHnYBGHSodRT19J0fh5+bjpm3
AXgoXvZtPY2m5BOBUW6XkzPfX022QOUA9wY5XTSn8W6heYHEh9Hf2R4dhCjKggHl
7P8OV09UZy+N5kgbompZtPi/drBL5es0ETPpfbX02vXg4UOZvE1gWXk7D3v3eTit
iCg6d5U9E4CqFdyw3/baNCaVA5zyPNKvbEXbrfxctsHfR4GrAWdy4AV4eXKnSbCl
krvruBY16+TrsK5rMEDCiX5yHW8rjPmxFlOksmxXtBQ2zpwjvg0yRPkv3LI8izH4
eBVYX7VcvTIUVfVuhnNNSJuFnDU7B806qDcnjmIO0UNDgS/SKPMJPoh3i/M57aS5
/ujlhWHrzqBd3Wu9MpM1l8aTCG7uC0VttoxFgacpQcJdl9puXSjw/3LKm2gJxleN
oFi4lON7ITVCc9qC4wdyKrkXy/NuLtHQVBzpVYrHvuTTVVPFeanS1HvJ+c1j4r7E
vUUS+kKf4sUyz7Ut8axTDxSQ7ZWzqE1sq8AwweBi8j0TgJQ7SfhduXolXnJa0zmk
DvfQXrmGIWIU17rScEiPF9nM7GUuRwASthSMatK11Srq6XbyqgoADo1TXlYpjIXw
sbT20t80Px4NE2FzTPoy1Kst2zwI1zkKyIoTfA98fjH/67taodNNlgSLPnI+E9zP
787Qz7LEAzc7NFRqy78eVokLKpdERIFtshohvKPobtwyf0NlgpGnMgjWGsOdL/lQ
gNT7BkASbCEm1knWq4ZfpmbFx5eFqHZFR8f+Fm8TzXxpIRJ5OsQGkKh/xK2+jn1r
ziVlFiy/3rHEfOr6TGZUuX7F13p7u3NPb2U10yMHudt1qH7t67GRe7Opa7g1yi9d
blXponaaZWpk3cp2ELNaVzQatTWMw+SF56BM7MhVyY/XLBFhWEvMYQhRpVUg+OON
YwGwG4CRJIOCzrurflXBdLDsw0nI9uQCQ9dKtIWAWbP4+WSAoDKwd6igsE9f5Uvt
T1GgrvGQrNmWIMTfls/D9DSYHyjiS8RWdnPb7VprIjpxNdJSfHA25n4aRCAx+HXl
Ied/Ys2/cwuRJidMxE9XkQh3yJ5+ATWap3jaQ9MmLjeMr824rdPo0biGt5VSt7vE
Qha5nL8PBRSe58B5/SYm7H/gJk2HWHIbQ1LKh/hLic2LkGQBmLZyg+y3G/XcmdR+
SFF559PtTZYn31TP8cOuS712q69NLVzJCbOZObSNZTyGP//8Jh00QIyuPPidwxhl
lBQCGWYZrlZUBDGU8fxcO+m4VyZOApZqauCh/FjhMztPTFNSHS08mvvPtLxJ95GX
bmdlw6KM6yGlTTJSnu1b23A8HCs9fkUwU/RLro5NXTAdxtWYW9aylymn8FFEwdVg
5MO94s/miy7lpHS+QvwxuZewDVNBeGYYAPVKkjtcODTqaI50aTlOPY/EGshzcApN
5e8kp930KxE4ZSXje1ItPtW7Z+ISgKCqrhwqzhwBJzYsSMQGiGIV+sni4x4q2MWP
1IZdZ3R9/3kvGGpDAuwSDe86XBzk+hiam1dtqxdFjD9aF7nu++659Ra1M3PAV0CW
QxzTqGfsD+HU85pmTLiiWLQ9fIHducw/eembKTsi64Gh5k7CThcYmpNAaj7qT1Yt
wpJPe1fj0MmgjlpJ9ysjRWv1oBXc6UgavfXNos64EkbdzCGa2H2YtgzczJLjkIhW
lmWU2oN3HBzBw3Gq3BUWUvahfFjO5KfEVQ2LyXM2a/P9FigplNqD6vm+KhBpqA2s
5qCOvVsHBo1YIBQjBmhDmMKXW1G0UvC3sydP5unW2XLKh01T4mlrMWq20/MG/W3n
YRDIsz6EUNx/6hPtn+YMpJjLaV/MtAcH4YV4jXMdw7RC/neMV8iNFelAJZ+vX+wC
+Gwh/vdEQVoOARgP1lxzQ46zQYZeOcCWxnNj8yTErSPzq/4aGUkCpwEdHmHSpqo0
yXBvwbD67v9qHFKqON8IPZR3llkPrxcETO+d3p4HZeKoLITRDwrLyHzZTGbzzek2
EoQz/7XOTx8CAF9TWzWBSRG4S+/xOoh7rGaTrWmZUk1CVTDkLPVKbQAHM0Wdm9Pk
+UKYt+Fj6bS8lYB1P1hEUYJpYNMfT7CMAh7zLHXXyMOgEimBnWtWEtJu88lxQNVv
ebezLFUAJdl07Pa5wJk8toaVGisyRSqahnJ5xQa6SLjg/HT7p2gF5SLs4QhOxYPB
MSHCsIGwV9wDVswMLiEs+uaOHONjA098POdtNozyIgLI8zXQ7JflibtOkmjAgBvn
6EVEIeumW74EKnQiMvubwis/kEc+LFbAw3wXUFtfMdG7wIpAgI/1tViSkObiMXOO
BN7OEqxkysmRpw6S+3gy3LZRvZ5bey6MyYrosJKaOS1s2q/y3W17Q6YskqAFLbQz
xwAT++OF9cTXLeDi+LEQknwpAgbTKUzMoqeiBuDMCGIzpr6SOl+7PphE32h/o0LV
uQE4LVq+1PVsmDOTK2AfDZcXpYQYl8X97vq+XdeSaEDykLxANtXKdtISVKTDJwrR
75YJSgiNFTmtmoi4GuhVPZVJKbvJnfESf3LTSeKNho0rP8pPn6RgjMjuSgT56Qgt
LyoS65lluY7PXSHg5h1li7mHmCBw0+XeJhBgxyZ1D2oZBvaAou9UlE9mtRAO6I8h
w05V47pkvJki7OWyuLaUeAXYEdycyPNWSk0jKwdhWPP0GMujK2ySFNFlNjlCoh2/
S14/LztyYABy2CwZjU/L68WP8hWoqckMklZEdB9k4RYUD3Jwd7To4GXgjDrd9xHk
k2Z737Cums9X7WoCGZc/qSlO4MmSHB1axrOjQCEs7Ji+t8WJNN6VZ70C59von5lq
nqf3igXMqRvOC05VM4jWNdcDqGpCy3hFzWafV7CNgOKKo1W1ElaEgeNySMkqaudl
ZIEEd/ldj+dQYE9rlgajOlUbtS8VdAYPWP/ZvPR9z5qlcAMNxGlEMT0WE2LgCzIp
oIlPtTQkJlnHflMrJbpWP1JJDL4aMYrq98jbo/130CjiDi71ESNDf5FXAAzXS0mz
MhNWURe9t4YFcWtGRCZtD2H7dXptPWJNG4GSXfZg2wJlJUQSDcnte76TXbrS82at
OWd/cUGPf9JEJFfGpmDCk3imgOYbrkFdzIcJyYAcu/NcCXkobMcEI2xh4KSu/7zV
3TqQtt9lKCa1/OKgc5knk0PmM5ej6/xdXkxH/2y2U2rKeUnQlKssi6otQPGeHv8+
eZ5b1HgxFwNOpsJ4LcIIJZnPtGeo3yP0wSB7trTMv2EyY+7qvZ7+X3bUS993Ulr7
b+3N16PG0UtnN9ZJLQ3KcYhc/bG4N4Q1x+hc1jGb2w/uLhgbLJ6rufYm5B1SyNOP
tHXPqNy2ickTr9AEJnQR5eFQL0dA7ju45nOvRRZ7ulH1xiHWpYHHM3R8FcpmB4VY
JGaPDl0fBv1VhzDI09fq7z90DIsdETxpOYESq9ZTqtV2DIXbcJu/xa69xYKI/XYh
k3ewRZVPXBPeYXNDYex2AUb3XtPxOMGIj+MJQ8GuOrqiG1k4Jb+/hxzpYKDMsTrG
Txvqki7qqhOYjuaUSoJJoK10VNx2JVs0UtIql5EIvghMJjkFkPDHFe3q0G9b6+kr
c5Z2kUce6EpE43TfMj1vabGNcRHbS0B9oJFRNKjr+rYf/NhBsag0MT3TbYHafhvA
oHAdqxvF4XqYA8Lxo7eUtymJCHY3oKCTPZ/QG0gf4MEi0SdtQCk4oUO6C1VQ/tCK
+BFowqi5eWCSH2Xt8/Wq1O9RlNGhdTgKfbsukHh3CamchHWX/Q8JCn9eoH4f0M5y
Cw+cPWVcefnHVz7ITYB+Sr4CdcoXvSgOimcT8Fe9utlC8MDt7hFtrzF6uBOjQjfe
8zDrkV4xUh/1feTybgJ1KmrnrTv6od0ZCXNmjwY/+SsxrtoaZ2/cvaeT6oetZ5od
EcA5703w4p1f6kZfNEm2QulCPcv03x7OckQjshzFd2eKPxE3piV0QpHk/gzhOEgC
ik3JGcJ0OJ8wQmwGkQtz5YCLvLCGEDHCPU8qjpKz4YLK1X2Nti2g5E3jdmenT/Wg
1i6OfJUUmYVJFWyh7319UIA7hQXembssGybjhwaPa9i4Pgze//CI6zKKzgT3472g
3xAVpDkMOX4iUOUEB0jejE1Zfts7l0rIZTsrYPQA39atAiqiRyrCotYdgbA7e5SP
7tTg9vMUutLKTVuzYLflVsG/Zsmn3gRGAFg78fRV5LRkUa42q19/ZLxxmWWOXdVL
RIjfqXBeS0kEQQntqg3jQ+5jEYMK6bY+aTqn+HuTO3Z6CWwy+wMdcu+8LF4OZld0
PjzGOF4SVDibuf5PUXuMLhZhCjSxYzpFga/pgI9BT0yGulOEIwTeff5sgMj1HaWx
ZSFmZDQ2A4MvRorC+xNmTJeSsCZNnt0u3tt2tcrcBF5DQLZjohrdm5UDKtMX3sd4
Kzn6BhOaJ+FCBH5VifRyzrFSMGNDKVQONp4iSMQ46OcinrLRcOrWKvbA0/x47gKt
M34Hvzx7BaO6ME862UPbBPajWE6XUrQgp0yGHREIUTc+N2hYZ8iRsJjTESX6D7Lv
7sCB9nhBhcf1yCsh41kHl0fUH2RiKfl8jhb4lzznsOtn5Zq/GHCMtaUlnoJO/Ixu
XFyEospl9dGS688cmZFpQrxsU0Gs6cg8gRjr7K9hGBhkxttYkuYaAog7iahW2XPA
IIkhQVbQkS1lBI+0q1WP8pbwyFHJ705mgAw0NozJXZHNgyi1eti1+n07ZM/aTt57
rUuKNSyzKJwphyHRBlRB5cYOOWg2X1r4PuFX0RkC1ZvU2Jn6BoGSsW34oI13j5na
LLhk0ZW7lvevW2Ra8yDgkUHyc2jz/xhjGIHY76ReZ9hqbbMYATpqVoBb+Ji2PRCY
LUifHWQNG6M1nR5MkCyEIvABWimC9+3UE/Wt0H7ekTz22syGasRYD+ZP0qMGpLuH
kY6RDTeInoDGqCD+FJ95QL9Uo344MzuHxg71KEjvrgrbdEUQfr+/wmfUO3tGDcUy
9Dru4gm9L2E+pwJ/oHTdPXNb27ExXChpIZ63KXw2ZQ3CdAnGUh4AUymXBtSXTWTU
g+7D5G9gX0FrPBFtuNTAUL3RzllaB4i3jCA/ldFwzv2kS8tTw7sfNfbdiOu4sp2+
zjTncgNxj8mtqiHax7onClsn7m2E+GgzQO1q6xOlKiIF0tGaeK99cWNApQIZKvAQ
XYV8dStdDFIRMzES25SBKIRSQz8BpTByCU+PIfuOHph1oVkL7G8HrL1SA9QI9D9z
pSPH+OG/Lg++N0dlbeeVOQRCky7m2UdXu32fXZX3+T4tMcg3yD5oQd28WSZJMiXb
FliuLYIsGJu7aI05qcudKGnrhKVzL9wkhsnsgOSjhl3iIL0sM7m5An2xc/S4dqOe
LjFprdCK0IUz0iHgjtK4dbn4L860ahx1M0Bgw/rFex0dc3qcXoFkFTCN5KK/ygUe
gC9CogXnzRbjg58YN8ZZftLxq5nBk4wpYJwAsb3oyS4LR13wDAK0xTA2xaQGhf8l
d9p+nhREkv9kroWs5/pSEzI92qfdkGarx4v8NTMfUaQEmphBu9+u3Ol5lJm49zEP
NTh0FeYcgiJx2TAIlXWZ1GuwsC0JsAMkuDSLdcQKdZbVDpFLU7dWtZSfwFOzO7qo
Ap1xlUlZk67ivtX7fW0XWCCwJnkxnP9VyW58IzoXM0mDSqiHdlODeY6J+5txbuVp
Ma9IzQG+YOWHG3EktWzfPTT6YqS7jqxyqNx0Ib0p0ytuxcsqHc4jm0HZtrnMIC2W
1s39YY50oVR67WLzok/g308pqpBMxM6C0wOVNqmx5jENjVLq4XY8EiVD+nAWJksM
0Fzzq+jDpYfETBT/IDyhxO+qKip5jqiBk2X2qPFMiabAp2MGwt77byAkXv4X76pO
GttyZY434ZimsjlWuwMfS9z9+MkP+wHNx3uEKMvF84CeCKnOkj39YM2f70kuBUPn
OQauEX/aUcgxvkJV9buvm9IL4r7Mp/VuWjLiErOGkN1aPfx0k3tjbFwuBHtit8ok
VZoVjK6IeEQF+c/itWURrNqCokoAbUO54kr4CmsKOVaMNkbolQgKXsfYRyOl4BEn
OZk4Yn/ks+w4c6HHSeuVpZJ9UNatjdeDpvlpXkjJer/mB86+sOuVya5HshyHbqoE
0Wp7bYHVxUn6D7FXMZc4QBw2eWkUMpvmNHItZIxSiJt/sc4hPbuJdOs7ytWDxgX0
d/PrjDQ1YvI+xqaoBJrkWgRCwCoglM22Pz0+xLGA76Z5oweNn4ZZZiFF+zxe7NYU
Nya6YrkudLVueqxyjnpA6mOctyHpzlpvFmxqxfrKlkFYV5q9tYBdzLyV2eqOTp+2
Fu2YsRdIWmfx/mPLwcEUFr3iF7+0+3qeMNXsSwELpzfaP9/zRbEiMAWL3Ztu75n4
KbazQFFX40Tir1PYo36oj3Ow0j7/3CSjOHW+u8rqr8Q=
--pragma protect end_data_block
--pragma protect digest_block
+D7eUHHNvqBf9iZONTHgfmF3lI8=
--pragma protect end_digest_block
--pragma protect end_protected
