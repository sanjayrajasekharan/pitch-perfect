-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
RztnxyP80HbtkzSX3HTj2xwhSTJqve3CEca5nA0Ec4wNgTWMFuyv6um0AzvLJJjQ
zSvIzCwBNGxjrpm5gNzv15P7PacPzrVSoYJKijslFFWs6VELqqqSNaxcjnRL5Y3N
O1u0aqHv/+DByrme/iGMkYfU/HKkSIZ3vmVW0vwdre8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7712)
`protect data_block
ZVYjhDFr+PRIUVedPtXRhfRYVPjA20yb9q1lR0hNt1KDXGuxMW2o+2xwSXOdnBlF
PINP1URz5vfqnb7c/549K/BPVm5i0GxdwozuGu+OZ+UH5mGdqHqogJySYgdiPvkM
cPkG7SGgQlCqh1K/lHHFjKFPr0F7EGFpICTlwl6bK5NXTChg+zA1ofkAU7xR1c9+
ti+3+bV2Y/xAZxAuyei96dWUXm17rcWoh3IMmyhuZqTnJPwTiN3b8ekuJ3+Q1iAr
sAd7aZKNa+ZqhcLIv2JnkoWnKmtQ55S/gwyPb6NKfW/rvg873R/5twlprU8hiLYr
nIZpoQ619L202Sfh1c38OstVFRKLY3sOcojYn9g5DI+mQRiXq5pdX8oCb7zOkdZ1
PRPOFHKORBXPnoWoDgjy1TALrb2R80CnG5zlXQEG1rQvLJCFtXz0VbabnfBpSMX3
l75sKi2te9ThjLp6KgTBKi2VrYQ7I9R4iPChI8q/3RTC9aD4T5apQQIIvrRh7jRE
q1jwAe+z/ligxxgUF2PpcZKNuakQIZes74IaU/vG3ekN8ITdyYRszT///MshbcUe
VVoHwOjjQZLHIgqBEJsGh2NHMTHo+yi531sU2/qXbGtbi9cPFYKTxo4Dpdv5y2Cq
yN2gwWAe/p9TjszqFZ3ErF1/G3kfpgvbZfaNBgsxb1M1fXKsnHM7HeuxPlX6mqeo
nUhAP0dXn7qAd1S6UrDbDxQVaTiruxx+hz1RSi6OBLrxTUleSfHSHY0PwtgdMEeH
B+yEncx791NsgC0PdSERb8wBNXtKqKj7Y8JSGWqdk6L8P2JCbDOz7sPbAE/NRog3
SvbZ2TERYV9/s/hgq7m+IA44EZZBZVjWnEixnI85bQj6dRTimOk0bqk8+8XRmbki
781pj4moU1qHCIj8+j+eTq/PCd1sueKsa7LNNn0E0asbjCXsf4JkEOGWkon0fvCm
x/8JlXvaRSG8/trJU89CK+4hYA3EEM9E9XvLksaXAFkYpSus8X5GnoOnkCCrz1Mn
rE1RaK2TkW8BNa9CjMe7OsDjxkfPZDjLhbXeIM2R/QS9LFmaetX4bWTOaLU7CVsT
ocKvw3dqvl/8ULQdvS0hGuflDbR5Za828W3gf8bMg6o053xPQsopRYgLNXUG0QAR
OissEzUPEFWJF0lJ9T39ENacdgTU6uZMYT5vRyFPwSAlTFcIsE+E5FQUXwEs6/He
AW22J4Ml/9+7TulntYHbjp21P5X4YkL5ltzFGKynBsJLmOF21I2nyM2UpuOiYGw7
FhE5gSgODFDLM2Bf/rXDdtGY1DPf18vNBmCFAzl3TP+rfe1QUk/j2RFpAhyo5o/r
FTPZxAB75Yvsjqt4O/vO9tXHsd/qq4F3SuaY8qT5q+RjK04+nY6suIxkh20mpIFV
8qOLnb3dQpAUV4OCsqOo3T+zLLZobXZhrWxdQ74kiwW7oczGm8xxjnjuHaxQckB+
t+AWHIfHXbyTf4EKgzUM2vDK77G+C8KrdKzUv04BKGeHWxI8Q/41+Xo4xBvwFfPc
ZsJ0DjlPka/GV3wMCcG5+S95cOrQAUPyHi7YYtrNHbuh8XxG2tOotPlqk8msD2rm
N3uWf6+Ipl2ZJpOQiKe9JaN4/db123kjUZoxWxbsiPC7oQQRav7gDYRHeqNmZcdX
nkObz06eSRysy79Zvl1vLfYLMK23NvdLib9UUkkIq+Pw3pT3oEJTIl6dhrBufewB
y0A8ydhZLie0Jksq4wcc3Wcwwd7nYwhrA0vVuRKBElCDkavnul2QZ+uf2cDdNgiS
OKu5qE0N+5bsiRCAaUCuM5aT/VErc4pNjkc7SUjABYHbat7sN8d5QHgQwgS4vocd
ElGSwEPGAAaO+RUWNNtX6spyp0Z7hbDkFKcsDv8gHTO/By+y7pEX4T8Mxaq9Itiy
mKPaRTAC1esQKcQJNPzqCwGwox/2gI3kqD+I/81LbBP62t0qw74ir3at7f4+nQjT
Ejj8P2Y2E1hY4ltA5opSIGDMvL9qOWMleWDdLXjy8O/RjzxIBvE+t5S5JchHu/2B
AtN27jcxLf/RYttiBAs9QV4jHtIZfG79OBUrhUiCc7K1vupKsIShUdCvkhtfgf0N
d9Vm3CbUVQwDqJz1KmUUcpON0yGIqOK/XptX0t19bxBGklJ/Eldr2Mlk/SnDh6wr
E0CKkSnLZMHLdB31mwKQM3SQAg1KUuFpQoXhftOpzm4nkdjbwd0cy9/c8D4XpBW7
0qoWlTckVNex5lY1pqedn1cyDI7gUnYv15j00LMMZuo6fOxp/JSiRQSo0QVmzej/
NPtFk108/p1pJqdVLCvA+jk9PtUrbcj8sqT+mXOSWLPzABg/lms2Kgx35DFXv3Fz
55UpUGpbo24+WG8K0ljVcf1r9apJ8v8vapVQrxKSRtv71AHqYA95hOEjjOLeAA9q
H7Va9/YBkYgDTeOVpEKJk8wbrldMfiCjAzlsHzRt1fGiY1bk/I06XG4luFxPh+pV
l143354o5aWGOuF/9RS4YaVBqDncFZmosO26biE0xhiHanfDw6qshB6afPlVER8+
0yRpap5ouUD++TZQ2BBSHiPJMX3yW+96160MJm495YrnhaPyhtmIKidBftNv4NMB
L/EOtBvKsYgrzZN6Gd/5kzJV7cP7q9QEkB8UHD21p+vjCX0DcwrZ2ifh62prBmUo
hClj56DUCjE4lc8iPSWhSgJ9gsFs+m+yLSfpRm4mTUuNDIi4VD/34m89bN3L42ws
XV/9GYCCG2OGjRyxrGF0F6jmnp40m6HuHmTki+j5BZ7ePsUfzUkKPSVyq+kx8snQ
OCStJyU8wTPFRwNfP0XlOZbVmKmkmkWK55NUwmF9dAKZ1NxrrUcdNZnzPAnIMMEM
DvPj+CANfc5scqdKse20A8YHFOHJJStUMMS+pYKv2Q6wOy9TwdsU8tThjTMwMjQO
Ny/Of9m2YfnNiUnJgziXldHQ27H+dtJTqs604lquK1bWtmcaId8TdnHOFWruCZ82
9jl8LRTN153x/e1eJ4mo7itz9Kjw4jmy26qJYnc0ccd4e4InXUk2EOT7FCHckjMM
UTL4YiHkbb21/5xOeIPjJWff7Hq6AaERV5/GSWTIQEFlG0GM2lVpTbjGFmKL/V5B
9O9mKmxi96BbD9V8930xCZFEfD8r7J9raAGN9e2F7aIqVxYwlK6RJRaBVp9R6u4Z
zKmpA3Qj8U0w3zB6XR0hX6xUgWPapRcjgndXrwPX2ay5duy8KJyxZOSRvO2RSE2+
36CNofxNS7Dw/KGM/13LyKIHxMS4/PGY+JJeVBiURUBLPJ6c2Upp2+fFu9J/1Fn2
UXRbdmHlU/wUIk5jT+ReAB6SyUgD+vzOyelJsDK87hFq1SbuwIvD9wO+4A15SnaD
mPVx8x7W+yq9tz18TZDrEmz1qCdrvtihX/v2fpf0bn+TbK2hDAjZ7aYS/LLqjvRm
xNwbnaZqtZKo9a2cBTi6iDU/EE08UCN9P9XkmHSK9g495Xg0dxR9vo0KSb78eJH0
MyH1i6tgrpBEJfUHlFhm2/wVskj8L3A6rH2Niwf+QnCK311Dum5Onxb1DA0/11h3
2fG/fcBwJlZ59S1N/IiUM6gkG3N4EIkOSHQ+vWcOZ7JpHjRaJ85QJBd78tX8TUcp
h6EJwfhiw/ZFdx1+EKuKm+u9eBrZW8eevTxXpBssjJUD4NRRBeZVI0jhTtw3G1CT
wBDhC/BNJBpVlonnI2c6WPW+RKZKp13ecJumZfOKj4ZkQlbj4/yfbjDdiv2r4Eto
mEnSJE2v1PfA30+qV6Vnce30fAQ9LQOXNj8tYEZBDvzqJ5N5oVwhGGgq1G5UpcIc
XCN/Y1c/QZkNsAUYm8dFgEbLn8Au1K8FgsNF0rvFH+7mlrsueUFAxgrfkud8F60n
JUjanqzUvm59MTfrtTqvkZ8dsEXSePx5PP4etHEnSGLKCBFHMmq4dhT6BQyXTsx7
Idq6/szm4AsuQwuzpB4OjbHfSgEXx4zHqXdqU5J/nlwsTUA/p+5aUzq7XK1g2O9v
+aORPtdiKshxT7p+zM/hKi4G0nPW30kFF+/cvMPv0jH6um3ODx/ysU1mB4mIJyP0
FD20IIeXNWAGWg7QgA3MJDAek46ieWHvDW+yXc4roQvRV0Xg1JJ+XLNoXPkAApVt
wpy8nF8bS6sklQlALOkHwJadjNAl96dH3jMyQPBQus74IppW+BNb6N6R6iJB6ZxG
9lg9ZcbMMbggIZ49K/306y1ESTjyLNEBNSCrWvpSK3dhpupbEcieHNS2FkQcvCwL
dOzLEO+a4LBSG2j14wcRAYrmRNB3uGPCvYhe9HPpigE14HAxN1pCBEB5S8sFz3u9
4S2lw9tpGDnTtpJt7tPvfpTYjALa6Glmydl70OgsTZDKmIPu/jbvdKdEqAtHzJWt
WJ+fNgRREV6/0lg0sRRS6MmE9zsaCYY71lhhnntxbwR7WaN5RJrKISZCB0ifmpeu
6LR7tCAhan5Fx3r5AZgrBBAegYN0UaUfIb33ekrEvMsH6/FRou7BUHDKSCQBk7HF
9OPkcLFvvXi0ZVuK3xyjBzxABL4AlxF3bEdIonKK2uFd2rs5qdakE9H+N3gJZAO6
XRhFAGctYag84qfh4VPSeiCvq3KnxA/Cd4RXL90k3KGLl6VtAz2BZIVQKm5bXW8m
3SYPRFAXP8XdSj+B2pL27GGkkqbttpU0o3TCDJtgKfhMkWAXUhS7xhjiDTfe3UGb
XgSVCO5h6UBZ+N52jwDJVcl/iCfyW7jmEX7C34oWsevRDmTajAQ9nwvvERT2jzYS
/uQD3WoHxGnbbHdn44lBqLk9jTg4nqKUCxwBBA0z63iXkyjEzTcv6471b1PiO5Zg
f+0ly6ux8LyM1dL0OCPxDCZQL0tkGgBKGFCx0uEp5VUyG1clq8YzKNXtgXtHX2XP
GhqHj3u9euKeVb0134ISu6GjdgIiuoqursEOroD60kexaZpvG73V6LRagbUuGFjD
Gkoi5w3+BnFuVo4W7OuNmONwCRUC87I3dUlWvEeq4K61foF/xVvCkLa9B3UQE26p
zaBeCGbII/zoz+YcCemK9lxRubFGVjW3tJwHa7a/wH6l+XhSx5MiGjydvxspM0vm
4+DukUcYs3tmdG9fCvlzWqZTOD6EmgYcPBdZajRl8PsH64btSblsJTGhsVqcevIv
86BbeTuDQgX9yblj/83BtaM1hQsjvZploBwUfFId5egPGFw6mADYVXN2VSmWWq1/
uL3qSmbQhbCrk9cKB7mRDIqg5RwL07k101cNyJ3N2WNKlQ3a12N31Vf6Q1HJusnv
GNZzkMOuzIs/2dUZ7AlszLjml+GwshANV9/CELrA+d0erNL0F+ULsPtrx88olZjg
eyPneD7Rseb817lIIx91f0x4Vrjh4XweS2M215HUlboqfZYkzD4gKMahLiQMHyAp
sxtYEkvOIKuRwFd35K1gI+CCUBtzgDqSEszTABnwEVZvPWoX2vfxIbABnWVE3wqE
vbX3BuVOE7uQLpw09Qpb9D2+qfIcVsNn+yaImQ10LsydfN9U9wIrLrzMCiE7bRW4
CnlShzVV5oa5jyXRfBre0+z4MiIjMAVZTFy3XZ2pevKs4hvQGE9gGvnZBQMsAFBW
3wuTL3RNtKwQ3p7CtIBoMW2o3Sx4ftdBSJPm+WOVWf3TMoVeILmvo0sEaspsAPw/
egiLYCqfPk39l6rhaxakOIu5yJ/HnPV5B29ER2Y2fbke3yKaa3e2ct0XJ0Nl/fYN
Ip5AYnjT0VdVHC5SwvKEVWABPwYoSgkDIDYOsSSGFVrtVZ3ENMpxYRX/xrinOiYs
Zd/PJsYkSoOe5IN29PwhJf+3ZTOhNaJeIOI7CqpQoopP3uGI7r37XD7ybavk7pfd
CPk+Bw6O1NE/3HfnuU2RkVjFMG9dCJtNOyn/QitAbgIcTvanbrHsWdImFhKaRh7X
EyU2fY3EcgulwcUaDa2ZVamCwhzsVnpmpU5EEYDsFKa3V7WCtv99Oy8BsS0vdId4
VGev31At2NFSkgJRRg1OyGl5VDEDYTxGiQxx8Hm7AOGVLkRhShoKqG05xwdvocVB
g8rYefoqjRJPrYlOAA+s/cTUJUQAujnNsUYKBbi/c99GX2YBb/BsdsozSku54tRZ
CmWimHdk+zYhJOYgHeVHPNTE9oOqJUsHe70DRJMEH0JuiaeuQfMSobKmsrONLfNZ
wTLjLuWr37BbV5+U2NEs96f7//IzK/WnWnQ7gf5QhoSklXvdouSd5e2lZ46IsmZT
JreORjK4IQuahd6QQIyaI6tSgo4s+JtmmRoUP32NuTEaKmBwTBP46PmlRyktnPAS
s+WAU+SCSuw/QBtuXhFJwKPgCBSjQqUSjW3D0EvqgGFaHdpbjg5qXjbyq5O73UhL
PmoPdKuqRSLisM+K85lqVv81iYaW/pArNBIxx5gxNl98dbutxKsja/L2x766BQW1
DtAXZprNmT7SQnX9o2XXo5RJQags8K4jQXA0pa9OiP2Vpa3cw6/guoGN0RebTS2w
Z7A6j/MaufpHN20m+zcdb6/Nf7BeWLz8plNMEnNVRXuoTgxC6/chATrZwlzwNUWH
nWhIeh9tFQAb7aDIowW9aIHfIPhJzlvZThIaZFLWjl8Bk08Q4hZsWDW8fnqcmpA1
sXdkhjKJ9DHPVcBP9bYXTraELg6FXs6bRLfHil4ccMRoyag3s36BkCVA0ExmUmWE
oM8MZVM0CqnBpZ2F7Ygpq49noLOq98HM+RYDJ/jwNApjdLIo0MBtd3gZcTSnqcjn
nQ+JF8fWvROoLx7lk6rCN7w2/+bNzerQJ2G878GRxQLlxDs22pTszls5R7hsrJii
SHwvimyPb8txVhpLzi4MAph0clwt6DL8naNk3jWF3XZae5ijXIPpoifqnA9BKCNJ
Z9toqVaj8g2Ib/z6I6uI3eORD2kQf1Pxnv3GxetFojK5s7NJ2gX8Lp6nBc1ESGZS
fantVYEC64e+xe+57lAgDCC9i5JU1uyFbzai6nn+c5AFsneQdZleww5Gh2mN7V6V
Ih471CmnBKYEa1U03wiul7+4No0CENCEvvjWGsFK/U/HzFYafA4ao8jDjGEGvwRR
BHmlbKXcgjVCNPjsg5RuOIatBwFj4UxkpbxmQ+SOdLFzox4jun/1uhwUS5v/Dscr
7AG60xKS93/Cnu0bYCfVDgJG5zUIVI4x4FJD1cQx4P9z6Q++unX2uJyJiBfm7SBN
SImlQ6BtQc/CbuMZ/6EQHx8Fxbf8AiJswR3PjBhYR+4duMSngCxHth+76pt9bxeT
2lZK3o+/rNB5XH176NGD280WnSNPwgtgFkcWdcy/kLrim9bcIR+NVbp5sHrLNlGG
20ZJJcCvVhX1nz+aIarxCqBfsp69r+Z5HyRfyyDWvDh5J1Y5RcZch9Nzwm3sGqS2
+WaeC4j/ImLu+G8SE1PxzTikB96gkmCKFRTHucWOt3E3sJplhmEvn/xWOX2cka+b
W0B9IGRknsnGAe8BCT6zwqt7UW577Dni4dIHlLh+62mb1ItnOg4ld1pmzUxKvDBr
bAO9h7ZH2YbfoAvM2UlomoiaPLb1Jvim4zbbaXrxm73wvVFSJSjBJh+fNnQWwops
5xJTKlTzFHCJYhecWzB9hz9/cxEnzVEKcrvyC+ipfqlcNKXut/u2Gu+7VyIZw3Fi
AUF0DR6uqg/+z633pG+LsollTcevS6j/d/ZrpP0Zk47a9S/cIaBdDsfw/WemrMa0
tr8DupaaAUdmyKBSu/xBAIQC9V3XYPe1TiPa9yyP17MalD3JIqinXFTDzG0+oZLw
VF9xIane454xliogZ3gPBN7EnT0oB88wYFgXeHpnHL0nD//6NT74Qx1GWifJf6Ty
MCTrYD0pmTUDii9nv1vw/+HRaJK5/+13Az1bkoG8nuITN7xUqvoA1qPD5N+DtGmT
f3GuBaJW0hH1gx/7HZU88sjG6FTeVpUrrxDLuPj1SWjRjlaIHDGAGaF8ILzstTnB
AWvmC8zj3FpnMoitiJGBS44cBf/P0zfrPCwaFThwdeZ7TX0V1s2h829IXihp6xMk
LHlGpffCwf/uElvk1lBChCbved+M+aITBPCJQvkBi5kVu/brZZ658B2BaXTzTAl6
iSgUlImAC6R2IABsSujlzkAp68vVpicW41Dix1qBri1Usbt1rvHHwjdqppHrnYfU
XGDmaevz3OHYC6bbC1eF/cJNBvGKNokuaQYavac8ekTGHekoeFf6TsrPtJRnHJoq
VBmiBMS9c1mLX0ucruPgzD0sg7qXfNyvMwnGjyYW0UYpM38kegcWg8pe3JV49lTj
7dPFxAbL7V9KQUGQBsKxf1alCv3y6GJpGcPg45Xo7AKC5wTxrHA9i5UuEw1BzPAc
YK6kQ2VsVfcSYmkY0KcKiwSOff7t/Z4UKYwLjq7puA1bFdnu3I4Yg65PqUFkGW1J
0LfWIh73c483NSrFcltNioG7QmFVuUYz91qx6TsMCRCdUTbuJyW8cmeVT+E7eHA/
+ZvncDIxsvNBcGDJVhu2G5tU13WbPsZk8vHONLN6XwDXxLghB/KpCH6SskTutgb3
l22PsXpoCzkm7HMu4y/Qldpzt/Tpj5kMS9+Rd2iNQcSZb8SWcZ9S/xNvFnfLwZ09
H9gTAFPd3vJ0OEFP579Cba6q/ENMXqVPN75NHX68Q97mUOE6IpxdT0tHMjnB3ipA
bkBQldIjL68emFYhcM/2Y44VK/Tlak750D5GBoitlrsuI2prnXrcI4EoScczNWId
glpLbmtmnpZUowSdsUovtZIrkI54opid4ItciBQ9BWlT/kFAiRVwzhkxCokY92h2
aBfkuQEtIuj05t4Ts4hlCqMD3Q9QdZbc1L3HdcjbGBqvMAJ0mDueB7tRjwdKCcUM
ALnIJjrditrm7+W32c/6XQOGCuHyE+p2E+2YZpd/Dudifcw/EhoRqOvTdsAp4eXp
llM1u9e6KJfXDEGCzdX0vWSqXOG130GcWuL3LBs3UvCc/+yxXsA3y/Nd2PiTA/Nd
y6zz+k6oOB2t7yCqV5RpIz2ZaqJgdNBgD/p9Tor/UfWjgMrPpnFjnlIqDszEqwwd
SwK5ni3Urh/+w0dU9A7mq9fbVDgQPUNN6R8oes4dWuK+CdV4k2kKuaA5BsgKTfP2
RRTdWtRPebO0CMRHZIa6CMoxPKKC5WCKYB4rLR5MDHjgOGF/pQ4tTCxWIj+E/nA4
mHCgCPCF0EuFmL5NZdCOmW6OkaA14s3OYQC1OyxOu/KXl3kQFpI5Xw1yT5NyXrtN
i3nPR72nerRebOhCyT1vNuady8gYhkl31LxpwA0bBxB+l9WtnznNJHu+ppVh2gXP
4mm3ipRWVxXH5RiFIGxUUyDfD2xgekOZAkfrISYfszMd2lkRg8ya4E2/IXNlqOLC
izg7nBf+r58koYHZ7yurKBY6E+kIALCXvTGGzgZ4J8UFxTRSzMbS/rBDpAVJwMue
8MskQcj1Mk0frniOmx7adzc+mYz1EzMqPhmELEb+TSyV0RU/y9l5QvhMWiMMOMMf
U68TTiql5iKF3XSMzsrh4HW0iYqHcP7va27Rpk30GSNyBSq+1eqkqqFeTtHiHbr9
H9qZ3igbrBJXppGlCP81VkrC8uc9axiCeklfQAgzpknxQgW7fymWpNua7sMGpJ6z
iWPYS8J4JmzUw9LicF+Y47exwZDz3aRKDhjzyq3bzZcIFGsGhLOUlj7A+s7OwWUz
C7yv8uvXU2Ol40V2wrvCWjyqP09kf5/2RVTSalEIPYBS7V4FRxnQj8r8Too4I5H6
Zs9hGCnR2uR4MpM/iMnDQ4lTHn4u5ySGL1EYKAsOE+t6Xxz754pP4UjXu3C/6Owb
45FCE/STUeWXfxN0hLic8NQD5hsCotAZ4lLvAOMHwglpQdNNu8QDtGbRwgy5NJRT
ynTa+ebH6O8xQxssMvacvIiXBIoGfVxwbRRPgcfG7XCYtLsG9szR5HdlXyoCGDKA
+ilAsnDZHBVhtHLDv/G9I8itqQQbGBRj69a5o7F4fH7KDUJlwbilBnN7pkKaI043
RwKRLY7mC3F+unhVps9DlQwKE1QlOcITQ4gc7Lg4ChHhOxXlvABLebQHs9SWbB/Q
5r2WudM/4kMLnOFGL6wBbue1XOg7o7xTCMSbHtyAuSnaodtcpa6d2i/yltuNWMYG
xia95IT0i5eOeaH0K/uzH+12t/mpRLo0YJAEvWNaCeo7RTMZEAqzIt9bh2Mv4ZCS
7+9P1ZUMkal9VdMZiZf9RbQbEp7vhuU5rSkzVwT/jjg=
`protect end_protected
