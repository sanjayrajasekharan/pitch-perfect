-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Bieo+PcxBGz6wTFrnBp6hGUvPo8vUA791uSOrZF7cCNZLjIKHXjAJKpzKal7r0qpKb6H8aL3Xw7J
gcwQiohQPKSElaCADKI4zfEJNHL0PTRkDh9PCOmRRtMXEOZBZoV/ipm5gjHpqhDVi+HowgyvrCv5
Iw+ndTj6gRwMv5Uu+jD3C/hEk/YsUtHrYn+9myYr9u3z8raODcdDEfUPSxjai+9iz7HRxnMaRyhz
B/zYSbg0wSe05DqVpz6EXDq+sbLBRmxR8dW3BQ5/jIPbaKAjndGm2o0xZwV/4y9iJ2Ue/KvNN2po
m3bc+mTIn9+STK+j2T/UsTUsFJBlLCKX8q3Tfw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7984)
`protect data_block
e4csC30ng588gy/pFGVD77ZbirUnHzINY/cxJVtAywShgn7GnzzMq+EPldo69+yGru2fSWcdjXoC
H+g8Ww21RpKOadCTm5vxkUWqX7A0ZnW8KW/VBpy4slACV7c+aygeMuPQfZjPk3TGV1cL0tikvEQ7
BHaVR/6GN9IeOc1/ABS5/xYrbY0D5GPc3ijXzQIJi5r8rUbKQUyL2Yujdnzeh2yhKxofBV0ysZs3
ZZFZ7BRX7nqHl+nLHkwd+I3D0hDu3t9qJCy4XTozf1OkCZftIPKUNjG7a3/O3iNPjM2yC7f/XTj8
0z52xtBBoeKgOBc+ZmbcsM1CIq8wpmj94MPqGuS7bwtXrAJvEh6ox0rPVpKgygw76I6ZoHyLrY8F
CUpNbwIz3SGhQ4mngpqmAveOXpNuNbIRnBHStNlgRq+M73l0xh5bVgBYMEJSBQZhGpkz/Jpg129y
H2AbcSsgLtrsghUMrHEZh20cXFlInEG572oVbJJ0xGe7Qz4kW7d5Y1mAZWq5s+ODJiWerEPjuwp0
FnxqpadUt7F6ZtbHvrcSgBjUyZ/HMeOBHfpSjUzz3Or4Y1PO+IN11J0VgVv9TlZJ5OzZgF13am0w
3DJt9lEi79NIQEwO6VFxyoTLC0zQuBGRmed7418DhjaRS4vLCo47dOslPfNQ99+eJ4Jj//BQRD2w
xD1lcEhGYRcu3RnpbZhI/Egc2UYpk26ayVMZt+PtJHAQ0fkSC+3NcBBM9bD4E2qIMkUo5dWKIgI7
4LIJsBgMIu+NWePGZNfB5TZctKxsSr67UKVR+Vp4a1jFTT8+mXUp7pFNExpq7S015Wb+WMssFcqC
bS3DIbYwMKaqeC6Vm77fkaOI5Tx38UXJ+hVBLYRq7Jw/y1PfjOMBgvCaghYhB79muzhi9vfsqIbM
0Xqeu93zL+JedJyKMWDBObbHRg1k5QHaGnjy560tr0fbrZf5DF8Jv2s5FHQC24DYUgn0pRHpQ/Hd
J5FfmleP2O5y0D5L4Xnlo1IrXoxMaQcUza/DA1zPxoLW7C/k/j0K8nI7vYuaidnjSnaUfwS2WTgX
1tz6cOjYPXtynMzAooxqjbaMqMF6zEy7AR9zajfbQV5yvdKIlwv7NBOVKDtnLBGyGjsGhGATfr/q
JuldBJd0gVSEIKZO9/pbX6lj49IiZWZ96R/z+n653QEvTiJBl2b/SghJDWRdf9/OZq6puIDo0Kf0
QK6XYRoyQoqe8tN6OXMcJJibIFCNRbadpW1X0bLVOi3SLu4klYL3dr1onQt58T1Apyupk/s1chxt
ACCo816gIqHSYXjN1oWg9BJGZZbohMNH0X+DAxfkrPxRkC6j5rt95VD5onQLzVNV7Z9IV71D4t9w
4rpshmyIK4VxthIFvnT7QnivDCagmSSl9TK9Vfl4BFe0wHcWnZfk/cST5PhCEXLi+/3NGv2sLHRh
2c+UJ67xa0WRAJnVbkdSm+mXAv/kU21QdnR4WeK0cRS/TmM2+hKK4MrQ5DN9oMw2pqOB6OvIGH1R
BABjnZYzTLAu72e580qPSc/UGw2P4AYROWroOjrrA/MnLdj4g59HReVVfwBheuj0Xxxb+MUOpEOe
s3BqSdZTy0sAHuaHpU7lDuoe9CaI1PwlSsUbeIPUQMwvWSDGynbtTOCobs80B8Tk4LZQNg1EGKZi
hV9DaO8hggwtcDqV1LG2kRLohZt1duspzji8itv3qAXVMSxGZHEKGshXaC7iL0wAMw8VVPzkGUBs
qaLMDSWQA0oETtafE0I+8zH+8y69rdTFEe3DSNwYoQnHlMz5Xb4Y1DkesqiPQcygHsmy+eS+sPQD
9bEMcZIuZJhFp6Qm7/QSQcMQ5YDsWQa7nXrtVM0U6VKI2jtgUH/i7qUum1uQ5P2EssjVOf3FR2Ov
SpjuKA7VWMIHTzrltc8eFN+O2ShH5mRGbwB6zhcdFUiEdOnPvOp5FxtNMGhP98NQ5WzJTFRlcGmP
QzK0ahi84J801/X2FCa9mQcQ0UuBopWNknqz8f4u53M0rS/F15QqPAu5npv9Q5rq2jPixPhba06C
LMKfHLwLYjS5A0Jw3v9DCT0Xwz2dbtOz5Axt5eFD33SnMJLejtn938GlsiPT2GRgk8s6oSlQt+Mx
FzS2v+f1Yt5q47WthJUlE007uuah1kJ9TucwK1V9XGT3MPSJxvhTHC+mpDEj65+i6pcyj0vMn/Is
vZOGUhddD1ZVSdDKLB8od3/YVTw0Nw3kayTnIeQm0gEliwOVpSzLqyDg1Wklfx5FdAFgFlil/44x
huTcU9J+cNTwad51gLwvLZoEGOcEaT2OI2v/IOFncCJMxFE/kEEA3fJdchgyT92DgapeABuRLafO
cttf+y1rtX7brBrQd2iJj3AoEEZjJ4DOwc2qs2l9lSRvRk1pbHRa4gIpGnUPrtWwdxkoTjsRxwnL
IKUm+kAr+7BFjrH2mgmAYcbrSSNxRTetgElGsiF2vpC0obzElwMYE5cZOTIzQjcAikUogQ2fXB+y
zL10QZuoi9bN9rSb1DP5IyTsZzOz08VFkzVxDusbbFjWcFPgjXcsWcKPXpGzGHfrEXAyYJ0N/z0g
5fhwPp0UrwvTm8Z+fMqbW+Q0VTkBby5i8ENJJ7ZgTgcDv3XMNgxpt7+KGOnFcRonRmmnOOiTdpVG
xw5c9rpoZvLoL395esfr8qgDPnAcfB+NAmnXfy2zBdK9STWrSco1gKN9ot3vxSAY9eN5EXwJ8vkt
HqtCmfNR/KC9cq0/5VqgiE+t+9ixwp7x3lR/565exbmnIM0Hq26rMDSO/0CW6mimV2Em4RQDHAxI
oGB3fJczrBz5U+kFDm+68jOmmn8wqdR4cr1++hT5jNDK4MlKJUhXUpf2Yj5MHJdPwjSEh4FXRDsV
/knS9uSeTq+8EJ8Y0H7OtxNzypCg631EuRoB2OC3KxNx1eb2kiIQcWBhFE8YOkcFAq25anEqFea3
hDt6F86+C1IqCg2b6jNUI92AYPdPVFkRvJL5fKkRn5H+YRJp5CeFgqyncMMbGp+GBYXXaG9CMMtr
zx67DLD/s86ElzEEnUlyt9H757btXjZQcdZz4BQIphTm+4NxnZM55xdDppb4DCTzOtI462fk1MRd
1Vi1YLg2RQHUz3KinLrLEbs/dZB8ZycR2qAtKUpgBo/SftRh3AoJ20mlYSDfRB7wauzNu8Sz92QC
AEAZlRQf2aRM0iBrGccNmAJCz8C94/r4Y2Ut1t7TsDu1/hzoRhaBh2+v1cojmjMVrv1iPRnoQ7ed
Z8RHVh8bWicBPU8Fnwa/vE6iUI1/LuYH1aeLMja+4zlyXFchSW43BxjwUdBEPJCNLJqmBY2Qq+Ct
kdvrHi+vG+mCjcmbGQs++SjQVl2C8DFMY41Bl8wVVlS7X8Xsm5LnqZDmhseMcvjAEcBSgamgJ+6q
lNGeVLcoA8YQ1H7ZMHqE6l6A182+HCZkDyA9dkK9gfX9s9gywxjs1hCwkc5Bk8AuqSTDS7DzFG4E
KvJZbQHnOCMJSRwbgbtDPCPRRM2qX+PivUve3097hlknbCpsh3ihMAZ95G9xXmErherJ1Lc40fp2
2HF5XVBGNdMOd+6gDQrsbXpnwoVm88pwC97gXGnpm4xK+adNivzX0RzBu4HFgPVfRSpDVxPfja/j
eWzwAKQylc9LKX+vQvX/Pi2Y1PJ1v8P+PkR7/XUuhoMQxUF9+faF1jvF0a0Datm0DCQEjcE+zASB
HeMAJ6nKvsaBjkXAQUmZQWJOEN7HRVa6ITzokH7y7/1pBspchvDDucnmKysL+QwTKE4iIvU0Znx6
erObYlnmr/FEEpiR8wIv5pE/AuHlIomCxVjbXJaklHGMwyMdmZEm7SHfuYM2yTuQPVX6PEi0HhSR
teXvPNM+1sndPakZp2v+LVMV2yVlxA4fY0qrC+vn194kdGnYwd3wATlRmp56V5XVAWvypnzKz/cg
CvI99R639owB7fFsQukzHXz2L1g58xi62ygzilvLdyOdQ6oUNo7f3pv/Au76upNKeS3ZSrYXUJyB
I6vijAi1CtF5M87Et2fDCPyzAaHdZMhs0Df5N2qIBeA3CI8aY5yFYfgMBSi6rrTk6XYuoSuKC3iC
z/SP26bgs0r5/IrQ61crIw5uR+ocmm4Wn3HWtdfJIK++jTZ0roeD4zmiyBFJocPuYM2HSYvLk7Eb
S4YjIgyoU9UuUl4Qi7fqD3CX805DSaRud5Md2Y272OY/MGVrqJb9NG1IQGgjjGCBQbAhFxa62p9s
BQl5KhsQHZXQmgQbV2NLZh/VRVmpCAlUotk6OHy14Z5/2Z/baB7UOfi/h/EleV0FnWyRAqvtZDTC
jctMUCvLEiDXz7G9TWs9zx8J0xF/n88nAM9pn6zPtuItBVtkdwrmwwAyE5wpN73SJrPLYhrWTHhF
NQNkHJNLjBC7/p9S2wwPmMkZkHKHn9lTZbBtrVT9x4OeXd2jsLLwLKYfXGuHxa4E4abncwQZfSMg
ESFTc+t9wgE0XE8A7CuWHhtL6dfNeyqewGG1wG5xBp0eLnqN7GSllRc7ASDZPFXHn12KDnl5A9O8
sF+UnWxzBVazdbhub1b4JTbP0JbN+p41b7O5Ydees2rNBsrPYBKmm2E44/iDZxWxe1JcXgG+EbZq
SUnHJo2bVisaYjrs0weRY5ZYRKXI310brq6rDf1MbjRhcGdJSjzUWluA5E4LAi7O+D0AiE+BrAhL
Hhz/7LrSAPUDA9GTFk7hEgVcU1tUvqWRtdMZOrTbdp+Uh9Euujn4xS638gCpTu5BDq+IChhgbyI+
DdEBfjyjZkZunDBXtZACPQhEQv65EIpQYfa+sJuw72zhrJYiZMljGJMXF5iCeG6JHVnkgNQYVN/0
AzpRyXAmrks9vEah06pzyRfCLpcIwvTRr/2FMxmSyEm5SuptnXMfjKt4hApvDlg3E8Qfv1Rhksui
pVMiozw+dtC9e6XIW8OzfkvyxdnXlXa7OwD9HBoQ1UEyf7Y4er/ZNwOYPqdYNfM21/NzGNI/rIxi
+FBDLHO079QThWdmA6YPCYOj62Z8dBai0AUUAIhUm/qp5jyuvUtxouXnKC1HlE+p8gbRjF8nZ52t
MvQrYx0Wgs5zdPbDnsPnjpQtwnAyUnAxJE5VHf7Xca8gMPPkr0MAPXhXMC07FheEVG4k6UOigS5i
8drtwH7lNmwUgp3VrU7/Bw/C25shK/L91plsy1gtfsmdX5jU2JMN8m8GMBP0IpRHeTv6zfrF/8Xh
nu/Emi4R/JrwzKipe0LCzE3Jk828FuYEp3shDnuvWJCzkAzL8r77I/tLsPO5d82VtWkKRBOnugEH
p5XsXkrjeM/LsaV4vremOebQVDg6CG3oGb8WSZ5kx9tdI9HbfUxC7q/FgwbIHWDJuZguzH6rgssb
Go0K/pSJARO2XsyrSr7ju9DJ4I1ePxRt/QljiunITNsF2xKgvxSh2JkYZzJzr2sDt5Q5w0sJs3xe
cxMdBO1eqmpIhDi3C0VWrxdo8e1JuQ4rBe3P7j3ciJTgKHGI2zGN01Pi7OhayGf+AQFSMNkfvIZF
u36RMM+MXmU/2f3G8HnGlhZVaXt/0GWkHoQ1UzbFhhN5YJuex2wo/djurgPsttYZJBDYIHJ9dDwb
md4Izf+RyDfI6FipHqThfijaDDxp3EfEHwj0tEH7WxVBHOuurWPUzgsipTOnE5lNYr5UxaMjC093
6/chtCtPfuGRCW6OZDlbaYh/1mcMzv5M8NNx7gWnTgFWnGCMw3E5MrGpR/3Zke6JbbqmRsiY4jEZ
Eauh09ocE1jNSEHwr42CuX1LJBNIincMem6fwac9kCxL2gJARazZwK+mnBdM2Qu0sL/X0eRX5Y0J
MaKplhwEtibbFx6ZLK21mtYbYQ50f0T0x30uzuw/7RuNIbjIQhrDZJ5op4BlqULNOQdLMkwsm4uL
ZneYQb3w6b5UqzDIXh6YiFzm7swhmZiumBCHsFX93UXVeCne+lcGqIlsdAa3aWSWIUQoqiaAVFLy
e6hdjXqMDWcUzkKO8ZyNjOkH7IH5d1QsPX37R5DqlN0ASkfCxsWo4TINBr68Fo1Cg/yiFcrUavTK
UR0IfrW7PtTfe50XmhsvTbf2v9jHJJaEhXzrGG1K7FG1v8mkFGFd372AA3sUMkRaYC4+4P/RuGK/
/xJDQTTX8OK81Pqc0RrMrMpMrVSMSZyFK4HITWBqVjvmDQElEU+19oEvpIMVKZdxM2tP7iCTox74
7ZYt0IFGbEbmpWMJMfboc5MWYG3pdFAbS4lwBjOkifrKCi04bXQUHY4/It6rAHFb1DmnX5bNycMx
/XveCwfpyqKvlrq4DrRzDKuZjeo+H2/rnUUuNSdg4AkzHoF0xEbs17gztgKpljxtrkAvWDit7VjQ
ktIOWLpoU4DLJJkWYxKvhYXJ3EXuCc2shQpOtqnJOv7tI4yrus9j7pUlw1U0mF3im9wYkMd2jxEq
L7bp2htutq0J3hU8D4eCgNs1kLDq9o0d2RRiTD7zsD3Jg8lTdi2tyaAX40XAUCHAq96/hH4BbJ/T
n8jgBFY4/9ZzGFs8kwNE6o8sYqS2rwt1ZTEE0/JEeElVhvIS4mt7WVjsdDbPDEDJjwlM98coqoSV
uKrGe3vcoZEhsWzseZQmvcTl3kcPaKNgpyaDL9NZk0yVy55xfCuXLDiG41u1g8BzlzPQ9IEidbM8
2oW1JKD6PbDnHtC56/b+ITw2sluJEkLHOe+3DvFReZ6lYH/kc5ThD56gthci1t4XeaKJMsRBjcT6
RlYrKBrqqhW3iXYmZTgPw7vKFUehRtZrG27kKttKoPTzf7gubk1LppcolbdSMuowep6GxAif8e2n
PGPJWnhhaZk4faRI4p7NJofzdnOBgLViSVv4GLSa3uqxgfRsmLVw75GMJ2aHzV3qkRmfVdEPeRwK
q9HDxQ6sT7k+9KOJUjFKyiYuwevKIkniYwjSmeVislLAySHyYrCwXQZG2dz/dZHNH3LDWgpxcofs
MgtAbOR+DU4xw0C1wWBbw4XfVqyXxf/smiRriyOhRE6tNM0XPY6w6NUVqNmkxt1vhsFMPnbo5k6c
2Nu5obB+mCvECPzn21e5lBAyfsM3Im/gWIHH0iNC+NXHxn4EBLHp/WGHB9h718IuyFcQiTA2BM8c
OJXSgdINmZhgrjej6A68a/qYFzI2hPm/ytIYvwSV442HjsXBSVOLcgq6jBF+D9UFpeqVUca3a+XF
ubYdOCpO7JWN++CJcoyPaP41Agvw3qfsgkSU4yHtGbf5nzVUBn8FB/iRjyhbffm6jy+62+H4czqG
NRTVDsyqZf3FZ0p9EkpCUF440vvDSgi22f3tQfIX81kRtzmAmZd+FfrNqldCY+cFUEkxbgwCYsqv
/+P+nUIAy9yFMu3GtV1W1Jf1PotcQ8uh4xVDAtow/JqdJETQRKuXz01kDBqyQOxpz5c0AQRsRlt6
VUiTWdaTqHghsFoOHZGHx3C94Py6cENDPFV9OTUrV/D+snIi3PCy9NQpYWGTnQVk2Ce4T3sC6v8W
C1d7P8KA90ASp/0v1MMiafdrkoRiBDy36XJ1KBxe0Z3ePMMpElik47DkjvKAc7bDLyl0N2EUhAcJ
H2nfA6dqzpVrSwLsAqKZi1rwuoIHJGM2NmR4SY3BqH8MlKH+e6DOpqsJ5fOATt7ZPpCTH1F1TbyL
Pkg6wPauiO9HEBwy2riWPcPQFUcdkjxqrEBVgZScbVh0bmMXd/dGYP+G36WVR0KCPpj/ofgiAEkO
IksjOtx6ZAdPp2X83LY9qMKmqD1e6LDxBEupho91TM1TFSqUOa5sFfv8QDIVvZrf73iLX2jqufsz
CnFLPNsfOgXQLryAX16J/0Et60kf6CMFtR3uRUGkBpjpXMkc1W2Gbk4yf7usewF98HzkZRpiMIbU
P1uen2HhFIFucrXtRiOT8mgDyp5TddWoMsGGt+zRgah5Rf6pSxbyuvU+xDcXgtaCTY0xxGFH0Thc
X2kKrasRuPY4Ww5e5qQ4J1DJWnzr2zWIXYIU6gJ7UsqL3au6vwIfdmkJIz5QcbH2C1oh2Sz6G7NU
CxaMuGzF5lSxS7qpTQzcBeJZ3gEsBtwVOg9cuvh9RO219fbzxj4zGttCLmTgtkaDKxvF1UCdXAeJ
GulzQuttPQKRoouKPAWieg3Cb7DXG6lLaf0m0m6YykZ69vfmQDB36yrfSjn4O15fValdpQQF0sJ3
p6WCLg5RSZIrW4abII7FkNZyEjaDgbgHl1kFO4MMDNk8x+VR2OGIETk3Rnxb8f+CMX5Yg6EvZH9h
puakj1IE5KmCdXYmqFlWRK6+zvsXWHAERWHZDbRuyZerYrCUhSxeqSkANO10/Knw+0QAD0z/Jgfc
nh/eSs/ShIFZp7eKDY+UCl18SgaHph+8+S21FluvCrt6Oeb5a5yT9q+FrOLtLrwhWU5S0/axr/Gv
FkZeJ6nkNwrreTI2HxvOcNFa0CXZI4Yr05GMVP0YNIPG8tcJNWn6hFlHjqO0dJi3C2Dx2lu34MYZ
wbWat+MpuLW875XrXkYN9wt9QLUeT2gn6m2bJJrgRfTQSW1Rd3FJ62e5QNpC5yKSLeXA0vbU69jx
vH6sAuJ4bd1w/zu44UR5+s3JscJinD3CHm8gZFYn+v8ZeHJzxM9/irgY16NFCfYLMVIUG2yS5wH/
qr5ua+9L3upueX9x2Buph1yXOHs4c+LTXIb6SF/WHyExF6xplsjIK+sYPBY00PkJpJhgpChjrH4o
Dcy9HZ6oGawAIinaZ908nb+bjg2mqYRStDfhMapCFVVhGWaDkmiEu/EvKacyN/Ahts0RXfjPVWYb
t6LUM+quL4CDaduCNS3YQQmMr8nP0C8FUsoiYQiMiEqrih/B3KbOywrIfDQUE3i4F/lHD33TQcIt
S3xDeWddU6qwq1I6WFCxjC9flDrUAdDK9auBzoVFsxfYOc1q1DLjTn44Azud1zSa+YFyZyPZcfMt
3Oy9PnsTJpRb3XoiTzG48Aq5CwdgxrJiiiJNyFGedrYHa4E2UGKPlvMfPUHsklYhUq37RRGJmZXF
aGV0IUcnSSDe8riGzdC+1a0Ls1eyXSQDG8Lrhd0/31+d/SEHH6mdmkbonsdH7XAPYKafdizFhJy2
FkQthLO3hFkDqcg6jVMXUwoXAHu1J/Z6yeMb183oo0IVhjDOcnv42rr5/ayZZ+zucbpvE2Zegh1X
c5AsTwj7y6qE60cC4Wazma3bofvak17qgvMGjwUNc7SlaLWADH8f8u14c1WtkuAoKkW1+TrimxVR
xQu94gwNeyxdHAboWfsQM4T3zez3bRsz2Xa3c8SvmwzDY4jqeem5qRcW8lvbb3oq1gDE31w2nBWI
0MavjzJ3uwMr+74z5p/4bwXnRIwH583ZG/QDHUAoH7ObvcMVNSou/ZZWx+JzT6zhUhF7E12V5JOv
2gcRuxb2caYohYQwk9W3sYhVUwSpfiQRGF0zyXe/6d6Fh0TbuO4rLHtpQTBiFJassddJdTaXNyVt
nyr1HVYmqWxxm/HATof0z7ORoprrNAYRqbuMju7M0No850cPfYDzGf9tuCbWR0Ok/ANURO3H01c+
fvjLvJG68e9szA7VZmELXtV5ncUJPbnF8jgW8dWV9Q7G3mEO7DXiolTGNucu3WCbyywqa+whEG57
/aOtbB/hJf/WiBPHlrqAkGkTdvgOmQdMUq0TVRnL6fciAdug/NtfKNLcJ2TIY4B9mTtTFpjobsX5
BvzKlSJ8/kS8mCIXjVTN3wRJeUllZnOjWQvw2gULFgvNWg4OTsVu6D89s5bQu9y9r1rUMaALaPpO
awDmwVtIogrnaXwixvICOiTiE0As4JINqgEVp1NI/TgtRMsbxtE6hXZCsb3TVmT41OMPlNH2jVx/
UYf6akD/Q2y3mFYTRoMUD0fZmg4t8rK7a7f87n7ISbTA/PlnBNQZ1MZhsbsI4lFNbjw2MNtQcM17
zxp4DD+HccFZr8+Cy1LUGsf+reS0M6eG1MdEkYM5MlVqibD+aqKDPyeRZWJ0qML6b2AgLjc4DPuf
Oy0K91t9GmbtIFiU03MiEicXVObc2phXkZ6Kc0hoaUp13VvkCG/2yJ0DC7rQxgeTER0tZpn/ANDC
jQ60bcmxICodZHJr8ppxR2csC8s4MkY+R6jXmzS7jNZdYvspii39fUi2e11BxqTdHuTk4fc2VZw+
kDZH4MJNQTvjzOr8tozHtEznyAm4BPkhFH6WDk4tyQ8DQUH2lH8oJBF9JyRBDuVqdmaZuOYA4m2W
DcGoFmKv8tutZvBf1apbQHVywntD4mY/QjOXGFClc4XbxrxCKjBQrx+lI694cWg7gwUH9YnxUA8Y
t4CtNj6/el7LFccoNYB7Y/+mqNvs7Op/LTmoJadkP2viZHiI0RZUqARO2hID8arYHPoBRQHRCe2Q
eFM+xuVJxbD7pg7jarPMsIXLwvKMqqSE2hl8NXyIbfQt+DtQYRaE3AITyAqyhZODPQbG5J56PJg5
hmdsZvtQbMQPHKJjx7J0zb6TCAXbkWhCJ4P/IizKtTe1XVX6y61l4TpeF/4FY4RZ1JLy3Lloou9r
1pvQ8CSoZbU4HrDHXWkvY9HRykBrhceG7NNHTaQzVE8qDupsQJ1cjb2SsWMIjdEiVfOITIIQWOn4
Z7f9Ow==
`protect end_protected
