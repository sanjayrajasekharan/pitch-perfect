-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
kD9e6ew8QoAtYD1lBK39LQe94eUz+su7GOpaBcvpFHi+fJwIFTEDnLr62eeo7JQq
8BpXq5TnW0d84GhFmNQysR1t8effzV4vLMRUz6DSSQd7+HCFb1qrA6SUOlqjWkJu
/0RQMjq5YDln7inmUOt3PXoJ841H3u4j0gc+qDlZEaE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 34704)
`protect data_block
nhrgKF3QgZlb1GRyIfN+6Ynwwr/CeNdoCjcMh4zYUI7Nrh1Ey2TY3l5pkzx8kFuy
Zzrg8AqY6D3Gv8vAPi2Z2w+lp73AjrklSP67nf4iFN5DpG28M2gxDF+6CY18MrWm
mg8KPhUUGZc+Yy2i6H1qczLds9hS+Wvme2p8WHgeNdN4nFkk7vs2BSxjHGFpOnzh
p3F11LD+0J7n/r6w++z5+M0mmj8xELc6sQJQjBAEnVUvwGZD69ec7W/9Jomtbv7Z
l6ehfbUuYKnd13DF2iOkN9128Z5fU/vW1RBeLY+vdHbCutpXU9Wjcs+o26reUXHJ
knjK+BuFAnqGh7ZRI9HXNSmmjf2kBF3aTPZsUX5E0+12xKr7texImSOProUNXdM8
seoUNXLgbmsCrr41t9SamiM6txo0Adn7D24nJbrJ+l9eYi5HpiUYsw1a5SS2Od7G
99OfF/jBq/j1aKHojyr+waxZRQ7QylWJsC9kDq/j4pnGtJptNAm843gliX+Q4++z
bUyWtBRRdqGzvrJJreDzh9yv24Q5/Ak0Xispvxcs3hXSoElXMux9A1D6emZopZJt
2poykhLKUFcL1CX60H0lv4qFJdIWc9yV0VfNodam0Puikrcyg3MvXHbujeRfnpwJ
TiGqoxPSQOcvqyAzqGRyVUtkYkT3Dsmls3DZTha2v/TU91oVfYIYma86a32zGB++
mTuA6mCKLmA6Ag1E7PQb1tc8FmKviaGT+i4xj1yDj5Fo8kFXCiQImMfR/mUbamkK
5yYA/fOWNhgOvGVyrX76BR1BHGfux68maCxFVIImtMSk1RRxz5gDl47DTwEBhFRf
tp2y2gh2xUl6ZvZkRvjbW4BURsriAGbJ0c4CqX5ED3JnPakNF34y/pB8Fic+gHnw
sTZ+OE2eqMSlfqQrJ4ZHaSqm5Cwq4AYBnPyRU2tSC/FNAOnt9RUzNbdcp4UeQSFY
4UIhfbggkmeyjb0IQgKdcixOLV8b5XeJK5Sl7AoVu1SoNsJNpln3gqZgXsR/dgfj
F0TzO4C78MCeu2SBGgmgHJxdXpkK2pqNCH2wRfJ8CUnrzb7OCIlMhKuM1S2cgtNL
xeXdBxStitoQeQVcA5xP134cwz/UPd2DLbBG9ozvLJF43z1+xt2/D1Nrcy23OnWv
3ORLkFUA6K05sPtWHbxwGzMjDixbJDSKirAhDASb/J4/HTm7mUt5iTGJKGxwMALo
s+FhbwjJjmuenS7r+gVVskNedT5SrLoAP90tGTY7mPBPngPPa6/RCIMMmzAhu/5/
l1AyxnC58eIK3dN5SNub+kPTRe4arau2ny+tIL9t4ULLlEr5AV7wW/GilJlOhdG/
0NeOPygcz5OZQ/jXPyfnp2rDpRXa7//JLANpjP8iAgaRzWWDQw7cOs4ELjUC5og9
lZpX6f8oZs00RXPDPvZ7JZsE8FkzcsDvp84alJZdb31bDhbXJhk5fE1EKVDGziOa
z1LMIxeDGMKkycYJliwNjj2WqMmcIRrax7pwvBoPLXjpl6jg5cYSBkwlqWEr2bJk
LUcC7Chp7a2JcNYLDhu+yvH1Q5PHWLz5ESYnn8cccdWYKFfYM7613Ycpn1GhpSpp
JTgdtoIMW0cG0r0dEHEEtjYvBTEzML1Tw/v9AgUOdwBfKHFTtkOduPOyzRcFEuPq
huZSmJ77sTGXq8iQnqzJPe0wbv6bTAA4EV0B6a4UtsGjKzJfLw3cG4ldP8RZVfM0
xoi1dsZK5Gdnbex9E1gPExNm/JAHMBftfK57W5sMFvy7ucB//s1Q/5w1iUu0E5UY
UvGEk6gT4nyIHuKcGzwZ7nk9/KvBYAQQFuuGCKP5oLmzHxXVYQWCa9M5sliLPYVr
tZxO9NsRselH+MXCWeN3UwDHjQxNDNyjtNSn2VUGprTmO+t/zCF+N3Tj9Dvo0wn/
gn+u5Fj1MstDQuYVPT3M7TOvVPXSN16F7FWD7khIJXemzw2DDgSaH3PLmIYZG4RW
KuGKl7kWJ2WHAI0XyFtL8hNlN63YqRuY+fP3S9oDQy9gcePEyezn8/+8kWsqoTe3
YJFA/M2MAuP9TLs8kRRCZgTUhXgxovrw6t+2lnAufOSVamYKECA1BxPM0o1SBcEr
SHxYXovankcgFkCPzHPeVlJVLSJ9KPe5hsbT2u+C5Kd7nCzJiOTcEW/4wzGs5UVD
+sgvqAXmy9scDGvNwt1yqXpvrsJPhz8GtnnGKp6uB8ishV75UBJk7RW8+2VP1MLf
X3XRv6TQfEEfhtntpQhVz3hCkML/OHbmGz9AuXrbHF97jdkpcPtR2GTZYsEuJFU5
fZB7TDvcQTDzg09CGhOZtEMounVIX4Oeu+gk61a5ZHig230+5H623JfqrUY5aMk9
DLakdMrXJUP5Sym+yyyJdGDVI50kTCTKt/aQODxIjpLAFog9m4EnNhclcI+xH7cw
191nTl9DYJePcsdux69K2DtIboUP1C8P3whBvomX0neGpllS+HqZYuKpMmKDVS4B
G0uGCcxMKaMDiG6gVVGoSdB94WFULpD0yyxhYWjBkEVBnXT+VduDTPeI9TdAs7s5
t4cUFBNDJcFkwfpS3TBuz9a2CLNtfL6zLudRBsw1iRH2LBCVCZyITAMK+ADsuvEc
K2z3gtF9DL21sAHCYAMNly8Xo2ULujXLxTlw7qSgoQHrAwcZS9dZVSplmcBkMXED
ytS6hQi4OxCEzM1uXp4kV/fBgS4IQGeS9nYYJLurRus4sSFR/cWmf4N8bgtBTM63
i+l0YzLLciYxO3Wquhi2AqljZV5G886WbVXWlER6XNCOP7mfi2NASQ326SQ80Cmt
oGnXNEBcqCwEEQNzDekvMbbxaeXzMXVf4NkXM1vkeCqUSPiG8zoyZf6jvw7Uz+as
MA6ZQruUklhrcbnD0bc29xwv3JDY7phKJcjls/qsIE9DsURAfgPj+ZoXNEYpmsMY
By9Ij5kVZIZ/2qmuNQdyrAWYUHHg4encBoCQA7wU1maUvsk5KlUtU/ljJ9Gae8VD
E2qbdz9U9DmK9YZWntmpjykefrFL5snUIdsRdSQQ7T8v+p7hednEJrx5mv5z2PS+
i3eo1UAFaxmmhWf2FcPZ3r+DRqyxx96EHkqtuZpQ89KiubPtEvzQV+txab5pZxlq
57sqaLo/2dF1hcbO9GlPn3yfVcTSVNhWzMYPbndr2Zbbqv4LjmNv8I6uP9mpE5Sh
BkbDcNWj2HBh523zOxPofS4g4O9Nkx13es1uwxZ+t7djBuq2Dlzpab0LjSaHpJsf
kzaQvNZdYS089mA55EOHm+L9qT5j50VKDU9FNwSfWeLGBe9X+u1s7Mp+lZnURnzy
vVAf6u1lRTKbVQuO0nS1lUye3qBM3cNlPDmBebqkhz4W9ZJ3h4gsirb1Ro2SsLIR
UtR3DMnn255t9Z531EL0zOXgC7Uf/RMOzK7t6StGwcBWGIzIE9WYh2zVOu8XCu3k
rJ3/oNYvqqGHu/If0xnkKnFXgIJn6bDunJogslhLS8U6/uEhaKFDlAJTFjXWQShL
sxY1GZWgW68P/zwbNLKHub8Tj8N4cYM4au8gu4YsePfwp4dz45pXvqepOqWFucIr
//qvwwWJYqVYo/TDYYEy/IRpMHCLMfPKTk9peTDe5oNRTkUFcomVaLFRTjRZSGQW
Y8bldebF+T+BQo2fW+prsc42bxSX1o7tojgAQtGs9OqUeqDTwkg7Iq3NCZo5GgNp
MqCz8s17p8mAMw+P0NGsJ7F6okiilSIFXXe2IdMPyObosVQ+F/v4Kw0xHpfe/Byx
tYYbiEPgynTodwCMyq/nJzDduhK8zZ9ld+hczKWfeczTSULbSzzTGEkNzqLTHjte
q5UlkaqireKlBZtU0aedlDPRZFyKFh8Uoj4jo99K0LzPyxpmtQVJp+IDGbiF/sGO
TAuYjMCBW5iqIpD5OjB5AykxyeSWDEmgTi4H7sqJzwGg+G9VQVtfHi0PFf6jTLHX
0zUEfvDOXyC+jqzTHNNmLbWy+awx0Ovv94PNlpL1SwLyseZdYsCwd1IfZj19IpVP
4gcHQUD4oTBaNN6bmCgHwNgtI77KSwEGOx9nB2vC9oaFBKNKTQ53p5eoYnjmqw6b
gHPRsvXFPt3yRDQn7/Ko2F/UY5YsL5HyLMMwJ3gVhGLI5fFLQUfKgOSHhtgelRIa
9wR0EN2A+iURsbnr+nPqkSP3T1XYuui9wjuu6TFff02VD6999qWHmnFM7RfCI+Av
SFSaIAA1A5zQvU1kj/B2IR8J5/DykNPI3nBf9Hfgb6xYyuqYqubmk0Pl6M8ZkyMy
zXgLype7XCNNNhNL8fxPBZlbwxqejDnhtYM0qlzmn0pDZWY7jPNEweQ374w7v2Xu
KzhWdOrhnwXuE2wDAdq9+MDHNoVWTSYIgYfMrekR3XvAqxgKYhkRRX8+0H1KSlo8
JkW1NPKSxRjGgxX0neveBqhAgST0bdDpd2574VtY7MZkS5ebBJ6xZkSx/CW8cYzK
pD5vFUt2di3qk1dImoDEqt4xztqo8gvDl1dTTlHq3HqxxufXJZRF0clAae/plvvT
ajF2VoJE8xsbO7AAISBlFoBNgVPiBTbhY6a2puorV/NqPVybuobYNtQcKuLMXJHa
6APkwpsOxyiQiT0co7QMQNpivCxOSp631FvhkfqSmsFinwo+XRK3GvhUA42WvVxp
rWDcsME0ajePTJTHkZjULMFAVV7Oat0BwKJF5GqYoS6Hp7/j6z49TPgGTLCbl3Bo
iqsnURPah2cD+NIMj0r//3LDtETOay/7sWD4JFtoqUeg4iqc2G2fCmS20+eEJwui
8hv4P8I28C+u7f374W7TdlZDEwI7md8qcIE4RsKy1J8QxiGyuVEqdqhBHJIL46+t
t+PXU/HqBTXY8MgSsphhB08yy1hrC3NJVTSbW2t14eLGJhlebpvRgWFuc0q++j+D
vSq8eDefrw+LvLOoG2ulQveer1f2T0uZLKmZQzOmngGqPb6Md6WsI3DP01rVHHc0
Bo0osqcgIbrQH3VYUMP13GIiQSjZXSouynlEWYHZAQ/N2q00nta7eTzX1itdY9XO
4ZuVy4gGO1RUJs20vQtw/+2lswJS5zjP6/63dd1wLe+71TVOI0K2RCDGvm1f0dwy
phxjrofFZsEnPw7+OnwnE+doaIENH1hKSz3t6G3hUte42zY+Rqpzj7CDhZwXq/fv
OJpiCfl6Ze1/QznHPsAb5lfB9bn+/vlGNrUaB86STUJ1OS9qEQ+3fRTUe2spPRJH
joedpgWhXdwn+agrnQEjMumCBLPLcIfCxiMhKpjdnXhExh5C+hYGZg83w8ezsvAz
OTFwBEarWIxn4zvw/t558Xmk6jpSj584rrugmhwICoHi8XP6tJEeGdRCEEf5D5Ep
BgzmqILwTCdVaSPcT4MfKrSUMbrcqj7NtLU5+v0G1a1QYHUH7jmjH/zYRKHkvqMK
YVH+A81c70yt093EBAoKsoQNWFXYhoyqRggDtVryT/xHUKllLEiNB64tmg5A2JGs
1TS6xeBBsJFQwsYsDoaxXf57S0oTdFnl6Jh4hfWdvoAPJOc42heCG8QNu3hVymrE
7zgKqa3TyIDv8qGv4rhEuEsJU7/PT2lvSV6QoZWtxWY8S6yFGiHsLPLoI5pr66cA
4KG7SD/4QmyE0U1gbMlrUncFmtzvl/yvJp5hOMmDW6cZJCwMxLQ+vYDWJGrdYPue
Y7GLAJoxd/z5Lhoawj+kcI90ZoTq9/Atg/SIaJHPQjxEJy5/1wifXXv0i1RGMSd/
BAwUPpZYGvobz7wySbZtKzTNyAIHkKpwHsQYxslBcjJCM5MV4EeMAgBwGUlO6Q4U
l/4Q2+uq1ymXK5dNK6WNqo2kI2fN7aONrXnU9zHMgB0udQw915wNQznrbkXf7E49
h3A4YlxWEevNJSMGFntBsj1l61PNWUjXVMsURLkU2Gcvf2a6Eajt4dyNz22PyB2W
syTPgPNDydPHwsw9WrAIKwKP1wQTSzMk1kGB0lu9kDAAwNV/fll0XmiJhF4I72Ei
Wi73JG9K/H/mNG0paNAlKp4FwaRsGzs0U8suSal4rGGYNEWhP57JzwWnwNQoSpxR
B4zk7x4Yj98M8D2mam7HjRnuMUiAJwEocvNy/+hvglItpOUxJHAxihnbVtfpJYLi
J5WYPqpqfiwBaHP90GOMyGt+cYeDP4cCSYmFE9oJhYNIxVwFQCotuO3CkDMKG+8K
mtDHlZqjaTAWHeKMiJdYIptdDpZPX7FUY9N6lp8lCxaAOtsTd7tkTmv5OrJQK4Zv
XgqPxkqxXlgnmQS05BZt6yTqgUQJM6a4TZuOubPA0+BCFsOe8NxxputhpLxqc6NA
JV83MyNh5DuRamwWtX6d9ytrPbpd9Lec5aqktrv+X01xE4j2mqD5Y6Ms/G/Z6b/g
+NfF38lHOlg7ur43TaghwKq3Cqvn8PQGUVnQNnT/5SzkwepQqPa91UemcIWYGVfg
ZId09LXJUJxouBv55+OIlOIdAIolfrU8qgQtp7ZvZTvHftWPQwXExfUI+M9ifLa4
HuO6tCw5TuJqwSLEwJJgnga+9EDJp/DpEVe7RDMQqvnSEZ7vX3AVGfjXNlzNt2+R
8mIkJ8GxjLow8qo0Jwe+tduXgm2IrEVciPOOtBc7vOTEhi8gr16fHnZa1BbNqBPN
THQYvicEfl4IMKDRrOcXoknVbYz0//CnOPVSmsYia1KGHPBkzk2p1vSsUUWooAVq
9C9KQMhX+JxnBXJEr+cHMw1QqFJ522J4d3Kph0fnrwOtMPpStYaO8tzeCQpuWv0q
G6xQ/8aeg+RLzlk+eaXQVjTeICHt0vqX0FSXoTDf2zO27uCo6z/rEdKbO/6NtGzI
JTgQKkYcdRJtz3sPi/kB6z9zCbHRdXWpDH4k5MwSyqZ/mYJqs9HBVlCL0uu4xKSR
9VjzyG/muRSGiuWgqhM1bYXzdclq8GoOJ7IgNKxpM9MMWWoPq7BreLc3syFYudjb
CjTUQYqbTXSY4sD0hI7b8FwDKEsntJieZJVhdEOO27xxMus4VIn1EsjFAgnTcLsU
X+mMBVzNq5jEKOH78djWPmlfV+PXO0t14bS7hp95DV+ng34roBPUogFBVC1MHFhb
XYz7ou4W0Z3CLvBunOM/MK1ZYta4eOVjk6IakyQXpGaygRH0Pxu8qesA6lAK6qh0
5rEPjgrqZPb1pCyJtSR7RH9jqKm6Q28t5Je3NlEWZYRqQgcVbt3duYBUndnVNnO0
q6l3AtSsSmPvPNdJlaqlkfZm10gs/aiHyEiiNwnaQFVJJrMeXK6iwEhVTCAf9KQ+
JMmQFNOSeu3+QZEH6mRKHEA3G7XvZlMsbCVzBHEEN1KBEIC2daGRfV4P5X1l2QNL
jer9T9GAYvYwk61oMugDBnM/+ipbh932kTQJj0tn4/D5+R3IsDoaSuRZXXaayiNL
NdL1jcBcIzuNvZi1QbWtEQvNeTjxbDjXOu0NHicgg3FqrTb8GUBBz9RO+QvP5R1Z
2VZiPmrETzXbKO1Y0ugMv7WTnCsJy1Rp3k+mDCHlEQW6e1Q3V0eRhj/C77AwXmB4
d3JoASkkPIwulzddxjxtLkr0OlZI5o3ijwxl2azUM/BWdlafeuVKvYVMS4D0CDCJ
50o1an/a0agCcasUns6Ecvqg9B/9a/uHhqFWk5idJ6c4chWUcrMC7OHcvRvpSpWU
tFfa23kpMVMu6pGYKOL8uuYOWigBOPdNrBsirkrEk+LtBjXUtGO2NlY5rKYBlB0R
ecf1GoNRRa+fAcvKstoi78bpLQHJIuFwfU8cUcNrLE0Of9XeB35njrB0oGsiSZcF
sIz/Tsan1tudgLelxMx5ChpWxohDDSUHVQi+Hjw7jKnlf3wAuaM3vmCF0FoiS84G
8xYYfeGj+llrmZoHqdsHeVgnowac75jGaZUqIfj4THXFbB0MzL7jdqqfCKsJfK1v
FD8HXadbPUBpiErfGPwLdXcwLF+wwHDbkfSw3xLsGXYQ4lhuGC9RBMmd4I2EsUln
eHnXw85euqn1/6qAQexVJT1ALVWx+5Tg4HJOy/dxVgGzcH8oYPjX8wTDG+ANmGAK
71+p+XIN+K3QyQvjiOSoCmMcS5X0e9FWWe4KInZYSLDjJMIu88uooiYNFxVrBIfi
8r8pACEbZoljNavHlr/Z6nms6038srMH2dr6pcz8wF3tfyyKSWZJGs0BqR48JRTf
es6QEQ8ufnTsoEgQOYmNjz3LQnCSkXSBEMvxUvSHeFRqwn3Qf9g+0pCIgLh67xt1
7mpuj49rvDU5TcTaDD5Vn0faV9+gWUs1KAnne6LhghP9skePDhoc/+dYWTOb3H7B
NrDrVFVDdnd3OzVlbkYyCsK/UqVf+TPNCHhpLzqwBfIPUE7Beb3eb1ZkR6S+n6jJ
pOoGjYtdGyWGyD7d5tJGZC3lcYio+VaYwkp/+US1/vuKN3v/nP1b04LlCqtUJT3i
wAJ87zu7zuGExzgTDV4jOB0qSyMBh6a7TVgJB34YFFkkOVt9lpAfEbbeD30CVRoV
cT5V2CeCb2+YUNi+2cJzr8PwIC8hez0N66v3Vew0ttlK0Rzhb+bb4UAr8CDSOVYC
aGHkzo4zv3ZqmbkZ2Pj8+x0VrQNQlY54NULPgDAKRqYtSi1cU0O9Gmzdiem7E0j+
di+TY3MvECKZMZ5F2e4G9sdeoNiFPshlyRQtv5flb/S3506Yf/Nnjs6B6auW/747
XxdLuM6LczUA/6FVKaY1NW+dEfb/d7cbKeQ/A3fr/s43BYH8ZjDnWE1bV4rSxg+c
Jz3UiJDw6/Zn/A0Zii7Yalv5lEf++cyOIOOwp8GAJp/qJp8kD1xoeRrJJBiNIrHw
1PJZZARpCsE5CdgtneorK15D9XJ/n6DDyERv/C3LWFnt9kQB1CL9icfH+VQV/8Un
aLPKN9DSigGMsOnbfSmVhc56DH+5TF/yRsIW9ldAM4ecXzvryZkTj/lixOQ3F47/
rvgFetg/4YVxA2KaOpU5XJMPBfOpjRFPBm+cZeOEVXMePx3B5okEqr1UBGrJJZtG
0RPOo/eFp+IJmIldqbJ1BmWTD9uu9YIFNCWdYZRg0uZoYZ2CFT8D/RGcd/7M/eTs
cjS9fFIMeo11UcYkSe0J11f6p9PJT3r7vRcybLSu0DVfa3LZXCHN+mMpumnM293E
9zcB4vc2FQXGoyiCsagQ4NRcpxoomvsjSZhiIRr+Q0e86JGucqTazenPwcb4wWbO
1SE5GJX6y8Gh/rDT5b0W+nSgLgFYykf0FPR9Tf06IU4++BgdmSBgOUzI3mtd4sID
flwMSCqZyC1l07iFANF6hOQdtbwZxWX8Kwmy04ew7debser7bQkyv31zm2/aZV0a
nMKJy4h2NkPL5kORwM14k98qHbUQLoTrfrqLYtwQNnziVRmRiIRQ5UXdQr0ZnKlF
/coh+hPBG0R9Elwdxo/VOE+gNjj+haIfxW8wTB60UCAfU3kQl6tzJwroHjoD9u1i
yhLGjYlGZ+AsPH5YQUhK9T8VV9FO3yV+g/DPji5hOu72uraLU1E3Uo1oGHxkPV+4
tfo9t3CBWslxxbYXNIufCd+XdqfvnEVHKfD1eJMfi35B23VltToQTZy9b+9u2FmW
UgtreKAChW6ULrySgnomKRs6NLm8E5OxcTuSpl9iWZ+y9DrFylhWKdESRPT9ix7c
4ihylq6bO/O8Xl3DnVqgTj2ouabjKvPjA2EcxUxHuOBBtyDKc006UW6fLmSWMily
DPdxomP3X4GTdXBQu3ps4sd780jZbzUz1ypEULAv9p37sdAvrRr5nZUWm9WsKy37
Pq4FOwfNfZ+MB3c+dA98CEIY1tgL3X0tnmVfqSZjB0J9hrlMp/tgCG4+KCva2L/g
MYwntJ+QmGrK6UYOWM0EHQWykgtwHsK9oneq4Wewq49I/fD3NC7XR6qC3HHDTxHA
3IUKsMvh5dlWoLWvyRNKkENN+SryYzF/lwkMlGxFTqZ52QkA0Ceg1q50r+L2R/KK
fE/keyARzp8RciNEHtfPSWTtutVJMr3MgY+eKiof3TO4Logoc/2lYq5v+LnT8ueE
Q6w3FgjHfNvZiZZQQYm2xbR70GNaQ3s+kUgOamRr/pmiZAtlMduZ2TFfKmo68mG0
TInBP9Q7GQejTSR8+PaJuzr5H18MqSYPf9lPSEICnvyMvui2OCUXWl+XAXGDJvfc
uMLVVr68gv5C1qGCP8PrW2WJT/7i/ftH6424ZW4ExQAGdtkwfHdqE9FokURp/1XN
UZeConuKjbvJGNQ506rXRSz6cU5kCndQzscPRg2p1H0iIUGgXuIBNGzFau9nqD5Y
M9sO8kr7CH0Uivr5VZ6cxY0LxrrAWjfT2pKvff3ZPeqOvJ3rrl3oOiUjYI4zD1T3
Zypk1IsiXguaAC8IAtI+vFc9sfI07Cm8nqoh7mq2gN7M7SCBZHUGTt9VXJkcUrhQ
DF4dnItcePuNvrzxtbd3lO9TVuda42k6yDO/PuzPgz2fj08FXDguFzLWlswoHbla
mIwwl3SsWu2AiMZPBWA26mdo6VS8eTc3o4u2cTBil3mN2LdFB0Ys28RcvJ3YBDAO
2Tb3zku7Ubk0xGHwJ3ciwTkfhRH7StbYfRjPVQWdxFRrmdktIfHgssErwYt4igqT
rRZMYU17xKMEnOIoahLrRka5+GBeBErkLwDvN7MFrhmhb75Pzgrjq808Y/4wKNTj
qXFBCx1eELFIBH1VBNqHLsLO1nL1FrQmt3+CSNKRRdO8E1GkHSmWQKD+8Gqz1038
oxwZaB943wWQ8O2h3pFj9O7LOkT85rV5Yt+A+WW7mEtdDOZ84zBDIgwOYkGGDmjL
gKBFsfx4ld++cbLIrIkdFDd+x3VlIFVPvtk4u3kSFDMgfDAOAt9GigRu2yKXNIoQ
lFboLI0dF/fExyn2CuK+K5+gp4cvT3HlwNkbJ5/gakL5Vc2HWZA28HedwslYdpbV
RCGJSBO/PFSZrbZjoNMDZMdU1sXSP4z+uzwDnGFWuWZkBZKqwj0VBLnpIDwxV5tR
kSzTcer5+R+tvmCgzQrF45zTo1LlUKTPfMmwpCqBWQM1RmO+8SuP094VZkM7qFZx
yPJ/uHQheLXixVBT7AxjeMr2XVE80g7la1i/XMuRTKaGMwHkdwFy8JSaO0aAdU07
4d4qNzS+wEiBuVZCRAzMjYw3+w8M+kSadfDbWBu+voDZg3SaJR+odR7bVm7eDloo
KD1Tbg4YEtkNLOFeCnxHXD3cUs5EA4+uVTzgHVX3jyw/ump5A6bkDnFHXfiWimH7
QOAmjj/LKODo+mcihRBpz+X5bsbbdu64On24d/wC1u7pZ261tpStGeJpM0YG7P1b
C89aMSlmxwTBowX/pG+8mcWu1rSrUWieIMw6XwJXCIZQoQrdFyxK6fJwLCufDYGI
VXqRUgedfgw6rHVL7NgM3P6CCnITgTe7yaAIncYHPYffuPeqCq43nns1TLrNUzcC
Fz57S34BBb0/8QQaxqVTwUodbrR+UHTbZTlx/Oa6AJvGghjdICUyQ+5/clTOqwPA
QLlk3w8w+coGWO6TEo0xrkuyVk7CspbiqVrmVrP+uF8vqDcBZnMJdAjxfwUzpxqT
4tHuaFNbcqUeQVgPib7A/sc8BKRHxDETasmTQ2LuO3vmhSTv+wMl5i3EjJe4A93k
dnXS1hn3OOhJQz7X7MtzppXpeGBweFPc/PAJqJNwW4OJMtSG/NkUOTppZssxhNPD
/NRY/rZ1iX4AeliNOz7MB4n7yjC0x2FCiZpCjkTAE9N2o9cX2f1p9Q6Nc0Y9WLQu
r3hrV81MXmS/NHpIYVf5bRF8RY0TJqA6NH9BocVvlyiL6y6yWO0vrc6mor+vC4HN
t8trpQcoR7g9t4TdiI/qk6tWhTUAmUn/px4pbte5l9Rv9NhBI6janVIu1o7hDWck
zUHx+DBxMQykWmppFHxnw1mMxKrWwyLQ87uv1t2HNOpa1rL60hwEnmci0JJlbo2R
z+timqA0PU3+55MK6/CjmCnyu3/WE6nUr48UeBnD0tTsek8fUoYrs4udUE24Cs1A
8ovEhCxEmTHFjIqgWrhiIU83ySPwJQnwupjPuyzO23CWuadPuOyloIIiSOh960sf
rYz6V31PeoAKwI8qU9/EhIw+eU4JD7Y/yzniueAGEkNE4/ulVfBSMnlVMruJOr4e
03dsKat0kLYLyD6Qf8WoYujJ0DlwEVWHMJfgdDNcVEpZ8xyaS46vwpx5R4jD1+Pq
lUW7Aesx7klRInROgVficmujSG1Tj6e+1lXoO2PptCrbuVH4Z6+6n+Ta1qL9fMWG
Q2u6QQuXZHFjRCP1SGAbF02ckBRyTuzRL8VRG5sPERZdbGU6h8gak7jDQgGVqlT4
y3wAGxuip35LzBBkbWF8wiMrg1dEhzTIDuWIHo9ZnqSp5Q7gPuy32Ne3ug2iGW0P
A4AjAKHcNtfHWIcCJhJIxbnW0Cw4/5ekemWIdDo8mPVo7X8D4T7iw5vHUy7bZJln
jhiueXE7+RrdMUS4nqgXGKyM26LRnvucmeAWQOuv1xqE0ajDIkAlYU8CJC9J9r5+
ztHTjN0XlFHf3YAHrRHth/UzoGH2UrJSNG3S2Ct4mgI4nL/2rApCIReq4bvbmuCt
p16uT09sHbAqQatCfWRPiy75LvupszmGZ3x3AA7e7Njyj0jUalWyytobPZzdICTv
Byhd9x/+6l0Xn0+PckMx06ER00nqTOjeuHcrj26ZAr2FnKWCXnw8MVm68UtL4Q3T
6bZbSVl6w/odK9O1Cmbhd4Rd/OM/g2hwuYjnUjYZnxJ+xcAS9ockA1I6oyyrlOSz
Le3qhXHpS7WwQYlt/QbMv+Jw4zM7Q4kwluz017+QDKVVYqZMuS+wlSb648GbcuNS
8CNocJP794azYzRkd5M/vLOm6Tr2zkzPZBb0WJmSwlXUOlqg4U8cXOz+VMqe/EQh
6A/bqnvv6PVvm/x9xUklcrlI5MMFVCAFllSdIEsginmVihCiBObMDo+OB6htgHBb
nnR6LbdtCzTrVOHcKmZDWsfbhLlc1Fso3iTFVcTHHZwFqp0BLELSTW9NPiVfcCwD
q30s389oFj+O4h7pZQlKOiVadCGD5HpWrB0nEu7FRxIBx9b/f5R439Amvv0ZvrZ3
CoFstS42N8TZjLcaaqPiUORdb94MRIkBB0y+N3eqcmXLd7J0jT1ShgExT04cxFjK
7aUJHRqNywI3fMhu3EuRIJ83N+XLEadOb44G9e5greHdoA4EeX19WZDS2ySeLhKV
Q4vSrV6cdIVjQi0j+FgGlPfVhCUvXnR+OYH90KOAZM6fAfybLP0/KvrCaGT2p7Be
AHrFAZJFduDnKnJm5NyOEnOj7zhY7If2FTb8xsrfqDrnYRkoke0pAjjGOXCtGEGS
fKyFGKz1srhpJNAt2TEHdHLImFqKsg5vBG7nNT2v6C6ddcm9lklrT7MxcVZ3DJUB
Q2xhTezKBLQd1xoIhcvG93+yxp5cdiP+GpqU1Z59pVp//YXf8MyJFW8IkE7/m8/7
W5ScZ0X+RUIwz088tSDghCMb6I4EuPPwqjIYBkvt8iMjZ6XEN8PniRNsx3aAb70J
8UPoxDde+c+maIPZyOa/WrzGiGwdyZlRo/BtdgstTWXpudP4VMFeoJEhgPZ4zjYV
9sreTvIyeyiU8A9Dd879t4I4eZxFDvcsotgaXcMEVH4dzV18h5/2xg1rrQ51Y+uk
qkYtuY9Aemk6q3hg6DSSK3B1Y01tt48G79aX/Yz6NuecFsRWY9Tj2EkGlwXJWmH4
O1yCh3aDr7u05Ghidk1YS4K8VPk7UOOmpCi6i09nXQyHkhdunsRQ3FnBqXhxFJ8o
tHWQ7nbRHFzbzT6qEvgrJ7wXxgtpyjuk5jbICD9V933MCrKxL+hPedAKWwgVBV5t
MbHsTDBaPY/kfZs3+RcgavY6nxVL6DE+2NhA76qLc56PxGOjkAq/6IQv+6m4n3Sa
vRFP7xOYZyVyori51BvUmsyGcNHBnNVrACxUyAnZ0HZVC4Y7iI1LkHEB2be1DXaN
67ssziC4j+1nHosf7in/GcGpbkLMvcbIuxFHuJcZYCWqeZiJd5Uf1oNco1OlxtCj
3e/7M2XAUQlzRm+wjSTiYMUABLQNdWwjkZ5AuSiqJv23jdMR0mJy56vSIzg+ujGY
Lmr3R6fszTpJtTXvmNm9P/rs8hbaixUYMqRiejjBaVsrhIzWNDb08j4YUwSNVIiJ
gxAJKWSuInT8PfJEBVOldPSgatF+0hAMeV9TpUpbciVXdppqBTiKij73KznmvRLy
szdo47r5WYpsdVcSysiD46nxh9HG0i4CI2xoLnCTlxd9JTUkBf6fxaIq9lzHSRsG
fMgRrxju1bUhIdv/dx4Pb81L9exn8CYtCR2OMGiawpEdkMtin5Oj7in2LPfrlgdh
eTA1Z//6wrJh/PJzdVCet5v9PTxIwVQPKcCkZDzRPMDp7ft/ekQmyFYeCX9vtIEW
kt/SPMO3XPhlTggUY2/E0LoswT+JylIpd/L7R4dlPUjKJfHGN5lVEWH+H40KkzRj
+K9XyeNYypNS2DFnyke9375L/jEJtNoMjNsgL34pLoB/vZGyUG+Lqarp3i92QUry
/OseYKOIX/Pbr/6QAFBdJJZpL6J+oiiIOiXaDBcMmY+i39hBwuSsrNSRe+Djp1M5
8TPUu6H/eRVdElowgObzXVmkLdrJ1EPU6C9RX+k5LGrPMt1WW6Nnj3wxNReJIehE
0KRQNPZKHhFvydDy824PocYIuJLSkHxXp/ZG658JdzmYDXCq1iaq3GzrDuYCShpp
oVSfqqgSS32D49UFKbhiNnJBNFGIHwHc/jqLV6vNaSAfLiT4t2F16K9mFEg9TJbZ
czq++y7b4W/Xhex+wRlyZb+Mxqsne/MpjFPgdZNSeiuLrLXKx/Xbxd39unFYbxwh
Evabt5rXbOfYNSpzEQxe+a6h2G9OrqKKAeTL7a6AaaKEkpSNPHbuSgc8rH/EtD1D
ZCNOcCXXHi6RTImnTQm51WUTy43XnbcUg8EkQ4Iv36fDAuXeukl7dH2WRXCnXoWo
KaAuAg6JUPEMt+F6L2JSiMgRBfOIh4sniczpx+01tNnao/31xGe2CNgfUh93jlN0
PaBH4D20toXohhJzQqAuimuy47aAUlT33IClQA90eI0pJoFQGI1KhCho5wVNxGIm
VDmyJ6gZ8aZTEvbL/9a0KlPsoVGUiGfd75HQPeo56+f5OC4St8cGjvmqI66KIpyc
7H7tHb1hGXH9It9okLir5/UP/BPX5KeZac8VtQiEpvMzGXFhZWvutRR30XFxq1ti
iK4qs7RVUNdJMErycPIN6vPoHnThyONM0u6O/oKBqCKH4ri1CaYNbd/d6Ew+3oIl
hnLcxV+T/PViHa64Y8VxjhvQr4Ej8EQe2+9prs1S5GMHOBN132C9gxD6j0usY9tz
0Pu5Dnk51pqf+/ddqh1BJ+P7s2bz8AnDgV3DBcDXpgmBB8Uds8Dndgb7Hr7vhZVE
dpbgSvJOl5IqEIApL8Eqn6TEuMqIOmTAqPiWjARxYPDInGh+3toeEAyqSF2yDN92
BlpYLIB4mRXdWGgKYQ1Sr2rTAlNx87FxGsZ4IbszRGQUNqFr/H/TpQOdQBexClDy
cMtcWA4pcLhEQianpHXoNTleM9nFSdoYHbM14XLPRXIH5PkmQjQUeVgEYdM21MlD
LOPcJWIieT0/yi1Q6lBU6mdXoY5+r9+kklnh/lcZSzU3MY6+YLl20dClqi7PQunf
CwCl/04Kqh3RK76Z0oh+XN2RZ7fUI5XJXFgVT5poXS7IlNmvkobMOvs9Spm75qFH
wcePJr9OqbaJCmkyEEjYvyQMDCMdMOXPKBYNyWXNHDL/gN9HcTc/9siTbufsvgvz
AYfdJxBdbdBK+FaFcdO1lsSbJmg2xL3OUXwwgg532cDO57x/XyYqYF6780L05MxE
1napPL14RZsuccPJa3Dvkz2Blic5vB+3G3HZ9WUsAyUjwJCeRTAcZxGFMtnnCTSq
9YZ0Qpc6eqCpFsqY3QezNxfrIQvhiNxckRguaobWpKEkq+l9oBiWyPD2z30i7TNs
Retwf8+egE6S8yi3XOSv4OS8w0sl8fwUZCiY4CapYpxZfqChqNpWJwSjZq4c1XQG
c4muecxJhQmyoXRLaxN1HEM5AQx6PlB5BlZsJFMZe2aFEWnXf9TuGKewyCAXuflp
5oJCdgaN2iNa6jgDr28IloDwb5LmnlaVs7WKX0Wwn4P/h1bsovnx1Poz+3mC190X
XVv47wUVE8u5ao/aL9jaSdCjcTk+6KPTvteBdn37EfBFFmJw4FaI8EsEV9LaaAwT
eUppuOmQq59ncXHCQl9juJ9fTYUQNqU+HyFmPRifAsRIHLqPCrW7X2ZZwzt41jA3
ajrCgsm64EuR8/4h/HJQhhlMyV5YPOHihq+T8CdwuNkDzwKtyBDGmzVA5FadV8Ss
opH42HC0fOvy/ceNMBjc3fxTwUJl8SxqiBQ7Yj4G8q/oR6M+lFqpE2tsKZarLO5Z
40N/WIMnSWBo1L1AlZjenpfSDFTLhM1/pkZam+MrW+IgbjzY/IXDlM0M5LvBgtgI
EBrzk6ID5d4/uxM4eiic+79pDrXPqh5AEb1qrdgJzxIk0uT44e9d3wj7KWFRGn6M
SOM6fZX7wmbr7E2GGM5bebiP3pP28FcakqKfBsbgoghHNqtb6hyQduiXFOR+kDvt
lKqgo9KZtE05j3cyXOKmT0iJ8u9SDu3x04Ew34JvP5wOmTXfAytmBUKfY9JqsW7d
KAfR45HbLdIkOooD3Efw1D4rErW7bwRPYvCQqq10KBw/tbFFlZVc/ZqxsGtQL72v
2mffHf4jv94bEeA/amQ/ARoRzT0OPabQ2rw713WvAKJfJJneR7QMunl/g0lItBws
6pn9hL+Iaj1SsUDUtLXRogv/mGS+w8/WOqExGe45or2b0acOCHxDXcuKqtXkvls9
4GP7X+7aZOEl1beYvYS2hCdqiruHXqkM44YKJ00k9nbgk38xVp08NW7jHu5ONOPZ
Oep2zarUPIGSg/kIYNsbCR9suyt6Vr7LhnPy1E6NkNTZQaZ9x3oOLVO9IDBw7/tU
x7XyK/u1hIAg09v1osbLAG08GFXDMFNLBkUisPYEJ/ifWwR/byNXYcVMwMXGqM/z
uUKiHG4nUY2ZdPIN7KpPMMEmgRnK/TGsc+GhPUBoQDPKgnHhNQ+XiKe3jeHjyu0Z
W4x5F/AQxl/S92Rg28TXs+BWiRCPM3+WH2THNjdDeMEsYNogKKbmyi4ztjyU6jD5
GzswYTryVZfVCtw/QfgXd4I8vRq5RqG3yEKnU2uQ0HW9McDE9ZP8Vwgg8cA7tcQi
fGn9KAHFakhHU8HkBLz+d5G9SAmpcYByYMFOuFu9oOQGXl913E6DQUD/7r6ciJ73
O7xn0ERrV5ma+YybWniyhjOH0r7mu8H/DM9zFrGI2b6gRMMmhvB3aAWnbhPBMrEc
RGBcvT1vx/bn1sflosrKGssNzRT6tvTzrJXAAYlrFI+EYCOXSW1OnAAuW8pAdAzz
gHS2RymWHFuoMDdtRAdD9bMpRJCOy3ns5GJ8nJbjMQyOgaXjdnMVWjpYYXRcgP6+
yzwk6YReiDQm6nsK/4V6WyUYueMFZ1HlxcUhhkDV/kw5z15DgNeqH6/isFzzpmFa
ROCpv+rFNkbx4hdm57e1L3z9Dg7Mw8tr9bL5JdFcDFDgElNjiTrhYb3eTp6LgipC
fgBtkD99eJJrWWiROffxpbxzujHlkuMgHizDTZV1vZZRJZjhJ2aPClVvfYp4iXjE
2vXYyZQ/U02q79m9dVNIl6E7xtlcLHScgOZL4MuWwpM5VC9YnjsNNYKpGHpqUYex
A8Z/MnoFhgJmj6VNsGR75hiiqt69zqIZ4Z/kneJRgo8Cv3GV72pVktRyKjsx4B3C
859CIaELugVzDJvX+kfF8R9MW3giHccfPQCTKIjmjXjC1O1IHhN8yktrCflzm8Jx
gAFqqzTz1hbUO2ztCtPsgehi/Cdcrds8YCpZfpvMACARMpqq2QslcHwQUxepqYhg
EJF9Rjkd2y90NrXfOHVqNqaiy1rndzTw+zangNnXm20hPJ5f21VT+FPkc9TV52IX
gyeSKy3E7LJEHBAsa4jywZQ5d0nSqXceAWalViqteyRVbTT44Kpy2JOqy7kp3Ztf
vxevOK+DOu5cYFxcjD2JspBc/XtBPjPxqu5gAPowM0I5tipO0aj1w5btJXnw6r38
krNyov4zR6noYPBQaMOGAaHIOO7j7jAUGhwyNNF15YtHchoa73ZExEsaLtrpqNjZ
meRX2g6NXVUG8U4geEujEr695osqbXKRe9EZyyKdvg34FIFWE8ltbP+5cHLiyq1l
0uUpt/6v5ZHU/NaqKXqgSgYtrBZiA086xBf+h/qrXsJC7Um53E4D3F7ZvoYxnPTF
aK1qMLIVXu7t2C2lNgTNQzOt2hGeXpRbuwLVagTTJXoMn5sTtBG573v4f/TEuoPK
qOQ47O4wcu4E3eKNozEqAGM48MJOfazX2vcPFV0XisKIEZWr21EA2FfKf8pCIVEx
0WbmghiPjTR1ipcMwiT/5o4v4B57gpGD1v9sCEPSEqGUdc2em6b4GYhikzbcncX+
djIcfn2riw0ExMddBeCkOIREDHCkkr+rH1WhTbQQhIUFWi4D+HhcWNiQLS7RONeR
XzbCHNokKDrzAFCR+4kcyo62Yr3rHOd0lClIdZmm/ED+QCsnoEfhhXoZ4siJUbOw
S77+Hbic3TBf40en9gqJ+Q+uvhkUcM3d+rERvZPOV6RWvZ31vzZfbmVh/RqWKS5x
lwtfS0wSm8qnVB29eXelBKiSRYAi3vQsPGJZ1mw8rrWNgGUT1EYLqo7w1CUhvdrD
NzycGaTqFGAO/+SGAbYdzHK3arTCQIqVNacZwQIUbcfiA7CO/jAcTzr8lHS/pxV/
ACrAH3/+rLrEyKenOlvuI0gYtrZCgGrzouJLLtbWNtrxSaE9cUuPNgjwqIlqKu4W
OSUjRYRg2w97tSCObar+1FiO7wK8po+kq/HFzXWOrvO8DdjANeOPxgFB2JWqMC/f
E/ITrTKJAmWpQT9sfMT/wRdyXxHV1+NnFEXiT1100r3PAQ2Jr8zhZiOYmbKRlY7d
EC4ZXtF4FyamoylwMyor3z4LKKhABfOrNc90VEn3IxvDwpNERA1F3AmQJ51HIZYr
67fC+8cLToYQd/fdS3Os3+OQfbkzDl3yhRiDf1TaZCiViRsF4yaCejxnyBSuHoeT
Mbop5MMpeDR8pCgXTZ4gntU6qj7/gnMjObF5uUdF2KPYoOa1QGpdxBGxoc0J2+jv
F6LUqWvkOk7Km/+A4PyLhc2xJ73xg/pusuv/sqRw0kTiKEtkQdUSIhjhpuRzxGQs
5PBlhn/Z2Gac8Tvi40YFpbV/UTWJmgeeJRf9PkyEiE7wxSuVTLeOpd9vKUF3hb68
P2wpj9McxrT9wLvSG2h3dVk0SMhvhKbSJt2QVH1Y0Gx5fFxPkUS8fNQwh5ThpiiO
1YLWccu5w4pHztHB/AzdXwtte1NWGeWgSfVxVO36qc/qQXRX4lwLViAD83qn/0tP
dMOrTse67khCxgbBLro05wAvINsDXYMoctNrOvgNyyMVH0O5oPWTVXj5aU6pom10
XfnfOacVE/ftWWdJRaQugaF5Zj+SvnZF+xoG5P8akiBg+ewNvBWE1ch8aytPU3Id
e6KvzKmJDX5sU+YoUzr0PQE7KDw9PFQKsz7AWPrsjDmMBxzT1vpy+f5pmenCEocm
69U0BkneIJnw5VD6b7FSGL4x4fb1B3dAZf9sjKFKQytUN96guWobAa86Ub45M1we
2L+DoE3O2GQmyRNvd9Xwn2Fz8Qb9Au9BF7ee17q/SBt/5iZq58EmrMTkFrs7a43g
bXJ4+dLOwcULJ1I/osMyklppM63XVT5SWGgACf/6kfJSNmF4UmE5ra67gRk4onUO
QvDpK40fUANxkvhnq3/4oa0vCNg60sWg6efkgkpVRV/hoWzdmuKZCfQQlEQeGp7/
OtPjSPyyL728FSbQUUKjXzwHzjGvDCpV7EAj8qLMyfDYZryUWCX+/rX8EaV+1oaX
sebrw2azWvj7k2AgBBKun/U71huSTjETOvVXEriWkOf7gX+CqHwE7WWt9VrcXFIs
Ip+kvEINZw+LPlaaHFPcVm9AYGVRjrjMyEM8GOTad0tM+AuqqH0O5/2/uiTAA9ac
LWjEkrBI3KpE8ngTjxaRKrY1WL6CtCyhNGg73CgMJjxOuzQC8ynUuO80XOoeUeSD
xjLYSVEugtkxrOgYZPN+RUoQNnQN8Fl5pf6Gu2mpklSFzAyfG20f6rFdfDsERg0v
74nFommbhVB5faVjKtnCLJOvKF5ZsmcW1nR+nHK07t0hpxjOhd9g+T9ZRS/Yw2Sg
vq/vMK0W6ALzdOlksMs3awPbvCqkjdSkWmXs36HXFWpLWAiaklIz926hDBPjfdGc
UzikzubWjN0/MjKLTG7pNq19dcz9B2zvxNLST2P0IWGzUAcJxj1WXrDSiqlxZpHu
WC2IZzVGO62ap+mahfEf+BCUhxzCLWksf0WCPTjTps4oyyZNaOrqr4ISHAdVPpNY
t5pKoDBsZHXJOosb8vkJU+Qiop7pH/tzP/2RSxNKv1w86cQkOGbH7rr509bSnzaF
TZmA7bcY7JW+7Puyu1GMBgfWDC/1E7y/FRBFRWhp0OQCsmsPhWlna0vVJEKHXLK7
AxyFkR1dXz/+7HRCSA28vAMRH8k6DGISc+BtMWkCWPrfLwTIAipzjKGUzaEVT4zZ
xpobahURFW8bv4ipBcXGEf34Xti9shO7zzgmdfknproMwv3zfzzzc1GRZPdjtTbV
LzaV7EoGKFNsHUBHl4bhOoCK1vS/rnT6YmpJznZrwnQWP04RK2f292oBf6q/vEFL
bNH9KLlq0gZ8blxO+O2cElPNStVdbvU0nSLPdk5T2YmkxRBZDUOvJ/GAt+NahKdU
8ELg2cX7gZDopgPH1Ks/h1g+OSSeQheQWxUezyyckPvaqC+nXdc65E90H5Uo/gK4
1ug49/NOx4VZ2lVrsBdlqMr7C9CTiHmchVVSTrAuZBK1CBVqB+BuObNWjOAm41hM
tTbnklMCeLTfkkr6HVxYAFFJgMR1wQoBqx/OpSE+G+sVvhcXcIS6Rv7qLg2gY33F
tOFGZIMrFGNYe6pWLCaoHtjhB61GBsy5mfx5hB4B9NvFIEdD/VF1zEzux7YzJ5M6
Gy+qyCqjnyOlsRpocptCTVCsDzm3/h//RsgpQlDG4QJU1CH+tB6vAynksBGylfye
l3UukA8SWU1dKVNpQl8IUHI51lC20HHwGy+cJzyrKpyAaIkx7MAv037PLdVsCqtG
60L1n5fHtcm42qOvQraLkZz5BJra3tNPn7YXq/xVNabvC3R06lAAYFxh8PkL/iq6
gRDRSbU8qHppQl/u2TJo50MHPknsNONqo1INnLbN96mxPsoWMEv/KyYI3q7pc82P
d7fumJ1FCVoEBB4/OBdqyJA0fUwvNLwcbhRQxOEZHfG4v6l2V8rnaSQyfm1ZWqJj
BN+x/LVG5qwDQDC6yIZQ1IkWFEGCdMFCsF25kCHNb5K1NqfIkEdFpzVqSferR5UT
9fzIJ0M4PqdAn46xE7gdJLCPxBtkhpBHWG/zZsuaYVs0WNed1eC4zELjcJHoQYcv
xFaBd5hHVS6AE4UoBaZxCvhLAK2Gx8WLGKoUjsFNB623KfQ1RZy/knkV70K+Hbs4
VN+1Klpe1Tx6HFhb2m53g+qeTdBLaEdh/i6SJ6CKld5Tt5yVWB4kFskGekTDEMoh
QLVnbxYrhMyY2Zm0fqIJdpbKgWIT6wnCpP4JX3A9K5czuY4+DMC3bW+vhIlVYfp4
mBVtP1C4wxWsM7iGiDcrRedU8AseVm2ZAOm+Mgo/xlWR4/2i+UNagp2juQ+k5Wv+
z2Bl/7w6+P5ijdonZ1hDXpSIZrXfX/dV19zEy8sr2rQDr8Xo+tR6VsNfEq0lRS6z
WLRdf3HZ++eF/Yvq01bhKJg5ULJMJbUdPul591cHMrri+LYv7vtMacKPE6avr6PR
JV3XbRvUOoNxOCsP78sXE6enIKLIsjWKpCkj7+TxGWd7d1mOT39jQAqiTNIAXBKp
oFUFhjIMm16iNyAL4+x+sbNrGY1RVpqEadaAiNF0MA3ZicDkggzo6XvklqgOt0Zj
XckvEsLGZsLp21yqFZCfId4w9ggLQqBlpTcG/qZVB3f7Fx2orM5C7Fcm57mFiZpF
3DiDmVq1o1wbIzr89S2PM+HY1+rZ2FrvbR0YTc9xqLm1go20b06KKxLkDa2oC9fu
l+JTB//ur6iw6O74131Z1tprrvTKOR/96Ez/xSjhCZOUd6VDSDmm6Sh/ugJNF+Sf
UOYX75siv7yt8FVWZwQwQ+w817KTmjxt8Pcdc3o6zcYq9IjXcb/xv0IRowFuEu2Q
ek3rivgj/qp53AUojfOLloXIaBvASKWiHY2lZfRStt2LGTO6PaPlDVVgGLlNjs3Z
2m0RbF4EoPv6PT1uTj8kPYKey+QOnAS+A4NOyxxKPvY7/d4it8mDFSZ6OySveVyx
O8PuKFOSIdq+0tLVZXoo5SxmmbWvyprQ6yuWTxX27sj55tUrZ951uLeqlGRIZ2uC
wxJ02BkFV5AbXWspPm6JMsDOAd39FSMYZYVl1Ud2BR9Fa5RHACFi1I7PGgyy41B8
M2GgHQCWSvvm2RDQ+TMr4/g25lbgjS/7IL3ObXmNbaW2TRaPV9aa4XUXj7eQHjdq
NS1HM8ruvOcO9B1qNVFwwM5k7N8Xt3zcg5uCLtHAohSIndgCVqXIZh+Batl2apYS
Hh8uvxFfe57PJ7utfzHY9lRrf1x5Vn9JiK5zjo02NTPwjfRcTtZjtaipand3q2BO
En7lrH3mEiBjgAbW4nX3P5CR6h4piyJ/F95wercTdehdj5BIWroJvsWeDWMbnIle
SOjVHy4+/q8ZrvXeS72/p+biw+MPErln4INyiryi1l62r5IAs1FbyHy8KLrpL46X
RyRKoQvU1fzqNqdl5RTL5+WPeUPUDcJBt7sbgjh+toYtMWujtyGsQhBWh6v7YJEH
0v8LW/99FLIXk8UyT4HnAFxiK5o7DTvN5pWXPWgb5YxT5ZlxiFylzwz1YuewfdOn
zVjPRKQ14TWLpDBaZii1HokDcfrwCspbbduYJldAh5AMW0Q4jV9AOJ0278fbbYUd
GQnaWAj2dlUZtE1BgsOrBhi78yRAhESJ+gsMKv9otULfUIa1vsG95kdZz8TJAFRD
47r11BfmKvBWssGoQVBGmTxKCS+J2a3gJWXLf+tlIBOHCEd9ApwycDL2tXUqTsnB
SVSWr+E1sbfQnvuQ2pe+LQXvj53G5Yqtgo9Ju+p5oyKkcE3NOmbQjBAkdUKJ6Acf
khKoD6ipO7/QNP3rpmeqyFX60fL4hqtYlJoC/UFcfrQYHyjc34IKG9Fcqd6FN9QZ
XoNK6KH2Pi9YFWvItgOZCoqFVm6fQKEsL2pw0/Btqcs1O6troVUdLZoiSDeBajPc
NK1mdKJW3bB/jMqHFBA+tzrYFAknE0VvDdW5/x4f1ltUm+8XnejTthBk+Ev3jM25
VVwiJD7M4mpEkOrKVxKXRPb/uRCG5up39YRx07Mqnx/wLqRWyqjBq8w5E3uUhz0s
EM3/7Ehlw+APpoE+qWling2RUqIpJj4g691kDEMdzwHFAScjSxRfGoeKSMmEexA/
0IQyi11Cz/EWYjqOMzM//CCyIVQo4hHnpbclpjBNMO6kBCnZQ65NjhVsEHZjyXD9
lGfV9fCZaRpiAxB98wWP3wR69GiqRD3RS8hO0UQp+d6uOfZy3yfbKGaR56xUjM7o
8dhMJ3pppADB57iFYXUghgDE5x5zH2CZccjwj/gCsnSXRC1YCHRPaaq7MTYXiIJj
3P9JR9G2/QYraRy1aBsOnVj88wig+G+/Gn+R+hTTxm3cqvockOniTFduV/dXahIV
9TN1v0DDWKpyf4gqd0LVoVnTAdtVZ5r44mFvRyVmhQpOMtuxuohdnPLinb8tQ4ah
XqqDSgBv3QygcRYlAvAKh3a2/7dNz1LYSJlaQ9G7AzB8Re5x3BBf/0SC0cTa8F4K
0UzK878osJiHYzZO/0OgPbBfwhf2qwXZ3SjxPRxptb1EeD+MiRNeuQUEFtMkxOvm
N8SBUi7/8gu2jJpZCxrIp9EGYx6bwHwfnf2aGWNhIvwZZlqQG8WU+NuXbgyx3bv1
UCTTl+5RdrAN/5crqTw5uWEhgqRXFcub/Mnn/vgCWRUry1mBiM34ebwP6aO+6Pht
JkgoegygQn5qYod1AdUOQB3opzmL5yO+h+YschJfdfH9jso9GE1KloJVJe7yQcpE
em/APRachxxETm3IgAwtCsHPj/uv0MBerYRuSGR23G8WQWTYsIiH1umjThdRef+S
muVxaTQhQ2kTvmJBUH9+1KKoz2Hsi1bE/+66wajYoGokZzIvmTQclsJZHAF7flve
BnqoAVkxwWUpxWCy0sNlFsgRglbG0JA+UW+tdPbnr0iDZ9MbqSIA3r8FHxBFgeON
slWhczDkp291hoVqEC9i2khZaYY82LVnbDruX04XEC5+Swj7pZ+4acskKJMpSeka
hpa9CbbRF0UipD/S8KiBPCtwIJB7euWvGsKeG1eBS0VkDVCzZmXpOtf2bea6m2FE
TMVhcyaD8a2Thbr9B6zKz8O0QxjozpqrMXbN3F1eLIu05NonFIFbQwywr+Nc+H/j
OEBnyOzxkj3YXfc+e1vaQGsG+4tW72/i12Z5eHahU6bY4Cbc24tUHLbb7RBpsEs8
NqlA+8H9rgOmY8hi2j3+coV+nvVxnCQUyz68hr/BXwA0ddCn/0XZVa+Csa15dthV
+/p/eDQ6cnsM0QqCUSKUrPpltza29KxXIpe4hpOFBDcaN7vzhvy7qPVLTYCcWLlA
rUQd99RVaVvicKBFpPpO9N5dnhJ5CDzYLOnPg+7CGUg9PEDvwVBFI/LSEyPjKgrV
LQMzBk21S4TvXkNrJk5jk+8ZBjt60t50gIihepXqjHzAlP4COlXoHH6Z7n1UsbAW
2yHIl4BcuIorGtc9hFD9UCmbnXkCPssWAKI+KEhPzsFHmHZw1ihezlTy4XkNNPm9
Dl6cD0TTIjUixO4M3yguyVkE6csVQAc6EmFncK5tUJ60AGGQUgCq1A7SuAWpOME0
KYbu/10IQqxwVIOQQm1rN9BlfGQ1EomxcLwxiiRsCoufHvucuhvQOT13sG3BOLfO
Qj9DWDLGDs2FAQlPvTjxjq3lT8M4c+8lvGjs5G3BAmkaPQdpkKpiGv6C7IzQkULz
4ttxVBBjMJCWrXJa+lZgat6+gh7g9jyyLNjKkxvQ34M37UGfgLM4npf17Xm3ZYrk
8EXXw76F/+KShC3WzpEVFATK+kl7rhPTl8cvQnZy58RI8NPDEwfm64HKr+M8H2EA
BejgICxc7bIvnK2zltoDboSWCnXmpdTsgyPbQ4dgYMpHYnLVSmAOAFgmrJiSWTCs
tiW3S0zBqhPBmO3Tamt975epm+NeQn5t5rcBcusg3OEicDINATGJa2fyprqtcAHy
OIMI3TUjG7MB6cjEegGI1AGnqJZShP+BaLbSZH23P62jWKsjVJFdR+6pLLAoGhSV
iWEoAYUedg1JIBfsZdB2TyFaWeMPdPCyeLhlIdEyvvaFLilj4RbXM9z0RxJgE4T8
cKuwlaxAPva5FXJANEHN7Xskwep+nWYpVBloZG/vVZcTo1q5yuNiAsnifdpb35kz
JgftgRCwEXnbOvw4J3CdqINq9nvibXsN75OxIkYBKjkkQj6Y645PAWJAL3U88TAL
KngVnT71/YgQ+HtSEh7NcfFTYEz3IB5NqfSvy5dedvaPaHZQoPiZueMfWJ+PyaiW
7THs03Ig6rVqb3Txi2Jq2UOU0j7c+rQSVtZeOjlZiE3bbtNyc4WNLGBKsLxPBV+6
IGnvFnwll2rT4zj67N4pnzbTGTd23PC4rqi7iSk04lyoDAtj5RiEMOP/fQ9iQEAO
e84hBX4tIJvyXWiI8CtmidnkTAKqkcoZ2ooXDBDmHD3DGh9R6+DPluQH3adla3Fd
h59VCm1Y/TFgmuQ1xTdqKXNXnw99T4HwsKLy79JNZpBEk+jAzjA1AOzswzNVCfkx
VKORbFORe4iY8ZaKCSFlWZX8621IkAgo9JosRAarx/mDyHMWeOJOiygJyciqlZ2Z
qoj1ArvGPAg6D+t6yZ2j2NmEujO6fUGC5moECwaqNryMypv9HV5bDF4HgyYDBiCc
BMKG7iRHpQrCO0iALGTDTx7jVXuTXnyx6Sd1e+FUzDbXfrqGU9Mjyvvqpgh3zJRy
1GiO3JDU8Y+0ledZW2ozLWyLNx6RtWbHVWWBpaGwm4uLIopZd3YdVxwqGdyZodxc
jKCKbJHJFcuvzup9CoOyhjxWe2x6PKe+7gs2XHIcR+c4xA7/cdE7KR4g9PYIertr
MJUs5soW8NeaQ8/9MLaawjqRZR32z1fqrfLurS4PCAVQplrSgmRXxNgzgrbHrgCj
0vla80FMPCNNALTS17GSirXMq5d5lgce33bJwsUjQu97JYtrq9yT88OuKLqW3b/2
K41DwM5Ew2j79/lb3Vv1vHjEt1McFFju6FdB/rBIDHRjstXT2Pn5Bx7CYibBJjT6
VgkYZhPukH++RgRRtAmym03pxg9I962Mb/6Pb4ffTNGugk+C8pG6v+Rp12Eag2H4
BBsJ4nt8MJJWHaBO0a9aU2nt7CtT5mPFWb/npx0HVEB3D1HTx2tB/q9pPtHFEx3v
ivDDBiuDJmZx1SbmoB7L3kOwGSuTFcHUwW4g41A1yf1mt7JObu4Y/vxOCtqulGGc
WXrySOwvwE06VZlsxo93NsYnDPUdyii9UjXOEPPXg6NYE+dBg2kZqWvgyammSIEG
5q0WEcrQV66tX0L48shU3leC0LkjnpGWCsWBvYGy5hxAo9hv1OkRHWicmwYvelDr
fDZA6tnXPi6fQUWCnegrb2TQhVnkflAb2DBbhIXilbQtJYe8UjEDYjbymfB24HN2
S1zZtd/ON3vQNpqorGsFeJVeXNbaofRN+7KjP2ryEBEQ71WVzrLakMJRCYuoDt4e
u1gjJwgglC9waQJIslakX2J15zkQIep3txsRudWYuWzA0i0/dLjIJjuRNfiB/a4z
dDMIJ23OZmylgtMxzt7bjKDph4Q9y3BsdUc3NSb4j/cmNSm781L/9o0dUrKL6Ck+
QfCR9FrHkJUEejRYWEF62Ca0gqcV0gPQFKiBM/AYR74EOod7J61/0ngQB6W4KJ+x
FLfLbHjyvuB7bKWyiUz+/cbBVfanCqT47bZKenZ5SfHzct3Ru298bskAOKgVpF4Y
SoJk/2oShfUxmUGFDmpe16NwvxXx7TdLf1IlciN0QGRYtr0C2ZdWkGCmeYyk7kLE
v35JJiC9JJyzWtLjQicEZop6Mhqp98/mkApRuQ9aZvKj8/ScEj8Arb/Xk8fnqb8L
Fmwa72ig39EoHhOviAk4epiCUWBRUx1tqMY57XdK1qCBcxBYtuXZCsLYR1fF8PU6
67BpSQYpc7VDpvDMZZ1wZD3C3v6X1of6a51/T+2qrvInUWgzqSH/z+Cp5iZ/v2IM
WWuaLPnrhVorMYAwd8/UYYr5vP1zpArv/oalzCO2eJtuGwcxGxhZ4pP9PQwmJqln
DMP2KxiSaINF7yt/Z6N5pxYmVWssaa2BwIGSk7VuUpLBiKa1CS3Bn/XCfhwzgRfC
RXGY5kYRiOmh+f9/qLTzBLAvbuMDbsQ3D1b9ESHXdeo6GNk3G8i5TgZgl0wiRNYV
+UYkIM2/4boZ7PQIQ9aSQcywnxQowGSyKCIPQ8wySf/g44zLrpesWXsYALkjXiEz
YwLPtxnwPjhFu+qoWfZ/37Oe2917XuCrz6va6MoFoUzcA+MWcEILLBNWOeB74VFh
pX39C23bhhJODnzmTR+6Zw6WTq/Q9BFLRhf1ubHo93Kpse7v2zBaVGY+BaTa1Ssy
cxlzPviJ680waWu14EcBZOft4rZf3O49EV1gPosf2yKDBQRSO4gfBXN3de9S70RD
TmIUzA2r6lYiWs7CrwU1Otb411390EZF8R8GQC4Q5DzsbudSLcgosWkC6OJzC3T5
h7CElRbN1YtqGakecZndjY6U+0LpDdlIGOdFXjRjeVeg1xPpHcuewNAcOFoh78qG
pmqpIPYcbYQmrrIjSYHSu5jaG1qfW8hfgQcLqKkMmRUGuc1em0HRu2Iv4lPkmpHr
wjkErsqckv4+ZqAHYxqqyo/O7FfK5pPf95jP2FTieekM6iGtJ6jKfrcTyAcEMMLp
pCPbUnOK640bUTIU0HfORrgMMJQIr2nj6OjjhdWWi+mleZ3i4NLHJz9hPyWr/yfA
K+GIhKUSU03hWJo38tOm3vQKRayIeXNwNkmxxu+iEkrzHMI4EAxp21X0egmEsfTm
ymSoc8y4mImbVxg/0XlWPxnE/Ags/w3hJgtyut7y5hqUR8E6nvxLpMLoy0C78ElW
vKhB7tBzGuOuXHmWsetLG/Z36xuwoFGWsHMD1cb53ZqkMA/RA+rGhcjcxiCV6SR1
2at4xktKBYHrQ14DiMEy7mK5QnSFez5zNdbi2tZ7U840Xuwjr1K8Bw+1uZ/4sIvW
lRhmiH+c7574IrcyPQcuoHz7P4L+8Ir5rA9Boc95QfBT30JERCn5WSb4jYRtPoA8
bLqhSYreGWsaxzzE8Wl/g9jDPFnBgv/77Q206SqTabN8mIUWEmU1pT9pU0rM+I4S
+1jUgXVrGgq1NnciBvdn/yM1WK5QEtGxKXpM6QLf0WqW01zgnib4ZRfzvjV9Q8Pa
CpWgtk8tsB5C3z8gh64HlPgEWpHoYwAg9Ix5ohGpmZ/Vw92+U33uoFBzTKmkdixy
Sp9dnYIz+Q8sv+SsMIfI3W8YrPRRjfDsBzu6+KIFvFEsNoHqtQd0vX1ztrIj9j8y
4HoEFkaKnYJ/Myp2+TSiPutptd5a7BpFJhMaTAS7QFiJcmIzFfqTJv/2XBzAGUiI
Q+EzkNAK3O53H/mE4aVeIlR+w9u90yl5MdAg3eUt7xfNSTirDi6tq94pgh3+JDYf
9lHzf+3NqsVLavdyKzMFgVmfCDlpZZSoKSpKoP0DxIy+9TzwH5PWi68kLHuhb8j0
MXI4ZAxl+jbAV64s75CZBWWCcwCyJHROxhKxEsSxipJstV+wpmVuSmFiKzlu6JJZ
tKXtX3RuqTjAz8uZVc4y+bsWQ31T4dVvco+YWQutSByYfVsCqs7b1U1mFHTyDgGb
ye8ep7fvRNc443GlAwDKeOPm5q5KPcf8l+mFS9wPZ06DJE7k3GY6zXS1l0RSTnH1
nhUfvqqyhbUa5z+XrOzUl9h06N53TqglLprsSTjn8diCRDdtUGNNQfib7iQK743s
URoz3RKglIbIxTdGZWYBtmz4bW16YekcQvwigq53G4wIaWhmspNbYXEfzs2oLaNp
Jqu3M+U4FA1kIP/mGnK6aua3Fsv3m4vqXKv6xVVNvL0fy7fg8so4quedn4r0gSWp
o3B9540Zsx9ebaq+3MJlaQCgWcTfV7DrRa7YJfd/WXqxQqKeQtNrOD6T8/SNzbTC
Lctpw97dP+D6SuhdZfOKFEOy9cKQ9rfC4oNZKbMLRMNc1n7b/piiB6ZdOhlGgzou
WVhlfq+0DWAyxaipLOv8NpAhiAVxWzy1y0w/Tbr9pdpmxkf45hAT4tlWS5qKRqDp
T0GbfENd5F6yFJ6O+dvk3aDovYKtNcI58LMX4zYKiPDPuEBs1SpRXCIp17eaSOFB
1otAN4IHvmAz1IFDwbNyLhhsA/lgL+1K8o4BJ0dPiIIPbolKVp4FH5Gujdsk3l4Z
MJUrXNGhDGce+lmx/hLwlvHoKadwLTYDuy2jY7JbSKm+Rx7FJPYxsdO+qgIQOfAb
gsOYCe+sHS+FyV5vuPl2FIJGZb72QSQuE1dwsSn/VfSJSFYlfkKTfXmdjhJE/bhb
PawMnMA57EjG3CUtrcaYmqk5GylxYQERDko/8WpL4Plijj4KXoHn6W1+L6z+5guZ
UONv8GoOS0WDBMAE2e+4/gd+JL9SfnKXrMB6cSSHUMVR21rU9PPkGHlgSeosaB4g
ivy9phpjl7h8WH2qjR9mDUzZHBXsV/9OabkfclJSgHvSmZQFsQj8TtsE/WvmxF0n
dpsdCktjVd7wb2qRJa6E6mcb+sNmVkUn9+HgLyMUg+eH7IaXcSyJfZA3LUSUt5Hb
pdClT0fR6Yelz4kFz1xKKftlB80H0M0+VEC8npIMqt08SCYbZm4CuNJA2tEeqmBu
5y5mL4f+bnL65VGDlSaG5jPJwvAPFbuv+YMLQwpthKajfEKoTtSOSuqf+n5iO2q+
ksV56QNJc3/Bc0gmoidfwXkRaIOESJMsWGsAjKGckanZRTz/G5mV6onqXygymBYL
3wzUqlnoqqdJXj3V+C0+Va+E8TzpxT+AaQoHGq1TDeaGHm9Ac3hhT+a6MHDISXy3
87U/a/dEbrCR9a99+4uZVKQ6LYCpO464DEZ6NogVBa+0JGAiMMjABu7GaEa9XbHI
AmXs5Hc+hnTVN5Br9qExUDLIWFxHT1iafGjZo46G73FwuAhhThaPAPEc/ANpSdDD
N8BVbIZYQKvIoJF8D1ohbdpxilCdmxzpzSQPtx77i5baegsB9Iz0NRMt0uoZlsWN
2lDV3ZgCjqkERndJx32PUv9gSbb6fk+mgMyn0XVeKHmqEDBEXl26qBr0zn4dlV1e
nlE7DzeExT59NKBZbMmVW94mLiXdr8FeavH9byVFiBxDY7l1kkaVrIVY42yY3EL6
lnKi/hmHJCUxr6Iod2mHTzfs1EoQ4vsTtVHjuESPsX5kpQD5ylvakruY8ZkKmt1g
BMh1CXiuE3r0090P43yNWovdb7w4jiANwsYQDrNzgIZfarPYb09M3kW7Pe6Exd0L
RBnUfSJ+yOvozctxS7jNFyy/fWZNpozbs4qcsSNo+eoBt5i9s5KAWoFOk0Fj63yO
OhdErsFez6jlUyjIIDfwX452LUk5T0GtkFHLGn4qRcqHac8CdQfhVg3jG3yErGrc
2j5Tsm9gAxHsDMvD637D7ZKggmJhEJfVzEd/oicqFdTfmoGYhdTqCmdhggOXbLz+
QLebnrFEYUHKpczkZ6KU9vRFVOx42EG7+YM/fRsQntPFMO7KNNUtALKsddVaZqdS
P5R700cuQuOGIYRg+j62hgyi1cqZvqAmScv/adfu7OnjvjLYT9P/TUTwwjdjhbm0
m85Ef1relhZ6IR5ECJTWV1pJu2IOcUbndesrQSNAzOqbUTGFJdFhL7pxk7fyuHDy
4SP2LqB7BRH3QRURWu47tleTtSyxO4Q/H8hGhFKZOCFazWGcm2RkBRJj11xDd4YP
LPeuMntSlZhmMplSacwzEb1EmcLnVDi1+tN7UwwGyCxOSIgWkViKi/WLrRBNQUJ5
Se77KYoKnDe7htFNtUyWB93r+yLF3KhUATa9LDJ1nF7/pH9oe+9JZKNZ80PqbHQq
BVMKv/VwSCaOJhYmSPItj+2dDTlhs8mCYq3M3l8O+EPPjv5nzKnn4/6jGlER3OMV
MYjnzCCczKJk9oqS3X1T3++F43XTKjxx6Z5CkWPegy3HQQc3kQ0JUQM/PfPDxDzO
ST1ihBT0RCyKwcF+JFOYym9ugFfdUngkdUVC39AOdSFthxMH2yoVPSJ6coSzTuTb
OaRUaZo2YEBcuJP4YKvgPI5r02bxjH3lZqJEIEBqNnpffCFZcceell4LTvZP1iWP
DOS1H81cE+5dx8R1ALhuHUQ7C5Lw7Fv4U3F9meeFLkVc6NUd04dqSgv0f0cVxeHd
5T3xEczEYQDeGFZBVaAhdStrGdE2FtpAqOmnxwNVZUuOCHCZVtzrA/jukc+AOH3+
yp66DQf+xZvrosTaApwgJ97VQWljychsRS7M1IJjZhJm8uZFrt7/evKBBsF3YAQy
wi+2cBbCugz55OntseL0FFyBvUIzN37caBpi0Mm0qG/6lKNBNwbBFvVuybJLVQVC
YdllDibKKYWmaZOrO8WgpF7Wttx7EDNUYb8BRsgl1pVS+bvvZp1lVOrE/gzv5cGI
aDX5hmcl6F38W8E658bO7GjXjpwrkpJvTd/BgwYII402UMzf1OdLaHWuqP3HNAkQ
BXOVcjDVUiTu+Fh6z7h4ogC+eXnuA52Hj/JKzzJJBT6UP81yZ2mo3/KArsT1g0T5
xjui+JaBMKw6aP6Ter8Ju8oN7JeRbHSeLerSiC8L/GAX7iXQ1EnTj3aFmUZfk19K
jWjQfw94Wr6wZtWMzHp+9XuHKAchs6W+oAgV67fdDNNhr7oDH1SEKax6lhN5cwao
/aWrqvKXXXFsIIIlJTKnvp90nXMtIVvIZKPDsovLSyifXQdmfgOfJzgPagpD6ov/
sQwgozGSEEkuDIMBBsC80DNcN3HXx3cyuyPCVNUOijeCGKEI/pAOX+MdmvUybmyD
vUX45MMCglh7KypO9ZCVjknWkXCzJd+Nq0iCMeXXRYnNY6Cr4tC1bzMNG5RDSmLt
W3qTbPwbAsyqOduPnUdZEnWF5dCvQEOoeqZ9ZAPLXD1Gap8K8+H37YDpPUbp25td
GGxJesmul4yGeMvrwy3jA2LqITAQWyeiOLhuXYe3qasA57+t/ZmWLlhji1NCPOzq
cMJbg2ldA9j1KP8t8UCv/IGa0eGIkHt5JMHkKKWHuDgZ48fBsEclzcrTmBUbzn+2
Wd6I5L1VbOjvPCV+wUqWgB5gQ3cY4utStq2sRmUJoMwAuRGR8KA3TaLx4z8LHBxT
qZMw+gk60uY/pXyCFX7YiBJCZymuLBoLBlWGVaIQyu3OvCbeNYIjawpOZ8ifJC0s
iWTk5P/5rEB7eFbc0X4EKyFeC6/OQwcx+PZ1neGJF7kycdl2v0owLQAKxLIP1n7n
R2So/stfmUvArnZC/ggrjKJq0m8pT+raRGd4RFmmqFmkJK3Ab6yJoM4Iz4HEqU+K
TR8Aqtp2GL0W99fofN3CoGCZHBQTkfWpkc01wG0e91FvDXF4lSlQ1gvT3H6jbvhX
N7lkWn6z5b6laWocTcXogzi/nzikwVKp2XwLvZ1uQQnzLMGZC5hhCtP6Jr2GIYg5
DSOPvcxWCzP19ZAZdWT/1092WWFmmew+nKt1wILLfJ99+zm8raH7RM01nBRkVFSr
2Rl6ZKZqpQIQ2z0WGngDDTIJ/THn5ngK1RZEPj+6QSeSQhZuoJSxvdG4xgJsEHbx
gSTjbpqswUMIczSoMHEYKkmr9IczGknNN5jvpfm7wWseXIyTkARBVFuv77BniVJJ
ey7iSBv33vfoKbE+ZoIi0PQxttQ2NEfJgARfC+GERpktyrpyT2vOA2N2sewi1Wz5
QA1AS5uofU3wtlaE5Ei0ZGiapgaSCZ6hJDpblJSHrfTDhbpatKBG+KmlR0YxobQU
WLSQdFSIw6cqWHGXl5pKcnC1BBZDfj324aTP4ed/Gpqth/Z5LFBotnc/pfu7xE9M
0yKacSG44lNlOiNVJlqaA2odnIFBzWdBITcZ3Suybk0rB40cxIcbfJJf4H+R6HT4
XuQ8Z/7FYxODSqWS2GpK8CY16jSTd/pNF4SlmQWlDGG6kNh/qAyzVDRmCptDKrNW
GfnD5b0L5phooenkp1XhIyU9H/cxYDLBeOdD47guXBteYw3CneHD8OdLpZDjy7zb
tiQwAasposAQDI7G02VX+A62KYMa/veIvOV2wCRUPETCIXudklac+Wn94509tvwK
kloQOzIxHDU60D6fq5tZA/SIQ0jycoNiGkoDCzMQ6Pmr8JjUqU6vyaJ7PLhR8Mn7
oSgGpPNCjU0+L3xGUoGr/0XLWpSlZslM6sVt0qHJmu604S9o57XVh/tideEsj/nJ
kXzGZQrtzZ0zYfugk/4WZRtAI8UUdsFzTXPX6oI0DluD4O58fSo2B4/lhmk3NqrM
kgjuU5LLWLtoQZaYUI2CfdDat48RLye9bsQLxC/IPz0vUeKdchInpIKzODMFrz+L
hIgtmcZ8VNtpqGH94CCjb8wZGtEELyRr7sJtSKcmDA0d8nRJSidF+7Hml2RjRp2x
SNcYnP7deFNa2rIt1SZEuBmLvAmCAHtUCU7kKecVIB6umKiXB8Qz9WodBh1vHw74
6c028N37+yLSnHHK09d6U9RSalcxicP9lLHNBEPXgBu9iqJ0hYyLPRmctTjrrfrp
DpD2qb6XAjHUX1OgEzYE5dv7ooyPvYDxzylZ5e+kkhwcm/xbn16NZN8rGBp+Jngi
PfzoGeMdtGZ3ZdnCZjHxFatQbJmcef3ficGtsGrfP069eiTok55KXk9meV0Kuke7
C6gHILnpCvxktaA8PCntcOiqlzG/nyJDzvaupQEDsMdZgJhSfoPT10hBdVyehzTK
G3+j0bzOsDey/JyWycQuwgvC77KXpyb/IusWS1l06LALeOv+MuP7rTUX/Ua+n8Ga
UZIwouOItqgJaxr8AIKAJUmmhLDyGa+yQdvPtuTpf6ENNtCsgua3/KX9v3oY6xTZ
fbIX/WOe0CfrPLgNHtvvL+cWHTpnjdcjCuipfM3DUqdTxxZMMvg1Mq1zoWIHxOiU
dAlqd1/YN9Kj9BN9qwDwogEvTNwnCQR1UcTv9cvoxpB7E/aehHtWeTSxcty+zVdA
LBYobnIwxIk6o6FpIyCUiy6nN0F9kEO/V6Hz2hQ+5OEEODC+2GqhB1KIiBaAZnfF
pVVE+dcp95acK5TG95t62+ZicZ2QunLBmSf/TQAexZN0iFQJwNIy3t05WzUUQK/M
KImFnin8ghpr402YxMAQkbPbAV/Oc8mRY4BBHAJXDfJaQmsj/++cSjtKOCMLelTI
XRw2dzzlj/agIJi+17guNwA5NTIpO8zy+GHdjHfJMrTD2Te4F7Ik7qcXlo3ri/yx
/qb7UcNoravjtfkjgsH+3LdvwDYoybUMf0ItR7COdgMuYBOXj0l4+1RcfVc6GemQ
8LNas8/mtyz6Hgc3pSJOJggHXgxI5huvb0dbNUeFymS08pGm5rkZLhB4pNb/IzyQ
0qRRTw/Y6bEH63R7TvCUtfxpXM/mWvw63YIkQk6pO0e8HK/mROq/VRr0tWSDMzjx
ykfuFOmZICqe+Ht2IMtc03wzDNLrcLZgldogV0sE/e6p9ysbPEB7bY4wIAtbITmG
No2zKS0E7BX12nlUTtUOB3x05qxircfZNoCtLt4N+/TxL/ZnEwOgZtgDSPm6W2cb
a8A+Aq40QCh+/JHJcf2q97KU3I09oOrDq8tQFUidLfx72J+hY+Ij18n1R/0iagwq
B22UmM2VWoWJkl1sWtZAHBHEA2BG1iLEswR9/xrMpjCbucLlH7sKo4eSOvjtSV/e
Cz+y0nIZI5doDk9QIfD/IZbiKzk7az0230ixLTLGAUTOThqs47YX8nB+Snp2kBL+
9QLNl+hi+E0l0hqjjeyK9NMGm1FuYKLKrLX/WEDghLEYlp6djV9jHOlGtgNP8lJG
FMb826a0ZE6cVQ4QKg+zKORuja1bHmZXgCoZUvBr1KCnTLBbQYBCcC9U2ZYfbEMy
WvQF5OG0A2jYG+w5f+B0279MbCpX16aAscFFbiitEg240BGuir7A4XHyOYh/5C/q
Jxq98CWY9DaAYHDZg1g0ENubYP5+4/OQVnVV+M1cnOsCzvH2U6NnCTGTtoNZKd4F
FvFtrOLjE0qEPUbbY81znu08MiiJ6WALoz0CAWkpWTgF9l25neF+HXiig8u6rWrJ
YgoeqMfVRaUx8LrjYlx/l9dpu6l7GVB72iRFCCwvgLHxnOs7nsF9ukkuXVhngz/q
xn+gZRvA7jctLyIcvyWxY/LD5Oan57stt3ZkLM2ERznNMcPzcci+WNA1xWVV6cRG
F7PbUijo6yy3HliSZtphTQcNeAwL+6yW/ujcncOk+sshMClDpbc+ZS10QC0dCCGB
AhS1hH6qjw7PvenU3DSpawUyxQId7YWfv5GVwIHvkKUDBSS4HM301BEZGYiOFvkS
0NALa3/e+TvZYTOPczYmCx2+2dkPmCARCPQ8YBKIdkNONaUlzNtU1G9euYgyG0ki
PkufysSjfN3VksVQe3rLrJGqvZulHN6Pwg9f8SAKd12DxZH3vljLI6SX+FlHv/30
STK7VInFWJDgoJMylDjlzoeJLR0uou0lRSMzOYV+h24Qw+NfmYSo/kSHlIDMrTGm
gfK8wv2L8r8yM8Cje1GZ+NERiZlVk1qagTO/UVoCyjSK8f+GTWJMFrAaO9c4jt/g
fO/9dJJOJQJjYRIA+EjJKHrseuVt7iYVSQeR4FRoicq77ZWkkvFHq6QL73wMMi2m
guUSMiZiUNHxJ6sLQIhf9nsLkYDMYbTAtpgBlk+8NkS7aO2DFvCA+XUMCW0cEnvw
rWivMUxiWFVCgf6Z1dlLdo7OYNYVn/+2eLXcODivV9o3kf60kuuiaKaeFvavgAHJ
kFpMrfceUDIAF5cKaN62785l42hRZT/b31am7D57k0BLvpwb6/uwtMMsyDl9SOcK
ypqPfjvYsXVTMOFYq9gbwYhO4MjfGZFQBeGprIkRiLJKiDYSZLdu+ejE0V4WENU7
F3qTy6vxsYbNOmk0jV3ls9kLKq/LBelcLj4tk+K9BvW10FqWgG+PVuesnLmabQoM
D+c5jfBwmZZtT4jyubaIDAvUqkir3G/iauidod7iJv00awsWPjZVqeAUFpLecVHQ
vwnq+I/SVKM7TTx5KNW1A474dQILsWqSEVDA+ExbG1TGgCk7jHo/k9dI0VJZeYIF
gYXcuU8mVYsEpUZpS96Wg3kBFUc1S4oJfv8gjTRugoAs41XDfqOM3+NmchFBcr/8
vPOFO6+Sv5t1SFNfc8jKgtm+i5ug54qUWue6B8zf4BIwHB2bVRBgGzDmRWRJvWCb
gzd0CkMmXMVlv5Ddq67WwXx4srHO6QnIm3p12UVUR+4KwVkty54jUcRAjsrfOeRu
tOLl974mUlEBAvIS9bY01JxvFhb2mU5srLX7ei6kNSFHfcHdEHd6LVnWzCzHr5KK
aez26aRB5ea96dLiiMGS2pT13L3ux6d/JwSZJksm3srg5m/F6699fTyKysTKS05n
CHF0EGiUg0Izc2W96mpTdk1bW+st7lmePrilwl2sJL1/oOiawubrYWTYm26PnXJI
0iYV6ZeSlUvZ82sTTKhuoQ/DbFAO1mf9WfO45lVkTTV4x/MosTau6Mvq47FxK+er
yWL9IQD8/QiGd2ySczUV2Fv6d4FaHKeucdQ9lRQcmQDqjnOOoA5llsfWwxvHW6JB
HYLdRGFeq9kz4nHfg9/Ed+1TCYB05JE1WgAl2nwlz5+LTFf5YjovMRGsNzBlViTU
/xgFc4+aMtVuny36p5k81An3KoLPzCCjLuh1GfkbpaSH5Cmq5HjhSJNSrHjp0INs
lVuD9KVZLSfFVd6qBKuHAIuEWSmbvghekZGTfqT7tMs0QhW5/1BFsovSUMySiNBx
LDTSiCL/JcuFdaOGK4dSsNbLxGgsv4ZbkhGA4dVP+o5rFgD/0Yg7xoZEWtZTi18e
baWcX2HkpRz0hoLpGxoF2w4YqSvgc4UWZScKw+NDBO9fYzCX/kasrLumzE2Bhfjy
GMwbqBQkPKSxi/bOiZtvXQXbAupmg6aH55xN6Ju+d3HysTNoQyP/n5z4/Fu5gbvW
Ab+7dNqsnaN7ZL5Ut1am1XFX9NplnVvUoFkYIYnhCHfCofGI7NGSYPr0dqkZN2+I
pstF7Mslxqhon4yxOpamdgYk4g4IVLKV/io+XcBPgWPn9X6UZT2qDFL3bz8cX+K/
wtmuD7NyEEFwjao4lDj4ovVT+CjRVpT1JiN26zyc04xmDrzfDBSUqVfOt80bMtLK
VIfFcT0nCj42mK/suQQIsxOlQyM50kkA8CotsSFSNrHhLo/SLvrRNtLNxO/G3snj
CTQQxVCIkCt8flFfaJmgH46UkrgvykiJBSicxbI00QKYOXV95QciZK55phYvGbKH
Bl3BbhFakQdMYom6QpIFhAUM1SFe/4szeRPuMMNl2mSbC1B+gxE6p0Ldt8S/oq2k
T9/sOx9LyFWCb9eq+Ldqt2FibD5ns/+kUhTIPjiEE9P7+VbtuhkaEcEg73UZc86G
KJqqLzYY2oUJfL6iKbslnauHyb1mn3M7m3MEAJnNgRC6IGRvrrl2otXkI5gLzTvJ
m1UultdKyYC24+2rT6ZzywKm41IrUfasCGUlHQ2AbhIIz1zfq5PInYwRCcImweds
obT1X4xC7xdKJWamhAp5wD7nKlZMZsO/epsYUkTaKQSD73DWOcJxuM3IKcYzU+7K
rEOHXwfHX7K8VNr1+HrEPpoT4ntQ1nCTlZ1jnTylEJhAAq0HTxANIKay/Ca4M9pg
jv2V7uG/SZFZWbobB3WPjIPgDP5uoBT5aduZFnOZxqZqeURrM/bkXCOKNT19hQHH
7yClEon1gUyQH5p7OaTOhtS0P68Ui9q9T3q+zSKy+W8VyrirJ8gCJ2SVjzUdiECj
mmMB54Epm+yI8mgkuF/bEYxflCLtDBL9E4TKAwRazAJvJeQjom0b2kfV7yhlSVyp
NW5hAxLuiaNkZ25XCSbNcADNYjwZSF/NlIhl80TPGxvvz+NccC08+YH7R82ZkwNq
JL1xkcxQB9HABa553OhgxyPRtBfK/XYTn0H+aYh33M43G6n+H3TcxbZY/34X964k
EP7nOv1EMUsg3v/uxY0+620bfueK44bb4vHG02Ur70TP5AF/VyOtWrGqqyWbdf4/
7GMPcMlUC/hgXPw5iTHiAUAzc4AzbuQcR+uHB9Emp92bcZ6TnOjuY054ZkTrnc20
aPRTDpsFys2Tm7O6B0zq8JaZyanvZCFevPu1M/s83IX4reEmYmGQSOqBf555z7iO
tSVNs2JYhIWpkL4W+3OSl45KOniEH6DxcU5FAQRPGmsah8+y3S4OcUVJpKaKfpdO
sJcDxl9TNzs5elJOWjHkeAhZLUmbyxOyTm9hAT2VShwKAOvHK79rVu8/VaWgDWk7
CKlCOLSJMDK536vlYHjy36VyZJkboT+OyNeFNA4TmfsKm7f3/PNAUsDjm/0GVjSt
eX/9jkYqKKxNS3RYMN4KeSbPFLilonMUIrXQ55rhQU9Im9kuITZJt8zJwm7ChEVp
+nM+KaO2Q4C/iE9dyp8/Z9RC6/o9ivi7/bcujDKYojy9eKNV+YVEYifvhlPhz7LQ
ETpCTj79kuYhXPT7e2NQx8t4zAI2gF+m7+ETujY6JTDCuAUSFU030xE8AO47SW/C
zOqHKXDJJfTrE0ieHAWTJIRnLs8yhCfMuH5oSICe4qt9ehezH/hNk/a2fHe/Mw8G
MjjVsoyagjhMbgW3UmzXBUqG1vLE6I2E4wWamoSTfJujeV09JVvcAQF8/GKde3gM
W5A1Wu2xxZAXet3TgRPKDE4U7jxm+VqyaxSmHavYqOpjgG7IPL82rAMEGEb5U0rb
xqaUj823VgGSlb3BEpnWpcwozu1msxIEQxcndlsAkb+bmPAin9tzK79BZT8zF0Tt
OcB/V7AexI2yaPyYPknDxYEYKa/G7LA0TwwLlcrZpN5hiT8M4z2NwhTzOnOHcPb+
np/BA3aPWx3213T+ik+kFNpbkK51HX2+XsWlRRc+yIQqgGZyrhvhsrniRhS8NvqF
+hTFhuAWkPQlhXnpZk0lsL6lnWxvm+QOt6qXjJIIOjaSFcZSQ7tcYwXou3yIZjAy
6Cicp0NIf+gyetQinxjaYAuHt61IHkPO+vQ/oqZ6kpjGo0U/XKdjOza4ldDZ7Fs4
nGqSW7kbbrGivp6JpJemiyqw1AG74B2M0sbfQZBMPbgcpbaMlcV6FV2SE4ihL89p
YENqN8eWPkZbnHoxK6TlabFVdAebfkf6lrI0nTiNHTsDovea2yn8+L/J+tYUGJqL
12Q5QpeYZrn9UtpPUVbcaD1XlMBcwaiRGLBGnGrLCq41YxKXHJQ5Ah2haVDGqSXt
r4L8zCc0gTRPkS8OT5aNNzDoCW67U4cKIFC1rt26QbQ0VlXWjMZDwtFMHHyslFYC
uWM2VdKHEHsptv1HyByvVab4exoQN1f2bVhy1HYm3zbEQ/+P4ZiFawG0PiYqUDl+
SYdJocAmIo16FRTnWpHVgMpeiOam6abe3KNMy626pNKprMNqjSiM6LymEKRzV5VS
w+E5ktmfizD8ovsFM53H+GewwbXTQu3r1rIZQVXYngMavcWOXVpdFkHEISlhT2KT
37MVelulxy0IYKOabcoXx+6gibIrPBbrGe6Sk08iA9eI6VS/lgVexmiLNz0WmZFm
bDbwtf1sb4JZAsG81WvedRqVpajr9NvAzZAfwy2WeuqATV18Gj2BeFIEKfLUbVd9
i6sEd6dIjKZrykW2x9vtYOb034KvPlagUjr1TjgoYUW9T4MZ+LdsouCPxF1azTLp
//Q0kGJhMSlBPyD3yNhe22lx2z0KWoSBwAurkie+3QyZUGOv4vikCHVfRJNQXliO
wZYzPTB2uWHqgOp4Js+5SsHkgwW8kPvWkB7rteYo9YMbC2RQL4hQY+vkHDEBfHPA
HWL6LPIA37fE5Zz1ftcqhfvpNQY6MDRomkyzydsTTGqnyjHoalFXHt2Yt/AggIEi
ASoEt7jSmOL8TPIGFsxA/9EZ92iCGx40vvtv0XYyOAGulh9lWfADSFdYKn15jl0X
NAqzJNWVOHWQCbf66D59QHJVZn13mZCKymIJ2hpTD2wjIrBaj/nsHanLaLTxI5zn
ETgevrw9EwBewZDAeO/CrtK/+MfbqPBj+96YOWG761F81lWtq9fO9WDKhW6OdSuX
PKTxDtWY+zO3X7SVoVHhTOL9m1t95WRm8gPi5jnlLnK6PN/WOaXJJ12kmdV5+Utn
xDdQ6mUg8ccOl6inYL/kv9+1bGejKbunuT77dZqj7Y+fIYzmgXDvR6emHeVtvPfm
sJNhmCgIFyG8Q94uf/SVwBYP3/aaiuark/S2EjiD5uufL4nD4GmfZKI7bKtBtbLb
lcPbeKeN6UuxTL0ap/ne+3iO6i10vz1bJN09Jtqfy+nbXPCyXmdxqk+lXgkrYj4h
QPaoxSuoYAvWalawnlWojldmVpvoDxtstqwLGK0DC5vHun723tdtAe5LB+wWzhnw
2l/0ZhPNMvtmGUF0ib6NgJI5/pDa8ePkvvxAt09Ubw6Kvnt4nZXAzs87fDtoSnsD
xMjuWjeItJJBOK+pFuEcu5JCxpwPSRAmQ9BLsVDap6Oz/IsRx1yPvATyYgeMTGlI
X4TseVPtW60TOpkQqmzjuTpnFqalhhiE3HIVgTfCPmJPjUoY1pQDnXesjDDUS20k
wgJsx+QgnnO4EmN5Oa7xYCK9k9w6k1MuWorvr/2tq2hIRjLCVDksTwm1aW8anSm1
0GNH8ZCz7/tD6n6HaSy2M/gomRAhZdSJyzPK/E9JcadGIEMn9cN0xFN2TxDsgOOI
1JmV7nM6njMi5ejURBfY530YGxu09pgHJ4FCruncaupy9UcV5VDDFMK0AYau+FvA
JhgfaQ3uLMGI3kOEkuzpeTER9W1CwOUTEddkRPcKC0/QplFBn9OdC8Kua9qlHp4P
ORI+gz+5ZcYvypKzIBNLjGi4QWE6forfHhhwzz1BBiiIhaWZvyWuHsGikyyGEF7X
nS1PKLEIw6biRC56gulePiVMuxpFkbYRfxXWhvHkuSGXnoQDER05QMBbDV8MpfBC
VqKs61/L772wcE1DtImraX7/pouTN52SPcqoCRx2fYynrwDYuMTf5HjqFtlvLQxW
X1zjqafWGnQyfqRwRrIvcrceo6gXOSyUsHcfUTH/XoF+MNbnia+LfhBpmxohDHHc
4FCk5vbi7jO/x+ZD8hPTScLzE3E1zWPAYuqgOX0HGGDRNV/ovfMExP31bzAdLaUB
73/z3V3hWWJtZ2Df4Iyzh/y8TjAdg7FMUPaTIEop8DbZCgJzk331cYA+cquEZ0Ub
v2/1U+5Sc6HoHUhwxoj3MJi8RfpLPXxx5YF3z3ki6N/2uPlcIfbGXXJPO07dk8/g
yPtNHY7nfBTWzlf2jwn90c7ZpRM30Adn+zKwm4x3LEhbBKG1ZQ6c0tFKgqiEFvUj
3JMG2b4gNN9G4Mh820pgyQolZ1/Wycf0SPktXZJG9AuBIxcuUuYufKc237UtEtxt
ELoNSvjA+vP8L7tbrUr2Xvog/PAcxTAmQGKypKJi5HIE7v59U0UjW01fqSxX8Pq2
OopLlc6uENhWvMaC/kFiov/J7UCX3exOmMhaoHwwqRqowwNZNqtaC2cQZTNT0ihL
Ejy1lTVp7Am9JtY/BJOPQrdM/RCCjqKpvjxEBfk0bal+bFmyFNGpAU9xYJB2lWbN
fDJWnZ/L/FSjBSbjiTFvDwQ0KVlu9EgyHF1gEh4CF72+sg4VFXxwPfnOvIp/TW7e
i7sAwkeKnKW+j7SmxK2fRkJiI76aVF37FeR5JCRMVZpPOUNyDCUoMHrQhSpl4mvU
uWCgCHWNE/Fy61OaRZ0ImHzXovqRrEqCf/CEXmk92peQoFBdKX/QHpJ7tSp7/ai1
TrozTpLmxEHhkl7cOlbKZbd2jJOv1jtzDQMyvcYqZo2gdoruOhMr8A8948u6RR/r
bK/MPht7gMCmQEP5rOXviGOcGtu4i8/VZc+yzHi5e6G3BB7SeAlUqfrm7b5a4MpR
0Gb+XJ5tabDJZxBmVAknkBvehIeX5blIdHWlCHgDwGtu6VLjC8cC2ObA79KuU8Tg
CYU62OApC1a0Mnr0CsxEaRylFRasv2UNxMdg/577j1mfEnL9vsEZiLCYWvwRN4nZ
hqcIfQPKOIn261tmwnd2tDIa+6poOPQWe2tvBg3HRK7IYYnYJzb1ehvtt7Ma42cq
qXo76FAyv1G3EawQQJ/RsGSc9y7wFAPUXRitlSLHmbsJoBFQsTUa9nUURwAYZrvy
B6xZAOuZkGY8sJ0CHlRdulx1WHqn1lV0EAF/5hek82eUlOhIGmm7WEqnGJRy9+zm
F3fsDG2Nfo0UlYrj6B82paiM3FM79KUlDqFRuAHS4J+urGrBbVj/+hQTEpruTspz
yNPedSpYM1isr64fuRO+huCQtehiMwALi+bXmCKS+RLZ5D7abhp00aOeBnrX197e
Ci0vs3U5OwbWQSz7gNqF4PbOqb4BlJXF6AMt0OXKAONEu8szy9GuwKCQanVCZZrw
sZSgsY4loO+Hi4xHf0vzItscoukgtDzPm/dsMGV083B1O7eYJsNW3Syo0zBJaq1a
JR/lVnvVjdmVDH3qqtYYyPEPpCHfw4UaKsoHYGbxtRdXWukZv+WnikiP9C6ojcgF
u8c+Hr89BzsTQVUUwD5RSSnndKv7cJ68citVUZMnRvU/ubMNIwxYqQlC7jNOg1s4
FP7PXlsE7jhzKiKXO3hpzTP3sPoN/zOMAeKgSt0zCBWfPTQ5U3l+rrCw78r9jwZF
FzcfhTQbTzovOKwY3twSWYEU+NxrOUeQ4l3/CFDMxk6+J1/0pUMSLW5om8mM8FkZ
jJB/ieMRdCvCCLv/+2bWDA2DhbLHPccH1xKHrtFuoyO6FnR1LMiUSAKjesf8fMRK
LhM0mHMkS30tz2UErhmSfam0Gyiv5XvL1xA/tvkexXvUo5B/IG0olTNAO70HpXRo
NDdNsZelriwleYrmDGMCmS2AZk+cRj46qUjAx/JORhFPdA6/n6T17YMV1JdJd+hN
lMI/pnuxC1jFdxk5/dW++C2cFGaEPKwlAmAspiVEfiMuz6L84F9QuyrKFWPS9L/G
lUUPx8fkSBkW8Lwp3bTE90+eO4LxpHlOxe7oDtVtaX3rz/cOBwwJ8Jfbp25WDz9W
EzM4HZDALK+cr33B7sN4Mxk+l6J73RLPQkzAKO3DLBDUnilTsosywpW69EQeZJV6
QXewspdMQWDTc9IzfcMPPY2XIm09xjxAiOJYoojjTiOcUiB/OhUok6Q2YRvH6gRA
Oe4jlgahtzL1ccHIFymlUk8tNBrV9kdm53e8CFuHbyhjAImjOjRtA1qffLG4yyDK
HwW5++4tbDQ3vGy038og8WuiM3aJOtzEZ8t1EX+/6H23Ezg9fSwDIPYHJD4buxQl
TKAjuMHCivAAWHcOdwZ6zRk0qtylhzgueOjHNu+ii+RnjqYzYi8sN1irkh6yYCC3
1OOPxs511yeLQXXdZByqa3ogtdpxVK7wqeXyhQT0LpZZsub3ISHq4Bz+zNRFLIon
g0QvV0PXoHSQN94KHSkpCDLSI9pe+E+C+1CtE4VM1FaaFBs+Bzi4b1nXsAiJqWxf
ejb/rN6TKIlVTQF2Og8l3a6LaHIOkNktrrdXaGjR4nrJtj+VH7+fUb5gJeHJTnbB
gNNO1nyf54wq33r+G5YnIoiOOAZP5VEHbB7NeCyTuCq1Bk0/BKDXCMnqHmJEw0N1
NR9j65DPICJsWBsMp7d4cqZofbGVOlUSqTAEIN9z1OBD4Ix9RASN2LhwvpXrNA38
txH+PS4S9U3MPtGCeXgiqm4+t1PVOykVpvdKNQmCB2Z2WFaa6dq7dKTk0lYZ+XYP
cVuaB9U3LWukB0cZLmTQP4PuUA8xBy5+bO33Pks0YbEAtW7sJ+v/HMEUc6bG2te6
/inON/NodiyWWHBRlwuM79bYl6AhnhKXjDYyd+SD0PgkNalx+qa1hDUuQnqXZqQ+
NXaM+kioQylK8jsbMgIvx492PLe2AEvcqFX0KzxZWmeaYgbsnFOo7nVEkW20cbx7
8gLj5ShNEDHAmLiVCn07Ft1o3kwuFgSVwXSToESSjkt1V0V2in2R1XNr7qJXP8cZ
m0xzKk4THqvkAjql/SFAyVzDTh0kO0WfXO1vQZwDmXiqCYxoaY3yWFjcR8jYJYt0
QwCuszY+q50klrquSr/5RbdNKu0MTKtt7tK052l1X5a4YZTxiTft7bfdnrJUxLzG
kAn7bzQxsSDAc/xhvbCOoFW/d7GO70nx3rVrBUnr8hOGMCzLK/f8lvitkA534+0h
nyGbsdKUyB55V5TB1bu/5hdlpV8O1OOQwGSDTxmOUEgjjdgwGWANo94x8VcSwtIQ
BnKkRRUtKWm97ydTPaemGVnhCsGv4ohs8eDl4ksCBvOgBO1IMfPUMz3f/hNOhb+J
WR8pWVyD6qHPq+S0HmlTfyXe4o8wi4ysZI5CldRraWubXBpjRr7T31tPE8y19qRW
AwORG1mUo5EE2KL+i0IqQK0vvevPvS0U3Uz5nbtALz/YjI7hJcybOhsTmhlLxi/g
oY9KS3dkVWRitLhp6qpIxF1vWvQFcobSmmb6dZYtvBVgnUD9duuohCaRJVrc1l44
VhvZLrqSmHY8Q0tCTN96DDBK2/Z6PkS5Sxg8Z7MlwG2XXa2y1eocRUEdKfVHqC4R
HGsbsBzxdeFugL1b2FEwWet+QOjBEk51D6JBylT604vWEFbsJeds6VFxqdX57ZCZ
ncuHcsadbYvyRH0QTxvLLYKC2b1Wus1CQB/aUtbuZ1xJbmALqiLZ/PebK42Tf6Ze
/QD0/DtPdAoawEUC/13jXDe0SdT2+9SuGrgMNPDDEzYElNeNGjEZOz1kT/ghmEAD
l3fj0TpyVhs+76Bgxfr4RihKOUyjuDJPYD2zTvVvcFM9HXoUBkVd5rtjcSe4QeDX
HIrlmf9nHPNKUYhckCHQWbJtaN3Q/PeXmvyP2StQh4oR30TH0wo2if0W6s62mKL4
5FlNdm2FAnTHczrSf1gXduEOijkinRHvM2mpFVePP1OFU/bgfY4fwzmb2uYYtXk9
713pBVy08+CtAudwXvvfmx7cAAukNOSGZ52McpLZe+qntOcxQPuEF8OMP/Veq0kp
RAi6AaxE614PV0dAZqCu2SkKYOZ/oy7WSs1NxT4wgpc+LmHEog0ww8HVZACHoPyN
vpDunxCAXAH1DR+E/4zWboF/Xp5NGKTKKl+QU65/3aml6DeC1oLtq3cLHElNvkUl
pdyFqXvyAaK+o5d8MPMecqpM7MxnSfwmhEo30BfHbDz1ZdnphmeGQibgq7gEHO5e
KJZ1VnjU99dgXdcLEYCi6hwWuEffVBydBzrI/WTkHzSU+eiaRekflbA9B874R99e
GLge0GcHCfJTB28lgLHM8t5sPE1pweE12cjsnyNgOuf4Psmf+Eo60J59E39aQobO
hStgKsvW4iI5ca7pK70LppAOH5tFWiUwd4AG5yIuM5xW6/OueNxLBELlHvIarsky
H6aWaeO6hGDHfAkq1BfMsUsSZnoADZRCH3c4wclf5olZJzlFWjnFBcUwJycLFATy
`protect end_protected
