-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
fDAlW2uazN8iou89LsojotrLyw7GGnxXtoJ6ayhDVzmCUfs+1Ek+iD8A/s7+n312
3XslCiIuV6vEgS7GLDc1bCC9s9rsUhQuaUe8C+pQnrPxsm20o3ElqRS8Hh5mKddd
MDB9u/7E9BDi0m3hcTK1rKheRQspgLgzvQbFg62zrtQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 34687)

`protect DATA_BLOCK
h9g2zktf6apkH79vAAqr9Mt/9OOxnu0dUMyys//CSduaERpDWQ/bhROc3jOdPxYK
ACa27v8GwB4+3b3rQMokm9+3gbx4+JtvNGsu8Y3gxsZZm1F9Zm5k4h3b934d0zpE
HoJ1PmycoAa8aWdAuZzXkqpurMUoSAdUIfriBYWYAMoIkh4WCo5pYYAglpXIrxkZ
+Tmm04q0cCTvUB2UIJUjMXZC5791eGE7N7JNVOWZjNWyTYrrjLHhzJd3GgjZhTC3
KbWsaA+BHvaGMZCzYx0HWiYXvSWy80bXXABchEAvCqsx3VHLVwSAQPb5jSNbcpeH
Y4agbNSkGqDPhFKk0oxT8l9/YigqjONMKzo1JsQp4Xi/jTbjutOK/NdAgFF3IGvF
uVR1GgBhQBBKm/sHimjK6E2aDnMFGy2KFRSz18GkzkAszDA+u98R/fixzBjNRVpX
KgLFhrVPrcDw5jrUN3MEZNF/qGVRlo6G5hURjkHgh2Km816+R36FsnkhXlWFsEKO
TWQVbe+cXKI0oYtuykqzPZp5rhDCQCSL8CKUn/bmNfGqGL20f+GRl2XoT5vawZCS
a+UFAhIeK5zPJJrjOc1ZFMjShcugGXONV8Rlg6VxnBXmnyPOeIkvUTB34tyTcD76
TY56MNrzvL6nYxXfNpUZHezHjk8Jq06reFwSIZnGVEmW/OjMel+BWSRTqNcVEv/p
FDYc+eZYegFA4LZ6vbaEWWx+7kdcDmuVbyLLxzOYADCPLwk73OL8dyrww6geCCxN
nhIe6F3oaeQ5ceQDBMOibE98tP5yLE0mkLDMxMKCOWpHft9HxEW23poyY8wreFLP
J9/wozhrabX3L6u4s5r9MUBSHBWhHxl0Fx7ktr+wTahrEiuABPt7DLBNwLwnZ5vs
YCxkfH3W6sRdtxWWvMZMCwJR7HXrPItwbnEP5ST+TsOL9E+L5NGGmCgesqHdSsSG
x4wpI2unV25dXU7zoG1Q+D5gWudT/QctX8Cd8ge3L5dFlsB/gSJkmVvLlSXE1zyK
Edahik8tmTw3gSDu2iZcMHYkDZr7ubTzFP/vkcl1LvzAqJjJzDQ5HZFf5vP1eC2e
lQ1MuJ58bj5PnaYflvn9YjblKIado1b9250AbYj+AU4dzWNZO8dFq46eXhht4Pkw
3ylvZ81H2f3QCKyiYn39dajx6D26+RkzkvvcnYNNL/cJghuaSqayevO/RrZatr81
JE6ZVVz+mXXZk23fTTG6R5O3QTtyGgk5yYcFRVLVbLeimXbHafmvIlVGCieSKWDd
zNT9N5a/+6NGE3Kj6r/E07OWyZWLn1ywG9s5Ef23SxCN7e6S9L7csXFQUt2briN/
Qj47otYPcJPYH2uC2NZZAktFPcXV00Ty2QdEXUTJ1RM8cXL1y7issGWv1R48VMpk
Gq4IuFJYvTzpdelN0a96DZiOlSJ5a8CQtxrZ0IqORtJF8Jvt54qceMdbFjKa0BzZ
VD0f663q+GkEYawX1qpHrJgtoI+NP2YWQkOWOPPkBxzwRHVluodiU+qQu1j2Py0C
ypU9ieFDwxtGppUzZdEPayDvJlRQbb6if8EQxfJQdSFUa6BsGNi/TO1CLwQ/dYDh
J+l+lltZm1kLM6FcBjK/J/mijEo88hZdMDbWP9x3dAveacdeIgZNv7zLBbiIteqM
UM8zxauRRkiqXNidvGEXQ/cbVYrU4HIGYeRePvQ9GHUu5HdlYJHBC+t6TV7MRcOB
T4jkogIPW4u77Pa47ZgzEnzx7gL5ChZ45Eh0Rcyrc2k4u6euTT7ipoh3MwL95v5L
QqZfAY/S8JglkTBPfPyiVVtaS8Eunux7BdcKDlTR4we+3YhlcfsG9HtjkK/nxtl+
5nYkr0cN/15NYC3zUrzq+wzs/Djw/O9LtJuw31PxRzaoxBICkP+6iPUV6Wk68iMD
dVPx8ahuI2cPYO7r+czRlNRVNRpt+ffsLtXcBWUsdxHA//6urj1LCyJuW6UiWURk
ayEagrHl2hlUZSjvaiywDwD6BNww+obVlV4DWQ+VZ1yyqIOp7ldOcfcevIfDBuEF
WF1QZOEgC37ISroRucLAOckw17wjvAxBPwp4ONvNT02zCuVFdNWIhAmY+dMiNZ8z
mgYXdXUz3Y+lGKTxs2O28G8EuaL+Bbbs9pA929LCDOxnaBoFn59spLUQiVe5fXu9
OTP/dXmLWrqKqKgh1BVyK01a5tfOQDzd5mkIWbtrjj0m6oRrV6IxthJaZsnHmyTt
K4MJNElgFHbytwlHppsXfSfSlnhykIo9JE0koZ88Qg6262EqjIoG16kxNgLykMGd
D6tUtmiAyb78Jj8zUwVWT7188MGacToBkJlGOIO0EafCFoXIzN7g3BTRC3fo2rZL
Bgrlp5/BfgluOvOtH1KMv7PmKBeIuTbw9iM56GMKsaygHnlRxCXMSchAe+1bfSmC
S8P5svqqdHMT0TLQorAQXB5JNPEs5lpS64R5B6RIfsbSj1Nd9+yNxmTr/f18kngC
RHjkRePFMLiqGKRvicz95d5L5pyWVCCOOAe206UacNftpxM4Rf5vydyvsAtttZ2R
5CEsKyUwC+IvhnM1WkpektC5jmhT/SGNi2cd5D674cICE5Za7FFH1lXO4IuxCGiG
SsxlioeaCCT7zJPicWatsu8p/lDN8Kc9hAkXjP8mdeNkm+1wMdUx22l2Br3aCsow
CtkklOkZbh1FvRRRrxmaNZhTCNtq/8/6h5m34bclAr4txMWFJHEuAwdehynWVVwQ
xrrHtwVrIT5Pihy8CjuPGt3igyh0XocRW4c7ESFFiREFP2ZjH/kqpQ35WBZ4POw9
qFtU0e16TZNhurNkzBVphRelJE7ftK5k6IkUa9mcco+xlixF/N5X/1OEO/Cq8WSy
Vnh3N+vcxOenv7stLwYR2nlkWvAUc/OHeq2cOqlszvmmw+4zEH8nWnzC97Z3sd3q
eHLfTKv52HL/HK0YahXOlAZAxW8XmtAFcO3nsrN6WIK5VbVfa/ywxKkfbCiUsUB2
0Um1pe2pOmNVqVK0ETd4mzREIHeQTpZnVFlg4DQ0jb5aOmGIzw6ufBT7VH5FfSnc
wvDY4b90uIZoGK0DLgnAV7ydu+Bohm3/h3RcCpwaSaGArwpQTQUQvFN2inQeY/uN
Ua4WdbkacAV200I7IRJ2zjZjnKz8roVc7vXu7n8KyARpM5fggnI2Pe6Dyf6So6t0
JTgrtPDA2fuVz0tVizMwmXQtyPsEh3XY1gYNYl0lMMhMf0yuVDcZctQrxeFrPPgs
GSdi8RLbml0phICk3MD70L/EwoGkY8SLkbXwAjjdupdC5ieNshkH/AqRVryVXari
iYmIVppHYUjc+XKv+OOLpyBwVImYQM+Y3RZkHCCnM/z0/IsH5CgC9qwNUT4hYFQm
w6/CTez16IH0sqcdjTeXW6S7AqeC0hxr8Wm2OgqAGnzGH/gKh5bmrhNQocpTQqAA
cj99cHJPgRuh8xm8jotplhmrTlFR513pMJVRp9d892mQpxh4HbBc2REYHy/BlvS6
3uvPlOSrwj5nhW+ken5JFExwKPfMo7KfJkFhdjN8GdVOH8gi/2DnVS1V9ZNbRQ45
m2K19CZ2K8RlQun7TAirN8I0FXxUOkZJxTgAbnzwn4ErkYeWf/tJHe3jtOaSpg3n
memvABivjtHPTmTj63jYAGhEK+dl/LM9sOIMSvrQXvXpnBeYfN4hgmB22wdGDtrx
tkz8ct9YsU9lAgcV4D9wRLnCn1Ec/dyPpBxjpR+cACh7nwCbGt9uxZw0IowOoYTi
w4uoD7ePJgkLL/iwpDqec/MaXzXxlCQsxKfAKajdvdbBKwIxMJSKi8M88H0nXM7F
Sw1+QCXBETcDX2cQGKTmGzElOgN9QmSBSM82m0mis9C64IrNrxeLc0CrRuOvfb++
ijlcKLin/a9ZI4A34wDqPCNqv8hXeBqfxOR3j/y40/RPiLR1Y8Ra/vyMl7ooBvst
IQqWw0bpmWRIHmD57yv9R4BEqNsKydJInl1vO/34ZVndJjdHR6ylJdH47HnVQyE2
PEjboNCLwHeMjavnW7RoTCDGvzfR96shfUE+gqzIcPoMWCVFmBSfhCp5h+MsCcnl
nyP2Vm1nBqRfE5njOZ/Kvxob9rOq8G8nh636fhiuBxmweTKc9N0ee2vBZ2Arr2dT
1dl1vY4WzatkntbITzXfJzPERLEtQ7eQHAFKaC72H3wJvbL2REq0Nd67v4/B1W3Z
/pJG2JsFlWnlg8UObU9KEv14xinGR7+xmTlqeQHS58c3+TWqWRWMDSEBZXoLO4gQ
vPgK/MlGdYnbjxSapWSThpkMPe1Gbq/Uh5GvLyhTSOrIbsLsEcJupPKb7gmo5Xvj
dVPgZ/WvJpA3Wnb6N1+mF7uFSwTzjM72b17aewgVqVpuW9jNKzQWVGokZdDRLTYw
orY1zn2dflc6fHeRUXZv8LL3nZ2UrSkdT/m2OOGJox7SLma4qYxnLSiTR/GKo6ND
MO1sUKYFTNAf9XfHRNVw84aOwEi3WUlRF13d73OX257u1M+h0YegtYzGV+qPrltX
qDQycn9zKUru+TvDnfOKbK6bq5R5DxX69A0stAV+NRqyKBzG6oZ9jl6PZ3KZBqsX
I5kDvxaYTeVbw+sm32T33Kaf4+e/HKqIcrsUWK5o8mViJUu1uQOOGWjAKzBPSG62
TxsOVdvCuaM6HQ0kYh9i0GIhmH/APJM/UqygbAFpcsFUD7oxDSfsmplizxSHlehH
ssOZSrTwhhdhrD1ytqdKfomsl2gL+Nb26Qe7djQi92Kp+0V1zfylsoQL4zpkgD+v
vk5FeQbsnSsg/84g2DeXya/fUrwDg/DssYXIw/1xP5U46DuuZ3nE7h18+HkBxc5F
eyy3OQxx/8lkBixdqnZBAmM3MgrO1D7nguA+1z4nqLGN72BZN3mDYlN+ORnTBXWb
YtYE+q1CWPYooi2pQHIOwQP+s9VSQLIt37746nr58Kr+ivbdzRWxsgnF3VVuvxgK
w8oZw5ofCbA2riwH6CMaMabmTuTAkCiSOliua03oRRFZRCWGEQdBQZyjVq2gcPJW
HkjPMBLNz0/RKvJd15rp2UiNiOLtHUNPCkZxZucLmFNjt3jxbHujJfWF62MJUAPa
9lvV4cHvQMo7mhdNq1EBwOve+otKlUClW3j++kt0GfXfe8McUeDMgKJRenjHzqV+
n2DjFiX+W3/MiniJvU+uhELLv4uvsfSZBBWEMVHl3aFEGQ/tanvWzypNbyFor8yq
IXVbuIni6IXQKWBaHMQo1HCJckpSDTuuX4XmEjgQLZEycrvGavUNKLlX6wE3lPI4
atIO4b/IWErWcQ1UtRRFbHqgKRfYSmByHn3WEAveMGW4mxiyZVXYbIaJmZcO8jH4
g36hEn7q0UaCxnZqgvSnk6cIDDXW1X4xF2A1ClICGeDMPpikmxj6G/OKb/vLNWb9
haUZ/yk4/m8vJ7yuedRNk12yXGeJX1jMCaDIPvV3mZNUIdBcO0AxAvLPZFSmg6V8
CzrvAh/LHuWT0XDffSXoyUM/aP0TAPV/2euNr6xDc/0aH4FgonqQP9Cx+L2CyogD
DV17H4CebvhoOuUlIRxE/LjnVipkVwMRqz1y6+0+xSNrC3OO7tPFfSrF0vkPeJuu
TR9mFxsRk8d6U52TkGieFsDbSp9+vSK/x5wRR4DDmnaV3jfr8fzLdRTcrib46snC
9YQM48alOQLZnpae49fQ0ElknCXUjis6IEMjGFe97/C2zr1r8oPt3e75QOADH7Xq
Ln034WjAORYSj2SrwazrT4xv3mkXUjh2wTEwvpIS8YxNgYSec5N5ed80zGAWhzOV
eMnreYjAt0qeHPkO07DDWAXCVmAkyNPQ3JgH0Iu1c/SYjgIVrrqxmWC9+PSKjpJk
T/jbaAaDXBU6Tcww6sIZTPY0HXN5T06Aj2aygAXiw3e6Y1JA+cFDWFPs3dR2d5bt
mOD78kwFvBMzB2HVp/FjJxyvljtli5yAZbA5Q3uoNSnR/dDoUzGIAwzSUQDYmeJP
Td8GyMT403PePUK2p/CF7Tcm4szERSuscydPsQlPqkL2JWA1VIloFcimWd28eICw
cfGqHakJWZ4BwHZCLrx0nHB0a8StnUANGReYFiYUeI808Rueohd8Ub9cRi/wj5D9
B7pYbow1PrBPSCu3n04+AHDSvX2tmrzpDmpJj8lgFzcV1wuLD5m+mn0KQA6eOkuH
SR7AExQfd77DhCIFpaw8XwbXiR/hjzehJMxaTWy/May5I49rewJUn+C7wZ/nEh07
9mh5kxkMFNZtP7ayBIXdnO9EQSoNdvwgkzOB9dEwLPL2PQM9pOcU+ASMIMsBsZMw
mJd9WX4KuCQT1YhqQ6+iYkmyRvlvbCrEAX/rNJvmfkyK4qc8xjwn/XuWkLL4wduk
zTS5TOFSJ1TfFCLJzztukx1Pr5sYiijh2B8dAVFqKmUgOrFls8jDolT6tDZOcLGW
Zc2fAGggcPGQ2gHwnT0vUqKm5Hi4VJEF6K3Wc5DRys6dMJpsAizCFcgODjTaNRcA
1Cn52lzdnUrzAClHR0jSfjp6cK5w1RZHqszvt61cVsinVulCpswxw+tkbK/nNSv8
OSp/IjlKC7mikKhWJ3fYmlJ259Zw5714fvmhN8l1yyYQq6Zm+2Uk/dGoff+rcU5I
6TJxQPmEcFYJtdFMsvwbKNtgaDl08iOjcI9TDrzQji7vNttdu6JyFa3RauOyBtSu
Xn1VGwtMjpWe5c72QHb0phs6GCMuUtKOfdHC+GzlI+x3KAL6zCFMjkX7+uek12bD
bG/RB+sffLjdEMR2zfwytAw2CoCIJBVMMhTJf8CtyyGoSsz+E7XYiGBxf74RrVll
FuVmNLd5SUFcIAGW33+4uLGuNwkTAolIN+8I5AcJt/1Q6k4i5MKSGnXuXyS12u44
tYGW+WwNqFZbSsHSu7XsPy93q8Sbi91RVH4+3guv/kFf/047qwmNLCHWSkcMiH9Q
d7l9E4Ju06gJ1E53IGaZUmcgT8O5PbyUfGEJVO9OlM77QVT409xxeipvwOeIfikT
8hOEZ1b4gMB5LXMepFXU7nV1cfjCWelWlDmKymNv4fjPzkVFKk5r5ebEqSTmHLHH
bnn/dkemVTVO2CcpXwwiqPZB/p6EUhhiElmhmfeBU5ZyJlBvi+WwPM/93/QhFfbd
QdcpondWgcjsSzJlMDZAgABvvS0FM3RDMw++nh9hNPvKE7mNanh/hogcR7fUU3n6
29b93vr9autpOYV1CuXDuy77lEMwhDPfgiJs99hrqHB+/pdsjbJrYcr7343S4T7X
yXLCx5+NaNXQ/cOahUJ4kS6xBOMx0h3tyh1VObHWyZNmaJTlofVkAb5UvpsmWr9l
i3c1D32Zup9TPdIE7hZX3ZnRyEOhSjN6i854BM8Q5iJGZ+ML4ug/0zCMsaEMfrke
A1M43oSqIAMWtJ0UBnYZn4aXzGe1xcDaPZntknkOfCUKiCBJlmJCXXbNz1sz2TWw
Jk2JbkxSUKeeaLi5/9/iCfRmm7XM8sBMAovc1bg/YgmD2or+dSCHWDAtFxozaTai
c5DC8AvQQFaMB0UpIYSKEfY2/8lf9gX4MxZeTGh4ElwV2LBPNbRHb/bPySoKKuFK
pjNbtMIoaGlqfKLn0eAGW4tcvzdR6srv8H+fBmN+JOMjq+a0SvHV2NHmuMBgdRiT
mpVsxXE/e27rxr0JMZjSkdsB5Gn2md47cjMipb7DHTDQ4neiji/M3q0QcwqMscra
G1ZDENcN2cy7TrpPBObP1k+5baW/vsONOHPch/Yq/9YHSk2+T5T+gKvZUy10D9kl
hGO2auH+SuyudmtX7R1EN1d+maGBAxwSfuukzvKQ0pa1XcOGK1YllqgBzJgX4in8
KNPiAu3ywrYfBf1ZJvnGGVJg/S9oVo3sq61R6mQfRcjFpXhuVWv33A9CKitKF5E3
laaAValy9Ky+14FV0V4DC+Py5F0fRFhRkxHmhlDDsJSTPdHAepUBPDeDDatLLVuJ
wNPXoK4XRZ7JcMKvFRLSta2n8eWge/X0oiiggm1HI4nioI8CBzg8sJPyUVysrRd4
dORf4UIr7yfh0j8LHqXjBSMNcdTCyPYFOJcS1xXU5jW44ZreOjA6BLzTXP2Fcc1S
J/aibfXQELlrklBRcDtQrKwUgLVNiIF8Y/VaWZ0O0AUf/2Q3eZ96Oloq3avJg4Ik
IIAL/ujvVnahWyKNAoNNiJywRhp/1rELOQorlf7tFYVx8/eOrUrKBO3nrQIvUt4n
nS2zmnUW6wlUmtWSSWPT9Q2hEBJ9VN5dN8F33cyPNuQNHx9K9Bn4Koktx/BFDK7o
wX6wjwdkHB8KC8XLTv6AfvlKx33qFwzn6wFFclMmkzXX6940VsNumdPxDFmQWBN0
/cO2EbwMfFu7tqUEIPAotfDRCbbBGIy8CT0XpMfg7kizHLqDHtccPxN6b6PocCgQ
spfP7hudkRQUZi4tdbhkXqKuniMJCjFPxpcWRGg8PShrplId65eXypom1P6pD9xV
EFdNUTCT9F/clO7IouJ98sPcDmy7yJdGS/lxoOTMeHcd1AjBTSGosAyDXkngKaK/
2FIv3cJEV2tPFDZw8iBZISqOJRS63WqnaWE4cOzKwdh7bqdoBzIY+dXXLqJZXcbs
xeO+YlUV2vkSXwfMTJJ4WnnsDmCxFa81cpRTVix4BFXxwIWdzkFCfCHJs/7VeXVS
qTkEkOL9lFhPg/0E1+iV8NnRnBbaztvI2SMC1vAI3qzWqsv+uHFcU1+fFchcVIoN
LZ0Ek2dTi0CelCr3feE8wxjQVv4z3KqnLbUS7DEArTEwTVkhP7Y7fjgkLKvsah5L
QqnFbDH0+TGQ88I8ocXncwQKkLfxcyH5C5Recq1h96qMJk+zXWbqrXrLBTvfgUG4
zcffjfjNPbtrQnqJQGLr3Q28ULpTBsZug/6fyKd+jWFUtBKmahlT7UKKMrIi4EkF
elq5s1QnBvAsX/7TLWKdxvUYi7iVwmZgSauxfdPJYtjnJD2ltob0Eyj5lqzbYmXl
G4CvgseBojTD9cT8TmDDRHXa5eQTH7KDvOdpc3wv+ARGukYRnmL7IXMtm4M4UBdW
rLSuh9W9L4FDFhG29ItfAGOU8+v253jSxeJ4xR4Trz7uX0WaJtiLGEUM+a1Axwxr
kv8y8ZCA3Ihwu+U9Q7YWqGjjhncYL+syCB20uVPDQ1/E2TWhTpNUY7EkyVBPWBeY
tmFKWhDSvrwqV2XdfRhgcg+PFunQFF6lNax1rOkXXA7n/k90bdAIIgwnTVgSFCp1
WktDot3yMnCH99eCfoI6fXMz2M0ghXO6aeE9jLU8tCrCeT0Kax+aGp17Dw4YfjSY
P5ptS2lRC5vGfdR80C1DorQey/IOrS9PvAkGk7N031LQ91t6mnEYoYG2pCjZrwR7
134J+tBB0s/+p1wyvaKNgFBxSk9VqMPE5Q47/RlSJlgthUekwzbGWyhpWfOLCmbg
XEr2JWpKCk3zOKyGf9lGJf6aofVlIqVaooJ09YTvde4sXlr8RjeJWvPQL8DVM/E5
cM9dchGtV2XIJuiaMVJfEhCIj8ByIStRPHju1viT2ZfB0YqKANQFumeHmgYswMOR
qnxmYgKhfllXJXMKVyUOkYdyccYAlll6id49WcdGByEIHcbqtmZZh4sFG3YqlpHl
r/HV+lQnmdMyGA9/JeZMteJ99G8cjrSJoMy/xNjsOHOLh/iAI8R20Rthr9Rr+sZj
MhWxqll6h0quQyTYJuRf3VAF/JIMxqdiTssQozfKilQ9kCfE+74yhTA5nTclZcsm
Si6hRfCUcIPAKym2LIXcZufvhAB28qNMyIHPRjUeMICGuOzyUTHSR1cn72AnVvIw
18MZZ0xx762mB/Zm4DLGDnC8PtZ3PNEKmwB0HXkc0JBdROCCneuV4+A5H7S3VMpo
QgdSXoPVgBSU3JdL3wjyv+2XlcSspla0NemvRkRZH+FE1vTux7std8cX8WvRXJG1
Y3Zp1JlvIIM/n+fnn4a1jnqxMczmyIT1f5JUNln3lYFBmvY3wf2CoVUKICeMgLBa
wpNlmrCgaUtZO/fT806QW24D+eM0smmEsU1w0iPogtQ96puSb2z8+tdxtHU4yhBK
yJubawWU/CShYm180PmPUuLljjcUibHKQVqNk+HBOEhWWzgHFeIpll1HthzUCtS/
qNlqS3OgniwJNRF5kl2WYXxeN/Hz8XTri0IThwVpECfyEGi9YUXSbSzz7oTjJIIM
UdJI2fbT+U7zMCzPIkKzp1ifoqWmPtJ9zFn15XZlTEDAkYE6hFd3fL9yAqLIh4fm
maVJvYjYFGl9CfIOWO1ouKa+g1HSW0Zu1YpIJjIKlOjYV5/1Eaaz5ncC9JDN9DxC
0NvqejUUW663QNZoJO/Y16dWL6RHjzK4CLsUiVWvPEeKNEMjLZdV0oyIjGRXhC9Z
LjSmncztzPUv613Z+ItHl3i3j45hQOgVa1hAtW/NPQ148voV0eooIkDfMuKOHxgh
YV95SJCLMyOm42yjVfj6EeMAN06KZA8iqjXjSS/uNzq8bld+zwYhn3Ws6ZEzraDZ
abupPNOF+vzasToQ7/wpizCW6GUYaYwuOfTnHyQCKN0Lcwz9y1pjqYlEBybDn9Qd
YB9e8QXivvTOjTVebwr5uHnMPdilhvSyn4Aha/kUV5vU2qHdV7ea6rjlyKHiNQ3S
V+oBy5CJwRnvUUI4YSnmvCk1g+j6aXFLWNWTXRU+gEphXeX5+mcrajyJ7aQZFNr4
9vBopB2lLyw0l2OzVXpTeVuf2zDL+LlH/G+kH7IvV76ABHdX8T3CUR9bCPU0qIAJ
e/59RSJ/VgB3608n/rtwooeOePaL9FacPTWfjLIMDBbf0iuJ6VKehquXy10IjMsJ
YWTgdLf0G0bHcG2S2YBxT6vbUmypsri/wZXyG3CrbhtzQuC2Pze1U0kKhhQbVUBx
emUGSIWSbCSTA3m8KKGuNxnU4Fd3NSKwjtc8yY4Ud94h9NkeyV+iFEos8Vu8Qh29
s7vP0Kx1KiWdH/x02Bb+E6IRnzIVY61oaXuBtA2PxQM3s8g2i4bYW+G4nEydaQRo
T5Y3FotSYpRtY4fQFK6MW5zSDEn9SX05k/6bbUeKnxLCbZzDKXKvdDtU6XX3hqmQ
6TC/+5v7mzQ+NLscioaCwHNOdOjplceXTMDUHUXP2hLgaHbROPDIPsmLdGSlzvmf
OkaLl11jkSk+Pkkg7I1kGdEkdQ3dXbhR/7mcILDHv9JwIkwK7RItFXIeLMdkqdQM
Z+nh6suqTOUuARuXbApp4vmopuo6xMV3oKgDAdR+IpMaRV5JaKA0h8Eo0ZyI27xr
klFHCpI6uyXksVaTL/PRXYC9WiZqvO8Zo47StWYkPJDPOCLl1zJUiZeb5SeB8Utr
hYny9IRSa4r4EdIiXdjOoycJAVcnfRMhutQAp1hTERd3ZSdyUz8LD8yJrt65WQuP
zXfdZhz0TcmAU+MtI+VPiI1/+9fjkaiif8dgsUbMmARWxRnACX3xxMHxpfTGDcdB
xR2OZZcqjB2wdJizzTxcWvQlLfSllZGHjlH9f5hdhLtA0BevPLHjqKBN8tfiRQdo
k6t9CR7NGKvpISAQiey4FoG28+LYgU8rurDZQy1EwsbbByM7orUaAH9XrrNjlG7z
/o9QO/NDucWlz7B3cxG1W6T3m03NdYF7HMkDp6FGZKfsyk5WD2gT/0TzpzHDnySI
fYd1R7q7uPoUNSnE8ORAoqgXn6gVpObABrQmjl+9Qf1QcSt+Xd/Acjge47jxKsr7
datDe1RuMg99ujTdLsLAifOTg7MmPQj76MbNj6Y0Ip6/IqHPcfcV0RCK6sYX1Hm/
U2Zi1uDEyd1zQYDDzkssZNTV95BDCwByyiVIPTGnwMFzs7uS6T4tMtaMJ+B2j2Bs
XzHo1ivU9IuXgT8xYkidoC2VQL1+UNkhxCy0SOY52uwhzPAbzQTBcPCIzSO+//Ov
z5NdO1TWJFmw5ASP8iJzQZIlPQ30+ZSD9+Pp21KlXhfc4f/6UmAdkHC5G3wXN1Wa
NTkTPAiOft3mAxBkCQRP+QNafN+8jK6Up6APf2GAuivBcl8yGEe40pmri+4MJDyi
/mRNJpp7GKVKEVtTdvWwJX5zjVmkLaYqCCrdaMCz9QjgxwOeVMOt0wYLk8URPv4L
u0dM5kxzWQ4+bbcxbOira5Eo5ySetbNz9LlrLrz1q59JL5NJmUKOyeabcVB4mkjM
+bDU54LsBgIc/+YFE191RVjUtyBbVXUm1h6Ee3DFR+c5GfSjYLO/M2sOa37JtRAY
XZORYmM+wOP9UgTePiacawyusNFmCha0GHXAo1Dv8dulRgZtuxDnwzSLlbzTAYuP
+rMH3UBQVCTaXac6NWRHad15d3YiuNWjyxMkzoXcbbpd0L8H14OfygDWHYX/5xKg
LYqfU/GdKHH0c4h2RBIN+IzBWM1zf5w3JmXjb/OyYucC4nhFdp+rltIGKRHCPX6J
2twxoN4Sc30YyE93GjqTjguTXIphkCKJWb+U8WtL6AgUtc418jZsMu6p6wx5dsPv
33aQnXUv9JA5BalDSfo9m841dFnNi+XaHR0HW6oJblztHqQUoLzQ/bXWwmb8Lj7T
RIkiDOoPTF7aXFrcUNzsTQuJ9VPDV0gNq3XST1NODT4QrEsDC0hhZUuDjgjlxyAC
N52vYDPX0c9u3IAy6DVlMBrx+MolS8vuoIJuV+l/S0fxFJHzYEmdau0H8vZ1YFdw
zO6S95eIj8BO4Mu1WriWDq65IUf6CMtw/avVJcDkw2Ys+TZi4cNrt7x5j7SRHF4l
L0LKbpyCT5Fq6M28vDCh19uRd66X2spif3Vcfqc/1F5Mc51YOz3QroQhAaVLzrVu
N1bF093Sq2s52/ZfVeYJ1vKKz1btvYTsF4M6b8+L+9NmOZ+U1Zutal2X0gm/LHaN
adS3ZaqBtKf95/dGiferPktWoaWa/ULK91i5uRtb61S1AsEAVugVbR8PKtSrG9ul
gXNXZBud5xuIPkT7/RI1JX25gSiHEeb6xlxUMR5Gx+jFie5ovF7uRIqseEF4l1YN
JyGk9rL+Xg8Fm7MJtdDn1IgzNT892C+9BO1GOJl+7993j4PbOwPmh/bFCTeSB9AI
NAYrktyejSdaxH7shQA+iOth9Am0zfHErvMAbPG9HJlbW+skPbJFJHcMxpnQGWD/
vsCilSRHyr+uqa+TmLKOTofRjMBF66q0+im3oR5rHd/pYbJKKkyZAksiJfsKAx2K
2cGkMJVlHd6duavKbus/RgCindxSO4epyUnYpbWCJilMDxv/G/8Ienh/a4Waf/H3
asK7XXKjh4Ew/oijQWx1tXkCgSXHHr+n74Yc7A6Lhcit3pLyrgZXL+81UMyFVosd
O7Vqfjg8gwLK0U/9du5G8bvT2RL7HYn0dgOozCeON397PxhFXrrMzSGMfrcHweFG
mbKqJUJQab8Vqh7Nvf+aAynpxrTR/2QSapJ14xbsdSKjvLhQgwN/oV926ckFCDKL
U/6HNFmDbtm4/Hpa5Ab7lEKy9rF7omtPRUGZHfqCO7lR6Ha253FYZIOM6+jd5FMQ
PV29FHuhSlpt/vtvUb1LA8Hkx5V1+m/H6SCnoXTUloW3ogiUgrvDdelLDP/aX5l/
u2f3ZOhPPHRJkWuhFDlGg0jKMZuJswabbukXLqG0/Cz8HmqfCo5mAUMDKY3z+mdZ
ew9fQR42hNXnWjh+zUDbEGvteyofnrsb5di1BR7dGm13VkHLkTTnxEn+9M28m8ir
UcIOOUN6fJPcvNLcvgAsARH2eKDWgOSHJ7CdmmttdoUDuAgZdhDa//+9U0haYcGZ
A6bKJHJpdkHkyYZ0s8WL1wFhYWgbhqlWetD7Y6LrDRvMXkKPzedKojb5s8f7LW6c
Kmv36wM5o+mYYteePkB3iQA8Z4/9rf2/ayFozh15RQXyErDbo8QnHn60DG5jRDX+
KGl9F/iyUQTugwj/8ntYfjc11U4PSHxEKjzqjTQV2/d5qFTBHrogwvUPYHSvHWzi
LByyVS2oICmQfuwMUB+huXPdiipK490ZvTuNLtAOtyW0/0tHQ8H13yjVaYbP4nsF
LwRMm9fcS7sgwfHwR9Ik14dfChp8AhUsM1Xsvs1uAUqY8HZv6BEHiMC+Pjk1z+hH
7YFwXCfuOF0aLkRFsh8QkQUQ+oeIhw+tNFEib6og3OA3hW65F0rgR49IMG2Drfd7
ragmD3kr1T/KdDTYXRLnGuY+h0FrNo9GVaQKainyeGDLtffYcPHhY54XDMHJChLo
SKdY8WEELbv8WMVRCJczbxEtsBJ05gEIb7QN8cP8YhCo9fQ07KPKGCKg9k+TbwuH
WozbLZpI7HB1ry4Z+TE5ZYNOW6e84CoCq7KNH5X6w9rg8yD4RQ/79QHK7k65nY95
xLYQXIZoVAArKpPGXIcCCN+N5OkQZB5EBg92wIriVcsCtLk2YbJxVexiChmtqolT
xtX/ekv1NS1k2uWUJNII33SFrWLqARZNDip92GMdDyTn0HV//mGlvkSrJS9+C71N
n9DBMK9uKdy7yrCBrkf5tCEUCjZhqpxi+eIFILNmiIjKNP7KYlrAvHf4ULG65/5L
Bw3ksE5l1EvrC90WvvIbCfSl15anhbHK/rrIL26UbFiHKcht4zUox1/frFh6U3D2
pkUSp6i+/SYgkvdQDkj8BPIqBpn+eJIqnHXiUG1Y73CbtQudag5ww2mzOXywk/kO
O5fTYCDTdJ7pQWyzUx1L07EreGmGuNXf9hH4WlQqt4nBUuH2cBXYWgZOw75fBw4Z
A9X+ZVnh/hQZpHilBn1tXAh20J7zgbrQ2ZRF1qdmu3JgRsXSbrN9vG4enVKk67u8
TeLfItl+YBijGNuC/IZLU13MR7Ho9Ig2f+94Uj0DeAHRglndhKD2HdN1y7wvK7NS
LRZx/8GgEbplfe/vNwmVacfkgkPHmQ2Gzxybb/4sBhKs+nQ4b+u8qCa+/jBYdHmE
52Wgw7ZgKKc7YGqCq+JTDWvOyRHh77xP++7G1xtCRYQNp9T5Ph52NwcO5sn/srwd
rQvfDFL8/4A/tfYnpp1v0AAP/Wlmsi3dwn+S+JktG69a2B0EOnwPfid6Im2FKs+f
itxMbHQ7uYcKuMJc/ETyms8bagjQJFfzQBV1SvnzzZDY6mgvWimMIqOtMn/QMuDX
FwHrorq3/WH0kjSXE569GQoVCkOpjHAH+Js9j1pO7+amZAktV9Hg6SSDdF4eQgKv
f4s8W5LVBY9VUOvdpw1+Hz3zOPy82G2WIBe28U8xrhtgIXXa4Yd0u3VT0GJhLVot
iETVaDN8O1O7OpB85YTZBgpa+RzF/XSUHPK7zt4tiUbszZUfL7CP81CcD9DsDxXV
FOsA+UGCNCei1W7wcBSMcdDxfqy9jIkYewT5HqjoRtUvoExeb2f1dl8SUCQeXa4C
wXriN1Pd9VDVlr+RKgKemZ3QaBPD4cKxtSROdcR2YzBdmbUIWDK2npdky1LTgkwX
GrBGZ3E35BBVdWHQmOE7ybzf/IXrY+vFlLaxClF2o0Sg9+y3ZNNlwbo17N3yG4ds
zsfUJjjACFL/ToGas3kp55QRoA7swuyJe9+Jw0BemxWVWC353Lrz+ZRvjMiUTnne
W+Q9BmT3hKJX2D0JOo+xtG3wJL7ASO3z5nQEwfSI/QAzp7p7JCT3kCBTR7NcVkyp
eYAYo1jnuLPsjzeiuitKUwd7gpjlmvsHSEp1BK39/2iVfMPoSPpX0MrMzGUZAQ0p
t3Xxj00BvKkilT4cHKu9fd1MBN9LGBrCy9EV9AAuZCWlXmBruWokbWEhGCjej9M8
7bboN+jqBw+EBWalTRV06FCiRtQrG/7lR9Bf6O2hjPFiOBEG3AUsUPOgBxZbze0f
wNevSRaCSDVMAndtbcl7mIb0d//PCI4LtTIdbp7/1wfNECi0k198cnvp9rxShBxR
F0IahcpmgbHHO9As0k2gO/CGg4EvjJqTiPar8JJXf7FVYvZr8cYp+mHuv9X9pFDm
Hw6zMGWpygU0Xmyrh44708JI5Ya2To4bQugZNegCcWdixR4XiGuo8mrenVuFSlyU
/fqYcuGJQ2eSKbQ/eb798ZJ0o1QdBedgLGyzBwqa5Isvw6hkhIQsIILfU29nQi5r
+CWnVS1hpMD7pVz2xnY8KCGwun7iHoVB/ezqlyogtkz5Frw47CKZRQnDdJTEBbQR
HSzOPBEK2FDIeCxgeuvdJb4WygKWuXvSuMLuuvv3JCfSlcvtAaDzoYwQwxcbUu5M
8DRI8yRhmyWyM07bK1ZVF5RRsn8bb0a8U8zfnCYSQ/6/XvMt7RgzLt/sCE2+12C+
2oSbdtDWWSXfzjWGekmxubcolOtZSF07W8ZQhmdtfl89MADKerjcvavmNvhP3M6A
49QEiX5gAO8XNFfO9U4nYUP65exSV6j3x+4hM+XP99tHvwk1oL45sYs4RtBdSbXz
IBvTr7BdlUQF5TvXSRen+TT2za27KScWGV05QvPdOwawCZ/NUYV9dBp+VIha/vON
nNUDJsLCHSQGk6mZ0TL3jNauai0fPSnCJUIDR83P4HMOQc9d7TGA8SA1Ra8321tr
hMiGblgPngE+y8492+CgUKh3PDKkU3Pe3ktF3OWDC2OaFSle9dU36L47sQwd5R9m
GRtSWN+5X1wypre24f8aIxbyFTPHbCfYkYNuNhjR2lzwG5kUX9RS8nUSfZNmLGjl
z9ztbCx8KFfH7iukQRu5ZY0DhFGCjtizZEPyR+lJg6y1RusaogJpvHY4+CFqYFpq
rNvQnpAsk8+et0rV1Bkpsn/+1hiU2lADJWz+5ELoGqNUCOETH3Xh2QXXQg6kzA+p
s09CWj+zPscn7dARXoyJyWQZ9pbafnFzN+f/Sz4f8gEEt9IXu+EhvSqvNmJS/lXk
U5lxRuxVposSpaHHFQtD4HwSjoX9DAfc5Vv/2O0Lsff+RpmRxviY3CoS2YE3ctVi
jmRkIjb2tk8QhnEgJEVN9O4P4mnjfEJrUGuQ4OzLwNIG55Q6uXArIOb5F7pr5McQ
Ucq1EfwZoMpcZsie8FsPhCd/iyXSWOtLKcZEgqtrbI1baE+9n0IMi4ZwGxnCQbVk
Rfry4lkafAvi+ZhXPBGoUHWMEyLEwwSIllHmzaSTPqxGqRQZ/XUpP79lGdhigyOn
e8dwg0RtIPFRylug3z166YitKTmbdbC7wilay7Gect0EY4C+d2tfIplVoTzejF3R
IMRd1cZLFpiF4qC3eB9hMAp55p2UzYCUKqsX+HbV8oPH6mkpChQlYuruWgbrvuCi
ojS1TKEoZa8c6o+uLtft+olYLL4TOPN0L0KOPaQ+KCF2L/cxsT0W3SWLfjWV4+4U
mqmzzQ0PcduzhJBdnXZyLhGeZUkS6fexHeEfVGXj6ppGWMWPTGKuh6xtbSadkkv3
3PkFvBRWY7aJmJoBQCnPs5Zv/ePimKQd23Ns0PL7eGmDvvEvPnshOa58fukBy3bt
8i/EiCuZxdmX4e+j31fSjwTTzzpyhKw7xGfNvN16AiPLNLHDSKoZHpYIR79nMyDj
mQElSiZauO8sz7JrnRC+im6iQtumFIsXZQ0A/92dbso1FCZ4IhamFnED7CNHUk/Z
9jsQnJ8deBKG3gtvsUXUWCo8QjbbV2YNUH/bq3JCfJ5yPDrhiJn8NuJdDa4/Z9Ol
aPqX3ythsoiiJX1uKvAtEHEnEPfKNrlSw+ZEsywPW7ANdRZiApx6odEph3g/FJxl
MMadKSOapvfHywSf1nV9DCz9rlI1VOOuFsSttGb7ifYF/NsQb53a6vVeotwogxII
nRwtMBNJA5gbXVfUK28djZuzB5oZYyVGGh6m/AWoE+uqvMmzQ68q5oapHI8zfZGJ
7Aa7Qn8/4b07EGN0by0SbA1plv430yWcbDz7rKEEsL8cFX1WNI68OtC8bi4vn3eY
zRKD6Mi/ncg4EkzBV6ZUY3hXEzMhUC3vb3YC52wZ6tq+dqPE6kI/AsUR3ZZzODdT
632n9n2MGDSOdozx2W3qjeTWwi3WJHxBHmljzNh2/2UlUvIesB3d2CId9SFvD85N
6aarTHc4+bVR50DMR5lqsfmhaIqpfBXC+KOib0PKIb9f6NqEYAEZXvuk2YwcO+IS
tmDzovCuJQrZ8g/jEiMUrn4fg4ZF1eNg1Ezf24kzhyrAOMMCtGHaV/k/W/xA8edz
Sv4vLhgZc64WedehR/MbdtUaxBscgI9brqMNleur+ymgdrfqDxyioZ1u4D3F4XNE
yjDO+NFqVwmZReIaq7RKdoD00q1J03fl52r7gQzByQf6w33voycjVhLCJyMhZ/5M
PCqRzgrq0jCQyyn1M+NpVNRxoqJVRrIQocqZ5Qpo8W3r6Q2JGGjOkX8TMlftx/1z
i3emGkSSffV8E8K2vNOzicrklAte/AtWx8OY62lcrkgtcH6acyjtJ/r7oOce+Zro
ivGSior4NrNl+nL3SK+Snl9ow0s4KjFf/rBzVyD0ISEKLw9JbhrB7S1QrlvSAfQQ
pfW27E5iZVoBLKnj7IcKPcxTjPXTg2rssZE+TkvVLnwhhhol+XONI9S3DggnAEyo
Z+zK/JwC91L5X1aPLEImK9xv7jWjIcWg40mPJda9HpkOD9fXtAHdZ/BwybsYKrX/
mbtp7H7yk2YwclgBpcs9/zrBBnvW7jYRto9nVEoz3d6nbNj9eqzCLiAVMiBipOSV
f1nL5D/7uLBfGKfwEMIQ5c5dO6pJ4FuPjDXiv9YoSb0ndXXA9oUdvuQOLXHpwf+l
QM4OJy8BIiCpXeBLBhlE8Fp8sCFTaGcHJ8reDo9UGLaOPSxOd+L+RkmAHxaqBOOc
ZpqwpRlA09oeXKogm3VB3dmVDScJUMHcd14wSIav5AVp4PmfI/X1/ELd3FYbc/ls
LGNLoEtvTMe2HHErZ7+8tcPax+T9W3uaabxsF8Zb4f5/7mgXxTOL3vrVqqXRXxLQ
1X0S6iAiV9X5L6hXzGsSF2OSqUXzH8A3PHZaudJWtaoai9WdfceDahgUQKsvciXy
ZIZW3oCoJJG81dDJta8uGA3M/pTwhdDL+Ahn9c+ycA66vVkIb9NuABIGSiUK1zrY
tafcyc3MxohZ6yfxrNc90YnQqmmAZWarhQ2yy0mi6c+XrsNpiPSdrBtmBwemklPp
MRktPP4ZY+YyRdWf8ZEZPvDRNkUG/RGnJFunjqh5HFpAQww2UsbQkgaWZbjL/afQ
Ql/f1m5f1sr77YWmnUpRNtZzEkK4XNCOt1QDin6rqNVceLTKNcbUkaGLwXTHj8MH
z02H79GCXLR2u/ekEGvwMtUXJ7QyJL1VvqAcSvuckA5s2qKEmyBR6yuu9wSkcjvA
yikS4csuB8zVFdIiJGjI7YXQrDbPoJChXqT5ug3qnANLdvxer/9+Qr5smSvotr0X
tDjG3FmQJpm9E77rWig5r/551CUAavXge91yJ9Yh3mUHVaieT/SHViMZDmYwu7xO
7XVZCVTsQoQuOYEDEPq7lAtTyr29ypSCsaAxWIk35PQ732bo4zQCrSmcxOwhCdlY
i+qVHNC7x44yyC4fC0eUmi3BanqWbQxR8TKFyOQutT5d6MjDctGSHtABDpZkj6De
hqVdPz5sK1KH6y0XQ5/m5xCWNlGT2pEua7itdN9jm587PdoEuXDO9/a9quoj9tko
ZQhjH3TbS4tVl+IP3qVT9MyMp5cwgl30QDchaMsTQ6sL3wPw35z/GIj5FNWV0LTN
bbfTyCfSfd3pTfWt3Nc8HacvE47hIO3Y9Um34DOVo9MghGTTKaBbDBQVpxoTfcpL
7jMvrvCLc4DCyyQr7eRLNEy6IiNj4CdtH3Obb5fFJuvlTcyCVcFkM5BMVEajJbx7
uhKLCEl4Ac14dSt2Ad3R46smL+N8h0o5fJUm0eP4nr4WNwUfFPn/jcN6UGAxgcab
VBLwmPjgoFyJ6XG6lccEPCU3fIEdgmSommZhuI7o1mDneDSIFGFL1K/zFpa/vp+/
WWsuTgNXc2dy8tRzFbTMMtjCmxD3Mo6gV+jmgGNdy4KoV2oNKB69zDrHAc2PG9lh
s5x9tFQ6Rh4y+NZmLq7xvDxrnLsEuNepo9LOpyJtfyUPAOl5fzRuVeUzUbuQ/ebY
OwejF3/Mx+aPxi7DpJafXjKw0NcW5CGFpZMGrJ2ixmU+XkGVS2E9mhRGWa98loNX
w3mnRnxNprKUTTAFimt5RR9mjoKUQF8hOvxPzCvL6x8R2NH+sBxMI+GLduHUW1rY
51ROvLuyim9UH0zpB+fGAG/x5G9d6nMwVZ7KmuP6fmdiubKfSTHJELYFjF4gXMMN
jOeKLWNUfpTOdtFcUZ9AAP35a9Q7Y3I8lWUxIymCMJ0oAO0y+MvO02sabJJ9fvuo
aQNGs1vNfmXmLurjcdhQXeAdANeeXjGw5e1sPytuB8JVMnbbT4uA+ffUHsA5Ri/+
mkz0FY5kBDqkA5aouea/1vBXqsLVehcJxdcaX8jcy+ZrRz0cMIxqtxTUUQP/fqCg
5R/i651ha97CiqbxK1ITk93OBZAfyI6quHYrDxtYr9Btr1tniCQ/1XJxpKVRlWpr
8WYTP74u4kBlixiUOM+Ebz3LzATfSoZKau9RbuI0fNGrFk9EC2YBE0nugKS4Ople
NQyCg9MzBjI0/CL03FJqaFqnkMCwAf94TNG4P5zOk8MDFFO1Z9W9TwpqC1DjtZkV
8VfMRC0st1xygzMk4K9733cOHcfsxrOPuQKxExJbpLBtI00Wqh6z1dT/lDTEi4MH
5ZDctbjamfqVOeTFPSOo4xKnNSdKZR/KeLvLf9GwuW/UtHBRKX/0M+/oJm2DGb05
WlGgRz0ZBLU51vXjL6k/KY4ORtkKGArLkb+Blbh3Trrf504DzfyGj33wjgp/IW7m
q4mgUmIqVuaB3sKha6ZO/KcQZia4mlliUXsvetie2vhtAiSdtU4i1aMc5vAlDGFi
Y/+QOKtbkmtUsC1TxfPlyrQa+CpzjH7wNj7nQtUwyCzJo2wCZJ49EKjV8XClwFO8
+80wQrF8cAEBPxd0SwJbt/oBc89dt8FrYSnzCHcV/DsYfUtFQXg15j/SPyPiIqEA
V7eEsGuoaRLr9cbxMljt+Yjkh721FA59bAS/8V0R6BkY+uIRCHrx29HCfpbVhdPG
W9M0jwqTPFZAOIYQbacv5fFXcEmx4MLTwydtY3oR1Faw/rj4COLiRpUl+2++sKnI
7ElKMmyoiRaCd8gvwBIUfgVrrlX46USkjwTs7KRPdj2ZOM7BluRFHjENvI9hbgQN
GX6vkg590okYmGQS5vH9djAJOq4qiopqslvQWAb9l+xsLZlYOsEgW5aG+Klj7mlF
vF3r0UcKoR1hOboViFNOFM6U2MMTfw3hMKQyzO3LU819QtIJcARTIOPCGrOMlVWa
PY6cD+qSIJuAS8APJoYYO6bRMP7rfPLuVAW79eiPSIZaZCOJxy2qf7RG60mK7Bba
Si4CRdQZB6MORCvKSubUK+kpwGQnPsVZgKpRbMkU//+8bDhuGb6Xp4Qvg2EGUer5
ErU69cNd+rtNXiDWgTJwyVfVU+VDzAx9IviOBUwbsGbYSBwQAba7UxbfJEDYRUtX
SLEm8ts1GFMSCwJ79ZD2ZujVun1/2dvpfxnyDxlT4LdQvH9yPJLhjwh8/Dxf+Xx9
rv3PyvUHf5AI4eFEWRE7PC+FGIpjFwPJIIaUHHF8EB/aFdgS+xUcBaE0R4Mqrl7H
bayaGphJNpBn3Pdk4Zo27UBGfSRPtISZh+Bop4hDCF4v3YFNw0/XA5RlEi0IhQA4
w34OczCKKjMgywFkge0Jefu+ffaEG94ca97MHPAJnYAl0rIRo0XjqJ8/MKXy1s/e
IVL2sDS9qA4g/lpuDe93/F+jyhs0GXbIqOeDYyk0KpS4HKR/PqP0jcsyAA8qrwl7
nclqnwgOt0ONusFqWbKdpksgPmeTKFmxtC6LdZkPE8biHxN+pIcu7vctietallA/
+T6E1oyXiyCbGn+Pdpnt9iQ7DkuPPUDMKrBJiEqWI+3lF0UQsRdkOCNnuAF+AujB
qgNj6UT4hqgUT+NOO1oHydPjh14ZBteVSRQk8rSrUDy256cbPr5jMljgYKxhlqIM
9VpuPUt9PNDFNV/H6/tIDtOLMHcF6F0Dhl+O93nqAAyLuccj9MCngJGNZgboacRC
FFRp9ognJoZ2TdTIM8huix5Dzz1kpGFtpN4iQOkoRIQLFC6o3K2uhb537eLiB+xS
AGhNaXG51oFniEq1y5+1nja4P3ZncB5yiW96CSQaVALdEiJdkak6UUmSIG//qLSu
0yTmc1kHlGzdQWPjNTR7KxycKOIp5UKaSOlPKiAWe3frEFAwIvQfkbEbT08VEYOx
xhccNvigUCVy5iqVKS79ssY40h3vooJKVl5+YvtrRlwcL5rbAXhXKc75E/gV1uFN
0X/zkbFkjvzeApD/9YnVZB4We8e/+unW8OUWM+BB86Z28X8EUDSGs9kUBHf3l2fS
rG66zNfE7KE7sMrlNWqy5OU2gmZ3KIbgQXT7PZa4tWDObiLdMje2w3VRHwR+sbTh
fldk50s51xx6ZDQ+GmUYAfDRbh9Xl7/WiKsCWJZOS81+B827myxfeR5ZtTpA8r8v
QmI/jqM724spAK+7PX1xtCI/1Da52NdNjLsA5k55eISHzB8cUkwHYAylImQBfGM+
8dOqXNg+v7YjE7DRWif3QUBBA04eYc/fTElDIeuy0XKqjAYzMus1k7u1H0BAdpNS
3Xhpb6Ax68lr2JfcOceWagS8qcVLlplADkoJ/0DoVOW9lp7Z9FUY7ixjr8IaTAGj
LQTF8XmgHrFptVr5nnp1Y/rM07Pkqf8L5GDE+/VUVoWuDaSN0TfYWcGVYWt7Iuuv
eJrPZTQ704fGgMbF3o0luZ2Tvwg86/xNH+a7c3lHpwVHLplCVn0mM1Z+E6zqbH16
AZ4IMyA/SNdzETJ+Hd12Rq11VQNGtHv09+zWRx3jSpfJC1oo3HPynVLqkXTUjHz2
BTkGYxQ5+nGQnRXUCNPRk1UvKqkQ9LmC9hOE9RgISskUUG2rq//irjg04FDeHJbb
xNA0zGwOV5oodmIxk23QvId3LHHlaMHqEvnYoA+Vm+pMTo1LazfnKQF5zLsgNGYJ
q1/QgQw1Y/ZEAa/TifFDCGLFddJrko0Msj9ftdmdextwM2PB60PyJrKmpWUyqHX4
gIT26KN6lCdEM9J/kIDEmxqW0RqRckqXLa7kKo2ads47vlX5VQ03b4IYQFZMWRwB
pF1jA0SgEp8RaYjaOZUBp5R1MEkO0PDoapqr2195mz0XeCMLX9x3o4uvg3BMhShn
ltkslyG/JTMV7tUVx1Xx54Vv8ZcsoR6AjIxHjKipKrH9boxpePxFmht6FKH8G1hG
PSPxTsrPGNU7GSX3k5YDoBF/oNc+zX/AXjq7Y6ZQZ47EjDGi7qLkNfRsA4NK9VQ8
bLe0wOc3mIZXP9/aJj+x5AhxomVbqq7FN91/zy1J13tKkiRVjeAo65bNKESSQIg1
J2qkFZLqr/aF3q422XE8AoYjzAeP+GC9wqYP++vz8TYi02VN00rMJLu8ITaN4yy1
Wf/LrGdlwgz593ARUwKajzsIIEX572sIuFObtaKX5VpA/eCgWuM3HBr0PipHbTz4
74xSkvQiv+41Fo+4weX7xTjkDtsmbayWkYw3fXs6vTlLVAHr2UEm+X2SakDc1aek
ipZI7dH2gjQoh9SbuOT+BWjY3r707cmmB+/vEDXlfA0wA8CJsJy6sOOVNxmMb7QW
lVmNIu5dNn8Zq6xcY9N7nMz1xD+dhXys2sRl4C7beTFkjMhkOSo/UEGUTx5VCofy
O+/Np6er/ZKTrmsi7UVBlt05v63Dj3BzOfWqZCw7mU+1OY2bQf3zZhzp00MSlz4R
pYu1zlcSnsmMYGL3b0B1jWHtRD9FTf3VlZNV0QAtMa1DU/HCRFhgOIFYZE+SFZft
mFIfZ9KL/goN45B1u67QcZ8bCOHmuAXZs4zdppDXkK0/rE9cuLuK8KuOqwhsd/L4
R/nG7ydb/rWzPovEn1XIkUhnadecbqjqiOLumKkdQYZqKWRInYC+It5PmByu8MZY
diYKg9WWzc0ld++4qGj0vFX0nfW9ikwxybwFSv5L9WK7V4T1RQUb0KEWZmVaOUR6
d7mCutfaL5VJYLs+DMGOmsqErA6vEab2hENkBTu8kIBl/YdYbXoTpShHzuiLeORi
WJ8zsFM8dLVXl3+x34NyCSoJeODbE8pTV9HfRLpjcALoHu73qu+btrHBJlIDP41l
qFJo7uwDdCPr2OvVw402BRcOi9LeEvAMsq28jJIuS6QqdcvbSpDh0wqIoP9RizHV
FMBQ0Ohy2xZvuE71C9s/d1zs2hYI5z0Ess8B2Z99rrIvbFtB+pZcRUPOmhD3D7io
/UTPtE56e8nOG49JvRazAlFzTN4AB/xxgXidzygYNw1xu6Msgo9je63f9b7ttb+F
bbTN/YVG20j4eEmUVY5tk1GR3FHbiNBI3qzDtFVIUIuwUh5Ta93T6swidTl6NP/4
K31zoCp/D/x+6FIo6GzWOj/I/70xBa9HFodU5My1miQbq627PJsFPfoify+Y/Ax+
oEsHM9IxaJn8DuP1nnS0jTUqyAJr87v9eKZrJqjgiZ8Twt3ecpMR34SVWtfHjwvA
XG2zPkEyjxrljvJUI8oWHCBpKHvuHjTaJmSGiYiaLawiJeblh5gLcCqEMbR8Rs4e
iNiwINSb6NiX1mccEeCtIuwKWyo3LBNJZF1ZkMGSNzBh/9XpmiSGFC5Uv2fmderH
5RuUdJEU2G3gKLGyJRjy+DFw5eGqSOf8FoSQQR3pk74ndjwWm+8JRnYP1xCnltTz
vlcFDchmP3HuOictF3FBVd+CAO6mAuxg9hyXSyJ+anT69CZTCTGIpvgxb6n5C88y
2I3uJk7jyGNKFZ+cayrJWdkvKqnrACNG1R2MCFAUfuZRKOEQweHllAZas9jDw2r+
pigwODt1uarze7gybMm/RTVIXwItdu/1ErYPB5MgNkC0EQMKed4cRsOdGWd2zAVH
5WeSU19mE3tu4jxu+Eowhx1m706F+M44SIGj7SJGGtFFzBUC9N6aaWwUcMe/BbBQ
pz6J7XgpXNPUnaqEWC7VxZBh6z61uQM2CpgTxxnZOieB6zkWpwVX1rGZn26YzYm5
VXrrVLqlV6af2/iTfljBpaUYT4QDYjYN6REyTlxYHgSzpjj2PJfC2GhLI3hx7IJL
0qQrOWZWFfcEHcfvxAcq+4kY7HbEPDkxjvkpxi6gBSkIiYt90y8r0FzHtjtacZ6u
ZmubmClWSeZsw4AQ1vg8Sj6fgK4jTqhOJvkxB93CLcpFYW0Mh/obOux3EhrEPna3
0g328/rqd4qurp8NwU5NxuUDDd7RuiwTQb6jD27eG+I0WmEkERerQVp/7d86rxSo
DQ+1fdEq6S/VgKHjzPPdpimlSC5kieJpYCV8wPyOw3rxnmHbhEY5PpxdMAE72Cbk
vDj/JTX89qaj/E1+WI/lNf8WfE63z0JWxnQ58PJCt9ruszg8Inia2W+Y5xicSLUE
Tz/qDJJAan0OqwQjspCd02Xy/8CaLYQ2plVRReLKhrG7i7l8b5rtuNaWT+UNaOMj
HPeJc9/A4FYYX3tG/rZN7Z8G/yqaIFM2FbG5w1MLwX3pc6eJ2b1fFhWa08k1kzkH
SbnK/V4HjGbfgmvjX7hgnqeA+cKJMqsxSs2vr/IUOydp7xGsxU0q0LJZuWi4hAOB
a+DpHzyOvyZOn/srg2HjCMVXdTQRgjNQO+olZAk2SuPsdoHuKjjK1RtCEPD7zhDA
MOpFgSY50DzIPZHfLKr95brqpidCGsd8AUuQebNGcommEae5LK5hg5uA6U7qC1tt
83BocNuJVY6hGClVjD44CXFLMKw6gIknW4Ie4ObDSoLOG00IKCXgRyl74w2f0roU
joApXrrEpAtQSCMmEe8VDdephx1MlvJhLOCWjOPKRmKVpWoiHvMCL4GcI95UL1tM
/PpcNpd7BCvfgIK49hLP7ymhNuy9aFs+Xi6pTNb/o4JwWfBE+OvFeByHCw0EzHRX
xKD5asdVTGBVwDRtjYpa5hd8pVpdRn9OQAVc2v8OLV1itOx/9/zZXO0EQb4qU10J
Lld8qzc40mSnBaUhZ5t2LYiJkBYVUIKRIQS6hcEcxxMCm+9qW6qgnV+TjQC+IJ/R
WMJwPEbuLwkF81/JxXleCgJnhtolslezhjrY++/WG3+LTLbW9uVyjh4/9+4fh5Tn
WrGN1Jd1Jpa0ucnCA/DHfqn+IiwNY5bad34HGQLF3NPP28Jj6uw60LKkX7Szg9yk
jkH/ADLG5gWmuXCrB/WC/e8mRibUuEvyk/7ogwwM3LR6RVk1eNwRC8eU4FMBTzpL
XePghi4GEnRIAwPGnO2JxkHNyAwdXD8WsNOdFGvZXxq25ZBbkd3xdthlPfrV7tS6
g5zPt963Gdc62kOalhCPlIefC/TvgfXwIqs9BmYo3sTsIhIm8LMtYi3V3aGfSVcW
eKehd0NTTt5l44u9tyj2ahQp120qAesWy/xiDfWiedLe5LMrsSjLIquyjvjrRD8d
z5NIZqc2c6hKK0R2r+8GSnh7f9WMM1Oe27AemDHgj0PnUYUVpvq2Xb/if7qZTzVD
cuU1BIzTErV442SV/IyizVLb2YWhYg/tGvutoVn2KQoyPW6UOwOkY3xfqs16vaJK
KW9t2e/K0bRUu91yhjKxt/QOzHiym7dJek/2DZJ5SLWT56iyfnuXGsIY6r/0HJ8p
GrQzoZllM3XJtq9LlOGAtSpEMh8p5z8vEq0XIfCaTeAj8iDznOuurFrObbAz4AUV
YLAeAlC9kh8JK2W++ZcKpxwUTmJfMxZG988lKqTxUZwcn1Bij8XCCaFwe5hormn9
2++FTCqu95W3TcDNNu/oILlyhf+6tvjOgk3+inQf+nT0fQuY7Rx5cSAB8RQ2T5so
vLsKLztaRwskONs94zb5P03yfGZiL+vUkf0ItdNGSL7DEJcvfUe55pzUPpucauUC
jGVivFrhFoxdEvS/33dA7FRTWgE+B8A6rueNbSfVfRvfzcLPSDpwwV5EX5kzYbiV
p9KDpkI7GDVr3GryBIyMjoamk1TOEuTwFl/seUR9/JdSwz1eWggUSJjmLxIVU0AX
QXFyKCbskPbMpX4bqoQMKZAuYE+nLTrMYjlFTAyfTNXGXbbxLjkpuLFU+ItbFqXK
JuUbI/jZtRLOluJqamE3Fra4rOP9xsOWTFBAJ+XTJPeqiXd7P3NEhQjGKltE0TGV
6vAtnut1tz0pTM6CIXGYYBUgtMyTEX56jkBPnKs0Y7OZw1bWkliryr5Zlt+mCe8E
iauUpJ9uAwAIO2Ycwkc0tgK3AV4JeOt3VsDH3covown/aAr4v06H7xYOsT3mfoC4
wO7AjBlq9ZRpROIb8fKYCgiOFFBsxMtI82y24dkRag3R3v+RBmY1PrUVlt1QnmjH
zccU42DVx9TVYibUvbxHuWESNDNNOGLrksqyqZVoCcVCd3LMYCnhcYAXaDzuuK9d
Kji/Mxk5kEasjbLMLyEqgOExhHXjDDVw3YUNgs4urdwU9UvZy8XcFTLjAL3WX1Vx
EBy2FN/O/c9PwuH3oGFz9wCmnAmJK9bdByFGZLrSjP/aGRnEEZkAjXGCcvtlJ4RC
KIzkikkOeBI4cuHeMHFX/g9WdLdjVRENsN0CrCBc8+chuvfkxaDOu5ZGFYVLem8u
nibxylQBscMhSGq7rQ9ZaaJQDQNhAcGja6+XQeo6WnywUWigVbdmnApZSP4CPmd6
pIyOvCJN3K7UuX41pOC1Vh9CRXOBOV5gnFN+867XQWJ3BlPkhWxKPj9T5fW9qWI4
kAYlEveizHp15ENI6pP1PHz2Fx8xOSHxpD3ZifT34vNNk5LBYh8i+KxcT538Owui
vk5y8XE+8FGrVIsgTXeBRxnPBEdRyRS7hzyx/YUbv2hLmoHOQw5yCk1PLFa9mrEn
46AZAiGJzPeeE48TNCoTULmmV9MZ5fUftIHVXhrHZn6YcHN48nDks1nJyrZxiXWI
aUFEfetzykS/2wEulr37nNnW+Yu3mOscXPW9TyF9dUuPSg24EuWhs6InW6zq1jsT
xzkmdOeTe9lvLUO1CZkIRJVKXTEm2nvg35bVLEWnfZkbVof2co3UqLuw+xQID2fS
0l7ARd5yrHc8olW2DPvzSPOwjHmbWK2/Rud4SQ5FAwgmjlmNOTwhyVoZ17qcgLud
290okHFbN/DZsFU7wb4J7AW4CqlML79lIkLmta+ETMo69WZS+EFVJaBkebkE3lD7
a0e4AusPxpFYmmrHre4bg/42c5zbNKpYIWA33DYVfKnQbUzMQeg+JlExKayogbyx
yGPC/hWmGckFQPq2jaPQq3UQUPCJPbnDxz2gZ1N2sjWmCxBhmt+EUZBQPGDHUrLk
mpD+vuNqQfMXZ1dfQeUOgZsXLpoIFlNuS7eG97zVLY0BR8SOlqgnnj9mPa17MrK+
hhbfLejmFmQshuma55LgCd3yIUKvxSYb7x0Fk8A2spyoZc9HpzGgGUVYyHfdUWnF
tilgYEZ+E70xO7TIoc/3XLCUaUlXpRpid2o1kvvrPqLIKNc+mTZRw/nHcM2T6roy
nVhaIlV8vD7Qw2h+oPJeO8DPlZgyDTd63m1XH3MflbGYaYKw4VXmfGQcYXtoI36/
bt09qELSJzFuh8/wM36voKkmNPCgQaZ9ecMPor8cdF9DutfRerrXKsSpaA7q2PcR
LskxMJYy2kRWg9KKJj0qWQre7392rlXQdgUJJ3e1Tdklr62bDPM42Rb2PifC2o+1
x9bQRUyz9ONu6v7thbH0XFNUNElH0z2EeTcEzR1eV5cxHFU8V4oToqDGGmCFAEAR
Zc1GkNZi5z8b2CoeWgopcKP7mmP/BjNsGGCQ/RkZE+XIKzbb1N0uPIcEIz8SsMpm
ilNCeq7VGTc0IrySUcfUsN90JC+cpgIYsK5GCXgnaCaVY+FXNCwzkFrr9CXl8HXO
wnZVWyx6P87fRd80e8l/F6PFmFCw6KayVNF7hptrVzYXi7PX/NNUQ/ZheibucqKS
9Gwc0tZQzc8FlwoxgJcA4j7b6oLmxOJ8eGtFrD6aekQ1m8FRKX6c9gWL7HuzVzHX
BOwhGAflzspQSl/HOImMdktVOxfl46QLXEyhYCZHIe9kuWMum4wuf2OX6LdcHTsG
/VCDNxCBNKQAJVUaRbDFXipBjAJh9HCl18liXbrbepUUla+gDAXTJWp9bNvZnGoF
c26uBnsHqxb5r/ZFL0XROD6sFeyzOAL6WDV5qS/ddbelx3mYjJuwk4qQQHFlXHG8
xubveUsaASWr+lPD46HNzg3/8K4QmR/qIttJSnfpU4Fg0pKFjnY2685Xwd44VRXd
AJyxU+QPie6CwWuq9vfCYj78mLgHTvdPRLz/JUJ/qTMVOWqr2FqzYtIZaSuzhrpZ
/vuOsINApu7Ld/IBS/xvk3+Oyc7CS/iomX/1XnU+IfmW+/bm4RapKzL9FyLCOtT6
wLLbaXv3cemJieBehUsv9nYIYdpD+iVkG6dy5Pp8PQ9XIa9azEmg+aIdS4KbenwY
TNgpPa8wZ54o6+BETl4zQHSi+Y8qcWbsvlmRksxZ4TIKu4PxcR6zedDGtTKAGqGl
e9WQPYiHHbxfUflvkzNqegyiu6tmy6UPBoSml/9j7F5GmgfSiyyOIzQCChpRL/iP
GOg5nYN6/ew7KhqfCBVA+0r+5QSVCJ8cSmEA7TwCkEv+kKbeiU5nbs3JTivxP5tO
gmgS4hnjyI/h4pMC23Pt42+ttKwju142izEiTpK7XItbFicdIjDYNcFpPbBP9297
FB8cH+qKgswBO7DC5jrO+TDV5G9PVGstCdIxs4lotYdBIUpfZYh+o3+FhFMimPWG
oBhZ47emBlC/TEy4Ef74UEphWOCn+To93XeoI9nkRoisAPiB0XIBzvl2qILLryrr
Tw7eCVrMKF9Zcx2qBp1ENLunDWAcBjjmAJbzl2Lj3p9oFZegTjMG2kT0P2Jb/uHv
s6rPBdrwKRJ1YlYVhvE3SIOWxKe7htgRnBTCf7Wk3i7/pgoHkwbHs1h1jjfK5rg/
HkrvRUAjbGw7y3c0nttH2OT3xV+BRwm6HPtIq2O1l9XUBfQfLteqCNQX+Ar4OH6N
kEvXfAmsMwLchtWKrfKFjOKgH8LO0C3RBDh2zwhiW4iAHcVroBD8fVh9+UyMk6WX
YjWlOJLrRcik4sg3lIMj2N09CQ+iQBE11ziFLHAAjoqfUcVFpARwP7F6D0//1I+p
RVqT3VaOjLNDVxRNdj/G0grmsVy5V2mAnW5k1OHDzTv+Jt12ac/r8MALhadQCGSm
Yo/iMEZHSD4nSeesSoM0kowkT5SFBLL8Uk6RFpXSME3yE/PsreetO8JNYh69XPDl
dahDy9bmBLFfvM3AWk2XZYwm8pfwaCeEkclkKUGJaCJju2l7Rk4RTWBqmdVaN3Hu
CMbjVu2VDMvxzoWU4yH2jegI+6Ouw6E7ySYcPnvqQwd598CefPVxRwAQSMmx2DUV
xcdOG2IcwRHZGmuNeQrliCs6P5IIXR1sTSHFHjpGoNlc9XkXiU7IvG4kYOtJkmn8
YEuufhIoFt5VT4iyg5wegVlHeuob/elISe6Z2Gwqz1c0sKIcOscBAgndSd8PD+H0
j8BCpVXb67SNpHc0NmVSyKDe16emaNDSVRJw1AfsbQO3ToODcYFfTwN/n+NZWL+f
mb+iKNw/ckx03SU6MgQTxtlISxZYXXKopGzKAgDAH1KnLQqlMA1g6JQm6MVcdN8D
FP3cKGMK4kCfcwhzxObxBzYlKH2AGLDqWT07McXvcNeiV7IiBKk/xtNYdW9ITW9b
hBv3cXXPU3znbrNlBs90df7hPKLf8Zq+Na8jpegzqW556AAfWZIJSSUKUe7t2990
nfHKHqMmLEJ22phy95NEI2ep4U5gH3QcltM5nMS72YIj2i1qEI09cebquFjhHY+G
FDeKwjz5xbFfUtdy5PSNgySb6hhyGF4kciKQ6yqD5vxZI+mfiVKxcc3iMe5Z+vED
D2BiKD8Um/qKWWecTSJAj3kN+dA6VdyHIICEmYQayiVAuponKgpGRQzz9FPzJptO
L0SIAYxJXeEcgJVMSx8Dd1/eWEXPFBbKcQENIqTDF1dyenzMifRdQrZYjRnRPfWM
QrQJQ+TUNF5Jqi5VT4Y81/TC78GoVMJ5F19XnQi88m/cnxOvZtC0AbIpW5nmVt2g
V4c6/Df4APUvpEcLWlmhDEjlT3YTciVOp055n3npNT7mtD88oPU6Xt7PPZ4z3DGx
YgMFwI5jy8Vsy2aDLzH5BqKr6yO37Zi6+1RvFazc28j8v5m0AgtR2fO+fMOC2c/7
ZGyRj6/ncUxm0lktnQbaWQlzSk24VbR503cB6d+InragCZIcp1kOWMM4ai8F7gr7
7xxdEc3RbE6Lydlb/K3CdQy4FjsJ7ad/ZPsnGSudSQZDrUUnCKMlXFKAD7mximZA
KcGcb7zDYaEK6ljDFG8iC4Lxffi1wlgN+DLaZZxN16Rkc2WjNYexp5I3680gpJTd
tx39EWLuJy0km1tu5FirhB+6bIGgay6PFzTMaCnn6jYT1JMj8JNlkcNn04rrLp0u
A3TcHt4nwGsmCti5grGxV0n/oPruotCFZPINqoekW3gEOMQ2R79octaUkxtFNHCT
xH+aWXT+jxZFtxRy5Yu7uUB+3e27wqz0wid0W1E2Jb6tAG+9JQfLXv0O6asIgG9o
dbPnVaaMqRdEe6J6Jl0gC1CzBkucABImwCUmmMhC0jPZV511WzwlLzYcMRGUdaQU
RBt07YzRVEU7C+rQUxNGycnfXzHder1kDpwFSEn6YUbzIsV6dO/lD9k8y9mXfF9N
3YWhlxRt9Bq3bT7JU21rNeVC6QcnE8wfkNFpNug/Opie4F1UiH/7PrOVfWvi0jk7
DuhUvnw1YWZn410g9K6/8NqY9ZvaImMZEJD0oeGgWq1+D+F8LXgXYsZrkJKmNAeJ
9MPV1BDQQITNEHxjGX9P6ZTZHyiNQaFevSNVBh92mPkt5WHCJKjLEdqUmWeKg19K
vin3eEzlEb9IKCuUL/nAcS/gAH/cKiGmpNtpLcYm0nkJpb9dDdm/lIJwAPGb6cPN
BVZnjve1J9jdFMFdPU76S+q0eU03no4+M+cvuzaDvNnp/ujLoD2J3Ov71y1iY5vb
rk3THa05l9UdiRFE19Q4Hfro0G6U1FeS3UaXFaSgb9J8obknl9zIvqW5tdLfzAGx
S2eAiJgFDhoGKMUQWe6WB/EsdUvsailTcolDTWOVeWePdM3TvEWqMb0Wl7tfZ62j
NiBrF9XcleO3saiVpiADMjqBBLcc0PiHuiDK8bYvlfA15zqwShGQGZ9bbIldRyY8
p2Z48DF+5x/8auuuUKRudDaYPzPlLtJQv6aVLyCVHeqi55fwY6mOQ928Zh0k6zlV
YPybbq2IwhQzZBt0JiNVmxfArsQOIkSJOmnmt8r3MXOJsCUnPt5Lyc3xn933QYwA
YqXTQ6hBavRCy8cgHdi1syk5lD2Abzu4aDv5uMIqt8Nq/p4SX91H/WSL7pOw/5je
Lkfb74ku9rLoLTxZT+Pl/bTzIyjilxDP8a8aenn9pK0urmYj+tLwoBjQ2qG31YQ7
4VMzEPihvEhTez3AAadFq2OXWRgSN5wUEvidEt6dxCG/ymJRRXPvdNzuC7oVCUYG
DfDg0E0RjWXPI8uo9B1hUI8Ni6w1G57jyRmfYR6VgvF1TSHkw6w+g3JgllwwQJiO
3X9csNuwmdALhvykM2ph7AWQLzG5GMSXXlVfi9QJ/XB3/VN1HGbfcu9MXyC1Tm/K
lDntntyTs0dTJ0+Rz5GXnoVb8dRWOur8xqYInmzmKwfXhPg2KisAKR+FzIeL2Xuj
mzL1iIpG/m89Cih6GSkf/ogh6i3s/dV2WrfEqH8mv71Q6qziyUtSxlGE8LKY9y9k
X76fPsaDBsi11ALTuyvAscSG0aW1TUXDpzyhre7+F6YXjZbKqwz64caDbG5fRkGa
FPkpbQAizlG45IlaC9wvm9TnCJCnyU123eOD0Z0YpU4+1/65SA57jtqRyZm0zoIR
z3KJji/pDKA96drOsgfBWBQ0pxyroW6hPqIDdWS1xmutBXqxQUC4r+mb8JeKJTZ1
8V1yVFQJEhLDK7dbjgimrPx6cX7L4NywatSS1Aci57rpZju7Tg1QbHjrAFitYhxP
8ZAlybIkl8qlVfgrC3xLtiZBDrEtN7TncXwpzkfbCRvY14AsRiKV8/Jp3obVgMw+
cGrh91mGjJ3Z1o/rUjBWEXH/cZSdbgP5mNQ6sDhZ5HQ2JpJ5+QbSdi6rAxya7HN9
nIPFLdQBA81TNgl82LYb1hLAieUyyd1tz1cWx0KUvmuliKvV1w2hAKLKyvESz2n6
dDHCMxYhA/DY98k31PABzzSUmDASYkGYfX7recumzeIDBTgM8zCe6Q6Kjpl7r/Hi
f3nxBzeoF9bcHnTWq5Fu6qw7SCLWkWyKasD/+mOM+d+jA7xtgKnAFIHNqcZhtBpE
7QM7uI4Pf6dECTkqFiAEP03o7QgPVcAP4Es85+f1lZyfPuiReGlx1n44PnBFoDz8
CDQqsatVAy3uIAOf8n3uuoa33vjTYEflF0VRCcFLwZRgTdggIJlUd6FuSLcZRhjI
xlzSPq6GDt81UFAlcDao7qo1oQ/vkQDErcgoSLff8eCdXlRDoE7L89MM/zVc8Rcq
UIyMt97ufnOQNwcwZUIFupnE4JPuUkawuMQ/8iql+pdpZcUQHPrpSb/3XNQwk85Q
QKmilzA7V9iYInLS+bZUe5LIykZW9poeKLUli20+xsNerrR1W/RLzd/O/nmXXdPG
1/l+NcRG5kxG8Q092mrwX+ECcDn/6NH7efX5b6UFFcQ+n1VnDw6t0nV8eQdK0ow7
9YA1a2/TFJvrGZxtmPA7OtfX+2q1OQcTJC03chdu3e5DEVzYpe1D9f42taarpfdw
NFWIstjE0i2kUNiV3oWNWRanHeuYqTiecjI77MkPe85iF4jz7tnyaEhsoSVRHEeE
12/fT14mz0TczRYbRn58x7Ac6HcLT9QJueBqMebZv9pJ/cThwU1DXSmYa2+kod+/
WJfF7aP+ZQ8b/e4hwPhoSQRbhL/UJASYBfmvVnSySfylsyoFcA4BICntHSbGBZTl
bjuVMudb51dNeqF+cNshoqL3Eys9QVKTptLGmjbPwYg1Y3btxxCdgethVRZF4QOG
7cVG7Uj7RzR4tKjRnx/FR0yn7PZyYtFpsYogIx90UNu0qZOt0ZPlNw530Y4d3sW/
Hk+KH561M0HR6cdp2mW1Xm/vU9lMWRQARnZp8T8+h/QRG+FOZY2/2D6zg1c7+td5
qnc9ytsdPSJiclpMo4D7T/zfsRenJf0L8cmgMIdVn2lmDh8zwGp3/SgzmM3tWtUZ
kgqW/xQ9E5qAZyoDfv43vXN6fqvZV8amjfGk4pNJEq1/dozDbGjhnKDG5uF1VyDm
jSY64fAuTXm9+g7rVyjP4CE1FImqJc6AqS1+r08xe/u752uYMZKx+rxSpw4RTFSN
+Qgw8ZJIYqJVoJ0chnSrXKfktOEpJmrLLhDEksT3cyu5ynk3HpUDkPcR6BXqB1xw
5qAcw7Chy2GohklTAEmC6QvaLgME1b135CEqYiaG49khc66N0iKTZiCkp36sY9No
YU76npINytMDFfiSXzuXb3mDWxi2lMt2cFZdhbkrw7j/R2UZgPE1EnXCRQi2ueLu
dBEMC3V9hn0VrwLpiZow6r7DCH1/TxoI4JjwsFPPiw5Nftqf7HvbdI8IBfddZLS8
NkJIMgToHIlQdEPZtHXCaGV7GcIo6EQNXMK3fWdR30lWciBS5Ao3zzvAppjT8b7e
S+senlmn7/lnGOTLFtYophypCdkgDuR1Shicdtf5VLhqrIWhQbi0Hj2PO03P+eRL
2uv3vSGqyyyGHO6zrPV3ZIr1u912gKmqe/qNDpLl6zt8DJK/uAR8MxIi2hDPKmQU
THchDTv8pLOTau03AMThZcgtuEI+GgJxHXgj8RvanqAg5awZDVDge98V0lOMgXAq
m4EiabRtRyCdfA3ybTGCKVsoJpCGGP0dj0Ac8HpqzfO4gYyhGcxTMYJtyHnfq9Zi
OzODhqZ4zhtMT1IwNjOQ0dPuA0IVL9+PGpxGlUPxDWXTxTQGQ/uCqzbPHYXM+S1A
STb4d/4Jq4+i2bmo5yegrJTDPoegkFmT2NjsBu2jtWVMGu8ez/0UuosRJGnL8Pq4
vkhNRJfCLkHvMeKuSQ4fc4sx/oPvCAJzcxBIxE0szGKWy2J83cG8qICsstv3mDu1
fNyvuBowDcqK1/ja0wEn2NUXViwat3SuJqih4W2nbMpgMmXsN3qHB8TW9e5UKZOA
SeDnCOfnp+2CUsgJIaZdUqqsjnGBjV9+y0NzoRciJWj3SyoLLDL/WJp8XI3yR0zn
KGyn2lGbE94njW5doWVnBk9AV7gB61DlaW0fUukkAUc3Jc29i3Fp19ENu1AvuGdP
PReK62enZUZyrv+PXd0N3NafN+xrq3kON2tg+9p28966iF8ewcN3UXkaHEq+Neuh
C1wIRghrvNEV7M463jG96agKUKAu8tqd8MmJyCGYIbEL64f7/WDJnSR32dIEpXJS
1McYlROa+xEZv/uhkmbuTiFYZ1cTA9of6fomnFHW7S3Gat15gVs6kRsUG4Y/I0Y+
nxV6ZmNhm6jtwFSSPPoyPtYyocu4mdQ/CVH4JkaXgew2tv7sAjiPESqERqMa8tkp
l6cFivYJ1cw5hqz2wsV+K9snn8tLtVzk5Z6oueP6RGzm/86SPVANfliQOYyb9D8O
pIOahpDZcZZzLrg6R2nS0tSmKWnzTJWF6P8hkYb6kzT4sQYDR4KNl12EhxXEtczB
XWPTG+k+xqaKiENKMgJsz2cZlcPrfsPEZing2cJNdpp7QytiqlXdlT9Gd3B58AtI
Apn7+HDhTQyUxM+5PCrHfQBy0Cfh17FRJphvvw5psNL/kgqrYuunSFboTpIpjIvQ
+RdxMb6kupsXNwHRcIsydapk0m0y4+D7vZd/WTvXXMIKzm4BfQEPbZBor97xk5ku
3E/3h8rRHoeGSN9SCj2ih+w++5ms6rzwvVA/SCvhU4223iggVexgzTV962B7e6CG
ZWKZHQ7SR5KFkudjS/f644pSkIS8jfYzja/SAptagPQRZoAvd3YatIdg2LHDA+Uk
rNmSr6MW6SIATNrSmHxnIlv3Z1gqjROpNhntjSe28NTFGYO9klvfm+nWBNUl25zO
ajU4nkJ+RBkcWcHVV9tY0gKOrFWIl18RjmHIOoc6P7URAUtBZoYsVCbs+V5gKRnx
2oihHozKdZ/u5nl2gQgxb+LEQb1V+BM7S0q6I8WApdVEVAy9TdCRY2xi97V0LcC9
6WbDx29WVpUJ6UUGIwIdrnhkUFe4M/RHq2uiJRiMJyFvQZ/aGxWNdUjrLYcIy7jz
A+5xY9kt6fYrL08ClGrheZPjYX93Xjf01wO8JnEjztL6m5RA+ZFra5QOKSUZiNEF
qWgNvGpd7y8TCudNyBHw5IMo+hrEow6WzxKZ+5bNSNCpUARfRl2GvyS2bb/IdCfk
LGhofZHP/GXbhxAdjfpRGngnu31d11/1P1mK0hqNx6YBEAJL20iwXe3UeSH3o92n
JtFNouCvpqtmPV3r4U6DFn/D6azjGEgJwgzkbrC9oKF4YcdaXKqHF66NIGzAQ+ap
NunqHz5BGf0MLo0BZMwffe+u7Qlkwhp3EsTtacrKckrgTuL4OyA01ubdcnZLDKdO
p5QehywVLtFWXHN/RoVc66UZDINEgnLPMBPNhEHFDSLfvTezfcdwWGrxPLwM0ovY
I1rG/dqWcuSHm85gGEuRkyTbsCt0b+gC4vCA3+ZTqXPd23AwROrHjiiOzCA45/Ux
vcj/X2dx3ugvtx4rSBZgMBZ7px7rF+1sYOpHd5BzDAY71eHIZOUXgYKq0kYzgS1O
ofNSlmnG+83UmZc18LZhJRMo+xosFwK8pRY6ZfVCmTuXeM9ilq9sqLmT4szu2lBr
o9H4tW+qemvkdL5CYo2JoLqIlPshABlFkzkcdzKOnKPDZ3t11/9/f480sMciOIaf
IyQUio25yU/PlCuoOd+fW8TOxlIQ+E1usKC86kh2eOW1mTsLa0kDIhs2qLp7xBao
ELABKo2ruVIqoQ8+EnbKfGhX7ZBrro2usPOChy8k/RDnscWzwX2n+uRlk2FP4LMO
5vKt/CuNJvAidyy91E3gP92ESY8YRWkPdcobgHg48iPvneFiqDlZWjXd3PAZZ4Ij
wgmoFZejK+GOlZmGz6Jdpvk2WQ/B3a0xHU58UpjaAj3lOu049wHGBwdjU7fTFDEF
ppEVYD2bHgpX+5P41DuHSS3Tyg5YguKSPgXO6aKlE0IbaMTI5ZAp2lyoBqIXOHkA
lNzMPUqEOsgpk+lUkJFS6Nm3A72WLmSFTm2GHBPObIao1Lm1gOsixnSxqEayYbSy
aNifuldXYxdWVmrII52C1s76lXBPPtIaRQ+RDC29bYh4MbUpFeG34jSaaBUJQ43e
JsQmw31rDLhiPR5G36qUu6nXxATThcKreJBjUpzhMu/YqmZRbJvY0kZu+vjV4tDu
gNPfrw0Dm5+RSZpg6MDia6m9MJFgNys/7MO+oAcOB76xidlv5CryDYwfe6G2e99z
fICGOEUyby61AGiE3cSqRPUy6+AHaMEYtvQRpdxfuC3og07S6w+eIhbO43l/Mx39
eBwcY0HIpyTMB2TqfTDEe3gwPDmZ2rNptZmf4p2XYMrcGY9G1BH372FDrk3Qx6KG
Lc1UmlhLWHCce6+ihVUoSsgvr3QqYYaE0sJiliPTsqlvKahTe9xh9zeNfDdoYQTy
V953MFA4xhZ9sxjHjtOriY5JO7gCqdvY1X6Uv5u/La7wqjzCd7/mgXqClYhv1omi
LPCHTrAvR5+1s9po/xmIIeMHtUpd3mmRlTbapGJP4u2L1DW9b6FWyK8xNXbd2kmT
IOWx8prET7aztVBBLAUNPl4YFO4YiYiR6KyCFhJvl1k6QcD/Lv3KcNrQV4VosmwN
kZVAwNaZS/oxtfTWdY/dJhyW+KBJJQ66UxGmK3EQOYTxDv+84jJmPI/pH1Dmt2As
4kso9ubbhJR0IkGoILxZcEchMhCbviaNdWAqRycK1dut78n7W71yvQzh8hZQTFtu
5aUf4J+1AZrhyRTLeTUYVQw/khWZChKh9pOSxOVUMiC10km6dqnOaI6kTk6bYgyo
03Uof9xETm4YLJuU/rKmd6JMop9OQkGrQjZlWyW1ELgSIL70Ydm3Y5t/m5kPKyWp
UreU0bk2oO7cRZISaH1W3J3wOn311ub7oau39/cnw8Uk2G7yEC3v5Jb3Cg4FiTLh
ln5AHA/ZeoBr1cHx5+F36jmqhiVNyYm8S+rMZ3F5rlD+Qvb2iAmjg5NyoDg3NbrY
sUFnQu6KtMVOdnSoJoT0N7wvhQ2gagxm+6TpcmTQ4WFxhxs0IHNRuU2E5p1Y9j4W
3dbwkP8VkAS5YFo6ICw88QL3QSvcVtzoc1qMScyXJOr8dp/hzSJPyno2+Lx9GVZz
k4wnfP9iPmdIwySvC/bMD1dDF4IYbxCnJwqoHe7ggCNRhrNkmPJTkbqct0kB2I8U
7vhPT3P+ELPwrgaXiCC7kfrmtGkXLbp4bL+IwuF2JEpPao3ZLJFQudYhpTMPm4Ad
XoyHYyWqVG/hqOuu6mXqgOb5+ibinGzD0nejRRzlPUcqXvA5MCkNEZLKzWDv8rP2
N70QNcdlF0fP7Cp7RqAqpTEpWmjo8wxKYpUJOnrOT9K1LCvxRdIjx8OLXbfGvdCZ
Z7cgDyzsW280NflMKWDULkunmUswEGVdxutC6E2C855RNFvslGYytZCV4HVBw03h
Nfdp5+qAihQVm3yLwsQUZ0moPhX0gnuomfJPuTjkjI8bHvm3lOKDGPyOJ1t42s9l
BK9fJlVTOoOw+QRCU1Bf7Q9YHXyUeN0qwPMp4u+s4PYajpvshG4jivW2Ir/K/MhK
MBp3xmzyrPXQJ9VwZOmol8IkytqCgJNWbaXCAiE/yl45vzc++uyL490SaXX/G0BN
dKaseMWXtkTQaXERNqO9X50iK2nleL7Oo0gQbpY6G6c/teHL/t6PaXqJhCT9OGsL
MFmgFUHCVoGKFwNZq2o9L58DCBH+Fc8mPFyec/vrm2D1kSQni0NXY/Zdehwk2dtp
IIGpQpugDViL2HAMJLrzwXiAfVOw2ZkiYaucDDj2GMWbovo3AV2x2GOatbRZWGxd
i3KSPzsJlgj27c4TD1OWaYe4glEoiAvi/ND8dpIOdrAOxsdpNrLp6e4vN+UuF30t
bnscLIxuDhoEz+ixbGXgSJ2qWIElemY6nYavDW6+zl1lJrDIaV4ukVeSdOZMgEk5
aXIWMhDMbTV86v6mpskkqC2mnxitozPDEkni2/esqSeUySqjVKxWVdk6cCJSlAuq
WTMAK4qdO537eQHFmMJ3cPXmFEBmjEg2YCBXM/zlzT6Npi1obPZVjYrWpF55HEuP
94NIOgzMlbeCoKM4R+dSv1CTN+9x/iB7deEvzv+XR1b5LMOZOMVrDMzdTrngaHi6
axpw9Yart4Cw+QGyJB5pLKozDwKyltsTqNrT/79GuLuhWI7T8ICFwfu3wQMLRTxL
NJUwih12JbCeGPKdRDF+0nWTMhN6WaDViE3KkGLkNmFejDXTIQHUUiin8G4UpOFA
7w3gat3iW5kqE2VFGyBejdawmdkZ3nkMoMPEw7Xlgo+uZwiM3+KMkizDnfw5ayW4
QyA/QYIDSA0aVFykn/Cwr/S+GF/OfsHXxl4KWKluxIbcuevScfZuE1wFEL9R1lQo
8VBfO2bhirS4v0i82M53/ulbsX290r82tr/WoCQO7puq67El1x+tLZG9++0daLHS
k+tWO9nRYOP3AEHHIIzDPHXMrmt+C2ja0oK85/wE6onjduJEjcG9nszIu+44LtTL
YWeunj2iT9EKwodydzlZoqVQxJNBfNTkjkjGNBTKM6hSefASBlo5oSHu1WHWOT5p
oxuaNese+3zwnzLS0U8XHZFNStkaGjb+rJc3OuZWIR6wuQYbusOizkJ+w7j+ZyB7
XKW0lPZa83go8BI52ByZOtkRlpOe3iQzYXbAHOmt8M6IEi3KvCIMHKdlGzOBIuA0
BUBATwRmmn1NC7Iapt/SXAxVuiIFmm+TiGKR93WDZQVOO1zeCkLkJDNnkgx0fICy
kZ1A3bUi3+ECkmrhelpS3tBYsjP7VunzZuFipux3p8BYCyz6lJA1C7tXrwYUTWAu
XuX2h6D3DbgtYWhGroezv7fcKb/vEa1KmOX/mgGEYPHZrErzuKktf3A6DKcM+jUl
NuXxeI52G4bS66DT4yZ6gD/FrIR1Oj05SGY+cFBR5CSUzl+gDOvjuK/G+OTyobQp
fJudbeKnJVCCLPDcimvvEMXG5X2HakdUnyv4s7RDFXp+S7NA2kfdGTT2ZCqy6W2k
wIKzf3HEhdLgzrCCScAAYiPVD+DOEdJSbsjxwHfFD6k+qaOLO6rZf1mUlZJrDXpA
yHg4zM9/5kfKeWzXkdjzuLg0t587xl3/xYpTX11L607vEgEp9O8NyeHON3q39o8r
TyQ0MZastqcaFC9rS0f59aUTZlOm4dTEiRgDsESzolbFJem6DxNaA3HMGLhDaR3F
iFbKw3IikXDBT342jx4pfE1pPPooMzlnIxkkISrN1lr1GlOK0WAou+hhUyuZNPMS
UV/UNKFOx3K1xCj78lhAlFp0i2BQ+FIfp5TfnljUL2OPOxMfp4ZZ4KLpOwZCtjc+
bZAO0ND5W/RzwfkEPzw5m49sWRujK/APUjQ2THTyDoa/Ur19W62tW06epgIWtDOa
zJMH3TRWAGZvusq+T3MkJznh6KAJYq2R8k/WRB8UeeBwaEBo5cT1EbxOHy2MfWs+
+JoiHSpuK1w6d2fNO0S+fzQjfgX3sr01PJHf1Zqz9QnvOM0Nntc8mC3t+oSlRT65
OXOJDw7vXNLopm2eso7VW84+UZnPu1XpHUv7AZZzm0Sos1zRzdxzhN6Kmqq/uzj5
kfuHo9pjBfncsKer3n3WLFrPzZNDyBbqaGWbgiJJU53xXaaRYiaLVQkxVfwssnqF
EoNtBfNE7M4JTaTxKzA9jA7ng8kijN9B4Iej5z43xCHrLsfuPJqHUcXHGG2VQ/+K
nwhTl7K4xqM/Bq2RvrNzkJjU8f1iBuIGRwv9YGsbf7uJvFcne7C7QGlIengCaASA
4XhVUeqvhWhliYQXMkRt1q1mPgVw7s1YnfpHgOyBvNj+MR95ay/XlwFi7Qyvaa+S
4Im9w+ZDGMu7qhN/Se54WKR2Cu3d+aO8ka+5Wm8vWoOS5IDCfAs58Sy5HeydmLiW
TaPe631AWzE/qO/oVUwg77dMZo8/s7ERZzVvu4CqxWFk49QQ/Cco6Pn9y0fEmx2J
isu9xQ/qB4QGjrxd9ENqkXtvKw8ZzuU68rXkNhTYnGgA6fIL9RZyM8JnG0tGLvYG
gnBJ9KjZdBOWKgOImE5ny6A9E57ohoGr3db9BwGDLZam6Aszg4vWLtd2fLx6Sz8d
s8Lcu3f7GIc1TnwLy7KOZ2z6PTbK/VFcbSPmc1DXK+MoOC/dK/1Aeb23EMA+8C5j
KZJ+eSQ/hQQ6eZZY9zi9O+zncbIe+5HPpmXRaw2L3BHQ3g4mKoJlJ2e1k/t2KhJs
gc95/ATYRaFTFbW+eH6hZsiw84e9QOSRXE9p6jvMrDNdDu+IqlBEfdJFRq5tBetc
SyXycs41kwKNcdEKkr4U/mfXBasRtN4bg1zHP1eK/p/A6MRZ9eiXliS2sh8kyA4h
GbT+7yZy6kIZHWaI17U6gMr5bPBt3papsIPQE2S45Gd5R8Y9jIJo6M+cloBUiLLT
6odvsHerZTnDC7MEcKsdL4MLlQ1vyoUgbOzHCoBkP7mSCgYtqMZhsSRpMbO+yhJI
hiUrAb+X+P9XMb6Ltzuubl7GEl39wStJE8XCIqpBqMF2v562q+haRi+nXSlJ9Cr4
BFKVCmuwqblePUH+HqYT815Gl3W/46UwRwF31nWjKhrvuCxjBjGPCjUHMFdyxO8d
5saBKSPicbXSeFx+AfDwNxrHBpfz89JutBV46+gqXcMHw2L8loIkRqObUnO4Dh6d
XIQlS4lhN/IXL3iNK/Lri6HR5zDJMUJVIwKiVeGcHKpczCyB1Xd2DX9hCP/PDAio
JMpM452OOwp2xQfgJv8Mj3okIdb+1V26wz4d1FDUht5vKGXFzZvyYZITxTfyfpGy
Njp3DoCXOfLdLYDOGn3rHl3etME4hxBi0l2jr31y1rzQYe4hFhqu/dcaGz6+ADv4
nRcnvzgIPcKPej9EQ4dwk8alzcHUEUyO/oA5mdq+BKjPDbrTdgcfmO9xXNC27e18
OZ9HvcEWhHSDWsRcoA83LH+0nHRBkjzz3YmNc/T78fL/T7ifNN/7wiLVpMna/Unf
Om2a4oUe779KthfWn1r/EjwQMFiVrFbeiYhY3wycuaC2seuC/rFSNJFVNKnyCt0J
+mU8oZl8Wpg3TSZqIYQMPPdQqlF/9xG7a3bvXWGbHrmshclQmSr2mmKdC/DHoueW
oDpuDyum2QqdBb4MZW3rxUyhgAXPY4UNPG5PJMxzUIt/tbfiTppc1JhGrGqWIexB
0uvOczOVBzZwyctGclRYCRRso2XDJuzjSIlObxWGURrkqI8MvVxEktPmnp3t1ym7
r2kldce9fEToQCaOEKRpy0gdMvbATQ22Z0a9WRVQ4iQioYmQG3NWLQrTbh0pYS3X
NFLHWLrIXADx5AvbwZRPvaS2s3aclia+WCa7NMaxAIIdhFX8FP6+JQHsAdsI6bvw
rDqmmMtXmHxuG9oD3XSEwH4ekXnZS/AdlE4pc4Q6DUrssnZ8W0ZhMcylY3OxoQvP
YrsmicT5Dnqk4kCVAOYnTtoghqGg4ABWT4tMGOfTHH1oGBf6s8DKMCQ9prUutVQq
cBI6jxLb4sSUlD/9lC7eFfH6Bs5xK1fKanz+PUCV5mFEVItVNYtDH2Twqtui7iCC
rNbZLYsr0jqvR7t7rIwH2WCK1GT8Ba4ZrTryt0kdfaNFc7/bg9icXGKvm2DnUOO2
Zrx5BoIUrhAYM29CnQ2xIZ8AYOFB1GMng6pN/2nWCrcPzTvTBrUy1J6o/BNNxtLm
ktQASorj0MJES7cs1sosroTRLPkbaXA5p72RS+V1mUyPWKSm8bssnaHqdP7AySv/
oXpCxgl8YbCdR34J+XElh9qne6UfTj7rlNp0mV1d5f4rL6k1ElqrV7IFYVfLjmx/
ze/j7SNoDSf//Squj37d5T9IZFrs0Jpyw2kwt+hpogUZCLwEeOtPQUlHU9XgZQ6e
FmIu7PTPs/ZHuqr3Hzc8V/BvYTW4xVojcMLoumaZOxsBwlp6ja7FZU1tLPBDU33Q
MvDeCXQl8/3UcpjSgyJOZ+EzIFt2LnHU82PsbxB7/MoxwvAQXG697gd0XDsTO90V
6VIxEVfVdQ/vrWDSzxlYGuOeMNxRVovxUyvoXXlDRmd4nCy8r+xjxtNaom+7Lk6T
d46AbsXThqrUqU/wgo+ayfY7Jxoy5LmwMoJbS4GGnQ9HYbH3XAnUL/QyIBwk68tH
+r2fcamdGk2/BzGXTK6pZ3kCSeuS2z8BfvDnugrljy4zOJYRypVGxbL8ioonKcjN
KkZiFi5IxTgvS1PeBxqIcOEoVI4QmLbRJ7ZVRQthqGBr3oAryvLpYMYo8RlLgmNn
zvp9dgy4m6ihrw//Ih3oPqWCg8276xpqngkLficbEJ8HB8FqzuqB3TYqdeTPyKtj
2zk5aOtvQnVSdMJsFPFkC58/4wlGzl/Pw/S99NUNjhBkBcoEa00fiQoQ7PPEICb2
qBFKIsrZ+QYY1ViXotWvnKpc6YcaB6tR6o/GwYrsHwH3fXerilZSbAyH4nlz76In
onFZnCoVoRP5mNw0RGEIvFLnJrcKlSEko77pTUXs5cpZ3H2L4HvAb38iEoTR00gR
DEw39fBnrQ9T4gIJaflNg8zlEfyKT7BF1VGk/uaVc87q/a1TcOBTtWFZ6KP46snG
t8qeBAOG+ewYPnZxya1+YODPSKjjmLqbMGUE93zaGyMWkdtka/SyJVTfkpoHwGq2
FeuLK5R3uYJnAs3XLjyX+Svhe9iXBZa/GSye7ZLRILZGyz2zMkmPMlFaaQ6tmK3/
LSDhHP2U2hNaCOKCHXebBfnIUkObDfdiWXEIL4XRPg/airX0rdu/73u/URNkXwXa
XA/75wKyic3zotUJQCoHetV2OEWRib4fBZjWdHHAXR5knklrZ+DQT3nVaT6cWOQz
NQnaQK2nepWO9LykYdwcrYqN0JOxIaeby3mhcCjCUZiEjodD8jEEIl9DqKPVbeCz
503dKakRrXNCFHSxhAZu8j79qycDlD5DkxjFOepkz9EJHwFodL3Tr2KSnf5e1Ufy
DiltV5QnkQw3vzKlD/2QXKyBPTzXCVcfiUEmK2PBO1HO7IW8ZC6kNb6bVoBpZF+x
lEOe8S7JcB6kesVxTh7LnV2duYGxArkqkpyJr0HIVHiR4uiU04fgv1gbcRG3bfFm
h+umH69fPQLHdkYI7OlQr8r9ybF1y23i4+2sCePg/GuE+dbFh5eRRmdpaNA0wBE8
bhMHTV+UDtPn1+wuaVk8OhLuwTChS63pxyiDd7c5z88U09OlzabFtPYeuLdFcYHQ
G1+Jeg2hEt+nX15RC2JhJC1cUHe1WcGpnAB7Wvf3XnNc/A5srerRC7WjOQi1vXJk
5cHBWlw0vAa5G84RzIMbYkFMIoLfJEyQeKVvHWnDqp5EIMdkPuYG5oWZfNv39GP6
QtNyKQOIUgFW58tzZqJNFauf5oQameGk++wbDkMQqaLbVeicJ4w+Ez2NDYblghrm
sPcbO2PW216lNsuG0yutLftD1ZkBUOyUIAxiYi8rkXB1eXA2cah5LZpuiAMAa6gu
wicQfDSH3/IvU7GqLRSdiAyhb5WG+LriwtG7CyGPrF5xBnyzRhFmRdEz1rPiKgis
b57g2K5KzAxLfyr2G0x7MoL3opPUvgQy1YnrxFQ8Hl9JAyEPfc0G+BPgkdpDYQVE
mhQSQzp7ocjcyXyCLR2Dl9fI+XgnH5/jBIdRXDDJk2Zwbh0kXIzWYgtpaW79hjWo
j7BB1z/H/Gn+em7bZOMvt183pDbpoe1AjhQxECja/vpKL1xmdSm+S6wqEC7OB8q6
sYi+zcFex5RfotFU/kt6Ln7reBNhn2omKR38Erk7FGd0ixZVZ4jY6vh2/uDLyLaL
CuNQnd8Vh736tiiAXGM4gCqTFqhOgWZE/TuPO/8s3QqmAjwRdvR/XoAkRlHdtAP8
eAq6kQI83bl8V8wAmyWx20leuFHGLPteIISRUG8fPVisW0KdxKt/SMot35Yb58tO
wnU4Drge0ZlOtVB8Vh9ucURGBYGg1y1KtgDmLku/dZQ1fdmbSdg04ShBA5YdhG2U
MPWATd+6C+pxEBFpg/RCnLvye+DIs0WJqH3QyuBORjbwctoVjArV35DWcaAN2KkK
Dfs0PVey1YSfI8m8VCgh5I/1HH5bFxnXtjNq4WgscU4nfwn4MWOSlsK5Sj68VZan
qFPqmDYFU5VwR7TyWuH66CYuuwcteLNauuKQ9fGVi8F0EG4fCd/ohC0B0tOdGCux
lxE/7Kb4ISX4Ouv5ru+eNqhXVjMZqPlqZk3h94s7J6iHALhkG6i6VpYbxBAuilgt
K0y7dKU2So3bLafgG7YNOvxk3uUH3xFHT0NGZeznxOUDxZlPS2NXiMG7PAcSlOnd
Jny/+g/IWEra91g1s3JGpzVgrnO6Ee2PQFKGMPoDRmJAYzyGvIUXfyokEKhATKiB
4ExgY5fs2Q4EvklNzWo1/YcKL7TRiGUTDNBbeV9n6mVBGi6cV2u8RQQAUFAn9MvZ
qFhaSav4hiucIP8J0piFinCry94rr4wvx5UvA7fXwAfsx2Xbh4+4d71J4zX0/6yN
SMsGTpOVgiMMaixqn8UEAuKOBQSJkvy9a+Bi+gs89UYNhsLM2jHn6bd8mne5NzYY
Q04H47GlQCRhSG9325eQO9yoUHpFXeVx72eMlXOdMK3XTRKYy8yKnCTbaBWB3KOa
MFuwJA1WaEecvhSVibmmlgY8GyqWeBFXdX9TC8dwPWI68qpvEFmHc5wrcf6OKgo/
0NixAJlj0EO4a28npTeXtGLvWv+0AL1EOPZzTp9AV9laDnQ5FN+zfzLVcEGLooLh
`protect END_PROTECTED