-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Q9nK+sCUQLReI4VmvRMAosk74UYUqAE5OPIbbR3UOb/27INcgDorkuKhp4S6Jxmq
SFrhpevXmdjKwQHwOE5BaeV2jrHkwBs522TYMKDaE6iuTNSt3THO+toKtzCXClh7
GGUsDf7OMAqcHKPu3MTLIV16t9owura5siX5oQjRhAlDnxxinltfMQ==
--pragma protect end_key_block
--pragma protect digest_block
u/ACfcFWV65fB25u9iMdDwxuNsY=
--pragma protect end_digest_block
--pragma protect data_block
Ruxud7p+QDN3kCUFMPSku+ZaYUaShCk9IN2RtRUW1tn2SfBAujZ389kC8MtMHV+X
D1AmNz5kLM57QZhuyg+cJjgfFV5Ha3UNAwtHoLJgrvnCIkLi8idkciDgGCtf0b5q
r7TGpcr9ZqQx7K3oHHx6KvvMxwEQqMTovi2HWMKOMB2yrJR8ZZpJ/0khXOoJZQfX
9h0RZxeYOLy9TzTw/unW7nuErinKeTmRzEU2DJ/kE1zRIlY5f8IsS6B/fXtAKPCY
tvLB46NFt4Szzp67We6DYBNN3+q32iyi0lHVqk5xVYzAITDxfiNRmwLZmvF8iah4
wA6+e8e4CrBWbD0rjywTHdBEJSDOfe5S4p0RyPBJm6C9f7dufiIbNYAnqXJIHkHf
1hildK0qBS5v+s3S2U2ikBMJB2D1Usu5lJpdjjgeAqDQ6aU/kBAKhY8wrN+5DH0+
+3IuXjVzJzPISPrXUovaVQiS0fbrMkrP5egPhzeIl0ZQxEYZ+oDFnaNyh1Pr8ecb
qfUQ/od+y9MslhR5kj2naXI3jkwhvlKPkCJxGANfHckk+KUezjv6Lp4KBOviMDsC
AXj+mAJa4kHlISj0dIUHB5rOyy87ulnTa/KnXYf13nPQ3OiMbNFeyiQz4C6FeWpj
NhsImBkrFRl9aCbtS/4/g8tSGRII3v1jRSQAj9kz0hwglQyd9LOlTfjIb8gBFpva
mHDaBn2HmauTSq/d4liFkea+D6rG3leb9EabSze9D9SVyK8fxsl5LXR02ZTElA5Z
DGhf3EhNzj/ThG2Ccj/oIQ0qT1qhmRxQdyOe++gC0ogar4qZtCkfuUbd+QSq8FuT
TmkCTMHxANy/C997K0wbzGGlNwJGJiumcDU9kglRaclypSmwK5+MWLaol9sYfIoM
EpoFhIAulygjeK9NZ5HYLcBdXj3dRIBfst0rXlsBdsThA99UgC7S/EZfJ0Lat7Nc
gp4jQNdnNZfm9cG9Ua11glA4J/WVSkuKucEYjNVeVKQ8YFzcV2ulkRp8L9pLcMkr
XPkkiZGpWIJlmmLfOZDVAHutPEKZEHDQ569ImNRdiYaA/lt6MbQZkY9ISkTXjHdw
8JwAyNPvCil43uij2WxreyAnxRoBF3SIVbkZqUvpZ94XxRG2l/D495ubSfUbCISp
vqWf+YsdGAtqj46eEb/uY6I3wlcpmak8M0psO4svsc1UeGj4JVTF9wm+OuO45jgh
7vbyukorqg8eZaCXkixkNPuPU5ZcbI0xJ/f3MUqzfZYshMYxEZzUyXibKp7tWgRN
ha2dtcHxifTcqAoxfguMKslXTc63sqVZzubh70JGpmJ1bGy23SwHlsnhpWCk/KNC
kXtO94FTNndr/Ig8/X8KoDqpAdQuQag3y7bLKcFEADs2dTJz7ozxb6ypnSbTcTU2
+6Eb9QMaqTksJ/xcHkhu7dM2pb3IO4c6AZX1DAVecHqXAVOpiz32lvXrMMWB8DNU
zylxfcYZZb0WIJlxI2Kv+Gb4jlVK2yL5lFXzcNxXGVqYgul1yHuHVmgTKOuVX5Ss
aiJq7P6r7UjXJ2iNc4MIyoywx2PisFsNVY8X70cM0nO3GNyswLz3EAazL3fk6cn0
SwBo6IH9iWZY3Fu2Sib6Rjwt6iNxUtW1BBaVhsCrClrRqGC5T1WZ4cznn0IWt4Wc
ko8yOey+aqUujGEajrxfOOKV5sGIp0uTKqPUCxEJpM7QThBVLZNtH8OwEHUT2qhj
WX4y8/tHeOx9PyrbMSiLTsO+u7L5JTtmPBTeFobUvnMNXAyvGNqGBYjcrVp7FGIj
apIrtptJpHVm+JGYIeydHwE3+lJTtb89CEcEgSMRrh9f0CPS3qX5sJfr0qU9EJzD
adjdWNW0FeKKY6En5x7fSNEz3ufO/ONTANF4NG/1CtnKvuAouucVt95zQFYFbyuk
Bk3IfKysh6GSmOC6AGnXdsR87CI7RKHqhrg3WXtD2BYdtsm0PtdCWSmUAe7mtyfK
DEjfwLuI4zKeYbu6UBOEMzJE9RJetN58728DuzTTuJ0xpXYqzSoNqiWZ8ZS4QgIp
hJ2y57RqR/7SKtPQsonPLvlimbyxN8iNpxw/PkNceVTwwZXJhCRdbEUDllaBdLw4
i/RJ0WFBieN6WK+wcolq+7x5Yq0kUvarTk4uqi3tBtfmuc4jSotuE1/fr8ShXbWX
W6fQ8jTdwj3PcoRbsH0fWx9CT+dMIXnxDeu9L4naS7WIe2HHfU7BgpzV04gTHT8s
GYql7yjg9/n9P71hYoPjuuCHtSBmTk5V1pabn+EzLgI3HqnfOigGu/mGmAQHoOHG
X6RcabHxkGsC2qGFrpGDCUqbZeEy1IpFDXbUc40K69ofIDTV0RGbZQSCPQhMj827
PvbMcc+ZqbyG79aubkX9stCsrpGCgvmg2X/MipPoF4hqIzTmLNybjODNK6U4HgZ4
RgVHpTKD8gF302BuvhUaGSOY28D+ArOD+lJTeptuu3HaacFvyJsmiKGcbfoOIs9X
kEyflM2/YBhRkGai45XoZFLJfeARy0fG8WJNPkCo1R05Z0CAYPjk6cODi7nGHR2l
ii8Yth5nA5YunxqHGZqIcYHXlAFplxjliyW//qK4nspeBx0RqSM6aUQejYzzk1FN
diz5FW8aYiw5VyGa9VktBcv87cYqC2NJ/nc8zowLfGfe3/9n5lS9hlQODgAaWuhN
wN0uBJxxgwIHS6hEa+8ExTBTbitJMDkJCsA7N4r0zw56IOSAKStWswIsMlc5e84w
yVT/2+PcL2upAcOiOs2A7lVEOTCKkfIsiRh6cJZVwKp8f6RGWqEJkgEoWg1h/AoG
+Khj7YjBZnHRdac22rVL4Sb5aL+gPkdQaeq8jFlnNTDGqN4bij3GV5ZoRBEwBFH3
Ww38+x0Mp50mvNkx4ud/5y3wdWzAwkT1drwr2WrHj+uY5k/jP8qP+PVTKgFXyyvf
4w4RthqBE3yjy9dtyAhiBjFqNR5TuwuBKwjIKQGdFTUQMlk2Abx+pqT53NQ16xgz
b31g+yONrVpJA7TdEgUwWhY3/6tVPVa9BtXNV3o1SiTn8ft+49s0JikqG8I4UbkK
xQFbT5dCR3713WTnSa0NccRAUJah68wMSOR2QtVkUdoyxbtey5J5D6iuXAaY1Ca6
hg3Ycqa/XDwldg2xJX/C5HWmuY0Bi9KAtSvfFsJkHcJQfZ3eH3A7fzT2/lB9QmTB
MN3qbrIbWn9dePKkr26uR+tt5Ru6qwkfvKh2H3lmQDT/FrAeO+gzkLEnAOsjZzaK
aCT96HDtzcLfytZpvRPSeW9r6Z5WPjSNpF7qiHeMssGJotXr/G2qJeJiDtq/UdTV
gV11AWOvd609x4tlfvte4jO4DR60U84B0pXb5cr0zd/Wl580C4MXjxQcoLjGdicp
w2JJmBj/7zDqeQuvUzm6zwncOfkXwRs07ngjPpw/riElpK6w3d4NQ1jb5IJn3ZLC
7pVEe4zZ5H8/eUug5foI1MNNtv76Fiql00gBZBV+5eO3ZEm890sd5pcx2JPNWT1P
6HaBqEGBEA3GpTUzhNiqY7abyZaAPWEM/ww1udnnLWpuM8/vfuHcFzQ4hYO5QVD1
A+/T0qaeZH9mdZK8lJlOGlxucTW3sG0lxcE4YQV76BITMIe0tiAZGxPqdqklkkGm
Vo8Glcu8d7RgG9fwAsOEiH0297IT7HU5DF2XDyVj3Ah6M0dbu+UmlGZAE+0aPSv6
ZxXRnFRq4V9izMd9/uI70TuHVRF1ud22P6jI8Ihgox/utbFC08jMtRA2NABy5joI
teD7IrzMgU8bnolzrOcXvJzWtkMtOK90+zjjdAUr6ha9Z2568ZAxX+v0RWCb0xJn
pHqeDYJqBKqJZhm+Scn19IUlagUITfTgiqsgaX8VfQT3E/fykYkevgqP/GQi7ykM
8PT97TAJsLV89yTarU6iwJ1luYfbWis3PYLqpcm7T4z7qhZxQhJuqGwomit8cJfS
20OfTl70ycKxTeDGZgUG65HHxOgAmBzXJLR6pW7eQDr4yNtHLqdjxvwdMp3vZvHK
7wwAjlzO+WSNsh2szuln8QcmfA1OG7IW6X6LY/n8s+IjPGYkvgDyo9wgX5M5xokS
OVq4kdkoHU/BrJJi6MkZlImqwx1qOYEsnH2ItJvoS5A/3i9yf/oTwIVd2bBsBX6W
TfY4kAZRApilXDy51I1UiRsy7e6gWhpWxzVsKkAH4NA1jZcDmpc3LAnhsPJXOzHR
ObrrdalRKTtkZiLMvZ11skuKsx+5cZzgTg3cWav0d9I3mv4Bj28+dp980/gWWtiF
GqlpmgnVkD+Lvg6HvRvs+aDqmuWQcCbo33Q+E8ymuZx29DS4oXKLEfsgx2Zv2Akm
ldyMD9cTpedLHfF/vqOMeDZshVnKVtAFcDSMnrcKa3uOeZ01jkU2c0/BM1ye/ENM
cT3yXszpI0VfBkmT47qdZagflCJLTvLULTqBdZl9/LSJVFtc0UQ7vryef9auq6LD
+YHtBMLlXUYqJ7dXMCpA4F6E7IJnMBhVMNdNdQ0cWGUjxNkg6bbmmF7KX2e8km+O
lhcVOetvT1hgdkyq1d7gE7QRuLp4DUSAlPnrNafAvxKDtibl4U6FymMs1BXjrFBl
P+o0M57dQwcVs+hEwwK6Pgfcxf+5/mNFSKW2i5FYt5c1AMyvC5ik6XKQYyUwW7wt
Fe2zeSZYyYF9YDFI+3a4qtgJjLSCrZxpddO00I4m5jmfN2uiinxugBqbgKfpLtrn
0hOaCpm8aGo43pRegaj++S4B2LL1UP8K9mvVe6WNCAMW7JkftJgEMmW6TILOn3Hf
EN/zyg4Akya6LmWZIFrbPjAdWjMkkfJQfMC5cQMRX77nr7wCvaGo7o8IVRSrgKYN
grXJ3mqK2+llOHgiiDQh1yyaPgU/a4wmXdmQjsrKW53UvahEb11ZWqETo5ZfrEpN
XHuO8eMVjjXaEqq/+9+xaedin0OThjNqakrT8xkyQBz+zCju/pT644yCOMKDS52Z
tVkZKp2DbpEJNvlEAYJGiSgJDk1ld5GEOhJwB6aiTYsGjaCuM1aGfBX/80ycOKqy
dAmOvrkD/rVGC20iqAe2pq/ZwlB3Pw4mGEyDVaCIhSv8/4OoBwdbyfcGR4T5PIze
f+YVmimd2H/ckzmXqUJXI59wYXrTqQ8QfyVdkYG6WWVVx2LsFIJvNHzjxTGkMJTo
Le6VfuUBFaTZDDYnt9JsaOma+tRsl+cKFALA2GkKCvsdBR81hgXQTO4uJYGH8GEY
gsN1zOQwogOalakI/8HJRJibkgGltEVEQE4lzkdunenje11p/OlqbJHlksTDcGDb
ONNVeFvzEoKGK6ZyJJQD/fgt6g31vhLpI1Elubtzqt27b3NiMRRIiFeevukV0YD8
Ldc6Os/YkWZWAQGlUBiY6eWvsn+g40yKak/3C6nk3DFxBxyujN6gGbEH+fZZvFj5
OD+tVa1NymdSw+M4Q0i65RXcBc58Q9K8udrstUGWL8O6OO5kD/1CxtVMdw1aY75d
YGjMKtsycYfB1Mm6mA1fK8eXMc5o9HOG3SqZip1fWMF50s9FIr8gYU7fnaJaOPjD
G1Jhf9PRM7r6lwWW02vEtZfmABoQkfF1Y69ZY1U1Tf+osxu41lUNtv2XghUiXzOS
uNmpqUjOp+EkNYWEf+YAIrRtwNZXzUJqxM/RkGnrZxXI6CH78Xj2K5hobnx/867+
ZtheYtbKqnY8C4pIGEbJa76TfIUQJ2xAXiqpyhHdBxrib41eR9ZSuEzAwDN7S9eE
xL4B1P4y6j3UdkPpPxo3D5Jb+6Hsj61Wkr2ZgFQVIjyXqGQ9Udo3RakwD/4ZUTfT
RPAP2FI5NWgnLvVfig8GZhPHQ+Pe/XjZo6zfRUoT7lcDJ+lpD/MEC1UE9Y88FGlW
wOSkb0Vr82/81xgUTXYMwYMNYKWFtfZRpp8HyzJPu4MrBPKSkeU5Oxa+/2k14Old
mDPYgEAxbdDKx96Q2AYMeMnOJO0QKMgjuEQ+Ywcw8HiRCg/xtXXie2Z2bOnriNal
Gpq0wMA3FxfvPGk4zc73RlCBlDKVJsZOzjFmG8qbmEqJvMVLxVI7VpGFQ8+t1xsp
wiKr1E6rlczj830e0NiLoWVyFTquLfHb3EEJxGDyqmZwsPXeoVa4KgAULYYFQAaE
y029kUxwbbvajwuNChXeec+U+VQF7SdOsA5wcsE3SzbPYQYhzsXKGjVNG5cGNSjY
kkNaqUahHMu8M5dxaVANQgXQtFNsx1So6gNuNKHXfshRfnr9aqUHxSsmLl27KrkR
ZY6CZwHHLir8LOcYKMTzHsyaSG4dHlhVFiqam94HFox2NKjYoMoLxKOYsiQ2O0gM
pjW2mEGW0139VS2DfSn674IbKNgPl1rjatT2dhCsRLK5YWrnXmq0lKoKA23fmXhU
Us7uZ2rRJNS0EVUj4EqN0X7XErspbT8YvW1vIIzrmf+oAsGdgVZKaFR/+FEenezb
q24Yj50qttLnCqsrsB4dqlF6rV8Oh5dDP2Gk4yNivmXAL8yQIC0BTL18n8hT/Pes
sNgoXT1IBEd0c48ArV4Rl4iaizkzMi9uQoUwXkOonqhtWRKyEd8Ezm2cGWv48TLL
X2mvwCgt0UDcdHGvYNXzE0AOaQBJbe0WnhI7SxBmQSufKttKOrxgbzlpIZeGk3Q3
oB7hBo515axFdvnCfEBD1EwIezm52mhD5POk0TTHxLd74s7sXG5hd2NoxdQDL1un
DKmq5IoC9EPdGv4wPDqTT5DbOh9nJl2zRtReqqby3JiSbPJ0aXLiYST8jQbRmsy2
Eq9E9sBfVDIgg97Mr3j2APwo68MLvpj7fYQDzbDbXK8NqXwcL60iATR2jT/3SW+U
F6Plbyapd8uUS5vnCJGkG/mHuUF6f4apRonTiepXPDWc0Hi/GuSvpHTJ7BBPL7Aa
AzZObOqptLw5YGV0yMmEdgEhYzNGyCrrjHrkCwigywMcLsx8Y8frmJwDHlR9VthM
nHH7nsvTVJ0LkZbK5soOgrZafl998JdsL17/EeNUU2s6PR87y/m0Maq6I9nJDJp7
Ooq/A7WFzrAlaBNw8eFJg44igWrXLDuDDeOnhdz5mRgpRZ6SWT7PsvG0kfWP1tJE
85nY9p8zT/9qnht9PD7hAtHEWB9DgxTEtCO0lisKJmAKGx2J/0oeuHyGCYDq5CKo
B1CQ0O7aDkrmopII1n1WWFhs25iMy3tq0jRWlW1s2SA2VTYtwodk6eQZ/YbOz9XN
mzMaFbpxbvhNxPklgTp23ysStdSRZSd+VRmeHvMSHxMy9HWIfw914W0TDS3aVkhP
n1odN2KM+pjhpcxcxJqb73p0OVa3xL3N8uTrrVEMXnnjeL8Ar2lBUcHR4Wdnyhuq
qiIP62ilQfX8ZZ6MgNkwie5EfNi5QiApAzIIZh3S3kQm1mFhWLE/JCYR0QHiLhGv
aUkMrmom65h+a78XxPCW3+p0qg5nYZQFQZ2olDCBjNgxII4r928WA0Fb+WzWblsi
W+/mnccMAHSlWmB9G3oYIlgzy4wyfsimWjSGQWTvxzJe+i2oWrqHAzIs8mhTTJFF
sErQfT1p4F1ClDdViCL6e/qDnpdjGRGf0AE/+rdmsYRcTMxffxxKZG9OFxiSWOQm
5dITrLLVOVTQVR4crYLuaAEJfKgAijFmm4guh4cQJ5OVSDs7Kgom/wjPy2Kj6Q/C
bn4kFDPlWud/vHaHCRDLqY62pY3ZNobm3riUm3NTsmuX714MyfmOgmUzUtBojNyr
RaoQwYiM+tkUik7xProM3xSsFB5ywwzf9YDWfXqlhgnj9rr6AOHOh31bGpPHKCDl
I6qmRcxEQr9oHYgrbz0vyJ8/p7LrX8yEQxwM3nI8/qrnpjAaE2+qZsNhWZ35US5D
4xmQiAZZUKasa/xo3Dn65LoukBO4ZxoKhs9caK1HFXYXnYxVOSByGPaxRNBD3z8y
TNVprpIoR/JnTwOLdbUnIzqoYZOYHgZd1Dv3x2NEYF6oX6gw+X19CyywX/I8fUwG
UvWhqyYjVvh7J/cpy223aHAXj5O+fu3Cj1pr+7EETHufPI/5Vl/8uS/S3Vdfx5PB
HPPTRvaL4QhAzoaq+uNaRTrV2Gj5BAr6ze4Ec/TS9f3fM/a7kj1mhhQ5TOun+VMH
h3OjwoYtMs4fnB0z+8l8+0jPCGHC4kBkJBrhfauVzf6TsEqpV0dAuDcYMCvyTGi9
Os+BCYTKi4E6qBWEA3LIgCFfz/6NQMhTrPyI5qK2zt+YN+X0hJpfneelA5NuQx3u
bHvRaiUwl1WERyWZIGcc1ozLQtrU1/HDkOgXJ0z2IsbXK1icE510LHpRlNS4bPjn
l8fL1yKaxYAKlszbcFY2GflxfmxMG+gr/voV/U+DSHuw21CilByR7MaVeSUVrXaH
qmGewO5QfGkxFONY4qP7HMjuQWviKDk1pdPcufNonQWxe49knqKh5Rou/wSruAx8
gDbNL2fEaXUOUBtlG6/fSw89+Y+HZWTx2YFzJljUmvuUN9iN/SpqbMnbvT/6opEy
aPxiyckBlEXsaQxgklwmWhIA5Pwmpsfnaxt8MUz8nnYxtx57GV5XhE5lpAnuPVbX
bEBt2IQCHmuzNLSRVgFk3FVU51oJtHHyr6PwyMny1T0aosAjMSYdNL2DZknAlUgL
0/OxG1yKXW8pK9bHH3dnm/BWVc/qFfIFE/wtCSH3hTV3RKIP5dMobvZMFFp/54cQ
fRs8nMzL3qxC0WCOTPLbUysK9/S4kaZAlraDyZ6Z6+mcwmB8VRi2V6rwmbKfErui
Z+Oz2U/vP2ZeUdDbXgoHMAdf9SgHsk+T4o2g3ONCdtsC4EJWsw9xT2jMBI3a1z8T
9+Tbbf0VhKthQfSluoQrqrtvvO3W66HngYKv0lJuf81ffcqzZSrU3MnmV00ogrYz
OtFnImUVC5rQLfh4mw/QraGO2gOuKIaZQqklZOKv4fCDPb7q23dTKjx/fdAVZJaW
Nn3lvdOfTSgFXfH9w/4gIQNIL7I/rgvkxymnAs7rnF9SKbb0Ywz6OJObyQrcACUy
GpUlvDtpzeRVN7EdQ7usMOxQtNjqR6xA9OeFkEWtgYJNh56SfbMl2bMy6K+YZyEr
zE9s0v9nk9UaX2nlHas1oopI67mqmwdTgdEee0/qJevsvrdBzqY0BuNG13vvhw91
SqRRoUBMUOFogCIHa5FsMMeMVPp6yd0fbUOesRbKmH6jqZ/f6lrHV9bLi7ZA35Zw
dagjUzHjv39g5WJDAiJ3e4GIPWg+otXhteZ7O0S72IMLB5TV5lDQ/tG9ytgLYC5p
DfLqNLv9SF9SCOSGvSY1FzYX3DWEkNu8U6PfeKpWvU7ErVSmCLRVamHhFyPduQ6W
5Lx87VCs/RyovpjwBFddRyHNuAkMgFdgdtgO13XmU5uc5jZBFWnx5jqqRQB5D6vp
SWlaI9YBfhdOk0gHijknQMI2BzPc+QDnWMPiW+8G70RUaxN+GXiuRHGxd+2l2QdZ
aDdlhtDt9+Rq6pNluCA2/5Dg5k9kZradNWK7RQJupIBFy3L/HTP0ZatX/hKvQKNQ
03QaZzArZ8cRYlcXYOsjuFIYyOLps/5Vmj3nXngHT++l9etcQBh7DRNGtvR+isXM
+b9EEKRBDMn4EOvQFi9e8e9llN5RP5/9M4kAOxPL8Yi4cBxfgseeVrQ1x6uLwvyv
O55gcW5a4IkF5ozZgt7Rj3Cjr2E3wjZ2hgiwW0Fxj6kSSn8df0iZfUTFQOj/YOVd
7XV5t4XrM7gT4TO8p9IfOA2DQhUqWnQi5HC4mPYHsZt1JAVs69BE+uDLUGmPKLY0
qPPb5Gnwi4NWx6711On+ftp7rc1iIFSs6mYQJDGwpw92vR9AjpjzGb+P6CSFVzz+
a1qRT6WWiyzx3YVz/w5VwhH6nCywEUu1UEzTVkv4ccWkRWLbluVNZ4kCwjqtU+u4
Y3xvsh7FFNHSBkKjqXmDCt9MBYe3gHT6187MLrSAcRqtllyb1nrDtcx+tyfvL648
UXdpRZYmgqjS3TgQRqHz5CxI46vsZL2DZn1PwH73Lm6z0oqaMt40qpgXFhicbLFp
+8mRNy0smpBey/fiJUEFc62JuCf1ceEbVF1jBY/Vytz+uYdzfkxiEzMkAAUu7eUc
Aey85258cYz71hLlr8PuyT+IRGWIbJ2fZb8o8BTWRqGN2vN8QiEAVwmyyhE6vvHb
39Ez+D4YNDw84PSwjKjswGVOUNo6ksO2C34p2CEgdzz2vNR8twpkfhAW0i13dw+k
lxlsH3536q/UBVqTHob0JuJiweajlx+fFiGuY5ZsflVn0EnM4cf5klYAlR2FrKGl
wPu0wOOwOktQHB0/+x/xmwUNktKWwx79leqbH0t14wZyDqsTz1yuECxaHIqriF7c
eTVz64BpwL6l+bZx1rNyLAp90Sgppbv51X78WpostoPMRBkeF6h1l4AtuzXBYBnM
ioZ75rQN1yqJwatnwr7X1dWCcsYhfff+L58tO2OOBE8bwLVLULgqVRRUFFExk3FY
Hu/T9YbxI4n0e/118FdCgNjqfgxZ9PUGqMg10wQDcBJuSCHJRZemCi1uUTs8T78A
P3s5dny2yeJ6JTftuSZucfLDafCZClFxDXKxYxiL/G2xvWShW5C44uUSCh438woJ
e43tYOicXIxmjv/Eopouub0Nf7LYCIc9/QynH4ycMSrJn5lyae56uc3pqqloI/A9
MQHXn/qkhcMVChMEsjePgDwnL7ckRzUKcz0ADG9EnZei1zSWgjVfbVzGl726Lz4D
ZuQWV0J4debWdlt+jaeaVWqXudg41VA5xBxTS8X7gKUs9BRStDp/WO3jd8SiIDr+
PqJVI/YjUJNh8YMdiy7UN2e09jXbbREiqcbz9V6vr9GYP4/1rlRADh/Mkfzc9t+a
rXMBFqi+NXO+SXgdo4D0+OrW3iU5J+o14tNYSQl5UjIne4G9LKqpY9AS4T9hTww1
z2djgbuQ1I7cNYVhrPOTBRoTZPqwm4rWz1jdjCPWg5b8SZHFo4OunbFAAqeDG9ys
bZZN61o0s2rVPIDwAxCyp1UgtCgBLzs/BYN3rKHuDpn10zTym6XktGJ0vhitxJA6
oWMQA8ZlrB8ynSxZ44QuNdCLEjK3TNK3Yje8bK3+39mO3HsPmjMq2C6sCjpXGCRV
BCdf2YCS8X6DuowVdyXR+vkCH/m3Si5uEYh30jDFSScUJ7Ig5cJs98jmufIUtNM9
b5D/msnv8swaRofs5ZoBW0LzvrRmaLYk4tYX6GeAMMfMFtTiCVE845lJ0XBcvWCt
sAnnV6+uf2YXKRUUlTn+VRXq2sk2KzJUwb47rhE64XicH93a3bjcDiGNydKPkZJS
7D5nGTgkC0jqBBmSngEvEXB/UuFQrmOkYiHSmYeCXEPS5XYVdsn60vmOblcZKCBJ
kqG9gWFIRPd8ZhXa7ViSgXgH6+p5PBKczBVTcvUj29FHrzJjefwiTIoZnQDf7KQZ
7Fy0Tro5jdD4/FkxH+aVVvvhG7FviMGkRh+5asHd/Dkwh5f2bbw7LMmjQ/D6qgw3
MP3iEVuxR87hNECuE8uKvB2KXEOwaFVqWZV4hUyQ6mq+hamuzzVshGU264v4wzdR
rSbo+MSBBhYghh0hqWaQ8cSsCkq1P8CkDgjxO56w6ARfSibR1YEIivpNQdnhzEZu
jLn9Zn1sCYjIXmIC5kWMNREJJhkUjl+cOCqTCoS1ex+A1GS2+WvaXfU9Tyz7R9i/
MdYE05ce6sstWiwuOEbg1Lly+eBEGODswfVva+HiOII4kTurMzKkkiq5mN6VoCeT
1RoBjK401U2N5U86fuRUNuEEpSnZJTet1lTB+GQlGfNKNXgIgJc3z55YLChyvNZu
b5dU4LN9JR2Dt9i0gMuEWok0tQxEBhCmvR01BdBs/KFAnxhN61+9iZc2IFcC7dEc
+naYxX2un1csLpZXB84zE50LkE+O+E2aUH8XY55p7rH0wYVu2tBtiG5YrmG6Edn4
zlT0b7/wk8v1jsDfO5jKexKYl5l08LykoGmrfbgB9Pq1KE07RXUT0dHOasnvc6CL
9itRCXHaKTBIX85EJoy2X/1d8ae0GaCRnEyaTV1o+AxRogaElcrCRmsWwb4rd7XE
nDj3SOtfZiweNgz4/0XbvxgwgoWx8CQ425sRVuBi4k8SIkIgPQDODg2iNgqbFSC+
EzNf60j+iClrdh2PgsNQncQNs08plrTbcyzsqVqOCVQBcBF0EQlvz9dLEv8htXBd
tzxZeIqISasYJT1iSLRYzll1E86Amn5Iw5Tq2D0trlzoY3Jz0Ipc1mFXqtOkB1W3
Q2K2FFqy1j7wYHQ/DuTtdH7VhFUWn07O93tu+WJrHdw3+pHtK1JiflhpRf+h6cfA
xrJSyYCVaxMheyzFMDyGLYb88Et4hbPMehXw+gFRm6y31cDWwUbDbUPFEyLeAytF
5Sz7BLgPAoK4VdKueg0roeH8YBskGk3HtHSx+pIonyvGP3FEvzjuPlBk87aLmSAb
YbdcxxFhoQbAyEWJ6jcU3qyT1vct8x3uwFIRfudbhjCw1wCGUXkUhYLqaxOKgF5m
CE5J1WFnxRayZc8ec7MwfpTnKysloWlJCCB/lWQAhg+Pb8cqooppGehEdTiorqZ+
3OLbAoDAg6QbQliERqZ6r3On/mmTsGyYDfyfcksQ9m6BpC8YnJpsMQib+lLDwDxz
kMThbm0/UROAScELDddN6CZQ8AwcbkTMQRCONWUCdXHIHxzaoFzcW42WoNmFCCfw
zK9UYuV2RUTn3hFDpHVt+wAwbkMfZrclMXAKNZaW1rJ/Z18DAxbnrI4zi7OZCifD
nTOWRRor8uWliM263EjGjN9rVvcaif7f81Sf3mLXYnIOcoeFClG/1f5o0Mn/0UXF
OO6q24c8AuR6SrYuueliZBZEA5JqPSJF1/enKv4G/Z0GSE35KVozKwxLM+hrtYx5
tErfxgLSQs1oXGzROuI7ZQUl20O9yW3AwlCKNCe2tY7fc86MU4k25Hd5ji32TDnF
tVZeciMnj2/EgwOwSuu3ivbtEWPr2zxdagn/TNwVW81S7a5Kc9mL8FhodBG96One
kDebDEuhnOfQAmvLR2ONl3I8kFxE7ahA1VbWK3ZyLDY1fHC+LYasyAUbphG4yduy
odBby2wCN8CANla8w8JFm7lCXwym8f8qWYuQT/pJ8BV0cw4xLso+bSZdzjQ9hCyU
JTrz1k1Co5PepTUG8FeM0Qe2CfCtPhRd0SU4yju2X28nS9X6XJf2HjvFLeenEY8j
ctiHtIHI7+6erKQctv0+CLpYpNFitj6VES3bms3Za6Zoe8iGBFLneHvo77PaB8MH
0NNAM70b6ra0bWue8n26xiWX0GLWzn9qlfvrOX8vTemnmWwxQmD0xmp3Zs//DSxv
3zaKKq8sn/VY73Ez2uU+2ZfH8Am6lBetfffF2SzIKatHD8dpwaY520JRJ9IhTAzt
+pY6b0f4+iWy19DsyAERmwAkRHpT51CGju69kJSmifCcuR6zIbLHnB/f9sU4WRPN
rXc2e4/h9gd/Qybc0/Nh6MsUv5pbRHFsAV8jt1+8PtwNJNi29+4Ee6RazN42JIDS
vnS4dzS+gD5jVyBKUWnzdtdPkujfc4F+40Z0xtrKUMZdJl6TB477XuiAUQFuiRru
dLM+FCHzLaJxaA2KDsci2n9cs14TKyqlMNfCSNDvxLqeN+ZBdKnw67TPT+NFV9ZC
/PI1xDbcPpopCE2GRSsWa7dvSHzjfFG+GvtrzMV4sGGVlWWYwQbiz6Chd7aCFW+I
cpCBBknPqZyO/qbZPmlo7QgCbAm+yXgIy3zoCiokHraaaoz0+VVZImyUIu3EU75l
lUph4RYxarG1115LYREBByjkpEkYgJeD85pm8JhY7U+I1uzzFRxIICAAjtkYRyKG
LlpcNHwuPn/XYu7vjqc69T9S6BZyk0A3ovPIJnMcqoOk5IH/NtkFepMt1S0k5ECz
KoN9fmTWQR00UTOuMO9QFPPQNYZTL/Vmuq4/Wflb+o3zaIRgp6HsjiWFdEU8bK+4
AQzm0iG8BR0rK1+ixpRB/AMbXqC8IrY5lT2lx3j1QML00PQ+PPfLPAGP2bzxWgmH
Dk1UKKfwdw+P8+6H4dqUUd+r7H8sAD9o8U5+f3u2XeZ7F6nBDPNUw0Atph8vPN+m
nO2aR+djdLURsdJz9hnPwDfrOlWC7FWCHG0Wsqn6+QUEdrj2nl6Z1NSGqZeLQvJo
os5NaboB4kA29TtLUcG/cVNo/QB1g2QQPf7TQIVu6gCjSZkoRK0BN+zrXLMjMXk4
iF2A5oc4xUllIWolYJN0ZrKrr9pvLXb72HYNgac66LmJn7D8gjuL0WfYv1HnH3pc
UuixvGLT42prhIlzlkULhIYf1w3TeJ34kW2UyJhYJ24Z4wJcXu+U+FobpH6JFMCL
cwPuHJO74MGZ5eBuDrPzDeoBEIbxapVv1PXNM/LSQFNjrMmTEVNEpG591gB1EItq
2uMCdfKbOw+Y6WmO2s1WHAxY5O8Uv9aO/LngzCOYAccXlDyW0BTF2NrUx4yafD+M
EdI9S8r8w4MqzTXwAoW19x3pktm5B9VcGkQmH5/Jsr62ai2Yd5wP25j5C/75Q8fD
23/kNDDvg9bB2VB3Zt7jFUFGiqUd2gXEzRQqiok1D03V6m2NQVaOMEXe8uobrLq/
VX2zF3TE8WCVYGEkwD7VyG1nL2LEKwSj0EOmy/HjCgcGedHGV2Wgqsr+ux3xGwwB
d0eQ0xQE3UEBpCpy5cS4+2HHFSaWNzFZAPRq1IA82SeBS6/wK/Kp6xP41/rcwERu
qzYImjPSOJeiFICHJSc7CgqFfZT+9DCcPTera2s+WieLz1AXxia6vQPRsD+KEm/E
PZQDrWvItY6l9RfVmUwy1DGv3FgpxzrAxL+XwWAdp/wjyqbq/6lkW2BHo8vhLie6
1d2fcQwFLOnFX+hCqkvNw16tta1zxxvW9QdS8+NWpa9vbazHgNQ90d5Ci2j/0L75
b4B8W9lyF9ljRQCKzn/5BeMHDbt9tqrZzMB8gwmeVn9/VHjP/2IjNvYmZHTUo5C1
uoRwqhjvL7nfIqDTrj63z9j6/UbAtslGHYgPFg3vk5pBhjFEzU+ya1FKMNxVJpxO
JZ8vIw0iAW9qfRDjLN36iz8i6c0679jRiliUpjJ96ZTMsTRGdhRT4FsntaJNYR1A
jlszMe4Z2Voqp2ZxI32PwLzHj6/va3w8fRccFWG6a0x7CvL2TI0u/LrAPb5gQaAc
Z8/uF8uETVp08a7W/mj40Um4qv3T1y5e/9a+6II9cJKjKYOuqE1HUFDascX8QlIu
NINroayH7zHkA1/z/P9X8kEgDrRFTtRKsL7lKs+tHk7B79vTJeIcP9pyjkIwi+li
mpaLFv4dmg1ASvBgRIU15B2VtFxed5h0MfUewaNwJUwjEnqoyYn/LZCHQcaS2vYL
DOgcVldXIN+4JADKWkqEbRgqLUiKPQjd+wUuFbuegn7at9RTxeQ5RbS4quL4Bknn
zG9E5dxW9h8tOlaj+IMCRg+FA+FlJUMQvpthtL1i5bbAqaAmO5s1WRVrU8EiF/kp
VHyHlAAjAYmYm2CXUJdwsvjfqfJS2iDkwco71srRoO89CBMMjY69GpQLIaW0BQp0
B2hB59MCjf2JUALwd9x4elrYk8sExsCEdo8kdsbIFu8ZBzgKZFeYds9Vho6NzMR7
A5VbaFz5y6evzV785YURDRkqA1s6doUlZxdeLrU3bcwcc3m/VFFpbTCHiNGytLSP
ac6t3WW8Af2C3WYg7dBDSbzoicM+s4CnTurCmmbmZEm2LlwDTtI5lAemsE5hO0p9
clWSvDi/xU1nVIjAYLt01AoNqPXm140r6eRS1+lrzJBXRRVyxJUmGtWXkEQTwi73
bQhWjKKfqixPp9uQVRTlpTM2tYVk64kiEIcT4tq9ujxj+wj6rOoKxqzZVPbqd28g
6TCuc2Ijt+SOI9+Cm3G/4sT9pK1pSBLY6Ja7s7Gv+YFTOsF+CoJhlJkfY5B5M1eQ
3pYAaSH5oLfMnqo7tA9n+iU2nKIqpLK4z4Bqn4xVXH8PQSzH42knit4hmzpey7eD
hLO5ktq/+Ae1XCuWI4UJ3O61mm4CLKROzpfHohrwZaZK9OvcywwKrz57YBQeG72p
myYLD5rIqMKf+wz+yp45l1JwibB1KidrNGNaXkwkldjGv7SgDqPtFnTJf0IkLysi
OA5SUaufzFMueGMkZM2APCiqMPb5bvCKFwcbCVkENwuol4JJ/dGCz/UxNG5pEx3t
iH5woTTiVE/IGcNYwqZxeMx82P7vbsmveAZh4kPh5HrNUOCpDkOq5P8l1X1ZQxan
27hNIKrk4YpPOfE4WCBx2b/MWu03GiM51LJcqc6leApt5NsDSGST9L52tYUH8Adh
P/P9SxqM1zR3B0F2phOQPv+YZwO91OI+ysKd+3chq7jffsfyCZosl/i5lNxPJeBE
GneIxJbYnOU+FQWtyo+tScsmqEKPEUVuxdHJWBvHX+h/7FEK/OFqiLP1d88u7VM8
MT8stXBF749C77vyQ5/dWvWYpD1TgAbR/le+nE6PYEdP983AavMsY9PttfL86cMT
mjcMbOWDHBO11hOLPOEsQahJ9Vcn7oHhPZ4nOis5PRIFfGGfhgXLANlW+We57+O2
WSh7YjA3LARxmg1vmGeS8fLCCLtMrJ28epKUM20gtbRW+k2I5sy5/oMq3z7rSRTT
fRuwz6YVmUxnEzlDftQYfmLZRyidWkLOMc8dmEeryCrKcCuj8kik/zpixj03ZVdO
+FGifjOrZgW1Sz77O+JDL6JaDPdaXQvnGRAOKg9BaGGC4nheZWC1LVGhJBoQs3K5
XNNmGaMgFzV3zYbYbwAsXMF9r6owodmHRN3ne9jvFmGamzOd6BAlmtDexNqDs/I6
sK8oQDdeo93uu3ZDjncnTHFhiWSe2LWZkijtAxJMornD0iQOBuN/eZLSEvEZ2xdI
+aY25lIXJjlCzRSlo+5K/uxoOXXSwyNDHLsDNkBjdbkMv5p89qGJsYJuXYln+Ec5
7Al2arpRmG37BSUBaAh6ZBZo9junqGa+YdbJpFOMaYOBWpavyP24PApZwv2KgkOa
Wd/QIE0Uxu8HkM9I2WkVGw3b3qCVdHL6ivdkePpcXQ87H0CXEc2VOTPzsHn4q3gg
Xje+XUWdYpye+MPkXARrGK2hTLafasrR6iCTkMphrKuH5qhRLPHgrx7z8TSh8+EP
reR1mB9aXitYLoGBbSCHc0gxRYk43Wbimyo4j5uUhKCLqWUr+qV0sgNU/60bvABh
AE7/OwNNDquszhf0TEFknHC9aHPhybjwg7sJAL2lG+jMwfYMRly0AhZ7eIxrgLtB
S3qD+Tz2nSQhI7tCCSYKWBi/c+KSaVgXSvQrgH0d8LXpML57gCzxwWLUi25mA0WC
MeV+UqtToU2GXjrhQrsx91ptWOTgCC0safIFUHzxduRwhCjpxoPQCZZrITfwFMzR
+r5XF2VsPz/AWzx+T4qmSxlAmJHaaMFdzZj4TYAPdAcYXd/KBbd242FOtLpVakKU
yZdcD9sC2cjjBspKYUf6iva1X/GdCLOn6184TnOImdSApYnVa/g3+IsrYMw+efBq
z4JlnTz4F+0XBO3WC4emVNCIScWyof9isgStuiolGvg8EEDbJ6WBG/2nUYML19I2
2XHYHuk0Q4ETkE85coWFK5lLpDU/ZKThV8NERFWoJaLjBPD+jvaGmjzGyHj4uPHe
jDfxHd9Q8zjWm+Gu6GhhpMrhCoRUe1/f2XytOw2PwfZBJyQCPNZbJk8PLvaCn2SV
I9iuDhxTm7KiK1yKgoZFhl17zxDoAel2Sr8CuFBweF6J+kf7iweszvkCr63IUhdF
Fzd6IaCvEAO8FrprKhrKaPd0VEbIuntuhRj3h55NuwxDketrJr4yHIep2Gq+A93U
38+xvuMlcHFwnDPsBHV33+PS+JWUP5WZFUdobj/2YeK2CswnZqu2dTvlR/QpI/Rg
/Roy/A+dfmRAL7HRmyA6V5+qehR9f4ju4M+NvAPgX/UbHCTkAcXQ4Hp64jrMN3Dz
RehzqRTNH9FPBEXJjEKORhzCEU78cLF3no5UB1fks3tsnlzqEkaPWS+etpVZ+UKZ
Ct3LXHMJk4itlPATH0JRDjRjllUcsIJnheHuKV5DIqmXAbgTk5xSgXsoj7soMUSY
Jd+4UJalx7ap15xmhGLIYG5BzKeGSg3tJ+ij1J4FaewFxkITZruOfO/V8A3Y2HFP
voCFK3sDLoG200jnKBUqFgNUFq7dzfDj/yr+Idwa6AaitPiHbfIU6GR2/vxSJL8G
HnDctjvs3K/GYpqXK1giFZtYedFAOiKvJmijTogTWdd7MYPr2T3BuuSBm5FmjLp6
zd0YBMSrWHav+czJ19hvc0RD8pJAXS0O+YTrc80+tFxJaQTVDo9lINbN07RxgGDK
EWDiHZMck7J57z1c7VsB+yztt1Oh9ejj0JssWzShUQI5gdi1PiCezZMrcxYFfIXz
9p1BZI2ssXPYvENx2JRumsNpEcvFSpSqk13lhSJC7mEeo39LoXmE/KQgA4KHF8VZ
fF3yWvzwtbaDubpZ+vwcmMWwBYO07kgObkbSxeg8rMT6Q9gQ+o802iH9nc1zDBw1
v6OuySct/DQz0NqSkPToZerGDzuGK7yGMbYBSmzyPTiN+n880aDvuxObkMgv4wfU
crXC7Dz3W2uA5mMflUnqI32CvJ948XrB/JIy/OH0hGz5gN8CY8SB5vhA9kgV0rwR
WhDyRfkh0MqKP1F+qCiN1tpawazRZWRrLfiaUJyqVIhjX23aA8cW/ovecKPif2Xz
0oexy9suplKBehhRFtdFLNNkRhr4w8OrEr0SCZID3mCEHTxbaFc0hz+NwAYEubhh
9WZVzzJ3wIFblz8rtajvqaOpamVXuVhggFw/eFIBA9YQOnOjwE/Ys/gfUsM5Fg/0
FI2CcqzlRxyPCpFrfcl2N9uS9AZt/v9T5o6gaOZ8he2qgr9HLUEctipc1iIbrfnz
YeaW0D8K/wLqmTazNyMT0JH1U3TmHsKeVNgFX+ws+i8yk/GpSuI8obJFoKrVsI2C
a+rwPvopc31S/AuWlkNPMcEhoTCJUHUQtV7etSOnUxmE15m1/ul0ykWnynIrD+M9
JFCA/GUWiCqTP12YSwz/3lU6ncVK9Zq1kjb+nBL0qMPNF8H7zgk5wym1Sz9t90h3
iq0h0MFB04yyp71gA2jmPsRUo4eqsTnGmsGdQFx7nFbvEbPwnaWAnvYJiHz34KR8
uB/FlkW+3ZlkvPPT2k0NdtnThA9kbpgPGqR7ECXmFzzbx7iCgizVkqEWz2NZiqUP
m40oJP4TX20dbhWxej/14CCkKliO9xH3w0g+tk+jvLGW/vPcBtlQvVw4uvvLubTS
o20szUShToVDKi1Vmxs61RKAQikmZaod+Oft9+1T9SV0NeTzVgkyos1q7q0fXyn/
J7dY4TvPvQ2FoMYv4hWhQ463/hQDg7R8MND3oIhVAvqK4fxw5pqo+O6Fb93F/w4+
6QfVXdgqtV0kIN1NKu2MDA0WfEZ7fxIf54NMcndrva0ko4NfxsbUGPtw9+27pJfq
vdzlpdD/EZG8OB3x1RGeiH4s0BHCEMsc1M+Rxnht2r/Cw9Y9qBGx7TWa/ExlrJte
WlB1Co9vlRNlsr1OMwPSokTIy4fKz+wsE6ZOu4f8Rv4oHvn4+akPycDw3Jfbw9vY
BAPWbUfo/LVf2qo7sjMXhpXVJR04ocgpYDTX+fvWs01o0eprA+Ya5r3OF4cPemlI
7DQC6qKNT/SjpCciMYW0wPUV72s7hbs0Vsw3K6fojxPLwxn1NBl91UtXMclR3+UG
OzqeutMb0XB3NUcQOvB8NRi3c72H4oB4AQ13ftkdqhNtq+Q1slru++FcGCI15sK2
kHsxg2AkNw5UtqOuHqnP1bZPCOhT8gmP+DHefpPGi+vDh/5C0rO6CkpOxFgQsiTe
UsfxLdB+tqOGqpGoIDgcT7HA97LNwnUXP7gxjxYJWhTak9PcN6Vk9Cj+6sFMaoYZ
iK4hpbK6iPJitq4dcJ94MTg9qcDVgC2fs4BJW7/1/pBOlAH5doraMwr6sANA2MBm
MzPayx1LE8L5c/ynjEAsVDN0GDaFBTT5adMb5fcVfCfbGIwNbcG3CBspQnZvYz2D
pO24JV32DakWX8FEPF5WvtgAvgKcfbyfMgLACchabUvA3THU0Vsq0h5oBs5Jkbvd
VejnN+KQABHf03n1v1fCV/jBtb1MvTYlIuZ0zqjh2lU89QKPXrUfsnl8ixbWZAwD
rVSypPlpmn+ibh5j01mmBLeSrzPxAkVEYOHpG0XQxSdJG4VIkR2BBuYerz67Gw+N
ueDHaO/xPzqfQiD1hOoHb8ckGCRphpwFqApTn/Px9dZWQ83EGjCCQRsdtbMddQdb
6iIREAHW5mEkbx46rwsLZGNZKBV3PQ8hz1ki6autGSj39h8qAc0E6+fjGmQzCyzP
sH6DZldu5LY0qhlD8LuzeGmpO64yk00TjX0gkHPKMjW3QxKAlNroXGr6Oo79c0Bp
dTUJUciQ5ehKjusiXjuhUMbzxyURLs0tExGCKu0CPgqUNO3Ak9/G2UY7O38Ab7eA
EdEW1RMth0xxuCPx+IiKEYPliac8m6pVRjmiOZNlk3sm5C06viV7JyxhtSkwM40c
tGXxvUNQnXoKAiYswv6U5eXLaVioWwatB/BPQYoyurQvH1Vc6dscJGFRjrEsjW8o
V27Sk6aKoGsCzGaI4PBKy5icFQa6NXBntqAcBAkSyC3lxlcNe/EvXqLUZx6bzMS7
5du47W8IzDPqwCQoBmmrppxgouF0wXGo1XtAuup7Y5H4ljWXJVx/KLedjKvejGgn
r7cOmpyKqpHzxVetQ05rfrPFJf+FFG6G77sQStLUCvsIhuXZ2/QN/s2tAN+pKK9J
f/AuEaj3NMtzmBlUkLLpp/Fd5Lgd4BaCC/HoAbAYH/CtS8BEBsAy+VEy48MjiHxe
PXUDLPg21/N5Ym6vDdNT2/XYpi1gdSd3XVEYmX4FpAlwme9f+BZMSI5vJUfbuktt
RPS0vyGcv6GoYxwLco+Tp9MbiSBNyDkKpExGLKjPsfZO3AZ8n6+uvEsToYAy6Rh2
JsFAqexrimDpXNMT/uMXEauBchLjXnPhVcQrfSe8ReC058jSuNRXQQCiQ1OAqckd
NG6qdBQwtaV6R1Ji1dyymcNX+u77/ibwh8n5yFndAF/Ch7U2XLZfr8JY+c2mNOBP
zQ/E9BlZhY7GZPYguexOHnned+oLXYB5ITsIBdfFc91eFl6M6dvfP5TKg+ZQSZc+
TL4NJYjK3oyHEIKOSxpd+QaSw9jUH4S2D+8UA5HoCW3ps6sNqlNRI+iEv3nvhK5x
KqUgtg1AupivcGADxgALPQwV+wMVQTG3vmwPdorRorqI70EQtjH+EyfEL0f7wBe0
53hkjE5yx0NWFef5xeoTtmyBFuTiqKiKHCMkHGfMd7Thf14tAYCErJwJ89MFBTEN
vR2zSEZXIGZuk+dAji8UKRvQqIdaowYqN2kMrIYdvZuTbOG9GKsWpnkuDXpR025y
5c1YKUwavhkCWPmX++vsiPgYXehc1dQIUGMJFlE+2QsELxYipW2MO5jKlYiA81Di
cYcOF+justuc3AtAMeWdOEG/Ok9YwI9uLeWVll3ij8aX1UI/G157vAirSkLaJiya
y37s4Qj6iOx/SZSiuVebIA2ldWgN7mcaNXbnBFpvBxm8ia4uNFFPYx8VnNnfMIk1
ds6aqI3XAXV4w2BAvwSEjdPn1+rAENkY5lfCqlV1HDXzLLWpxzHFPvbXwi+Igp5/
q7CCeerzYwfn5V1I8NNy+HiULi1MVL/Dz+lGIoGF1qOfyoh+S8kq107UZksG9B0C
SCbVhAkZFYwi1ONa5GIiqggPuoM0RfXwIxEosFiYnEkibZQ7jw6+v83zz9rnlkK9
LLDrkv4+jRChpWpM4G7gb0iT8AAT8PejyevOF69nrcVljAkFj3QKkWenCYJY+XMG
L1k0cn2JblHeDXQFGjbrtd2I0IgbaB9DIxvrm0oqyUwASp8HoAtld/OM9Kt58Bjd
Kkw2WSqSiXDruXTNYQYXf+T69/UEaATsBRIEfqKdsx+WT9wBtqBPcEODee6KSkmg
nmGuVfLqwf5XS0MTNCxrVuSW5a0Sy+ALbErc7HsaZ8Kvb69cJ3myNhIeWS3uF4DW
ddjyRDWNFQDxyClmseVPdgzd4hsivnUOLofsCpwm806Z0TTeaBZ5W6uOv/+fze97
2YaPi9E2oRuitdc4e/uiJcTUzK1TDujNMUR8CzmQqzFBUSSgPLgLJKe9ZSHTn2vi
UgsXeCP/gHIX8iBAer08mCv0CUZPICByJiHIpJNDeBPir4CdEuAeQLVj+CXJfyg3
OvuFKR7cPOxiIU3B4ZfOHVdoet6y+V3zeNA2b8myYlSd6uA7XAw4m+qixkV7eF/F
3i4Aa6Fnz1Oi/AbUnNbKYCx0Ngczv1B+izalmQ9vbnex++YdaSpwaVh4n9jFR2I3
mXpj9MMPry3lvIbdMUpD0H4jvQlSDwqCNCEgNY5Yt3HRS8DN7taf81gL1gKo15D0
BGuyB3v6CEzEqSjfuNphv1PUmsvd0npSKk1V7OfTliDD2P2FwexUGdAnXyHY9UqQ
bYFypvE9rksn1+ZvsZAXK3fiKxejMz7D/62sblD27x0W0xoS9pO1dCCw7k6Cd16g
EVZuHKbec45uMMYxW6HvR9PTCWvwL4q+irkqHWmG5OROeljBGbViv2pgHy8ZEeeZ
46di6C3M2P0A7bJHWxS0rfM+YLYiUvalukKm2uwL+4RQDdwfthjruoB+x9Jljolo
ztB5IzFcNsTG9C+bUO7kDXXZ3PfDPegowBrFCfJCdU9JGVMl8kU9elPlD0+0i+i7
PGnjwACtZKBavhSJo8hXjVX77mJ4DZdWAZ4c4cc+sp3bCAt0cWCJ67ccGjya7Qca
orU77q9/nC8IKjYv+t/jTKdAtKr8iKIBjVTMNvHb3tPSnlQklDee8tg1PTTuLlx9
7Bw6Wr7r362zUjTdgPDOdMvnmxoI+IjNLr4Ik8pz4CQ6QjimiiwD0v8X8eRE3dpl
EFGjlJi9G7LvuJ2D8ISbQu1PDH6dAzXwqTHdbgSBeWP0bR6BDe5zsY8tN+Xf5x+g
zl3O/vOmbnKcbMqejd7ioZpu8kcQjS7QA84McXrxgfHpYPItOx8CfYCvf3/DH7W1
x7vyAl+07xsh2+rAUKYxSHLdVyfIh+xvTVlJl/tLdohuLnpzQUv74wW8pj5310R7
1+2PX96HyqOrxpctC/nEtPqRBDJ9qDHCgU7DHfPUZo9uhPZHExB952aes8ZaJ2Cf
ulcXkje+K5u8MJyzwdn1YU1VfEjODrWkwfMNnF1SA4MelR/Y0BWme2E8qBw3qRMj
SkzNtJb4jqndEOYuVnS+fCXnTYgE87+ILIRrEDSEVRqE3lYhJ5m1uAz5FvfyOk/l
TDLgh2x0YkbIpikoudb6gRfhMc+/SQGh9bCAN54J+SEXqF+HBkrXyge7comWSdlv
S7OouFSA0947LZSEYgDBCx91rXM3zdVjOeLYQJ/0FRnm2zYKHyaFfyW1qcX/lcVD
yv/Gaji7Nh04ucSkse4QutokDZCX1ADB/8PYndUr3diUx993ZhcUcPSzQ+gLpB+D
WNOm8O98+FC5g9qg++MUWX/RZTdHZ3qv7rSo5AvBdE+0EQjnKucUamnUu89NNzX1
rkmrpM/Fdt8ALhGA38WxCNjCgqVZdJhYiyVhsdIf0a4fwSHZ1gU1a9wkbhvo76Ay
TwNipVVdRbBY4SlLFbJC+RbRSfeu6qQWneUf6lisK5qjYztpV7OtmrSQXWmv6pgX
gSHZByXBACoxWleXOvtpZe25Z3IIc3hT5qApGauG3yzz/4UVpR4oi+f1YxyWXHRP
wq0oPNkeaJiTVu9XJ8tRRS9m5bSDNv9Yl6I1JkMfQrRUf3kxJGOh1ObGelVTddjh
pabbhbgarL5Rcs7g3u9MhCvggRtY5I+5TQPNtHmKRmrdvgadJlqSKzpvei9BJtMa
XOZ2HX2UV/E7qpNdkpKlHgxLedWTki415ds8pDWjDToZTVRW9tH59BwDpR1S2Znc
ZyIjwQ8ZLM8+mpoXTOQV3/TRj+JEd4POHiAP1YgIkFlSYDzzOTnznSkdfEkguadu
WyTyAcoZfM5UWCKrYCChmGI+WOy1XVtQbzXaM4J+e87rcILydjXxGKuvIdfJckAq
b653iePDaDGX+pqogvI2jA/V2heGoSTxvUKvuzaJdBIzC8/mnD4G6WHrZW8r00KG
jhjld2fmhujw1p4rExgxc/N6nUopBZcQyk/qs8QunXEBGFwjnu/DW0PIzdqTqtYS
owRrMy9Pjmi6VXgbWI9kwTB4rRRc7m3eR52T+KuzhraMBj0zc+/Xaqgr12sJSrdo
awM/fCwCBnWJBgBtBXe5Fb8zyTiQLzM4uU8uU98NXNPLep6T1M5OGGgM87RByYDW
YbQN9puia0m/hsTW3P815Sq+O/L6DcAQv91O7Y+1JutCFRuAeW4jjx9b28AFnfly
nJBav5wapUYyT2kGMcHVXKvqrNZ/eUHlFsqkHHa3eYUGodmnb3cvxxUp7e7VbpTT
xWDnZ6+2Kyt1kkwkEZitQ4YWD97SrtDbS4a9WVHbnx5ffOW5PwGHhakJKW/DWlMJ
MepsRn0eXIhm0AYgWBvpSL2l3RZvmkNuQuAqFQbs3hPcQiQSpaaC1dJg0lgkWKzb
9mfqscJ5WLR5Q8ifusxbcmrtb5YjBDTTI0xApSXuQh1QWxP0FC10ijCSkjEm6hB1
QAUfI6oROTApqbBTiPOPEZneiTm4iwLksyajF49ZEfjEjKBzy3uqQ6oSbF00U+3C
Jj2PSEV6Y0A04PgLrgOAuFF4M5fr2HOfZg9e9ItU1F3/M2vaLBFwalmIRyuM8rT3
yx3IvWEzf9FJUImmopmMy3Vv4WKmzx1jeuVAO3jp4lLl3h7iaSDoLBHKyjwFOnDL
oAF4wrSc8t4oEuGAfTbStCh5swaz4blPHw0en18WLXQCEVI1e11a6AyfRvoPkXZD
EhpXRC16DgK1oXWDwqnFlgDhNMF2RlawQ8J7zgEdo41CPkDZiPFhFFfKBdbfAQcI
D1/FkAFoaypoeiff4vhOI94BuJMaLlnAiVIdsUSjAat/jhCIyBh5BpLx+jjOeqh0
qLKzLiKfZUtV6q2hlErzLJfXCsEqXyoAmg1TTgfpoMxR0wnlFsBxsgTHmD0XJL8D
opeuw9M1qn4GPtn9xWrZ3nSSQmJ9a0MHXRdJJ7FTpO3VToIDVv7UUNVq3ai/Y1wv
s+1QWjf9iMA8UoalYwy/z2qGaXSE7AfuvskKnb2vevdYfqY8VZTPJIsUMmw4+ZJY
2/u/pRFKta8/IP9F2pvy9UdJ5yVDTOJGMRvscL4o03NjscpFdmCcK1g5KbZ5A7+s
VCKR+UTqpHQOpdkD8pade+U7MEDtSY84aVq/2RD5RAmPLZVFMox1lKrLPziUXGzv
P4L5LD3WtBEfOI7DK58KH2/WWUID95ZaPJsXtYg41/8k3YeU5mrAHzhox/vTn+Wf
HtvFzpZsVNHSRLnDSouZ+HoEnz4oiL655OjmIaTMEjvshfSNzS8BQQ7eFHXqD1Xr
pThT/T2J5409+WH4Gv5h9aO6FBAKpLyo8XtQ1cpLWapBJznFaxUmTpC/KE3nt80M
Db5HrzalU+bju4c8+U+1aFUPKCIYnlXzUpYSX7a5c9QLJ8UP/5y0MCp9kBHnhmpn
YPOFc2FzdhFQSDlFnjYQkGuyOv78b9vLIqG8v6eLUQ83/UgU4HfUFEX5voINBndf
ibL9FbGzCJRbqGzdBCvTIKBTR7eNn790muzDOyS5zTA6PrYx31Lu561kAzXQdtts
u0H4EG4IAsTZL4ZzLaNJjFhb3PAQ1LQFfxF80vrr4omb9f2NT8VOxFcyT1O1LPyG
m9x9s7NhH1S0vkGgUHg6WmL/J5jaVGKY4iR2V+D3NE2cPcfnE3GqdNXT61l9skkH
+cuOVQis//t+f7RdlzsCOxGLDx7tBVpqD5clg1RK/AtNaG21YnumrUBq6bpJKpee
uUQqH0b0LNWDYGoexBcIBppe6hZnthOu3Jo3jNkJSnfqOILTzNo6z1Rp4GWbsOXq
QanXAKUjyPMQcgCnpEoU1F4DrTYfJFoKrB0O0IkprGxAyfnvSV5nTP7/HYyBHDly
C+rU8EQiPOh+L5KmIUA3ipIvambbfPzOYVtokWoHnQQA3gCCaACkOqPlIfyyRlkW
y8rd4CaIbjGNYxEFlKP1oo9JlCqXawXv1J5MoQg7qaOYvvRxpLKMFj+3Ic/nVwge
IoAse34e+lX1mGR1LAIKw3vxMSdvh76tgXrjosgPeaR/7xkGKmrze725kkJXU/iC
E9zI77ud8qkeyGBO+y55Fw8BL+EVjQy26nU8Pe63idzf7f19g+fepVNpLOCPcS9t
4O5x+9rMuZ/oezgnxhy8pjGYJAcfuLlKc3pN/AHkIC/Ht9qvfQa3YR9MuyXCRKDP
lynyFmwgyorA1lmg2oCEggwRV9i7zXJN9rpCPtRKxcfTnBaQhMIxLZnyLG/HVM3a
tVS1i5LuZ4c9+q+N0w7XLDwF6Pl8BztE60KJndJxtfqNjjXSE116ZxH9T+DHouBb
FqGMw2DQe5h5+75TPrIZz9QZ1btzpBMS+maH72BcotpFmzlnJPZX798QRt8fygBR
uBjsYLBoBai2hxu2mNLyNB5GRqFZGerSgoDS9rHiKkqp0aM7XCWkCSjZnzh6yuxh
2KZg5jRvMdKthvHODsYmO6y/L28uf8l/UB7b3kO2llhuHa9LMhz2G6k/YasQHjpw
DUE6BlrnrmTSV4CXeqmtP9dS00qc6PFA3tuCxnACa7eKr/U4BiBgL527wXfRzrjJ
JHeZXYjE85IfzxC5VDUYXS+JSKydWWPf6I9IrV4HWlKSi+EK2UXpPZ5JnwMm7jgS
OXjw6pTVLiGCh7Q7LzKbHZk4E5aNiEfunVKLsRSpjn4Tieh/Jez6vFuaapZSWNSw
aLxcWjjRRF7VbgYd7IV9XJm4QMpDzaq1cPrcJGZojygJ0zYdn3+oHfW1pPqQK2UV
stDfYCulMzB+b+GVeFLLCTRv49/J1TbXNcMXE2p4r/s/kiMY7eWnIjt9I6O26Q9H
qJsF4f0o9yOkKJ3JvU5DKe8MyTxc10iQy41Jkx9jZwuO4P71gvQ1m6qUxcf+ZhAQ
gwgvUvXouksbxJw6g8XPuoxe1YzC2AklTnzEdpvUlxeXtftLXVdQUhW91LrfqHiY
Dr2kg0afkbuIWSDfRLu72ZtkAFHv8EGhsRn1jyoDjsbXF72YddQMn79S/xAuawr6
2cq32EubpO8768PnP6IhKhFFP8UqJ487tDGf3JrjWZTqMggH/5stdzuyrVw1jUpP
nt0I7zg1d68Idtf4nP7XxQpdXU0u2lRiUBVlbnJl5xL2Bb7tX2yS2S1SiFVqOcqq
HOeqvQSPKHOU9SfrGDITQEKD3HQbAdrGl/qQAgrn4GGQMhkOePS3KvRYe00/75lD
3AY8xesRTKL8b+Pp9/eFl/hxA50LvN4sZF3Y24Rkkm2QkZYmgbAkU/u9ZgToHEIV
AIZnzvL6FyxUlTeejb/R7Bi8l+7iasHBsGaVBps9lc2N0F7hFD/dWnqj4Az4+xn4
iaM/mrvbhv3BoUJudc+NKAG6t0L4aA1HLhNBslq4zc7PR1vJ/4FQ7fT2oOYCNEd8
wzCLPWNICg1Xe2s8syZbBOd1zcabaCeIxOOwm9FbHHhS2uklMQTSi1ymF5VXqwQS
blqxOS5jFoxJ9wWvFDfA7mxjpRBVjq35lzVu2uKtCZYtltkwbXUSYmfJKwkacTAv
42rsY+hMQyImbBcqKB+JxmeiOW9v4A5spCgGtN92au7Kz6dcUXDKb79jup8NjRz6
ItwFco+P17MHFOsjKhYzbfUhXrjGCZ+uexdGoHdNxUTnvCiHkHA6LKPoNqr5Aqcd
t9oRMnMD/PsNi9jqgTOAArLZ1iHXUMj6gaFqRhILKvMoeDmPL+J2t/atVO49Oukf
iahjX/dlgkqU4yNHsE18IJYOZVbSNPT88kbbxyYH95ckm9y8MiHsJa26box4s0MX
f1vwxltoTFRrUrLKueJ0WsLW3EbGMdzwFu+BzFq+l4Y0EwZyNntJDVlZj9JVIWbs
9TacaifyMkpRqxv0O58IJl/YGvt7/jC0Ojsskznlq7NsAUe0DL4NcIhic+iW9EVV
Qr2O+UyEurtB8VhbMIFUc3jnWZG9NBKUCAUS/OHW/mV2jK0fhLom5BQRBpuwP5NR
NGzZy8p0hb/T2Z9De6YLc2NX3ZHot7ThBEVfeNUp8Za0rJy6d0nYXT/yr0RbAc96
hpWXDEYTE57fn0UOjilsocoLnX80+rm6Lxsv2CMCz7ILGM8fH69xaILeq8hs3ReO
sxiAV15XCzKr1dfvuUBR8u1L/bIyiUwx2L5UFzgJ/Zg9wL7nT6lqQL3j8YI/FcQV
fwm5z07Bsy8wZ1BBHPlnA2vEAOO8VbUjHl7LV7hISK9E1zM70hLCAm/8x02K8gGn
rd1FK2cb9lNLVp+t6jU5OFNEEjraI2bjLlE02DLjzNeNWCGdNYPtF2GVm9phTFju
++U8mcz/ijr2ENSt5AWg5Mwn0g/7fbhFX7tlXL1BvzNfUiVB8/D1LBEsdl3vilGy
eljS9CH1lfxJjATb97Om9nyfG5g7Jf6UIwjJp8Keu+vTr4ApbUTpchDUNwI3TXUk
UDvEcDn3en7OCB/tkRWwy6k8iRxxvWCiL782fZviRfildmKdd80X7ZFb5/T/siBH
Trg9Prcz4Btbwwh859WrdGfj89m4aHAVftxUMDo5lg2B4aWeH6H6C2kX5clxFpSx
fFgNXPiOEeuMtyavlxGLJU4qcQYJMXD/Qu6tKJqyQh9k+hla8jBFfbBxeJSVu76Z
fzZwYekHYoxmI6gcbCeEPYGgQ9bEDgvGwHxAk5EugugGMc06fghmmSjOZ7NFVrHZ
k2CGz/Lk40YrDYe1n8H3/ZrAqKaYZZnzyHtwExTGRtF8QOO00f7zJbRCP0e2ctxd
Css2c4cigdfaYXsHxsJE/p1V3uHgQ5JH4dtP0sax9EzCKJdh8/sknTBkvTPJ3Cni
Fw1dIot3QUh1CRFPM2ORzw/Q2jD3R5mXyy91Oqjp6BD19o0qNczFFucNee27umTl
c6e7mhTxwnHp0BwAK1P3ul5C2gXjMWzlJKgANI33PHZnmT9DiTqUjV/n2RZBLzpe
6+Rj0HDlzPm5p2nOF80hEiGtu0iuhlVZuCKo95vdgy9jqNfIcBJMfOC9gluhjzKR
KoUOiA5+Zp8n1zzsh+gI1p/SHFdSU6A9Wu/nUjQV5hDSdtBIXvIBuekl1//nM2GM
iE2SawCCXTeYHpvThBFbiywaWG6wXE8n2w34PRt8q3Mxz0qCihRNV1hZPKgooNmm
sNio7udR+oMaE3Qn4b9/sTJbG2eDBBuwoiDPWU+7K+ljQdTsLDWW/BN1ikzfPjhk
vJXf4WWUCU8o4Ihr1TP6AchbwHaMLEuM1WI9DDAc0vF2R08Xk+hu2fLxB0kEfS1D
zofCvpLCZkPyGH7dDAFzxywzZ1SH8ATuO4Si+dYMdx+aQVbVifsOFdWsKicReK7J
ZxAMH+BWFk2J52L/QBhAqCZhhWzlTUSIsaagp7znDyg7U6TkBPrcq0OSglNrc51S
hprQn4/im+FTLk/hRZzrLoJXFVrR8lStd279TLKhpMOTrs56n5vMg6F7kQAIBjlc
xeD4eJRSP5/5RerVHng2Jp3ICy1AbC3jNViSdHbHc/+TxWDpHQVu8s2dpyWg6SkA
uGBjYGkufJD2tcsK75MKaLvVw481Uj2cG2uco0Qhgbg3S+bX9utdOJ6SXZF+8HHf
TxuTvauIWzhAptYrGeeMn9LlxzcFvAeFzmWrqULIj1EUPsm6/yZvTfeQuaNzolpq
juKXF5A6z2rw/vOqROX9dqu0+P7mpkieXJY2pkcgHwnAV8Y5G7JEvUWROJpUuJLF
5Vq2isi6UFiemlueVW9wTMmW0GMsmjhQaLbYHypAi4Lo0JicuybmqaN+ClXw3h5G
uZqNnOWZxF8FlIdAvoGQevMuOuerSb0VmSamyH0SCJFhFZtLzJ6Xi2DQhLofpBPm
9EzJraErdVlEn0dh+UoHzP38o9FENJcEDFKErDQYZcp5PqAXdW5UjS68KIkBaCu8
cr7aGfxObKUVmeu+KzXHLo6bXRPIaX67/Dog619E+26rlqJZRtsqOZ3ziHdwrcy+
9g11bA5oQSENEGsTJDKiGSKhqROCEgkkmVH4szh/PglbPHhAuK/Zzpj5nrtWued4
D0OfiDHiLong6UmXSDIzkrSua3+6IrlgmcIx/8IKogKyif5+8ffADayzbyOOITu8
ag6CQPusCN1YCJ7GCULImj8Nj+If8I76TCHpZkwuKtTNzzLP4ml7XMQZ4Hy1Xan/
/+DV9LMkrVM59HNULGWWtf9l5opj2QYSQ6s+PODSQT01806lIwZeJPy5KRRmGNYs
1KvGDRlwCqumGUVEkpgbMRkq/AOzVLCD65rRTJJjcqH6NYKU5xUix+YZd9oGDdzU
PGIN0jW2lEHRG6kKDr/nJqKdDa4wE0N7zVfixNfSnzuAfzDxocrQfB4QlHWP8g8L
t7AMVCvkEfs5DpqWatOmwv2qI/hFbVa0x5i/QuQ2U4uvrOtKTZ0ECxELSrnyxHOG
pBPUSbiP/FWcgBaUcCE6ui7Vk+scT7QrxA+YmABFCLwuFMi/tTg3xZZjHAPicb/U
SY4+tIL8tI/7veXbRr0nMsaxIsU74c4x4T/STzPdzv1LK98wYLmfZAVdOUXM/wGp
H7HjM5SrlifB373U/rasbRFCDjy8uPf+R/UvCrYHoKhyqca+DZn3n9Ofey1b+rJ5
XQT0O0E+moK5tqzeRXEx6XknDfxTvulEE+CD3PjZ8gmJMWwgaGjmUVJHSM7FH2Tu
WbueOI7qitC19xmjByDIuOCA6i4zIJZR4zSWM5nMcTwaRsXpUdoK70ublGbhbLsx
5EvwnoHy3ZDbwBYNcG47BoLqj7GBCfA6e/ixlJ/RtevJYoe1RD87EshS3FLy2Ptq
PissGjRcFAkIFctXhP0IqHckBcHeXSJNETLpi+0hi2N1jBffL1X2lzfrNTA8HH2E
CbSZOTugoCvFYUAaYvPhfrqks+iGd4UNDPdvZ/DpVeg2mZB+jgJTEDIQ3FoqPYqj
62OM/v4n3NTfoNv1LDBXuFlFxbuontfczPx3W2FVeGbVSDbbDxGn0+VQClj7rT7w
RxnBmATy8C9T1S9IAFmVak0AGlbLy3gPqdGbUwUSdreKeT1DvB3+jS+YJJydklJh
uGF6/GuDvBBH16CROHtYr50FOYvgIvDK6jG0ltGGLqFjjFQbds2Y9tRh5tzUikzq
KhNR3yURCEGwG38KHD6ETQ/pdvSJUsM7WnxoVfoRFbAGsjJf3xNcV+wUYUHU5bu3
GayYjbaEGFeQL3TPC6hFOLS6OQkKz3u8+pJUygkbBS8fMQm/h1rnxfz6iOFB9iwa
Y8kBV0xp6KSZpCoo6HCZFxqg1kMY9ClIr2EF44tGOo+5Kj8FQL+did4bbteQ8Rd2
Y9nhA3sSZv3h96snP3ryiHPXjyRJ8GewCKmTR6Avr5wOuWXa0y/uqPWBfljOSJc4
vFqbYF2INsquB9PIy4h8mqDOJsS9U5wFjnD7JWyRJbWNntXSl13t9Znl3mmrME2j
vfJw9vPhKKFIASbYglkfTgBDxfu3Nqk9mRdjvMfs8UcqlFXNAibfS7pdSS2vVwhE
+yOzeCCrzJzp8f4mtGT39E1fYg51phZkXq8A3VuLtuHYh/tYf8gT3f/eWOOiN7sU
mohKJ4cMs+QdQrsyc2ZwdH+sO7E6akgn9CqvlLk4OwL27NuVTcZHAVZCj/2XvpIE
IDMFDk3ZzLRiPW8PItAG74epToDAXLT4Snkgb5mUIgUvi63MOfM8btmOToMFtwB1
PEA92BDwxjKRXgydSJBX8y6t8stK5PZzlA2fePLI9i8GXmp8mWn7elel7/HQDq0n
R4AC/Vc2FGDil5zoB6M2F0zCYFXsQUD09dS36pmpmeZJD/VxRJUMs4u37V70P6YF
XFKPsh3tutyVGYUV3TYbrvxsH5vlXtUAKF4CVDe9zLRLvxnmW8/NcyIp77OwEy9S
kfwLmw30w53WrZTvFB9j6nm2f5wc7W13T8q26/eJ1rlAvhbnd9pbFZdYG4tiCVn4
WbNnOe86j2zcDnZdX0vd8XZBMV3MvkKKRgO68XHYaL45AAbMvmulsOIwrAe4Ns/n
bOp44SpI/ALYw1XVQRvkKlvmvVlUWA6A9qU9luA/5VsaZofUcBoRFxtgyah7XZP8
ippn53W+0KAQ3+wdX2ReMhQTEMdVInhAqgkhLNhYsWcINQ0O9HzYU5/+sDkytOmK
wujbXWkBdvyyKL/GxxIy9BzKMxxK/b0pSRD32ab7HC7/rxY35RuatNqYVhYFpVw+
fLq1oQFr23bR9QO1kpn+OsRhxkE5yj0DJINnQBdPPf/gM9GaBGxXgwMtA6jIbMX9
xkn5H0S0T51+EC11MVcO7h1ICJvhomHO9Hf6vdUMlbNW56INWpUZyRJtX8WU/LNP
lEGm8riWSPJbOpt5UKJqlMAwxtriuALPEITXiGg3fQVnZqdESkwqNhN0x6w/ubI0
JTv5AmzmZGWh0IIb3Hp0I8kGuAt5U0M3jPhjIzS5vL/Sh1bSQ29FgwF4Rj0RblBW
iujo0lyvxU11ZFqRljKJJ3ZwYJZl8jPHji31Aa4nAxdz6T/6Hs/hFKnUZf/qbWEj
8VdcGCD8/RalFuEk2wuTaZ9PwA9ALrZ+J//IUQBRqtULCExgaTbUZqL1CG1tBfAE
8M6achFWRbfLJdXtGC4QameRsf64quJQhx4UMGO6tMWVjdvW40GCyyWTSIWCYvk4
7YUAFQQS59rzg6iwzZTRaQWKW+3o0pUVnopn65oWGqfbQSgHv+XhbUm8pa5nDddZ
Y1r2YKJrIKZQh+IRwkyOISpTO/xJTrffw72WOQFs/0tIc7sJ2bvH7iQLl6nhz39V
j+YzWJ7kdTWEV4E030w6H/3bPHncGVarAtkWh5/Tlbs/mPvLtjkQxg1fn9xumnwp
J8D3UgNTKyT72nyCV6o4boea16WN0fm1VGH0LDCjKTNvUMadEBBNbFFIzjEoRk2f
JedeK/WOPIkvA7FqCbJ+JbedIfLEy2eQdfqn3ESlbE9wJb53gI63zCjV3UyJDnzr
p2Pg0/Qh+CgV0jC0URl5gD4QGHfbH5EONo4WsIlb/ThixhYx0H9OiOl4ZDqnrgMC
eJIk72QiN1yXwrNg4Z20lMhd36j4Ns7O+bh0+li7q9gzCBSML/Y1riff479geoqa
2wddbRW9LvvGZORHncpjgCStuhY0YFH6uy4yURDxKq7KCW0oyoQzNBKAjgYYtuJc
CSuZt0dhwgUnTApMSv7I4LK7oKcBng1rUj1ALKJ+lvChOfFSBBtmZiIyyfq4/54G
vxx6fG8hk/+d2dj+bmMpoYOqu0QpfTcSp3fXo+/ktZt0GUDEPoqBsHUePWrAoEJC
h/NO+GSHKCL59KXgmcgaL/wwMwYGS6bhFWV+CTkSflYjXtidXF4ehHey8hWy8Bpm
ExKeQDkCwiZcFoX1N6QM6nNCUSZq5LK1YPm+IwGOoYLpp8j85e0ZqMk+1fbmL2EW
jgfzAvMm1X85pZ+DSKhjeRaQisOrEtSHdn5DCFI4apkO8guf9T3yeIm+EZiRTmSA
wsREaSg/cGDN6UQSntMbxGLqSJV+7V1kcWaCvw068oIAG2OBiZp81552HvXLrWwo
2C2fgr5DSUelsAQ2iFX0uAR/GqoUiiIlJcEaXF8eEGvlh9mK42ibDEEfu0Odur+T
qXAJSsAQJa/4+u/a8FtjXNrfm3HZ2szKKetYLaQRyTqxprtTRhO0yXA5h/EsawWo
YJHysRTaFzRhlMRuWbZmU6z272rzalGscJlmhnsWcmVHcGae56c4g0e6efWLvd0L
tCo/HEBvhYhmMZglwHjtB3DSNQuCo0kckC+CpscDpRof3kYJ331l+M0V0YiPQ2M6
5x28KfdWdZC1B5awcl/w2oGdS51fptWbs41fvQt/lIVhzV8JUiA9IbBaLsqxKoT/
oYun+K433PWEOTgy9uikdwKl29i30ts/6uE/u8AicO6y4uTSfznxlZznBdzz/ywt
0XWsruK8WQjC2hfgKYjqTTuCuaNQ6RSQ+nDKo+2iJ6hEm88SWaf/rtI6gNuD1nxw
Xs1a4dZcO7FXO45RqxbAx6/G6V0FNQvx0zwVMPaP8JFz7MrLjIXzSYesM87oEi1b
g0Nj2DaG2MRM5+bp24IFPHaWB6yB3zybv9GNYBHS4KBXF2SNynxS7B//voBlOoJv
h8cI4XcdPT71hTPQjfpSSwTefPkUooXhnK70V2LlKlfIwtlxnNf/h4QSbA/bvGfT
l2yf7PbTd/f5yEDWBzBI/hyKJSVu+2Ih39+kJJorWkaGGLu6rnBaTA5f+bnEX444
21kleAAy343y0/jMLMHF3chDVq85qsE9dASYmXFMTPE95e+w6bKsXfOL+zRNTt+R
q1nDNSkjLH/wj0hnz722S4vBYoTKwYGhQxnHaBQs+49MOIMLZ81cWFYBb2iW1GN3
H5xO4fdzWHcBYwSbDzzL9eZZY9TU08cK4SMMGpfeZ0g7jNCfjvatvRtDPR3S9hji
T0z597oc2SWr7OEoykbIDSI5gd2CFo7YZIbWu8BsrDlIGDi/nV41KaO172WlzcJb
OCVgnYnySzjPkEb8YCpIIq4T9iDT17lxtap2qjr0yrGejTRIaHGMri21uS5uLZpw
r0XMwxMuD+GwNlFHkcUIxRbk/jhb/B0bvv8y8K9M0pqOIQOLVbRu801yHe5QYpoi
vdIba5lMfjljEcvsFmfnKCBD3BQ2zL/5iJaazP8YCiB8ahdWZkly7g9Jc5/5WFy1
WqSLSxugp2og72LEGlvtji9YyHMU80D+4EIANkBvACIwVJJI7I46mFBzEmC+Lgne
ea7wdEl7qep7TmACFXK4DWjbxYgg7iZLwBQGOem4vO0EdmsV8xw4s74aHCHyhmK9
HFQOPxINMdiK1aTAcSDuZztfN5BCoe137hf6EhYeyTCBihaS9OQMvidKt4bUw6pI
5qvZT5a0k+CMYK6pdt/fqLts3U8VpzUtQIE+IbhShep5Ps6oyHAl/52JrEi2P8Jq
uBvGKD/ilIfYzIgTYcahDwalVUYl9aK3E37a4+bouAqkg5c4u0TQB8ImsBhvIOeE
wRdRQbi2Um2e/Los6mFEaJzSAUC+ITs2lBKudj78cANnC+yE/XfCxMnaeZkfBpDV
Tvf98hBRb/83OUGAhlEJvtXgZzz1SFxyky9k2LTx1OPQDCGrmA/zssbjxrQ123qA
pvypGK4i0Y3BcHPa0r9BRtBjor1WT63p0YGYgI7F6rWteUdyw99gjV/XeE4kIdg6
QdWzmAjTCHFYs3V/72xmoMMc8sTQcuGeqig+UTwPQSBL0BR/hBANOBQ9m1fFtiWq
+EkBj4+OP79z+BNOepy/wqCJj5wcVSY3M6H0DGUHbP8PNRBblTs4S/+wpMJANxSX
mzIaiiJs39fqbfF2JgHU95gmYeuOq2RAbyXMVURc+HA1p2GEPrClXT/jlhR0QMtq
uPcVNQDELaDpa/LdCmeSdgKLD7/dY8nP+KWjdj7SwD/aMxaeqJekEDSUt19FuNiA
GB4bJ9SslO6CsP5FwXy2FvOlIYhGgRUb6dkxuaLDvycM2KjrhZlEZH9efJ4SHQyC
RTwy2A/p03kKtsYH0i/DgJm62L57G9YCWvgib3NLDMFFjXgJigWfKrpX7TJLN/5G
cHa6fw2CDAz2oMZ+ohxxrlOnetqBD5G9iuh+vZ21khVbseQGFU+9mq01k80A8p0m
RuYflTBHxnpRQh20XD4fqMp1r24OSQ0OTcSw36cNflYFuxHCTULb/Df2/eg40pFD
FSpMsu+x6WjvZHj4rUnynOheano+nT9g52ytYpD3kXTbKohYR0v+Ig45ixc/F6qv
K0rSNSiWDNisOx3Y8TEd1LXGsw9vFWL5Q9pGDCesgY2utyezJa9/caTMjWHrolrA
hfBp+d8rkyrgGTuFA3AMzJqycIa8hBHcPKHOtTJ1CE0otcbr0fB112CSQ6ysxEu0
3+E3URX1/sTng8Hmwnre19Dc2AqrCt5pBY2V8kqAPAehUoKVt/vOeoVsLO2IXk4F
DPlfN14WW+Imwih9ex5MqC1NOblpCMf3KAxhRSqxiDbuRP9qJYUmJFHtp5KSSlWt
tmQb96wT43fOiOuOxGpig4P76ZVGbJYqwXXH2FwGA0Fo1UgjYPUzULQwV7ECq1fa
Iaip1r8eO2nl6U9aZZYgtB3d5EXpD1Hjrmk5tJ4I5YoGjKDXJPE4PF4oXC/ps4AB
6SPsz/07hfegZ4hGHsptSW5UdMKq5POABJRvU6dC/kwNuL4nUALeddUFcm5swhZi
O5k6W6gtxXd+ZuoYrdhENaKtFtVOTo1RTsypU0uc7BIzK2v5OboJystH4wKTPZgH
rsV4vAgTOT8FJZUmsgZ4fkks3HGSn3YYJcdQ4gTwieY4IpYU787HHQ/CUH1f0TTi
eSt7j75Ikd+K13TVkCJ2/9LX+KM4X4R+3Yzk80kis5fpSRXa9e7GWLT9t2LezmJ8
qvLxxYwcyRAvrLbg0uOWxpbBAP6eSPugdwc4LuVTI92L9iblHrwcYsgoDZBY1oxS
MQ2g6AMsNa/YYWk5F2q+hkoHsZEN+IXYqUG8ht3tOgqP1Gg8N0uLEQy1a/htlfh8
Q0/f0X0NE6z9YdTPta1322DfhcrjeK103DlO/DpDvTE3P954Z2/xs0Z8DV0rpLu/
1xmJIn5UdmEgLJD1Y+VPnPXhJejRlhKtQaKDuT7t0pfFm2nr2J9HD5V9Z0JGi7Yj
Y8+RPTwweTk2GfBYSN+upVcKwNOV6q7/AV88VisY3EvLYvXqFvxZiGaI9dy2jjPH
tolkJh3w2dm4kb7w7ZVvykhRyRnAiXuWm0TOkbWmSe2xJDk94FoYQZ6ICY+E1zEf
0h25uhlnNfCM85gjMGjHsS5UHFKVt2tYmgATQer2UF81DAhBbYUZZlcG8Qcq4lSD
oHF/sfLxla0VGYqu0PbzFjm9Lorn5y5gSojD0Xosb+X22oaASfPLkrP38at5teeQ
KAemzVPThV2mkATzwp9GK2NGkPR9N/EDSdY9jbnBMjlKRNQ9pZdab3XatqxM7NUZ
xXdK1FoUxkQDGlj5ssX/QPhIeyp4cS/zDAU3IQRqQ6CSoYKgKrMtBLp6j+4Pw2bb
CjQcBoKdg9lsE8Fx0CjYs3xIBRQWghKwJwUFa1zsTJiMmaGF5SLYdIovTneI4MX9
gbIo1V80p0FMYaHBnChI2OaM7nkyproDbdKuuYa1Nu5xIzujETX017Hg3TIklZqV
4DBv53mr7O2XvFyTXW3yH8Xvr8ryYgCKaJArjwwnVKOEo8tq2jtvmqJbYxdq4Wxt
1ueGbnCZkLmUGm6zGLhtiS5o9uMUwh/KRfKGuD5DSolRswzqIZxxeXF6AcLMXW7F
tWeh9xF2rOykA8xN7o4eBUoLCAq43/IA27lUNzYaSwOcZZhDzKawOrfJx+HessjI
mBKSgebfqRUp/cEPCRA7gIY3RcKh8i3OL//xOxBGEqAMDW3h5sFQW2idpQBboy8m
32zwHr/8ClVclRVP5g9WsrRopkNkMKbhS4dtzsKyQSFW/WSugPbe+MrFUGqg0Fw/
vnE+GOhlLEIHETnHAN4lorlFK+EMaDJyThxgAlOHyoQ8WZ82zwAjsJU2iKng7FCd
oVns9z4ESCNcU0ru1B83QmPy1tV6PF+PoK7Fwypjiv+S1VX8uMdMQLj+x+KatXiX
qZmrjTHJZS5tojC4XbgqFTNtXyE78sJVzWItsi4rvX+AsIlucDrLye1GUB/P15Et
jhQGqpIjG5oqwPEuWG04ZmlUn9O2dIRupaBwhK1aDYPn7ePj56+YOUxbDkVuqe6F
8AAcvnj/UpRiiBtFmy6eOAeFO0Erp1vzAF3xofYqb9RQVeELvoYIfOXuui0IseAK
u64T1PZYjgHO78ckC2P9xLt4rNw6tfeHf4DuUXQdgXQpeTt1mkcdDjO9JTk+vOZD
qh7VGdsSNdMPrHAvWYa+QhAE6RpOSlZm5sjtR1LXLKv1nxiShzTrRZec/Edc+DNC
Wgif1eZ9w/dizx/ZZbQPUI9G0G/34cFHWzK/BLVQZLwy9DOzbAvTb5eeFuvvkx/K
zFPTKD4vPu8KvqojiwI/QFHYv1GHZHhkGyFjwyqTpIeTWamGmYL/R3zpijOcUam+
K8LIaOPvTTqzx2WG1DuhUS+NgLFZa/rXF1+nk1V7VN3HK0KFxf9fcEcAbdEewWJ5
L9Nh11wp200sMyEjiRbVv6ifij06CESlcrkANQZ9PCOHARjjjxSoPeuj4jxoXcEd
qhk+ecKT+pYoc4sFw0/wWd/NSoHp5M7+1r1eGxw7WsaipNOk6euRX1FPWSf5Ofym
xFORaCLNGhTrWfjkGRPfh9HCArxo9dvufkmtqAHRMCzKcw5ZMLUvfEYRf4GL5oIp
7KP1mGrYn8qDgfwy+A16qP96g85qR2243AZUXNQGSjFq/5xTwz6qdrCTlfuXOjVf
nbaeg+PsNKrEqpO+gk4EUTI4Bun/DCwnqakUHtAS4d8WQuW9KOdBu6H0tzStV+L+
IM2YxFDgFT3FWZtapDtx19NcA5kco9LvNS1MMEN7dz1/GELpBBQuZxZHoCnf1/fM
18HdaWItkroUEhUHWe0Ita3qzX89xo5hQNkk7bb/oKpPZZrb5bDWvXaMRTTlymY1
hoRTFGDe/2QdviU2tvtfUnP74UYgTWSky7V9Xf3eNSeulhq2pTVBkN7HV6jqb5zx
+A15k2HRpUOAqlf7MUV8qhdyoaiDMCN+MD9CNz7BZdMa3EdIPTJVcVL3yEyt1jx0
hHJ43wo7QB9wqfMaF8N1o0bb7o+pPuTOESylGBSqJexKEf6YCgwV1Hpspo3+Bgvv
fiq7R9KEOUDc5enpnfErgqNUlrZwDC25teKTtv+z+/K/esRNoo0rl2uHoUxul5mv
FFKqKeF3B7tDuo0LcdnKwgwhGA74cwIivyzgJHR8Lv5fnl1ZcF162fx+OqgtP+p0
0WJn/dIkTjtCO5PUax0YAt1Mkef4BSCd7gfwJtuq5SEnebHr+b5Q05Ct/7N6xXt1
R0QrwuNJzXre661AaH1BzTiAybifStHdOrhN3T1xzbxR5MxE0SRHBpXhrw/dZZ9T
ttRtthB79OCHLc6wm0Si4GCZKT49uu68MTBft1M6HxA2xZbKAR+TyZXvM499/ejw
HGQRBbUXnXN9T5oFvl6TJ4VVj/PwqqZn7JyQY+zVEWlHGPPIZkRkqWzb5zf8nJN/
ioURjWLu8QASS/6hV1UrGBKuxcUX8FGo6Z1unNXSIl1fp7Q4AqRARp0zWo79KD5m
tmj7AMYgU/jrcb6DtQ6gVoVg8pQGU/fOwA4XwwZHxdHnfzn3dRB35N+tZfu1QTq1
Upjh3HgW2O7sJogiUrA0srqgn9VcZ04DnLwzASNixlKHemQNJZMrl3expzE6XwdW
hOJBAhETcxwy60reKhMeNXbUzDxUoaIlUtEmhua3EkN8g6Pp9egk0KBaY9YfDwS3
wt/hiPvimLob9I9hgy4dmIF1rW5884EDPaqQ6Shpv3uxa+FRJ49hlHQ01hGD+T0L
o3utLzbfa5b9e3dMnWRHxZItvlujfane7pc/sK3kab1tgGh9tXw1yE8ZwxwNqC8A
ceo8E+7YJF0yjBVYg+zZ5SH1jNIVMrnmOpNVS5Emodz20UBFGLQvdG6jCBVumvGM
gtDTzAKIVUDrmI0mj5U9vwns/Ts//FGhKuwZh8sG4NRZ06CIVnLrdvobOnr4BOQG
Om9ZM3ozGEmXMQLXVvMiHzj+bJb4mAGq8BHA4zyyBHXBIxcTvWNXL0c1YwSY42AU
0871HVCEKWDiGfIUhR8rN39JUFvfV2nsiBxCYhdQs5IjjWebFA1X+5ygyGzFOabi
OkJXUN8lemQfEvsjbvuqABtlPSmfn2lLRuFlS008Va28N1waZ98qeKKHT7DrtLFw
glUaZlBCwKAqJlU4JlYlwxBJRhbHhRtNs7MCnul9fZCT1mobaO/hJjJDlCDCYgHx
TKxxjbjvRxRB8atKMdymrVZ0jAhJ+q/StSdW58UCXCrHKWz2o7nfrV0K/8A134Td
QI3J6eiB6PPk523dBhoMRJwnCqTWsZZmMzBp8YHpDupXua7rzW75kH2qwpRYydDv
is5ty1iqdlrWtNrT5cyBiZEbRnJ8DiLvFyPJffJlR0IyIwenCh/hkxZaaV5H8E5E
IYlKulH3c1VImsuR4OYxPIGUPknQp9SeHbIfnrL+rK7I5E0BHsaQURojcqLwLfeV
zU9/tbuGTS/7Rm5oteHcTvld66wsucEFEqQIvDPsHUum0hl31pv5sdHzJDch3g7n
NXNWQJuoJtQZfsHFAdPranCb8oIVhkBR5MSU7k8qahGXXbitVjXLBRGviTDUmbH8
qg3hgkzcrTn/FLC0AeQGX8BBpCPfsEYOlEGnq2L0dtA0K9YUcFmBhLb+0CXZwJCj
a0PJd12nQ68j4AN+6ypCsPNaaegDFnktevQWi50dbwrPTXVCPavo6FWNHTdPqieY
aj5/62q6QVClj/+uDKgIpkvAEpCuWjoccWjYV7C/zECKrZbwWaaVzI5SPDIH1rnk
ocScjV+Z+psEg6aBmrKyZzhuxBJZduB+nJLPH7QpKf20xHjM3hnOqMwCuWgsPTPm
jcBwSl6lA0nqPYfe7PQF+nT6FtOx5FnaHqaPBdwYGMmCHkOIt2f8DP8nfDES72do
7tnXHbpup+WJlJaBunW+W+yiSeYdqOUvdLuEHmXPf9QCvpqFo1tuQdH8vMIjr90B
1Cq05DOyj959+KiNqd0jVnun0O1VDySS5s2BoEfT1sKvLLzFDVz1Z3xPuqcYuhYe
kC1CJzoY5eEXHHfc6QBaetitdqZIhKCG5sLZjmV4ntolP4ZAzB7yN7CILT5A6JP+
LYkkXDb5lQpAyD8s1mKOnyiQbQzVCBLLeix5ssas0dna135vXj6syRXDbMd8Em1U
m6dpvmZHs2zcSQipYyEoWVPYICwv2cgAktecerywNu+FbmQXI7cP8PIzIx4/0Yln
BrbGNt50s8amroZDYiMjTGUsVNckWJ8TYygnl3r2FOtNkz/sUqv5ZqMhBxvsSGrM
PF24s22RooOfrz/EgpdDrYwIw1BVOwImCnlV82yeKbfgKd08mtC2J9OoqlXelBfd
Uer1y+CJUkGhTxVJykL1K2N7M0e10/p+jP2/cSHm9sHEmhi8Gw4fPl+6OUwCi0Io
sf0pxufubG2Xoq1nsyMDJ/NbbQ37O0RCIsfJpdfujBWwp6SpV4e7VxuIvGiwTEoy
lNbCGDtJ7nqI8SQr1QITHoOk6RQT++DYegSU3Sz2R4Z+GikxkbuMAup+biNzIZv1
ieVN/9Ouk/Nr9WmFgeg2cxiKGBQNC+RH7FhJHZgAsFa6lhSHXVKDQ9kDBFm3ySJi
fUHeVKERnTAHZ8OlUaj/W6i5sRfeBYsi972HAUYXMWB4Z74fuqFm9v6l8ZRwo6eU
VjhYI2IwVocFFXsZTZv4V4XxLUamP9PYYB85mKfcvuydFf9AvcsJgu/O4Us1zW/I
jB/6Xf1QYqfxAjEI5U7aBP0tQlARFkp81Fztb946r4hVObIcMJhp7tVpv/0+7Ef1
BkynZJey+FxH5keuzKkTYaJ7BVnA2eXH8bMpWdD1J6f2Bwq4muUDpYKpxdJD0Mkc
RPAAhrox8ueB98Wt78AecsE3M9rL4/vzwSFGTHdmZPZgX9ZaeWEwTvEbUyUl9cUn
f/Sz87RQP2mSjexkPk/tjR4DYdt6ZxPgNZzVv9r1U/9S31kMsJGwrZOgUx9X16aV
hddjYFyb28i2i6ONa9an/00nyxroiAs/LZij4Qer7/Ds9QNvI8vsbwVZC7D3go6n
MKLxnhnlrLGHgoGEKqcJtYfEYJ8DDDB/XBjzmqyJOTKVo+cUAdxpEmSOT+EXpHjD
i4Y2R0+iMY/A7OuZuKwzvuWg01alGJyH80WhlTLpwyKbWpYkoG91rmBGzxYOHKgD
m/ZMfyMDa+bd8FkBd0uc7K8Ix5fJc017bjHBjhxK+kcS3lboiBEfNb/Bqn0wss14
p6V7bFhmiNZjJiLWM6SuOoJf7LWsMie9PvTUoOkjxxe5gdYcLsTE79/m+7F7KiZf
Xoh8sZpKpsCaA3Vzrmo6ltnfxj9dkeuffH/GdjgFmv4eblDwNU0qhKCXs4JFTpsT
/KhuRitdRUeGTTDVbMj3Ntz3x9MgMvrf5t0BgiUP3SwlgyoPajg2372hRPfrNtUp
NFzUrgPrbAEH5n65HtmDS0WRBpdpqng29VvdyOnC+WuVw5/cJ82PV7s8bRgaQL9a
vDglHlMANyUx+j4G66pFtID9M2szr7Aa4wE9EN4orP5S0G+XwJ5/k4cjxRgHFfXN
QAzrA3cCeientcDs/zUIPv060YMOF3Zh2r7og+Sr+rd0+OtYjINNvyPqu+VBHZYb
XcxycLHVCVcW30L82PbMVVh7mHrOoi8bl5PErEOHR5TqEw9C+d6SpEodDSZf2zOB
HsFMFCW30bdxcDS3hw2ShXaQL0Gw4WMCYZoxwmbDY2dX1BJOuXNT89SZyiTLnIlo
2m3ioZPW9YOFdSmhCv7gVTpvypdbJRH9OxwmXSoICM5fccZGvXpSgSKE6mJDGUET
h6vF0/x9R5p8he5OXT2lujqrgnLK541Co6+SI/ox+g8Lg+5/f7DFOULAFTpTuLpH
FHxjhGG7GEqMo9XfFGuAIHyaCY8QgTTyPw9BKrHWNVJMmNeXZImWRYscFzaFNpxH
OhWLiQS0hus4RlpvNuGfO1TpYmQWMzFNsxVMIVIW8AFxEbXmuiUJ1QxUu2m4BZTc
p7CfUCglQ7dsWXpuyY7FjcSOvUmJCApLaVq/4CCQoMqO89315OXfV+hrM8l9v0m0
PKcNzpAZaMfE2NQCHd8YkDj1FIdbcF2dA1qtMviM8wLz/ShDXMxUqWIvNGsLMJ4z
MW6rheBW4f45k/8mRjJzoOESiJnSPK9TM14c7VX3Mg8HG9N1VWX6Qjsq4VH3OaFx
A1pI0tFNBvHulPmx3YQnQ797tpHj7CGkFwUPfUq4TJqRKivrv8i8jXLP9krMZxUp
cHb76+hUcbAoJ6EZm9q+6k7k7WsabBsUhnczOGvaSMl6Gdhu1QnBbKzEo2nxHPHu
ZoQ4MXkptNZoK4bn7UjwLWTKeM9kaZBwlAz4yi0r4FU9lddJeL2vbdXozDIJWuQs
7DX81nA6TjKUWfjWcwZv9N0MI0UUe6RSm1PAtRTy9NGCYNN4Qe41ifHF+OaEU8dd
+/I+ha1Ve2SBnbQUGIFV91y3b8LbvTKIp3M9KH11A+90vFEh6xvQaAxILiP0t4K5
JLecL+G6K3rREzNPY7HUOJn7TB/nqowSvGOQRlgLNDB11rIwzUo2Al9g7m2V0tdz
PCc5fYM2brgHjVKFFnAontBFjrO5fWIhg0HmyL95kDkugDPENdb/mX0bXo8rIHc/
EgKec5hEIq6U429VO8Q7uVjH/9z8SBJizzf5KTHsd4i9CwF2FW2LNxKflaIdKNMR
pkiKI35WgZzPLpFjzA90f8n058p7NfZr+oWU88TQygLbg9TooEyIz0XUUHb4cClV
+Bqr7XBorvkRENHAxPkvqWs8O+V5g2exMBdceefMJvI5P0XNRDJhmX1pYBP3Mekd
t9ptYqd8H1XXkQ5VpZsBigg9C3rP+WQdc5iRpMCpx3oEtGJqCcxiuK5Lh7vAJJEo
0fN0UxKktaiq5bixBKGqvOSsdyDPjEcetLr29tefg4ks0BluBol8pZGIyvcTEzHN
Gye+cUTA/ozxPvstWgw7dYjAKwgrZ0+ELCVqFyfDHU0+W3+y3xgLfJCM7AgMJ3WM
GBcCXtDS3q8XrC/iphdH91ItS58VINpDPENQZz4xJf/SJYWZ9yeEKVvJJAGKsm6d
sUYvKkX3+yjC2r7jEiw6bOQ9cgcxsmp8adzoypyvVOk1/xkvmWtN0w9Kn58b6dem
T6AzkGSdMn4NWJ6atRN7aPZJ3Wkdrrv+6XEg/9Zd7WB9rq2oJuCltEgS3WwKZF/B
3N9eK+7Y+Zp7CCs7899C9MiWnIOTlLD9FkXrQ3IcoCVIZVqsG5fPo79PO8adZe7k
suraF+GYjeri9VGY1PJEiasHkdAoWbzD3Tw4qUkA2yUA5h7dJxE8VWWLC0j+X9Cp
ZrA1mq0cWSXHPFeoX6w0TqgaGKfT9/7OogrzTBxAsq5d78G7tMAGdVM04EHsh3iH
j7gnT1hs02PHpl1o6+SgkO7rD2uYIPmJVIf8WIIWg/eL/BMqYkToEUPEISutOols
pN7fHaBMxR6HivoxnpY/8nC7oE60ddjk7mMX9+vIR3ltzTcTWROf4yQnMOcrAGsa
Lx0G5C9UnSZ4uE/gJKttynDdE6qEUd2pzZcTolc5r39ZsO9p6sqNF1RwD9ZMYakH
p1b7essnu7dhg3NHjKsCmnt2ZbVYnvrtetznLEusgRGvg8eIvpCDO2XlcQn2aGMQ
aHH0lDN1EdHWO9ITJGBMxk4k381CzTimvGZT8o9Ls5y2QPGzB29fKxU3yHyxdqgP
AJu4MjrVLp7G4QCPB7nNbkj8gyRAEYxFb7joadYX7p96ccaWZuq+TZ//iv8f0cu2
bGhzyz3b5Wvgc6FRe0DkCKo8XU1ENU2QDbdp4EUl6jgMfqWpUHeUovjA/USVIXsa
dFYhNhWuf02bWUleuHVUeiR9g+/PmY5d/nx4mPHtpyNViVaFnUBbzICIhCwNeWb1
BfOSC/H55MdBwTiDuF86HWQQOtMwZk1cL3gVzsjYJkRTL+pDis6LHJb9tZNgRJYf
nnhLuJkw7cDmkpiwVCLSXGEywDVdSaPMX7/0wWyknwQ0AhcQtFQTK04/n0sJ/0JW
S/6WE/TsPn7WqRIhxR+mhU920b5OymGQ5+Y33TJgHmd8atbOpFzlU1DNJ0WFYfFU
DimBeUsxNnr5KIb9BcegbQqZu+qn1PKibNms0XbkT/kmMpZPx9dx1e0a3X/AMM9z
Q/FIIVjMDWjQGjiRc2MtZhjX8YR5fBv3Nb0UlRkH6BoSKN41iicoulB4kI/pLcIN
26ThLN8JCnNdtyoTkUMaw0Bc84p9BBAPl2qcyxkCpNEpnCWZ9KJujJ9TlWvf327G
ls4J2YAvJuk0KIvtgzufQNaC969DyZ+kw2hw1r1jzAc6yySdCN7jw/gS85R/z+X4
sf1ROtuG/6GcqLs80QZ/0/6V6P9bxGNzSHCymdZE4AxeAaLovJau3UhOphv+cImI
X8dFcLX4FZ8xRw3Vgnr0rd8Mh5hwP69S6vzKevmy8QLbwFIrtIgc40WuOhRhv6/1
NyV0MyctyAQi63LQM4PL9jc2hxwN977MhABqkmdWA8HmqQbFFQjyy7uiDWCw0+WL
kv4XbPBcm2HkRTd75vG9CRj27HJdlcLkePLatAa/ZqJzULdwEu63gRN0pVwbV5Ys
iXwAYW6Mm3XJPlv/CORHFI26v4qXnbbFGXGZIbzSSdB3YfGw94dobuDpX1t+Yt/z
WIqrGFKSq3lul3extp0X7Huz3sr0gVzfjTRBIb36su3y7CbO0407EFZlbNhl18jo
ToAPTQ7AXHeArcRtvwkGfRg2yWfLBhHYkpmxD8VNNfxw2HThBA4BjgMVnS/KFC9J
bMwENtJCGmOGnfcrKxeVLMYwh26+MuNDkzRI+7T8OpTBlJib7GqhkbgH0gyDMNPc
lQ5uPNToxLXoFiC7WnqXe9OhQ0NDKaAd7cUGSuaGfePkBS+CIy26Wo2inTNuNGBz
InUjLbNQKLJY9Bknnz3Mluy5+lThQSyZ9qiY2pXtc2o7tvb4X1vQd+AGXSRqOBGw
6EP/jGbE3G417BzlZKf3h+gXLQY+Q+Yw3HkMuvG/JU/4RR/p99HSHjjSzo5N7iIW
QYbu5/xDZ/+aaWYv3Bavr67TUubq4mGT970VQgpwb28wKWOzpuuQYl6Dw2HpsIAA
DhFsUrut1ZXzKLH+yUV+23yBC1Uj3quUNzMhq4iPf06spxDpYdRhzfqapJ65SfjB
n+LXLQnYUEq5CDw9KmA/1k3T0BWJIJt9sOmRWNdknhGG2l/MqIPOx8+TX7rbD4pu
kOndEdSNCJF6xAbs0/ouX1H4bvl1T50GIC/dRJR1ts85GPipsO4fYzeklw3HACHY
I9LxORmxD6BvSbHmO5vv5vPN4LPAd9h7pZ5mpHQwpoZmhpf1QsqNkFfKP0kdw8el
J1ev4YsGumJBlg1OrMQ7GgbxXOzwJqzQ3hKkvfEnVKl/lt2XztbdvI+nKJwblGlM
ByDwZlCRJHCxwVP/WICYo4pzZ2FC4qCdS+i0Gi3XKEzUXlsOBrcEaWPIGFTtsK9C
sVQ0d3bNvI9T3CBAHk0AEOiZ/ANjxtpkxsO6+W8nkcqsB2PUyI29WqekSyBwPQNy
sBJ4sXgERQpo4vlD7VDWcVDpe3Zztlrk1UiJbETlwfFOsOiUIANm0MnhNT7oys8c
lYqkq6UFlf8gAxJyrtetQbMggGxEyLOONWoOrHAmaMiKi63PyvO/sPbII04HSlZm
JeqCSlbeS98JeXWEFjrfBHH2tqXSM8H0mApS7+YcwVJTQiepR+Hki+mO0SsXNhSt
pOSF3XW63Tg0YNcqpw8pn+XDo77KWHlmlRODlCA04nJnng0MDFfSXnZZtwqjm3Lk
ljab6K4Cg8OSfd6UmHExM4HRRX1O0AoY73jofkhsgdzBYpLa8niptWBn00+Wvpps
k9VLZmn0fZ3O50emk4TBXXyL5sR7q6hdPSdyOi0FLXXtJtQnq4VKGEYl2hIs16n0
sF6GNnKIGmgF3f7gpWQe0Z8tMK1hpF5ZAIAV1kWpURYV5W+X/YM4uDtdIBpmADbX
/6ZuNNbsowlvTVzrSZJoC1SugCmPmnKHV88nKHZ/eiSHiSS4Tv0I/vNJ3sybyCuh
ApZAMwj/CwUeyAKq6KbvK+RKy3tS7P+9NCCZlwl9Wbogfl/gK/titKvAnuLWgprN
WxZfqCgbLKfjdy9QaaoUyOQXUyuuUkwMRTuIDpSXi0R/KVrU5e3ycpumiCXJphjF
oJyOMw2Ig+o15EfGfT+sDyYCw7jvYa497EefHQtHxex39IcBde9LERO3CS/e5ceV
ajf/8T6eazeiAbRN8rqQYspwHuWCSid/OZ8OJiFgK7LY1Qk95fJYLenEPKCziony
AS04PpOOMvVysmUWaMX48tN1Eg5EcLxbVn0MUqZRQv3GXbB6g95Soq7DndFfV6zt
KFNAilaKIRNoSlrmlvGoM/T0IB8nQ4irmro9TFmGe4MgVVYJtqd5COaM1tKAUKoJ
W86I2ZBT5bf6Qtk8uh7DCDerpc00zFpjOQ2kZXMIfHSAxWakmZL4/XO4dbEUsPP6
sHZSxrb+2N1jVd9tCv+NNu9xnlBKDmDWwF1QYR07daggBskQlEqtJID6TnJLLL6e
DIu+rQfgkvIyvUuA5IhvIFxRSse8bZAmFJ6AKIaNpfIcbxJ9KcOx+Ykp+urJrRPK
DACNyDAlWju+EDiHef+zxHKC0XUQQ8MPpiqW9dj5vG7O8GAyCpujVw5Wq/82mqE8
1x5rBjj51ACjSoy2d4ZNs9tPVLI5AyqIKcaLWxOJfCP6LJqKWES3HEkJ3zVhvWvo
p3kui8y7EcFhsxUdxOa24biDCiEc9MYb9I+PCTq1ss3sczB5iWVSxrCOMPEpLVPj
a6+99tXDDZv04LXqRxEQizs9iW2t25cIQGSthfUOQ6wzJ9ZjHBmUwNcrIGjZiS52
V2lJEnFt589bpBB435gNA+u0HswWfJaoW+SpNlCO+MxNwFOe1d4wWt4/nl1hDWei
gmWRMa8fDXHwtOZtHzhTwDumVFl3p9v0KUGTcMgJ6qYjhptL1G8EMzVmS2pHoAHK
ST1jPJgwsbq2LsOGiEjkXAxpsVg2K5PGAZNB3OvkY+3eOwzzYjERv6Dt4XSLLlHa
S7cByi7BWvOK0iWTchiCXyfkYmVz+y6quKPHQ4GvVQIgKELqYtHLtx5yAGp+TBBc
z6/2CTN254l1ePRhBagMOrS1/KVzhqCXJUKpVvvg7AeXW0MGAOtcDrIh+cV5N4mU
ioQIwaWHu3UutDzG5pvlxYuvzLk4iyqIiMq1vZmBEV0HJoXrpWFJTycekC5iGZGO
UPinAnvDvKlFijHiBwAfWJEQxBSeaiSuF8hClfHTNZqlXDCGJBK0CK01aZl7m58k
cVzqgGxFc2CCKXpRLZd7pL1pw4pWuM5G+OYq0X2sFoRX3JtocaPrMCUg5pQFcfyw
QDtnzsa4f4FvrhAJfA/W/dEN6jTzfEWqnPyyy1u2kjjxrfQxrza+Sm7SBUC+dHvV
c0h3DfAj2POBos/MpfILX1cjilWXjrGJYozRNU/NbofbU5Q+1T38lE1NXae2wp3W
mxTQ1CKIl8G+l3+WDFdI35mrXlg1xCigtSx0Z847he7r1nYjjxoAyhQPHXGHWXcm
4iIA53kNXxyTlmWAUWLK001Xn8oq5Vaau++uyfHrkLz0GnecaIDiHSc429sdfIMH
qYcrB7qVmj1dA5n+jORy8GfaBNd0ciKf3SdnpQuEOGUxoVuRMw4L25CkRTwnGzp1
11s2oHHYEfODznH9k8lJrsfFXnlbuLB1isGwS1/beuFVmhIMy70/VNJCCvM8I6CK
6vJHAIiXu83qG8QrhXXFHL2LEeToRWeo74CSCgIaoLIRC3WJE4iwhWPIvo63qAWo
i8iUVghiBBySFA3sMc8hK9Malq1AZ3S12no22b7WLYI/343n/oh4XjAWpMYUFVPJ
2XF2hcQxYDNGI//O4kXsPFD3hAcYoLw18AENQuFJtRb5rcoASnHz2Xs7FOlh0AqU
WPJEvk5VJev154nozeAD5ce858h//SHs9crc+a73rPagba3eII83bQGi2tyiGPDW
YCtJyp1dmlYYYggrtGU8HiX7h+7ISRuC77uYdm0Hu8Xc6xHaVPHCT1Xz8bH3F4Gd
iM/NWAaML22Dl38fDARK1BECKNnZ1eLJp6uy5UoJMoBr0gypSaI/mdB+aFLybZYQ
9kUUk0FxY/CSg8bLcYuqMAwQgk3GD0hlD9PU6MQxse2128OQIbTLfFVDhB6+YQNw
U+IxZ1l59VcpHd7h2I0Ui1CZJMnXP5ZpHF0F7EheyI/08PwcPWN7KcwmstwKb0lg
22Ozbr3Nyo8B1MkWKwmqjN4VXoQuky6mLLB4DAaQFRDOA6xMN46+Qzbk++uqzBGY
5zXa9Un6bf9+R46hn4zJQ4taaUQ/RGkc/RUcQ4YvEtcOmfChpkmOZy4rJiN/L5Pm
wwHcc65/2QjQ/3Q+L4QGY/eEPA2HmidQaMMK5vu55WAqb4KHzbZSk3lzAU3Lgv+8
X3Ih4DByTh+FaphoCInaH3DjaJRVITltcsVVRQpM0S4/Xf0CNpR3Gs5u97vSyQ3f
FZyWAbDYSkSnYUSwD2rDGjxJB5rUebJ3jWVwcjresgyAq4MVG1gWYA6mMfHocZ+p
5H3ut/JPMkn9ZySxYbs6SUCa2LdmHlzxNukS1g18eI5PXWX6D42fr4zYdnKP4GrZ
aoWu7Q54TPtvqzkgN+ChaoZDsh8mrDPipjXji2rgqvYgv6S80JwPHr6iR2ZkeQQM
8SbO4GiwwN4i0PcXjNMV49WSPoPEIkV+i0r/6z9kO8NRB0dBunsDsmHPuT7J7bKF
fGO+FC5qh1H9LVNmD5XqXRPXEmz9v01Gi8bRBfbKVcSPnDwiAU7LR6dHrgXQXlgv
TOGxgUo++lfD5GlVg3rjqPDqdztqHPpsImPMpABS+f5PC77wfeATb6H8G7yIocyc
iIAquNpzu1Pu5n7RKet9yIWsHcUwMHPxv+q+fazugforEUx67CH4SkiX8mqVSepn
TG3dZlCrxCpUQ5hXLOpV+F+LLYoADLhHPooU8OepUFV/xR71zb3eDkWUrYpDo5fy
Pm3YWFmFpSRGBmw20sl3SL3tJLSnyFLJxBSndc+36s8v9e1DYAmBpo3fWcQEetqt
WkyOjpjumRTj2Hm96dFF46YyXT5H69DeG+7YHQKy0TsAI5jHUK4IJ0iWvif9bEH2
DlLOtV6zCOhm48sllST25YJEVIavxUsmlFk521/L7Vag9lHjFkHhbrPY6Cl2lPca
qkc/ncSisPY76vmlicxFKlMkzEqGjaHIaJpQekGTHiO/Pn/mr2EubkzFTye+NTHV
e0/L+FTEos3QNGsLG3+WYf2Vv8FovyhJmVeNvzOaRq6L5FuGMMfu6ROImCCwAlLi
cM9K0GOAPDj8idTwKcRnAgC6HttkMGjrk2FMyXjRTVL7KkV10+h21WjcB6o00osZ
W/bfmjk2dzLxmsSJPRT359SJwxWISULB7PrFcQpVeQzkwExhjSQ/uQAa87BsGAv7
6OKojBS/3pP6JvEZS35tZXAx++rkcQqrMg1Y6Kb+qlqXB68uaf8lypBamy56dLPS
CpKm2voMKhiPO1P8hKIWROXuwvxwEVitdVy3EYrUhgXN1EMHeWug7xjKmjxVV0F1
iOOH3US6wDe0TcvHH5hz9x7qRBGK68Krf6kvaLkDHGggxuAAmsHwsZ03GjadHynz
hRBYF55fBiqV13ziWoGOdOWtned45YbC/I5jhDtdBxE+R5mEPpXnVumTxwrIK86/
hE8moZ+qKbAMiTm+0V00ID9yMrqv1JaFBoyEad1bkRqHcLncx6Mzwma7n1QmUHq4
mv0vN6XV4dGaDRBHuYS9Vaaz1g1V4Y030WOJoR9Fj8b+c/6NXSID2uSuaGSTdYeG
K3LXa7sqP2DMcAxpJMePgweE+ROinzHR5y1qIaw0jVuf8K3+MB4SV3TYogrQ9fp5
hmUblDBDw9qzPs/Bt3mHDo48qasVLedq7B99KRkc2VGcu5Gy7QUQMo2HE9S07phA
vLCb5JhiEAP0T6Q503fn+TDz3cIfl6yBXsCLD85FQ22x5iHQ3ZGpkgf15h6NULNt
3+ypcBUoy7Xt7amv5GpJJ2lXmazlu5frX2ugxMrH1pJ2KlvqPxVKmqlnFp54aJyZ
4LtXHkdhMWpGtg0vUZXvy4TteVWDXgUL43Wvbvy7w1W3Gdiczq/GvaIPC35pN9Ld
+HOMG8oX+uf8cW9esP+umHGiWLqHSilcZ6DREbTq27/bscDQLCAK2fv9R6g9ye2+
4pLvuAHOoY7kRryJn0XWlH7vFcdAbUN6GMVC8I2e5dMWPPSwToGhN7BnREZ3Emhf
XTbTJaea1WqU9FF4AtV97Aj5OIfe1fLttskop1dRo0MrPSmLmbd7DL61q+dEndtp
Vz8Ten2WVFUz6vcSHVLQlZNxr56/vsOxKUqhdiYmc2MhvNsU1k50Z9n4TjIvvuGe
cONnIa0AsJtNcX91S1iXK0EQZX1uhpI5dO58aFKCY4F1d+HLfkh9TQlzfHzutZ7I
TRdI2NFxUXdJ7x7lDQqqaR9WAjZKl6anEPhaPAntAv4MRTtefN9TBYCzLmwaqp1R
uLy7CR8a+cKWIx9GZhNNDtJaYO9+I3/WyGO1Y3ZjutXbMr/pjdhL/Fr0SojeLl2S
CJuqMhhmK+c9WYPETP1t/y7vPUJgK7xL9MIOMV8IPbx1z4bhO/N7rZj1lgzLDkPS
CboIMrcon4x45mx6smGSGMLSdXKcRJVxOnyjOxIw3CDPR6kYUvIBFdwXodQPF5sX
gJDsSzn2iIsb4/YbMRlZVB2VX7NfhujBYjOwuUOBQ3Fdk774YRqM+5rZcWs/FCb2
8/cXdNbfGLFyfFMMNK5YSrPQCorcIvXXWhwlHkHn+SrGtzYvTFwFcy/RWOpRGRTn
RfZewjJx+9BRW1Nj8113E5z/Xn2cWxWuZNIDVl+8aNV2pTjIvzKOF9q4heKq5rLA
nxGT2csBoOPRJAq9lQANsgZB/n9luGo0n5zjnsAV8xVTm/uRq2//fv9uxmJXDVs+
+1gl+zUgrBlF4VE1eL/vIxtzs7zUaqzvzs8tB7mKdUctyesRd2+Pu3yWtEFU3an0
+p7IqzzXURqGraXH+vaG+b1oA/sSxCNUNozzqOedS/2+F0bBdcVKt4rf288t4YDt
gLjGUzOKixhhvkmo79zYF9bhrpGH00ZgWOz07vC1Jtr0SwaNZB5V2HVFKJrL6xsz
2Zpm+OmC2YDntOVJrcrDXEmhrVUp3PT9gGhzJnC0G4T+T31iYrDruWOdR8CJbCDG
NA8xHjGzDWUBk9KsZ0JTfXw+sHnhluTRDUcrHmS+W6EGI+xcS3XQsdDK8K3LkpdQ
i9MS6R7IepNf11GczS39ztA/JZYhdromkR46gzMAsmCHP7Yvaq012iJjX2R7Lw0p
PPNQ+xQGaFwF4Mq1v48Wjs5up7iw2woxtmnMG/BQeKpzBRwdy2RLtPnj5gWWPHJT
f4L2yb+k3S/QUYebCqOpqt9Fgs6xFK+vv1jSDZ13ao3gE4vw949p97gaUJBv6sta
tsKtG/zvDy9AUOzyvPDBIv8IC9naG8OwsTp35Aib/1rZDrBZTY0NUrvhNGkA/2DX
WWS+aLwPkpIf+sYovnuEofM7bEtYpulwMfQP+t+L6kxZLGMh2rGZwTcRwsa5z1sa
1TT9quM9ONsJt457BIdygozDzUK3MJPYJb+SZPW+yL0A/Cc23PEmhsoFFv2LFBbA
4qmmA5zQZ5k2qRCQx2CtzSxM3eRr3aoVUa+KLw1pu3p2hE+yQopzJQ6DFelbBNg6
tl1aKZbpTnapwkzc3wveFSgQbNH1aIC/O5+6mu4NoULDc6vBKRh8tsDzo+bbnWZz
Brw0gFLxCTeCmIGUew3KcA+wDkqC7bOAMGjhjhfmvdTAWz3jQ+yRnk7O3S542Udp
lynArc46Ycjr9szkcCjAK5l6H56jw5z1qKntTmMFt/zvc21pRKX+tgMtfWDilDtb
kfE4TYobMLISnL/4ZarTlXZkiJ6FGerJY28WBuwBy822rjYWfh2sL69XRJSOHwP1
eiVNa1lwUxLLd6euFjnmcPAeihQS/BK85QldyacIA27ZmpK3u2bdr4oaejRvkUx+
elJOpREWuet82Otqq8aUqmwtqsfZvK3kvUM2nQ3YJqiavv2cE3MoLNglpa4iYl+I
V41EtgsV5A+Ul69ct/SpeN1+xXWc80JXiM1rScj4F/eydaz0q7rIRh467VNTcCvO
8odUxRlob2Et7tbYWfusxq2/t3l1qIjYv+FybWXZNaKNLABM872N4+dDu7BpP7qS
syPmal0Ygn7wuA3gWlIsmAnmycb71RWjAJx4f+I5ulQM+f2Q+HAdAGBmSylfMjFa
8e/vqqvl7mYIa972pfm6ly/PQB+uIyuToHR6wNf+ORb1/TL+NE9ugkPLUd9Fiby+
a9kHhgAvgGC1bYRjMReeMN6Svjv6tZOBc9PlD9JtA4qmTjbhH7P6tU6diB9Oqd9m
gX1w+M3jU9fCVGhIgY3KpH8f1EvffHXAxQ9yAWnVMBllEJm6wJkmyT7iXcSO5xVH
gxks0njwq49i1WSZqmD9ijOwN9Mw/lH9M6kdv43KJ9907RrYWZIR/5NHE2vCCNZi
Si3RTLGADM5O4LDczfC2VHLncyIVL3GSOM4FvPkAzApfs4j3qzzSrQP5YtVtCuYx
hQYbdCFVp2SkhSGhj1B3NyyiEalGDtSgXa+Qcd02guL17+Dck5B13PnkznyOp9BZ
Z2ZvsKbWS7GRA8lQrSJe2t3bQ9uTv4xTpoe0oJylIw4nYGnPVnptGKJ2DSnRU6Gj
qrWfHqh9Jk75dH0Rlcxa0sR1GO/a03V/jAqRD1X7mqcOwXk2Aa9AgA2QD7pN7WC+
pSty+kmAwTOmz8BNMqEwJlhu/ulQzPCAT2csz3pkup3ZJ4KzJQ1hLOnb7K9J7ShY
qoTpaB8yV3oACOCz1XtHekGPGGYwZ1X++fvMFXluljMs1/4qz33qeB+LBuIcQV40
cphwf8UEd7hd0ciQdOIbnUg/TLazdJZeMFniwjB8kr8SxH3i8weqVQ2j+vonHE/k
87Uj34Rv+YzXkY6e+9CJ3mZYoo+pSuI88cPaEZ5l5mAbnP1ubLdq4zmeVFRZeu1o
P2EWq4eLo5HTwURPn8R45TCdDBbX+Y4W5ZGlNHkMRw8mBnE72O5o5NOzh3Spdqry
M7RfT+4MdZUd4yv7MeT3hIsYnF8egJMeJ4d3V8DU8Pm4y9VrXCFs/N7CZeCpJf6z
uow8eTfjkCVHUmUhRo1NxNb9M8wZ0Ru6x2oDoq1APs5IVbQSTkSh8Q7W4JfXh4GS
j2EGMce4xKgIN2bNvcESn1Zq84a1Xr427RFupsRv3/4gTvCLGh2MZVcjiFTC/zVh
6Sa+Qwe7BlMZnq6x6cSUeP/0sTpxEQtm1oefJq3RE9OrArLYXJKzgtziu68VYvXY
HKwyyxyhzrxW1MUyYVnMMhuZYn3yb4AIpPeMSwETEVtTqV+ae3cHzQZ8REgyDOAs
w0JdHb97CTb0O6rW5Ge5zYKoUYH6G/aJb5ZMm1+ekS/qGagrMVru8xe+fibKhelR
LnVFM9Xn2E5q5BjyRMSa2ssov4aiRAqviyuhWeNcmIwYew1nqb/3X1frp+tSfvJq
P8WuMj+20gf1OuxPgX+tV35Q5bG7BHKM7pBq65Gg4jDmYqElVGSz7kzOPU+uH3pD
VpsVOG3KYVG/Y36OCJZ0CUqvBiUCc6hYYAPGh7lw3spkbkwEwdxQBzdQiFIKv+Cx
xVBXgQkHGX/m0hOZEYINZVo8oXWUi5+CivlqRlXsIOjmQ36ijggXosji6MFse5LG
e6mmwex+b9neX3yln2bnHtZ8mT6Ipdzc+4ekeMySIP2mlABGSWlyMI+wXfE6bpSj
LzLoOF+Z2z5vixDkPSTuMoUX2S1olpUU7e+WN1XmFY6x/ssTEcInl4Jjxr8WXscR
Hw0MBEoEYLoDmzbqq0Acx4jPNrPqMR+PWvznWalgckwRmprE/q+tI+vC+Y+BJbOs
V/NKa6+SYnMaWAC/tm6OYmIXZ/NH53ggDs9mkcc/RFYHD2pZ0uI9rXUR1JKaRxqX
RcZIqFJQsd7Dc/EUSURzs0toa1fT8ASpkHjjXy7h5X9mxna9GssxgCWQF9HtXIz5
FJn+HPHbwyCZemLUyD1SewuiNAK5ifIEAO3f/HUdslEoOcRBQepjGE5NfXsukR7J
eAmHclbJcHSbB3pFQrbDRjI4knX3CNrbJ5+zjgc/PutqcvoSdD3IsoddkpQ8juXd
jhcnqModCeor6a8HlXmOAHYzLvfHuZImCPdnysCrr8ZjL6/6WNtuzkuo0yAttxNT
EiQAWJxyxgev+qzlTzoerHsAiNs08vZo5aAhg+uXtz/WeXYkN0/VwrWqsehGQ4h6
sdc5BRUCArzIRCRQMuXq1vnJnAnllOMkpgWE9B9Y1BDjcYwjGexwbaFZfgziuAHm
Gtfa2BnnoFZ04nMLy8oAV3AqgR34Jh75yCHeuWeKEr2r+SzHkN4RiQFQK8sbA2tl
HQB+Xvyyogt+dMynX4ePtW97SHj6FbiWj6Vf8rz8RUsSnBsp2HyLMurRELoIovYH
Tc8G4g7us2/tYFbUyIN0sHnvhvBAEtbtgyXM6lMWSNRuKLsRME8LVwZmZf2umT4F
OTEyXCP3DZAK8PG7KaELdfM12uPQw4I3TquVTgsg3GFUlJzX9Mdr6BhWQm+9yzBj
rOmHy9GbwoY+P2pikV0ctnIk3jnReSUr+C7o87Hv4Bwyn5vhN0jV6miQXHftDuEl
Qg5dH+R/xlh3qez56WUcbyZEjk4IgG++Yd1j+vSLAODVFB8RRv35UFVAMLzsS7ol
XY6cXNQH+B2b0enjfMdfBtNY0WjsxRcEXvcZvsuX2zvNuaN8qaSC2S3hke/U6pFh
9TidGF97SAICt1RDdeg+nzkePT1BRlEY36PmmlNypfFJCFKhp8dJWhh0wdfZGFDE
jgs/E8WIkH+RatPSGZbq39JYR28BriHwybhSBlaGfheyQ4KvY6auZd7XA8t9k4Mx
rDvcaNyqFbB53e7wDtC0AqzhlSnLS859lFjZx9js90HrkfqxJD1C6koNXbEE7vCN
XrD9rrs36+E9k3xK1rmYRYntIsAdfk0m8MedWyiT3IQMYp+5vzGHTIkgeOThOxFd
ZjCmoB+pzbZe8wdl9kRXtRC75oTxFwnIgXQyZFj0ezuPGA7SLYaLwY1EQL6eo8QX
8+DCq4CTdWYdfBpuIgy/e4StlMKKRAmekeZ+/MV95ciBv69O2CVAaKtexqHfw5sE
tu0vyX0Akiubo1kfqdcIpkIrzMQqVJ8mPMQedIRoRSSYbS5f2/uazHpf9VwRxtmO
LhpSTPbk6zJdOXCLsF7HmobAlEhxATV07LypLwS/G6YrRMo1ib5BW64Jxbr28/1W
OZUvZ0shSryhukoLQzEJnnlZL6gD157KhIyq2+kLWHkLUhnhcFKi1hqxLNRTpznt
fqi8IizWPxA51pxbeK5YOG4HSHlvicegFMJwHdzjfzg0up2KmsKPIV9hi43GkCnc
WyT3c8CZjM0KhYZthW+R5SSh64aJP7mPe25DWW49xkXVJ/XnpTGKkBGDPi1ptE4N
KApF6SpYarBFyIutrYxEwtuzWhNc8bo4yZnK5oJlolSSPM9Imkvj31y57wR35DSB
OBvAODOmMVl+YHXLLKdjt7M4QQyxwnlw5/X3vWipq6Fx3eNgad2z60ltWZqe7L92
Gi3G9184yMO5FS2eJlg4BmdYs2M1kdKbKV09UUuq13F3DSZo7+T+wRlfrIZYxD4b
Bcej+DAHWKSZWZMgjFeYuJ5dJHux72I39eya3ebhRXFUeJBc0w9+Dc6muA0na5ZI
f6T9dhl7ioOqhUXCkpu2FD2tGl8pZkRtiYRCpg7yVYRA88+wFoLrS/DleOQcs55X
jGlMIqZQdBCcB14dVoA7W7BMN083ceMFVtZbgrjCp9SEEEnbu1kh5sL0bzWk2ITQ
ewfYkWVIFqgcDPJN2faJbuR7m5SDTs58tjyRDlYXgr/4yKlQnE5DWY7Kj/giy4Pa
L4EAN0dqTVg8TOc1oSbAfl+ZO12CS6ABid8zSDHCqx/m3BPQSSTCP++KB5LbJT6P
4gjRe0yknND5B2nn7vNhjPt07p38vCSaYQNJwmvDsbHRxkG967kaVKD3supbytxa
BGmrtX2yWVh6FasA4IK9pZx49jizv4IfzbGR7qxKzxlzPAcT17VUCN4EsrA4CWlI
uxyJBmJR0hVu0X2hKzq03Uli4NT4CerEB6oCVAw6cxTIyJdDVVs39eT9lchZ/qFy
R7l/M/UcjRh19Hcx2tEhrI88gGXbCaN2FDsmwIG5VHZIozkITbemLXC/gVDLN9uS
JOi2Atrh3anQHLZ8W1djtnqB2x1WwfjGc1gMA7Yc6blyil8lDY35E29l4Ugc5R3a
2evpH90EOnpW+ukOGqV39nyAG2yHFsAN2gepVyOV5SacN9cMzVZWzGxGDL4D1OHS
QCcrZ4OlovP5ZpjmnhyBGq+8TB+UkYI3yRJc2gHxx3eKd2uUBCoIgV6QK5yJNnD1
/1O/N5BURrhJm1Rbyo2f9qp7/htIoMBGGVN189tsiloymKXSQRme+YoK4MwjU5xa
xZ4glbJo4TP3L11W/ZSzMEIFVRpLNfzAr6nbTvOi3jdK4spaYPUtOX6XdEmj2jS0
5ObpZDJUJS+doL4ViaSVi53CEb3VryKyYx8PIOPgHo4eumNCPCNPljaFZQte+QQQ
6NAvV1bMnyM3n8yFXVNR6zFTGNZaVrT9uqy/jqrWlnb8HUNeHnH0EIxY6tJ5R2iu
ZzbT9oftlwmRBOFCHJL0I0HT+5Q6Tn8UyCSaiV23WnObg+ry22OFxmuzrdg6oPHm
+Fz3TnT0HjB1lHGDf5GuUk+2YzEJ3cY/uzpNJ1WNH+QsemUYo2IE0Fe8EF8tVMS5
nVx16i9yN8xo46yiRrhm/uIjYbhevYtbF+bd4FJfaxpMs7FVaDtcLQ2ov8lNZzTX
ck/yzVRKUlHwjxk4j0bmuDNAW5/vySTlDfiGhqQ9JsUkXABBqtYQuvfEys8TwuqL
b0sj36j4+X6o2YNGX0yPCZswVF1gk2jlEb9wIW6jSyxK1Pspu5ZZjwoJJm7Iu8dN
x3l4gUFiHzRa0sMIajVU0fvRSNa0t69H57Cqzz1MQXSqCZUtVdpdGx3hVHHhRRbX
FoQfOhmXt8R5siIjLYs29c4Q9OqBVvooojzGmLZVetWo+wxi3CbeVjpRZdlmen/O
VVf7/5sAq9bIYzKj54+Q2BLD+1YTUgImOmOYNInQx7g7D2isDQNulFy21AzS/ZuR
n3Td9DyIMnJaDBCD9TCX31ezHWjoz0NMqV6oUiGup5JY7ZBT5jPWgzqz0Y0fepxL
37AB64oHv7zIulvG7gLGnzCAY6Rh104i5b5TeKib/6dZXG+Z1gkrlq6JfwDIEc4z
/4At7kuCqUm3eI+SioMBMvjBhZKQDQNfVqSQpOn6HkKPZJRWOvEBVQoIcQ5CLHIx
3bhExZ6HsjCKsW/j7NjdfX9AOAVLUAlt2ztIakapbaxv6fJGnwAATEX3U4TJopWO
v2p9uLGqehNyjbSMfKTtuHu42I6hnJPUrp48otxNk1K4iX94ta8BiAR3vRmZKDUA
LVmr4MMvo9zq4++tsP4FOKMZbujmTF1IlPBY5AvqffAAi0l8SWbnK5yIqWUxJzdN
xfuc5A9cIMobqaqAHoSoVBgOIflVWysIRb/8XMOdrI46oOUXQaeaGGyzjHQbjfgS
BOevBSujeczfi67bk5xiJej8AOYpNvPAVc3wgeZ2Pi7UxICCK4rlYJ+8Fy9zdbqs
aiTLOyGKDYVZIzpWnwhKtQ1HNON8Ar6q3FV59kdV7IDOmDYwrVG0Yi/ViGdbx9Qn
t8kvyahCWqICGCOtTOKU6Qu3p3Lrcu6bNCwkP0s53J9UTalkyJ7x5SVNPe0jRPGw
43C7O1cj/8/ssjcPAR0acCV4+o6e5wnPu9GAudeHtHgX8wzV/JYNQ9j7JJ+dq5gB
ywsxLmfKeYjPeONTwJ6B9EsGKAPCCGPYjkEZDg+1wW8BfCg+PRrqm+p1v1h4Jp6o
S+4U7PqrQ4QtsWNp0cJQai2oNVUEoHEtxWx+4Q6uiOx9zusVUo7kvuZpZDxv3xPs
J1lLoPBI+Eakcv0kIOqinSd/JOXL2KDl5HFnLBsqO6CQeUvGxJUT3uokrVWJRHMs
bHHOQsKC8R6zmeoXheBXYIDgNE0SNI+RumtUkHNwH3P7D+tTPSSs3oUjBirvHirq
rcgeMaa4Wtam3k+9vapiJWStikoMbf3qwuQmEjbXtht/WrPv79P9ebQ2oZ4+0XuX
ivyYwJVG6dx6MeLWGoLBM9jC4Vu7jud7h261seJK2Rt/Glfj3nY5XRGr5XGoaMKs
MSiYgo/FTu3cR6MbqXAQhyWGOPmHJ6kB3pfjiRgXFVQ1BEfZ4CVCrXsKIDERS/b9
BPs4Kpw2tCcc29kpCxcwEPIdHlePZtLKuPKomjEeIdROMimMhdxBSB2ZWQ/KVBuZ
rdW28o4jMCQ2ANcRZAkb7hxL2QOCqfoFkYEzIS/n9g0vT9uejGVwJs1WapYYE66G
8XnxK2OhLK1rQpUoqRGbRCCDBhOMMj7O+NpQ0wfQesqANZpRV+kEEtdS6a8ivgxo
UjPFMxNlXV0m1Zkzza2pQbJNl9DxTEVwq2cJGU/XCS+joHcLP2IZTqD/PiqIrWmK
f+wDgX/o8vyfDngz3tqlZznitzx+8gG7w8EesKafg8eAxQsNzSZO4Q9VivzZELvG
7xqvYgqKhIU98K9Zl+IKdtdHz8DUNeUIbVEK6RZPW9agzsj0ksA/yYCkj1Ip3YrQ
v84NZJx8+7tqlKQs2AHZyjrSDWbL7906r9bcd0liM2JnIofRrc46v7aJkN4prgIZ
Zt2hdDivkxtUM9XgEkjqRYv7HcnIcml7y5zkvYi8swcTGFPlcF9WFRE/ksU+denb
I4mC05sxyaBfmObC0i5xu/aIlFJecM3AHKqYQbFgWxj0mLFEG3CkZToStL6haEDu
zupENj8KKn+vEmEN0mfnFPFA1pv87Kob9cfohSn9+yiPmEJAnDIOYogdXuva/pPJ
TRj/foqpOfPm2ZOLlPnX/6s9f8HsHR/lBmHNhnqlloRalrCcmBQPnHyytI+lXjgs
jiCkNQ29dnSfgITDeFueGcthoYl8mEAQ/vi/9F0bsEdGyNzTTEoVs1bskSoSsJaN
yxOK2GVprs6/wjKhWfe7FnKEUmjJ1N6AEgQKaU9O3kU+EfoxF9u4el2nbqYkC5j7
3gxTokLWolQwyZXvv3TvvEvWfFp9P2RG+PWd7rgxle5HGOeH+SNXeKoyDmENgYzY
lZSARQoMBcIicQHtF1tHglssNTomI3eAru+2v+F8V2t3X6X05Uk7RKz4aEDLI+qe
bC0iLz+fHZYqRdkPvzcnM8kNlVNLXXJPfsWn7bcbox0C5eBNtMELRFYryTEM4Y+o
LyAY6W6Dv0c0RwGa05hJapXQviunO7Gd1vwGsaTEnle0jHJDHpUAf0eKgusKYZzU
+Y/TQ8Uc+BNamoy+oPYfhDeXUJRLLdxs55ey4tzTvXtU6Eb9dz4AYoBF2AJE9EJr
pDFmORC/ispa4vpo0Ajg+ezSUJbCzJB/7nnacZ47zoLL9iYPRCg7/OqnSxg4PLD2
6wRxIU0hN+s/KmuX3HKp4OSrQzYUR1YXQImW0Yt/5Y6uGLvJHnb8Ltje8wirx6wH
zusUWT+sORR/adzmseLyxX9yQY1w+gFJihXQqIH00EUeLGlmnglmXrSpsy61IG2b
x7m9OoGUn1OYSoc67PtrcEqLa5dpm8vyDZXxvm2DHB9gmWKjUvkzM7Pa9vy9Uo2w
zFEcm4p/zR+FJRwC5M7seaS27QnvmLKbyZewu6lnVAmIcBtKyZjBJQkjUQbqM3MR
L4scHneAdzbpQ+6ABMl8zWbDrer4SkmlPqx/z6IXBU+S/kZZ+fwn06MGd/VYtgVn
3huXFp6KeTbkChw1xKpzDtgLU+CjJc488QjOZGkfho4wqZmzFYtIbss58xVcoevM
y4u6OF6etqurqqHXLnmyBQ6CcJ3cN6yF0VeIX8QY3Ezw2Y1To7wHivd4dFwIzZAb
wgiP6Wotka2z/uWpGO+Bm1T1RFzaFCYY+hqaaaUsV18+sMTSphATrnXx/Swzfb57
iBIRPsuX2H5KQkv9CbSBhj6FD8c0oifWOw3NY+0N+/4bVYavzomU2puAIlIo6xwS
tYexL46UlzNmNiGJC8xIs2HRBVFAvAFCSI/sQM0sm9nivwr1ek4g2NNnkSLHMSjC
rgtcr+w+XY1e7bWvVre9gcATdbl/5KvNWKsNKQ/rV/u9rZT1mqKhihhSZgtXs3n/
Gz0+lbeVCODtodMfeks+QG7ivQcqZCgmGPHa1ERH/pf3BjgyJrGUslK/RnbU4EXC
f4wSPtuvSIDUUhYjJ4nsPoJlzzILhZRedF/B4kGt3KdisKARZh7kto8xeu3PV9bN
sBOwfzM0dFqoShdUps5QTcwtoeh36Y3WYZ0pLvcs1NtiOk3+aM7k9L/mRclmtCD7
A746wcf8So2jDjENAl9YXvVVIsq3xjEwErmzbwoveWD/XS5x+1SvWbC1Npfva1/+
XgvNK+yq9Gym4L4XqRV4wrxHeHVrbKA71UVXj9uDGMU5TkvCbqRKW54daojMAXET
tmh+nnicV3ZVd5j/KzQuKwKfxsDf5SLJ0znJDR1nWhxZGGXfbXVSWYR+T/G2Z7FX
MHpDmBERITCsSEYN9Z2YM94uD98QUulL3dE5lxStTjMNAcmtuikNmjeoHhBkWJbD
qjOyd4JQwKRyen0FTFc5bY2GYBMNCdojwE+eZtEWgkVan7hZXX35JY/BFEF+I9Yr
dRf0gKfedZu/zUELYadcvblPgj2z75aVG6acBsBVETxIb4xWTyAPiSg+TPtuOMgQ
tLxVS35dv6pOax5ltUzFQFUK94ZLApTD3S8E6FsMigByqYH2zz/S6W4LAvR7Gq7m
L2krcWJWBsJvFuFph+kfDpH+Gm2BCZpmbNmkrTYW4elm5tU2LLL0UVcHEDF70v20
JPZAYayrMcEEywzQF5z5kNvs9ceejYpaPvt3X7BkIQCVmy7gFpk6poO3Z1os3Nd5
j5mzcHjO69eh9QxQjwXfIbnmMgl9/xd2vwKAD8RQe02NYmyDeQr+uLKumzPV0LWp
AThtZpScJw7IhzElspdvjXMGMr5Zh0R+zKCalGkWt2T+KjEMMj+TnmSF66NwUFwx
t2Nd2oecoKSaBN/EU35F1vZGCtDS00mSy4NY+0MgPBBp8mmz/gMpoddhMY9RSefc
WXJZBAJbu62VJeePfs1TH7PxGEJIFL5q/m355jMzwo1cE8Vrn4AHlPpd2yYsCoIF
YOSHKwuDymXpFZidXFoTQidecIz8JmXyhRNjo2y8mLhTq6bW6K0kgRZW7Jp5U9+a
Y4f8fk9RTm/1jl3oSyANIpa18RK1XwKEUWh6dzacQq+ZXlzAeVnWOjkgSYs+1vta
3u3+N/pxA/U/ih3yDu4PDVYGk4PQBS5ybjte+iKuDQoVS7y3WREmYJTTuRYs2O4Z
OtS2/DOzlC1c/zDIe8umNsQyo+WJZzjp1VFmxaG5e8BNG5iUjaGoAb5n1eLzndz3
G2XzOYvHz+WMzWTwKSvH/ZPuW0tIrhPjsmgv9lHzYols+xYXMmA2oDGNf82i+VCY
We6WZYfXNdIFeYzKiNYpnEF5kKcjdayjEN4JQsJeIdPX1/7s3Lu9cZM6xSSl10Dp
z1icwge+G9VDE7MxwK9YbWsg0zmH3YUSa7onl7n1P+MqX/Sj6S/AsN8waPKHvuA+
KrSA7PWZBfQcUGgo+AL6VyVCaXRVhg36NuowmawspRC+QEti/Hwo55HZJFvAuETP
hlzJYV0JDYgeN+iyTl7Yha5uJ2Owj0kGIpdm43Y1Bm05db0CP4w2DllF4J4CxFEw
ZQv0liA1cCBlD9uxLlC67v236pm+AqBWxB8GpWxeIkQu2Sxpz33YwclJnuGg+i5a
er9Gsvqm+WqzqrXp/Uls0dcRouiDi/1QSGOmqPlZf6FRMofjmTikQnFSl6hBkDX0
Oe8toESMiKC008HMKT/lhYhWJbchf1sZCo6xong9n2bjWe7vkEsgfFDXZeUGL/gb
KbR+9Km8pxeov3RxLQPHnuClY4uPdU286JVwQEqgYh1rwI0CZiiF2QdGD406jzF3
iP7GhaWWZ64HzSBByY7wZ5M1rRQGpY6qdkJkXAgxOo8xboYVM5tfakWNW5Ua3fr6
KRurj/wib51w+iiHT2l6GkrvoudEJ5wAZBF32GPbLLZQwnCAE8DuXyVHXqcTF5wg
3Hqlha7ffpwUyMoB45uhQL6TzkHafzQEjvD9voTWCfKo4WP8NBcY24hBctSuVwrF
FVum2LeWTWLW31vvIS6n1LT4a0y3yXc0bLKtW8wO8avOR2Wg4Tsepi2Kn3hmHC0d
cV+pifwRygn8QzYqCdnBP6FRJRhWGTOV4SCCUGF9TpONORlUgZRiL+4HJ6TA6sx0
L/8vWC4RvLo5sXfhPUcTKLXMwC1qcyHPp8OmaW/NRe5svu06zGGeroK3+B0m582+
cUMGJSu2zD8fyQU/nBwi/OaxWILjjS/wnh7RbTCEUfiAOc7lDUpn0WUDHswoIETA
rjm17koQuWWH3IEEn1yPCgxXWTu2jXwe3KqVcl6S6jesPXLbYzpyplQk+RIw7Xuo
HgLEmeXqAVMASU2Wlq+AaM9wwz1IZxE60GWtXoHyqPVQa0yamPc3kZVknwvenZc2
e3LhGE0+VB/5vUfhzT718QR5B35W3ico5xZ7DicEQlMXsJZCPAzXVvQw46bTyZSt
g9LO/zzDILKbk2sLCobF46bZL5sguNruMS/JET1xW9G+96+BKH2ZUpU0Ooj1deSj
+Kvh5b+WVKAvAusTHzFiRw+bN/n23zJJJTrDOXMczJvM+4icJi6PWmfB6qwXZQmS
PdBOFQd5C5r9swpGB9kpm+Ekke/kL302PBD15TgZDHvlLst7m7o1d9dJlu41Dhxn
bBaB/JCeCr+KK616BLZCvIjTVz7rkCmV8oWH+0Dj87frAfuQoCParuGBSPNy0xgD
PKJSXoAdmspKqYedCL4YptyVjd5+cM04n/2r7YqGt7BmPZAkgyABzZpY2cXKCJcL
m2KR3ubtPWqQBaNsNu8cXocUGEzFkvEg9EfxbBk1F8Na0YgHuR0xK/L2DN/x2Ozn
C5Xx1oyYsdvALnL+B6f7BXHfLFNvOGfxnLhsNBU1qaWoSyfjWLjYtCce1F6YbPhY
59v22wmrgrjHD5lON3RO78tpYv4rZ2prxhQnzYfJaKC55KO8sfHIjg3jIIjxye6j
hT9GfdQ7lQ8AP9zGcVSxeSyyVWUdhkXiQrwARjhObwn99DxyZ1H98JrP5aB6Do83
wv6UQ5P3PEoxUFZTAXInvq11P+uhrAAmrx5OxavYl7VlqR9GEzErWHXQt4/Mz2cb
4w9+Cw2g6AMGcMs7HyfqJRXxA0xQH30vOTBlqAS3+QrhE03mNkn2wy6V1j8d4JLL
brl3YFgjZYm0B5er5030fshVa05Xfimbni5VgsSn03rKYEKlJLzcnmgFdJxCeRGv
rHnPukJZvn2TIYbUo42oFHe/0gwxsz7WNv365yC5N1vRy715bkgACDnESciGCd/R
a1txbDFJs2ZEg0WnCmOeB23EmePrEGsJe6p4y2xSMXa/mlZmJtc34j4+O4Ri/5eo
rFpyC0Trr87kFlWHHwGcNn5jmD8IegbD8qk7YqRXi4SeWYCEHoZhBVuWX5tfcyah
xzKu5KnmbtzkJVMWdHfMA1Ln+tRjT9FqF5Up1XXCJex/rDHG5RXPzYL3fc8K8JHv
s4nM6qwzEADogxShFRiupk7Q9uQjoA/DNQ1n4lxvex7OZBqqIub0jQeaJ+h9hd6C
p1AvBQYBaqXLzhz5WHIbBa6IWpkru04l+1Qx/8zsdqJMPkmk5YCz2OPxOE0HhW/I
Ut+bT5MKRhRuN99XwvTlQmXjOl8HtYr6sGmyA9DoUYWUatpigzJiq6m9SEUBYzqZ
cvFsFvYP5sA4pqBU1x5sQRXzD2Yb9R48rLJXSxbGz2q9F6z6KJEfDN+j8yT5xvJx
6GLhio3TxC6sg/gjhcWHwFsmQVhM7+hrVsi4RqEcqFVCh8k95Kuur/ujlKOdNQpZ
zi2QyeWhjkufOzAwG1otq5IEGI6XY6ltDB/Rb5UrF7/zVnnnirE7rZ28UlwhMO0D
2Al4G/7otPJza1dbV03/xFYgbszJRYpVzR1dBwE0FmufBeOQwWp0ohTtBt3OuUW3
pp6SdvrzPUUZKvQBj0SPOQ1RO93sVCyq5iaHhqWVyMGVJgq7nWNgTbosNadDEfOj
XEGfxAuCPs2nrs7vi+GseHvml6vaCfn01juxAQeTUf3D/74YAnDxD4NyTnvLAkHe
c3UEmw4iHU33cczcIgm53vqkvUJWDBMjtJN4l9s9PkUwotQI7bJyPDXzkKF2pg2F
NLlYobMH5Xmhsxw00GMua62oqHgXE37ZmTfz9aB3kBV/h8EWxsZsTbXTvnIRSB9L
bV4aH/BPbJqOGyliyZg4edPGCFhrS2AMI1/u+wckgfqfwSlTtS7U3QBJVqAzx6sY
1FfSl8P4CpPMimzAHVt82Y0yiNmd/gdMJyrZoh8xgMlXu3FbzG4Yyd+eRbIRI/Va
6OYJspKF4EBNZ2AEDxsmZuMXKJmSiB9ZIRQbvVAgEQlkjIsL3kL2Slqvn4qOa6Vm
GV3FKz0yK1FSVYzmBT5J7lEGLMTJWPO1V6zrqmhEHNUxd9HRulMzAZaLGq9Eh9e3
KLEdFAzU7xFtjb9uP/uX1IaIWMXyeQ8EWq6PpTmTHPUMZK9tJe+68fmptx3E+ShY
qZNAPWhTDRvNPFkQoLtx40QueduhTLVKMV0QgfrN5rInTIRwvyE4z24jEcPWIuK7
1m8YsLo+T5YNS/yaSKvwW9Rg/Ae5w1ZV7OlnGz5TS9zFQYefK5rekeSCG+Nv/pJ1
cvRfsTOFtbCkZTCw9hDF3B4HXiNspw+VRXgw5zspjcu7Fkb0tmk9+efLpWu3l3jn
nF84OfjVbC4S/CCHxWAGq1VjVAeWmrY5BuhCnIukAxx+axILLL5vWlKZrwGmz/6j
3rE62jG6usrPaP72Wb5Ld5hLE0+KcA+vcP++mhEkJF10+cOBSoYNlFBuSsQosqIG
y0yLanDn9+j5MTB1iP5rvliSg3iDMpa8zvjZyCQD8SFE22SzMKzsvKRZBYe7hSz/
YLhK4cFg/35HpHp/mdwF3nOZOsVFi9zVeR9gvJPtgtido8PGFvDn2PzYqjchk3Mw
I00f44HdOOsRuG0OWt+K5Uty4fiwQqtECC44SAteZP/PC7xWfwnYAtoRVUvv6gfe
xpw7zokCv8N5qX5tCav4GjiSq6cz8KcvCzodfBaq4NTqvnqox94RXcuXlSiIw5PC
dCWgZcAG3mtaTrjwQ6+r08klrk2eD+cE7uxX0Y2BP+Av/uhh92R00Hh1iqOXhpef
AfgZWzP7H+P+42ZFDIBOqOBiVdMdl2CHX1zGcQd7YV9xDZlZvVGSuqbq1BVOuPv8
vF2462DKjVAiLppjdD7jTHYFTgcAuW+VhzdbIpNZ12cnfHst9E34gEFhwh8T5Pmw
Ds439fOFVl8giznjhJ94ITHXEaf+ag7l8+QJ7dOtIZ+7pPOA6Pze0jyWW2APQ3sn
SNqwWIJEwcDO7PkQDYXrmjS6Rbx5/8GPnXm8qPYvjjgwgAqkLIFmcyH8zJWKqclW
rHp74zf94JkLQGjdo9DJkIJ1omz1CE/TMv2M0r0X8Fpag7b+x8qp0kawKkqR+sJz
KofLw7ecF8AR9/mDz43xOiEfH8e9I2C5Lw0mMd83NuYqq8o9IErd4t9urNhyDu44
MQBzRbYZngUeMSE3716blkuwkWifiNl0xVWjuB/3z+MVArD4wU1QpgyUcefCncKt
ZY159cmqOIi2SrO+PqXihE44Vx20CbdHp091L8kiZ5lUipld/UfKr8+efP1o2kqe
OusnCrw58XmHJwHFtTw6Q5x1edoPHowmxCcav3UPNqaSn7FtnoMxf2S+Cb3ZrcmD
tZzbQV6kno1dvY1zqRDnK1ad41HUF4BMMGUXO7tUD4Wr2ASBCMpE/CADRK7pAw5n
QJobkxtXETEq1x3taMximtM8tJwT2XVVq9T5YUQlrAQPcforrYjFRphqfe2B5UT4
mxmc71j4aVOI0Biqn1CfOSjz8t8bW3YQqPkHnFoFCaAlaHO8CPdb3ZdZfaoT/ZRy
MXcoROcbqbU0fLlhsFO1wI+/QTM5jDt+zL6PI5tF1R+qik/5qmnKBEzdj3oJp/Tu
N6txueS9EnnMqCfkzDF1nVcFqVHu4ZJ4aW11e5f9QmFwK+6kHkaV8MwVSqpiBWSB
Loz82VHBJuxRNy44+lsqASipu9FcXJp08w6pvqqhUV4ugihlj/GKlJOtX9cOa+jv
rnTH3CWFymE9MvNn9+Bgy5debQokgLFUs/hQx4EJqV9cbCluvdllyKfbmhNajZ7z
FeyroqJHnJXaqXMjZtTdCiTEgp02KGSYkqqr8gxolZSGQqwT2K4yHaBRi/y+HO2/
ZDM+Z/oPP+BNmoy3c9uCgVvThLmKLDXqgiA8p0QhUF3mNbqdcj4hvJox30JNBaTh
+xRVqNYehX2un4HLY31/sYK9YmZojdpNrcPqNRsFATPYspTZA+zOoh1aUqGCBPgo
tmqB0Y2b0m8RSiG+A0oeYdzPA2WtPUuyOjBsvjBViiUxNdbAoL0ib9qESiNxe+xq
j1/fkQ1W+Fpl1n0skKPwprefZOjMV4ABOp8g+T9fQHZYgp5g4+GmYUSQNDLPNvX5
36tXfSx3J9WucbIKG8WsW8Vtexn+AqPGr7kJX6VYzGUX55lB2tg0nz1N1iqcmPuh
9xw+BhCopgdP/ZZIocCHcZ46bnLnxIfNkASKiojl+i1rYS/3nEaKRkpUSN+N3XU7
ocRY1YA52iMB6ocVp226khjp+b2+cKwwbkAnbrlemrWF3OerVNrBaviLVpU6pVzz
zpvXUs7K2MRZg+kpEnT9Lr5TLXGGBH6FAWr5AaqS7YEwBRN4c3pPJqLixvuhS+JR
EFKcXl6WQAtQMSpGGj5Je4Z98gDhCIjunzRwsG0y8HV9uuJXNFyOU/h++Tpo2C2L
bcfPSEJzPPXxfCjsy2WMZN3lLeUW36xo38Fcr8prqw8Ijt7vWhynYFe4EJ2AhkXs
mVnFldmU9PNgf7ZLUrx30aUvbkbFO4jaryo405F0QPBZon7vHGQV2rbZ48CdWu28
iEQJNPI1kUtgkczPWaNRvah4sxaOgZa1pM5RtUE8I7Wr2SmC7UcIjYvlPyKzoW/A
zjlsHq6LiE8UYgguP+kn1RAye466uC+CTpBuRgobZoAiwA2vS8bGbVeI5I589pmt
uRBM1nqPJztgOSEN6grlcuMqE2Lb5LBzp5SELgUMYLm6bAJ2WmBAEhYj+FHlgSo7
ot5R6NbNsLjOaO05u8Gq0rtLQGt0x9983dIX25dB4CvZH6tVY6BMr/0rpNLOy41D
RK405OAKiINQTJOfZJUbYqs6/2deRPo2fPTLi4XQxadVIBJGu+dRHWMxPJef6S0Y
0IEXbER9yy9DZUd4WN5eogxXwixeCr5CyQeMdD64WxMGxGuO6C3L0wIhtR/H7YF9
FyJ0PrwlVURHJvrpX16xbiux1HK0+CKzNJ3gFEGh28qxg/dtj9Kgalvx/uU/YQ8g
k94JsNvPa//Z6OGRbOsZwdXB576nBhGhf48rM+Eb/g7YUI2HDRNI2UjlRdLc7lCE
FI4p+PjDEOOH6ZAvRIjqX2uvrK0s/MfTLGE/tcdtWy/tNphRiLw4bqcc7k6ZfviW
v6dgdf4di4yQ6BN3t4SwOBrbTQgJQKmOyh0MEv2ESbTkGqANlNcVqoh5+vpH5REU
3X2DkS8aR5n5SB056sjMhmW/LZkt93JS2EimVyd4WDb4NckmfA/2STZItFZPTdOr
c9gmBkiB6KBdINBY6CbyIQ908MzxbGkUhPuggZ7CnwLDEnqf+BV/B+gp1RaMLChg
SSDlmSzZTHXQqsh6f0DGdXZWdZ3n0pqjLf/zvYMQ8WTyN3qSnWXE/Fx9kT+UfiuU
mT27I9mIl8JuFqNpbrDsvmnOpgpfEh66aHpva4SndKDhvj+Ys7AaMdFRs/fS9vbI
tTU3o8LQIXqk/D8qHiKETKgFf31guZpEnR9XCDo3lfrmACsL6SFmUIcR2l3iy5Cm
KMe2d8X9bt8fzy3Xi5U+iN6mY+k4jVAN/SOO4QP9qC6k/KNwiA8n430eGXpMRFdZ
SR8l5dH6noo5i9ADXTm42B1FAXy4aF9hyGWtKbTMpDqt5fvgEonPMLjVSdJTwFWs
+yP3sdcurr8xJyZYPMx1T4cFp/H1TFIQ4yl470O6e7esXSkh6/3SQu40iPz8cEQB
x37Y7JgvQ1KLWHOFeJkyCWGS4y7YtgWP6RYQGzm60x+GG81KN+4WNqntrIXwBEtF
T65ORpXsH6dpyxn3QI+fHa2kLEJQ8woRuv7+Flla71kVArFUXpoNj9A+JolwTXSU
BfctgxXBy6Siw0tq3j5e+plIPbFHIbUfuAHBF5gxAnteiweCzOWBO5vAt4aocWY5
w3uDJKA0qoDu6kx4h/qdoaGAfx3VPGHBiWZAVQ4LdfR8USUa113qhEbty2ODdBWG
QA/+tPR7iJn/8y50HC3WknQ67UDc8N61h/1Sbvym1a1nFWXzgtVt+yvdKaji6Vmi
O3dLP4lo5eWCUEGXqgFEakkoRphPqZ2AsZ9nlaEibmIX9Xg2qnAN6fejt1nAx9El
GS4GnIJFDyCUpheCnlah3vtJ8Ch/zCTZ9/PhbFYU0LgNu7uoE+n0o9qcU3vDwUCg
PSsl7ZIy/eZm2ofGBp7UhZE8xf8rj7EArWlndFcT4NKfyhzeSiIo1BUHDZm9jfRa
SWo0czOBgnAhf+Lh1/1+GFFseN2ECFbzSwpoFzcYO7p1jMc7En1wrttciDI7AQS+
50ha5kg6J5FB7gO778lwd+f0z/xULfEGqca8QCS6USQT5n7GlYp0/qhJl6w4MlET
Dkjx8QyMR8Sq9OEqo/7cP+CeukceMXWmkIDXUWQaOgGhwYahBAJIJzZRqa4Op7Hm
nBWvAgEZHhODVNjw7rl2DO/oWF502/pjKNhr0tU6c3MXrbG6eN3oqcee/JYza0vZ
C2ohV6VnglMJYEbvMWWzjzvlZqD3HssWBz8toYjmUxuWwO14wM5j0TtPg8bpIZFp
dOVaxccNnZOdbaSbZT0k8CB8Rdc1cA2qATM/0lXSjCyt8PIQheRTFksu/MBq5Lc/
cx7nK2bi/tKMw8+qpPLaeL9nh/0DVW270rqFmjubvNWW7+xRIjmlzvXPrgFtNiL4
Aa4rpsj/TIF1daJOXIhvBTO1j+PBkjM1dOpQeP4KKeX7kYnB7/r48lmm6BVdLLK0
HIDHrDg2vt5bXMVemdzVWjEZS8j0EjKfWG06ZOkaEg3nGWGgmpdlG8eh/OliU4Q3
KTuhJG8iPMkXrvtIjTomN5NTPg3AQq562o4ti6TzNf3Jejeh6o2yOhaMPd9X2Ofl
Wh+8cPuyfepBhSDKijcVsN7zPbSXkzn5BvlQwRQpY+rGiKywxT87KMq8UZ79KgJh
JsKL5zkxcGa7Sox0VuZ53q9Fc/PO4Ip4GiT4eNNc3XuVVdQDkKnlqCmyqT3JuxpT
pCM8sD8bWFATwTsEjBO/OC2lJD9KGXa6gC4z6VPP7bxTB8u+8mJtSXRHff3NY4I3
HAuDqn52Myob8pHXsMQAc7CjyqKcoQZ8PS4texPa31WJpXux73Ndri6ZutxXzUrJ
KG/ISnrvX/gnHaSusNIojp7dgOqT3shV2/Eu70oYrYCYC7oOoMK7ImFj4WPbxSgh
f3EuDEvHeQTJw+akbZ4TSDJuMoj+s4Ow/Z4p24A1jGizIGQ3Kr0u/noddUFimVdt
RNiVjS2j3dtWW/AY7oRMilVUOzpGz6s3n/WGm8xUJnZfqOg9TmiclBJgSvbXa9wM
/1h5/NAhUWG9tCdbgbd5ojnn4ayjwralKSQvZN5A/+KmlMbeDEJPEZhlaBvtv78H
budD8xUX8apo5UuqSS/JjGBLKw2n404Pbfy0qlwmPIO9bf7SWRoWGD1q2VEXc3kP
OSOBDQh0suaty2cYmMt+Wu0uzy6THoVspB0F3c/BayNYcESR0QDLhX2pbXk4LD/X
x+23NnyPcU9ymzJlmxa5eHp2ijRfgKALkvkbAkrcwF+SGkF2FbhLn7D9RxWxa98a
jecNe3lTVT9u0HzRxiNBGtCgiKx1+xLoMkeGC88NbGyEZ+4OaiyexvQythEIbdCc
uzTay8ubgpqsDbLsfbOjEyh9reZ4kSmew/gtm/VjtZQopqKJNkK4OiU7Tw+XbNAW
ErLr9vs36E4tWRFwmDefIZiYiQ2ruOQVQ/du0oVlTxppjPmBGZxupcGppx9t9xB8
uD+5MPg+njr/wg1/uh/dKKs6xPmIT2kkjgspx3EvQdkm+m37p40GwfOqeJkRGKft
/8d/1TAL3wAN1qrFCl8qFRL9O7LhyxRAzf02/dpZWQ3QMAXejxQBM2/grxu7/aKb
D5Zk/6DP3+Q9Y/P2Pg3RVUn7WYAbFy2chHcfhgQACfDP5S50JcEBw7Bn9HPCmTRl
2H0kc+rqgQqdtkBb9Gn/j9d8NPm9QFVlbnP6P6Zi8jR+Iy4pV2hwf4jBQouCgiTK
X/vjzap0M0iw01z/crHSLGnbUIWJIlgHcruldOEmoQDuox5VVyDCSUPCQq50lxKx
FOeA9fe3R5nwbWtygiQy7AyFMErJBX1V8ghwPxbwnp08unia1wz7vlQz8+W2aOHY
c3TjiqRcC1YE4k8yu6/1T1uw7IeYAiFLiXKaE1sWB4r/meBpXZ+4fFRYDb/GLmVM
rwc+5enEFI2PytMqSVOhuNGgR15zHTjOb62FO83aQ6KJcRVbOGsJ3hfliU5bIyes
5938GJ0P452v7kRgpo+LKcjjBWEg3ClZQqMvi1qGJ7d1zhvdao3JUQa4AmSmNsrS
Ke+E/i7kbHt/OOvRFQY9cn6feRlA4a7f+r+WrsSrN8gcuKHLwYmkkHZ1NaSEKfX2
RU/T29nuPxrnhWOrL+IXQR2lln/rh9q4lZgw0hZYo8UPlsNc2bvR7p8uM6ggkJ+l
c09eZEw4kR8pYYd40TDZ6fxwPEgB1J9N5O+qn1WPcq1ERZfi4iljMIS61SAJtW/C
SXp+W7TZMXgmQUnJZRDS8tEMXJB4KBEQMSXvV3T2FMK31BkpunoPk4HQNm5zF86m
qf3ECCYx9NpCvpfE71sAj1wOVrr8/CT+6b6u8u67w74Ns059y+GxobfUzE+HMUPR
mXVDxz4o5HGBKe7mhWHBpgQMFA0+68Jz4s/45Ig4H8rJSTe06Y5/JseRTP0a0PLE
g2mAuLuAUTaGCexqcuUK42zPQfVMPjb7szZag/a9pMm9/QXnghu4PD8alHjC0GMo
8+DHtMXlrDr6JGaErGeoPjLACzBAyJZt2EJ8V0YuFQNKG3yEQMGz9RpGwIUnL9c+
gJcDOtgVC1YS9Olooq32lo3cuB2o1aWMa8/AVXLYWYmZ84Kk8UDJldlAqVCMAh8e
Pd6fwIpLRjq3n1Yvd2//6mB+SEUpoxzH0y7MxbEsqVE19y0YwIpD/s9AZSASRR/v
CIFl+Y6ySiINhKXPKe/58t518IJhY4SXtulL/nOLN8fogozPSHz8Cq7r59cDxsZN
0GN2LGH2j+OvXrfoUEw4njcP8bOynJLc5ZxFJkSGg/k2MF5Yw9QMJQTEO4/ctDHC
TnCVsVDsJ09TIxo6SB9/qOXXk77OO/XmcyJWI0nG6QqEdOiuL6I4Cx9ocJ/kBIM7
nNGd5iA9L3z+kYfTX28UfMriqrEcSR96yk1rx3qLi1nGzKolwBbUuMj5wdCsdE6r
U+fppL9D0rXlvkRf6cjQf8RYQoIaX+xtIR3DHW0gx/lw6qBWZTsvlpIikWD4r2mr
12a1OxF/7eK5PKmgdeHAclHbklLqyh4vcqkk3VLOYxfMpPF9LpYHY2hLe2aunGBA
8+tK1hdZVFr+pU8N6ATwKpqxaVwFkYivBgxIzZFITC3SOnGFupEYiDom+IJRIzgW
chbjlMb2FiUjCk4yS0JS2ZdlDpNjf1A6p02tK/50IZkBDyyQq2j1IX3Xg/BSfK/U
ExJ5s9zyMJTnRCOHnBC28HQmi8ZQYpWp1Rs89w35g1SD+GBUgYjVtvkbXUDjih/y
QKcsEc3Ini8uvwO77TAB2314o3vegYUj4K2Obc2s1oK/zS3JqXlP4i5ZZQ8aBHiu
oS6TPAOgDcWEVCOquq7vuGOVxSfAonMsdW0vjjvNKB7UOE4S7jXnB4ezQsqthNxB
6SJycgnplZcuhyx6ogYSzzKlathfP4HIkaxUIEfDGjpPohz/QU/7OPocsW8XeepU
CJKJuDfvalUIhcQbjVshw+JFWeCG39t/LWXUQXb8NINyx2e3OIvfugVn5U2oezqm
gLNu1rhr5OSGVcKMwrskUghRwM2CGqZtfgUR0EBM6PD6y6UqvjjTvILEVBWsnGaK
PYDradf+/88vqsQGD5pEo5gPqGIcM7ixcZKy9O6RmbYlLtAaZ6Gf+LBu24/FNVho
0RbDM0I8uHpNGSuK/xq12FvIJ6cMkJVcAhKuQmo5Wg5WC3hWLRXSDP5/Zr7u/UjY
++d0T+yN9WXteh/D4zl9NJuJ1jGdLExaVnuqkRk1l1dXEuXLxQrVqa5uvadm7JmL
zMj2s5rPuqsYgnXI9RQhRdfeMc/SBGzLcgK60FAWp18HGCgI3eKpH5ppccsbWxvt
D/meo9LEO6txfSp2sYSdVMEGRRQ7NLDdhhFZ5jxIdRZLkpIn7kC8j4vF2cBm1bL9
0ZWEPhds2oGkxfjpwI2qa2t2x+WPvEkP37psV1gGbQKNIz2XpltkHnptgQc8k9dI
cDHSTOKbmLzXPr/YtGcNGIIRtMMZZAiKmauDBpaZjpvV5bpEc5rcTTE+algP8NB5
0IXbdB+V07TucvYLOHvxubKGiXNHhcbGTdM+oQqM6fxzNQr9ftcxh/IP43HpFV1B
sDkTNPrZuLeHFnnkacqqLN/CAC6EATTrdi9grs0YRhdpDc9GghJrq+a1c12uNOwK
C1Ronf74Eh5guvE0vceESC8jm99No1kyW5qlY2NGlR6AvDBsCDraiNGCVah0npUt
NAPJH2luOfSOuCOKtjLuvtRKlae5Jxf+9tA9Ui/WizMP0by2id7ROclTzANn1pW0
iSkkeKjrw0gxKqrXIOtSOKzYW7y8ZrBV7FUXya7o5lCKrc3NgEYlYnlnAeVpU5Wu
QTEuCPcItREpX2n4/HrDzxcnHtDs+ee7vYgX/nLCI6G7VSabtZq1UL3+YWlhxRE8
EVeS2QSX3l/ADeMs/gKutfOnWIVVGqICa3rTyZLKK0KOhjNPGnGi9cW7q8GSTHCP
9oeK5uLHA5tdnUX07IW0Wke9JZvOGUsSsYopjrl+8CJfCWEaf78BgczjCDC2fRG9
GjnnrmQnYY0S12Rt4PyDrD/RQV5iEvL0+v9/NLuuerSZ2nLoNNky4IAYmFEfUpPZ
TajpnqKfakLGBAB4buA4NVlvmyHGUd/LjDPe3iAEK9on0Bzj20IqcAuijclzvp7B
98T3KVsuVDjxQXmym6jQ/Qrkpwgco/n0IAnCyozOgltcU4Yk9Dv740v2DaTPsu0/
4fagn+jcDKzx4F7pTGgcOZpCcWNijo/1yaJqPo760NzqjfKRfSEa4qffc2s4N7HO
0u0YsCK9wnPv0FW9/BaBi9/1EhT+a4LcPwDPe3SipxkyHGWyylcmLMyraf+JZvga
ed0R4IjumWR2wD/U9YZTi9zxsx2gzm3YbDKDINSvw49bEbo+1g/l8fugr16x3SVP
ecUnZnHd7oh3W97c1IPY6LWrCEOxoRrmK0/U+nYAwxsh/2Cs+1l5BPxsKWvE2LAe
VglXPc2laNe9G81QNdj78sUxmhslV7NC3jqHSt6LNEG5QfH4Ln1gucVP5NPIPyVM
HFDZDO/ZLv5SjpVFltay6Y1vf0vAc+u36U0L7OGJFPWWT7fPCQSHRJW0Sg1O3ZwS
H/OzJhRbHrpc0lVBB4+tsp1Tl5f0vo4MrRLhUQuzhQxfxG4BngPrFkJ2kyOghXmm
8kw/kiEWsBgoWmCNf+YEn21mTb0HaiYSHbWcxQg9EbW6PcvYsn1D9fMffMgXrmtI
Nxh9DSNVc5clmvBQoN5fN30fTue/SSBtnUh+4nsQ9GdzZZIyJjCEbuZ/vXV4gxN+
LQzpXCmsl0lCVhIK71qEVPMsg7oNKrFzsb+rrKkXiidgdzVEPJpiRqUVovS1ynZ+
mCNbykIEwDezgn+YNUu0iuoc6tkxIh+9TnUvO2p6tWhdM2rlGTxg24PYQ7o29R1e
0w5VUkSB3MioRcfFCXqkOrUcTEatVGCKvBfPOzRslNOyx4Cer5tjOrbTZ7biv9uI
WP0PT5sahsvrgfTKAhd/D47sDfRX/csjnVatejg4bWQDppgItYtRgwdoz5mTtjpe
+voMZIYxGiyfQQC21vDIY7p8z074EUYXhvKSWT9VLNT7vdYTg1rnpcM1aJbkoHod
omGVRB4J+TiUmxMql0dOuSBiQuzqQ5nRSlKJSnopmOmgKIIZDl0/1AKcwLklYy3/
jqhGeFXZC/bmhJy/+90qnd97DviBUNE9ALDaTJFPyBgR33tohWlSa0qGi6gZqlHP
lM/vIOxCxNj2Trixmkr9QadNV4SIjohsqsFzD7sEKmOaO81E+iWVNx/51oyyJCcc
wT+eb0jQU20q3d2HcM3Py1GQwuAhjpPxkEdfND8PWZtod8Pb7oskpvbXSESc2qwo
RR8HW5a+f9zzyp2sS5Iyn6+uFtQztRYJyTn+kmhTRlBXDPUNldzEY6db3yu33nZC
g2d9jNQz+b4nHDmGikdpVXHRmwhncT3rcwsF7LiNp8oRlcYxxJaQh0H9Se4JJ31i
pCMQZds+WwimNM5F3888vxWV3tIycyIlSo/UAPR/1ic2gcGMJHquQkHPpdfTgVyu
g5axajvVSQ8kRRKXWEduuLRx6w1PwEHHzjQEEqxPqtBTN1xsQvxm2cE+jMkE06TD
N6kuMs3ODGdRA2asKA6hYLqGDfxFOozpQ+NmnFMIk1x9uhJ0Ps0FP+W70l1E/j/E
d2r3gFv+zBhpaUb+Ni8vaMFf/yNfmZt5V5I9bgmQ+WydosLYkKSyAe/wDz/s2Ljc
5ohtTzh5vJhPUAA5Aj0to2iaOdyB38RAuzcBUxWqk0TQrDAM5bSU2TWJKWjUSa+J
oTdB1TlZMIWNFfJiMo4ZMTRv3IAkRof4mI/Hj52SxjV8sPzsCZFTrj416XG68WQe
YpYwwFC/x4yw2YboN84cbVCR5uwQcikGOfNgOxoe2VFvr0ymraY+NSna0OMT/rYH
JCVow1Jya6sF2sD8ojFRIbxfv3vVxqLVrnWO2raZNOyVXzM/z3OcutX/0z579Cnd
UOd332I8JBuXN809ii+aRuA6VbroMNWn9dTD9EjXU3q1Kfww1ddljoa+3GzLhN18
sd9JoB5L5w3tdOq4Tf2+2vD6udRQuRI6Sc6h9quivuNK6duZeJOQCRQVnzzQCbzX
2dlElDKlgpmkWw0j7HexLzbzf1u3uzQtMSXoJ/yxNqQG72MpveqKNraewc4y9NqF
QCbJb4TtkDSQ0FlpMzxeDBaeqQyd8mbMhIN8t7RaDgpu8gkY2uyRlQ8e6wKtGN8h
L0BnfC5YwZsuzGyRW/MZMWsZum0L94UZWYVOodZLBIloTussLunWRKuo053FgAQM
GAzVi3m3WbbN/B8gENCBLUZKT96TmTcGF8ZhWFWnbL/I4kfS3nebdZrwbqtw80Df
NV/AaybpfnukDRq3vic0XSffn2lnPkuOhxY5tT9fPxTYHC9WIanFF5839oEP2jBT
2FWSwtAGnYB3aoPFzOhG0G6xsPieVtHUftazlrROSMViUYvLxOh9iCCP7TZNFvpR
ELB2rPLJgpF3722CiGuTukWNMucKgnoULh+fQcmU3K732Y3gWmaRZrD7THKp4AJq
5vVWgBV9i6OjOq/7F/R+jh/MDyrM+HfI13veIOVvNhL7DEnbUTE+iH9x1F/ppfQU
ztSbPU6S8kFj3SzcqB9McV+ah0N527kfPuOeTFL4WobRe5AYrxmBUIF/o1y1du22
mvMTXjZavORT/AFoYTV6z92j7TAGn9IqPGnh/YChzPSZ5nJ9lfT3pLd2clG/0LzA
P31fv+nRRP7A4Y99L2hXkLCGs4/zbXmKgSjh9EchTsiKbanG5WAqeO/Dx/Dpo0nQ
lGQtNkGV3uXstN71l9aLXYuyU5rzcIpQzV7tGGKk1gFw7XAFX76eeW9Ex3ZpS/n2
JM3UGaVLbkV3/8E4bHaiOWTRazgi0Hd0+FvYjFylfcoJRYuRpV8yr4ChB8lMXk5f
cGZ1Kwzpdu0zSaVDR9vKeN8M/5kCtuBo4RPDj4CXvkZhtXc2laaofXqxLTkro/xJ
ekQgZG5POWOVr2QZUaGiujjc0fpoGNfNbzWHDv9m47grr9Khf0HKtOIx+4PJuBYE
gcBM37V+OP/EZ+hkWfW+adgTEM0NiC9qKzp7PkAXbakO6+K6S4MPKTREFr3lU2GB
JMXdHqoY3XTDg8cNyX7MNLCKsrMKinX7sR2N1MSSGohLulbfFqINx4a4Zxh0YPam
7UkyOKK40CYocJlw4IXoUD+Jy0lVxJUZk4U/br+t2KraPhfuPYbEoy3UK4epB+jb
HNd9VILU0nh8f5+R/c8c0RM1swriCqExZc6Ete20VvLYneXxAz1coBCpB4ionief
16T0LXTbVy4587itbHCHQTkRovXG6n4jh3NHx9v8tNUcP0ABPUggvVr9O3VAHuV2
c1EHxAejOi4q7NBxRZWPoakhMmtwFKSKl2nsPLcFet08G0jMtOONtivLWhsXfm1X
t5xH/6TVy044/PIsaBu8OJwHNs2Na5fv/Gq0M11uJ+4M00rvQG0tS8lsHdAMd8Nh
HRJDCZtddcWRs+cYgNjKFsBZia7p+AehtqZy8R8iTJ/h8/PcpO8q2ZDTzzJWE9Is
rCu4yWyY3dAMF58Q9/VEAPmS1R7qIgmPesb6YkEoDC3W4nqqCSH2QnNbG9vD6R2S
Rl0JuI68iib7PBnJN2GV0pyFjDk58BzNtBa+Oc4QAbRU4CxMdeRRp43BTJt9+zsq
dS4AE7zkcuxsKxDdSZGlA47qUiT+LMj01i973YXjdoA8fcrzmhvcAUXAA6UO6hl0
fPlttph60IktDiAMPLPCpbXKcFNs+wdaHQczWawHw7UX7DYaZEwCDdAKIkgatsbg
HRvRFQhxkacRSTzRzlmOoh0yaT07DzjLdLayFWfoXMrI6eB1tqW8C/rpD0W3uGWz
XeckchRkI9oEdzdekF+EeS9aMZJeqQt95ocdY538hwwJOdgliZ6qiZD9hlM4L6oO
bgDcQvJ2PbDAYee5kJusISMrOK2TZ3E3jgN3A988zVXmJupRGOVM6/BNN966mZeR
BqfUlv95TNL8MnkNv5CzQKz/7j4xRTBOEOmnIMnlN8NQabeVWh5ZSGeNqjvhpdjW
mzZs4w8fBTkrpV05T+g/bwIu4zfodNHfU1cxqzZsYaELa2pV8G1DMXDMoKT10Csb
sv6xBN9Md25bRsXF1Ry/1u3p+UR9XIskL8u2HshHcgWEsfb9ZGzRE3A6F6r4JJVU
9ND4QtNXxvvvsO7W6r8GdT6Yl2y7vPzly3NLOYJVJkveL2qqeayGDr+sViF2YN1J
gl3CZI87L7BnBniLoRvzIeD2F60bzEqFztAPgArRVZfAav64pWBKXhJDLN8zObtr
5MUSaj0GCFvjVDeik+mlHlQbFS9GUr6ASYzPYFoSuIL028BiRsh4KAmJL0WTC0qf
yzhSpGeZAEufhPYXgRgIVC2OEUV3H1DWInqYv9JRaRQa7H1+8UWY+IKI7J6IWKKz
6yOcZ5/DmL2M+6u6JQWq4lVSsUqsRrZnjxMVZAQ1MZzm0mG7abu4UKr+IrUXvhlq
dDYTZYjFkWmih2hLEYJRFyvUA+3JSwYbPhdoVzNsZplmlbxnUuoVclXRN5LBjiuc
Jmr5kjw44+MYtamYu67UfEYbS+cZCPbVPh8yFSuzsppjfTui9/jo8J/Q9vZ0ORVV
jhfh4liBy6yHHfWbNTs7rrRVJqosvIWP4artyhU8txi5LY3Up/2RdSmbUkedk0/x
PXNj6CWnoqZ1Xa86RdO8C+ipNgb9t8hoGfSrA4m6iJiMIGe2SODinJa2rytcLW12
bCMWw3q5BBdc9UG4ZzewS3uyveITqmSH7dYyKCBC1J3E4+tOLChkgxSEpmTMpBTa
0AG/xuvTdGJK3FkSQdQUC2dN4aGrJh2itLV+ZO8xB5u3mdehUPbjg1vlrDVGYd1j
sc2W2wLFijrAWNLpoEVzK5qvCnzYK0IItzz2plmVmfxH0kzstQIFDH/5YlFiiq8X
AZwsvgIuoS6FlKHujF9p6soN1FKaiJv6ExrwaETLNzXbelNMdl32l1LrL33f7MyM
lJGz7tYt++7N6vwCTsrPqBzgCif2cj58LiIk+HNtkb3/xfGfds7BTlIcTdHcXU4z
WYQxf8CiGWJBoIyuClUmyoFl6IllVUskOBlTp0wHJn4xyk6aeIdcf4nbQ8WCQBty
6GeO0rBbhMNrBY+jgeuK3uPy0GkSioyk+0ozflCUzoH1YJmcvsua7c0Nenp8prjl
hsRCFZqtWW2UphVb5UO8AfpIoO1D7hageDs9c0MoBlePqzfbnTfLm5jVRb+v8R6h
EF1hkZ1Aynk92MCPB9h7X02bKn5To0Yg0DXMPo1DUcn/nL7woT7HNzd8BNTOPNDg
B11hL8iCLlJ8ExsOf/7/QUUd6IsYQYPNlPF/0+VB6XNF5szTiVYgvA9o3mRWfGPj
nIapLSJaFTlNO5xTKWjJr3BnQP9+U2hMfIJF8YB3TGVNB7SD92v9Qm/bfYiFN2iy
6vJfkYgrNEH90MfzOZc46T1N9jxwODz1a8Rd7IkTr17Q/xMiqzsGtQw+dTrRf0Gq
NhmH+wPTv6LsvFPKnLlvMJcYOgkBctLWGeM+IWutr4Rl8EptzeDGiCOaGsVwSvrd
XtzK54NhENR3KiTDxSGnIVc3oc98NX86CRWMGIcSf6Eb1NQ/Caac+OZFPb4sKhMY
6XjM7PWSFMlO+h+XFNyQEgbARZEASX80FiLOtLexUwYihyk5jrmw5taWkeAeKoP8
/O9+bUxD/rCmjwbG5BYOqamFsbldy0lln1pJwFZmyKWo6Jd3rBYeGWpYcZ7IK/eK
v0RHTGGP7ix71VxZtsTZP/N4sGJf5E8ZIHgn/+nxarYHpgqPZT7kqUSJfQxTvuIV
xJTkfAL6ZtNCyuV9KupcSqi5qk6alcRQLuGQFZmylrLUqByb6xyBY8+mFYKMhFEt
E4JPT6C+Di/GP/9mgdj5a7OVWZ0sfFzWWfZWU5PkdEC3I5UTqDbWHIJM5qdd+26P
+1px5bnljp2hJOVCqKUZg0hBvzNjlBT1S+pWv/XvFbqBwWyIq56iS6NfHKfPwabO
Is+cpnw0MZIKfVG7utsEPgOnyts4pnvPIRwVsviOL4DpKIoZmsSC6l4O6GbPRkvk
QJYFsXjtbk6C0ZjyGPDr6qkc/AWJXgVdwCdq8VD7Lb/sDAFg9oxzMiVSO7wLTEmj
SOWU0kvZLtuLqBMVMHKXambgXXB49QOBvnSNd1jp+O6cpga26x0C2BBFV0+ttCed
ZyIuy0/SB0jJ8OzB/i8ikNQSN+3RcQASVT+3TsBntSYeLgcMxXVfOXeSIiyHQCr6
piiF0l7epOGzzSzECeEI80/HcvIn7+jXXcXquHi0R1Wx1iQdbfnLMQYzuG7E3RzC
Mfea4yPK1ida6PePbJpbxQ0SrKkAUMs2DMf61Ye0A3IUhh5Rqthza7IJfaYhwKVz
+L9evkF0rgxqMaxVIKoTF7bEbbXDD43xasbmAZ4VF6bjcwdZ9k0OAS/4wSFTk/nf
hdhsfzy5hDSxePiP+iLOKAohXESMMoyCiGv9mukXGINqeElaLM80PsJRGMKGsanR
TLf4xkScIl6TLWQFynYV881k4MC3ZqADmYp9gxTxiGlTkpAAGvQ9VBs8VGFNZ0hr
Tt8STXEx+eVd4aPvKFLr5QZg4pVJT/fYYDLbgzRA+rq9hzQX6eo3nqT8H5VSaFUO
JhXPQ5mbnxhN2ziBUYVbJIfXzswMmSJi2ICyV7Zp7LaV6mLSlkmdENW5vee6qSOO
gq+DtDZxeT0nwCIdGJpjCFo8qeHASr7FWWI4tC2sfZA9xuT2F8CuwR5/Pl8+R1he
GF1RRNKFRV1lw3mPZoNV6k6nWSl3S7fDDJfk7Fo0j6g9dAFHaOdKGtieuBoq3TdY
izIHHv4slBc/hMgFuq38AlfHqLDXF2WRFf1diEk44iicC6zkFvoSC+MuwTD862yS
V0zxdgKf3EgL/6ZY919RpIFDIx35qov0Ny3DIJKQ0CwRmvi+H10Hia6E7ipiC6o2
VJKcSbBJG29xsQrj4ML2r3hoCB0csbUSeTqaLaLsVZxNjZE3DpfZVl/8eEmQwNZi
qBzvXbaaXMeMs39csCs9c0rh/qbcur6mRP4L+T+2PbCHwuhhkiKBIenWubGl831Q
TpWe5BDgJnjsKZyNXdR76NeKNjGkRBBONhADaW59iFbV6cBNrfrc9Ey5+Woqf4MB
oT/GI6N6VytH2cAPv7+hkWXfbFngCWKWUcDZKzCoY69hy/rG41YcoKcSuA2MGmhY
fY8OrKGGfUsjcPuPRGvYxABI7FdB9kusn9weK9e8SJtQc+gAV6zctoIxjeNZrclH
ALeobpLRLh27IsldsAlb97+2ydgct3gwbTGUqhvpvZfJWUw0ih5p+FA2mEt3Ji6d
4HkWOTC8wa+Of6Uj71/C985rHRM/rLOkoAfOE86/d7m8O/TNj9yDEWEyXCxjmCC3
97huguJyG114Kn04uIguNByV1MydxwZFUJaq7giRQjW4hutPv3Lw12TuNRjO0tMX
HACJC/JGuBP8A9wAHmQJ0UNSYSBWPQJFo6K0OLAO7vFgstogNx6jP35uR4k3VE97
1XWYwF+adydX8VevAlTsqEMJrk9MzAVQaXXsGnmGo0xiOYr/y4is0gdnxIsvhm79
AjVW8mCYsG54LDdByDAlT7CZ60CjfjsP2BRo0DSJ9L0jXnrPTpulvP8tSZEW+GUd
11l39dvMoPN6UDcn4BDj9wdD3OwGM8Eglvwj08tm04Wy94JGwPa9Y/z0Brdt+KmG
571N3g3Xs1bE1NPhutW5NkTey5B7HxnAXbyouozxgFFwqmWHzRL9SbKBLSyR8sWs
kDEERUFbzrfuJYk/XAvQEvbp2YvvKrLPt617SWh15ccteeW/D5jCzp4NcB1q/8xR
fxbYO5w1oISnsi7lB5rpOxaioFI5E/waN3Dj8jjUys8tOvcz1IOFJ9YlpOjfdzws
yVRexn25C3wRT7PyE5+qWByCLoFH3/NQufKQjt4e8+6KEhWeuSdfs2FpboVT+kMY
BIL/o5p6CMbrtU0vIK8UTcP4R0QZiAap7uWSiS2JSxIHha7vlekOsHi3FvMO0Ifx
36WXkwVwdKV5PsitNBaM18Bdz+Yqer18UTdr98RLt/3BfiTd4AjWb2xZtCUjI2SD
DAbHrwAvg+OKHbKNNypbIcw3VIQWSTIG2+QuR1egeo4LDEwMaQMdqhbODGFkBg7N
8tFgHFEwksVsp818A30bojo+Ch+8yZMt2qGn858O59js37UJNjb34w/CPxSgSmac
e1AGqFB4Ll8TLTdctFS25+U+8AKuH24b8fG6w4sLp5T7XS4EagrMd4dpBfArZhKa
aJEFC80ol3dOeQoQwZv/V0lRanBcarm4OE/EX0umKcq0GD8POpKPs56KgxZZ0Ihn
qceCkYRT2EL/07GJIHWA7hh9tdZl6dYI8R2oP8kevSflc23QCJc2vCRfLN/EBpCP
PfhDkRHj9kazdi95PqMjSTumSsUCmQeal1qGig69ZUSAQJp3sQyu7csx8ir8iQ1U
HVw0kk+H0Gvvq2W8vHWAMNb9AcYXSN1ecNj19X2Pz9gOYuXg2qJ13J7ZUuNw+Ldi
doxZ8WCeMm5e8EAJ4rdyFEBucjAHNPz06Ui7r0K4Uy8tOWG/qD9ogfeB337uvE/U
6w8btxcsnqfhfALsIaxD0B5XJAVZqw2KHfQ/mvKrUO6si2BkJmGF0wFzOoux5xWu
erCfPNYMLCiRSRo4h6o9SpQyPAwbLftC9At1w6u/ChGSfiAGPts3mAR681e3Uvi+
gs4nzBe5YuzF+Dvy2oPuZJXds2wo8rThoF+i9zXy1GTtq57dazXSsyfsd+z6p3vk
ll58NVTCQ6soyAJldk3fS7oPEeVaCu1Lgr7/UUm2opghg1/UqWmeEvz+Pq1QQN8y
3HfgTSM3e6RyaTy+mlrnY/CG5ovygILrJpij8J/6DG/uFfZc82zo1TFkKKOAvbrn
RsPR57kXNuU9UTicdkYliMaMhxBYTlm2wSEpkCKoLTZGUllBBrvFBB9lqofdAnal
NH9b103TocNDSiR6N4E5MERgOKiALuZA2loj9B3ZaXw2liaHltoYSc0GajT74aUj
2i6LRDpp7zzQBIf3O9YvurmVQYrJbjYLwXOenu1g2DAV71uzIiToCG0Dlll5Hkzx
PkNl9J7NejeGK/K+WCa8sYRkQ3Z8jS1Gvde7KXIHyqx3Hdxg1DMRyto+VQrGfD1q
ceKaGMgtX6MH37oIewSd+bB1/Mnktijvx0ObGONTLmWffV97+Qa74uT05egDJMXY
bPioxnK4VcOTJdhu6i99PHSWv4CVYAljDHTZkGOUMW9OsSbAQKgHNouGc8nDzJ84
37VCt5TYhESsmoexLxmEcVviSxlhV7alvJDY2VG1NPJt1pCDDrY05/aFGvN8RjWA
bcadNzTIcyqNGfknhThBR0cNzFfJ7yUzSf0FIrRWg0TnGfedZEtlwVneYlEyiSck
bUshEZ5ENqNHvLqN/vpQ/2GNwsX8kHAie/PhS0Cx7MIL3geWHo+KZXIZfA8aHIOx
tphh9hNQZvF31pg1rjcPX6CFug0mBuK1w8BONHquQEqWpLF2p6pTlqOUWfAvU56E
B5oWIS5wxHykF0vpeMzyb+Crb3Kr574DVRJNEGDGWY1T/LF6Qw7wq3bQvx7vwvZJ
e5FVIIRyFThHmdxQGaNxS9XzMsJ3amaqrlo6Y7HvFNJe5hR+sUlgHJwVkNqzJUuB
3Pu8cvY5RbaQYXWFB1NQZaVLqMAMM64GSz3mFChju8H1wEuemNvt7ws+dGBxhBvr
m7hi1C/8fFLGzp03Uccc9I1+Ku0XyBsyoNfUXGGBzxyHh5nrAWDn5wpvs+5HmFl7
P1r0/tDpgMTQkVQ9gv2mvBSYjPn+22OnHbXVBT4250GxnWtaXn1FQ2UvbrAWVdCE
4nMcVrAhtwZ4F1ZFwVczTXt6Nxg8+zumk8ErydmWqTqOaMRluoW97AkhdGBfWJaC
1dIDkzoVyQ7wyoMe3nKrJ9DM+03wr8J7EfuUbLGsie/XAT6KSZi0XJVh3n/cfDS2
aywrw+4vunBnsrSm7rcblIUdwlSzherzpw+snwwm7GBZJZdiqGZW5d7xYiN980xB
L4FGg8WesCWuN0xnWO+aPn1zIntmW37pjnLQc27aPbmWXeB+sDnFA+z31Ix4BYOr
RHdb1O+fPpC0/6uCpjs48IOM8zBwGPA17kIu2e0cES+JjoD3X5r3xDrSwvnVHW6n
xG5OIfy5Hj3u9kJsC41vAQtCwdRdUPQ2WUVuiZuYzeq2t5SZ23U2SXuQT2cx+8n4
t+H3lZHfpaIWWytT4TWoFoZePkGaapK+NYwnzpf86K9oCLvrv2+a6XJ3jHqGggB3
0yzBqljHQ2F6Xzh0ChGhOX7cmAqFIYCwW3qLcU6z1fY/oXs75EMwWnDICQksSh9/
9sF0OMwvt0tVH7xMj/7n5DvL2armjfwrAUYAJiR2AHDofEJCKbIlVpj1JDeo5dwF
xmH2ax4YgAxQJaosfblhGoDAdOw/r/DVopmk8hiEp0yHnXk5iWV7Y7XKVFUz0WNX
ZMGvQpWbtKkVUXjXE93xL3MIBh9p02haIv4W2AwaWLORNAU3OO7KWpXOW+jPWuCu
jYmBAUTADnJEQI+QsIZogFdo00P/PqFdiEO+zbM8vVkUl+j+8hc/8YoMo2SbovMX
iJSy+o4KCOo8QcQcgxd3x4vLx3VW+vvrI3GTCOk2gRQRUqJFI2pOjhpRla+W5CIb
SORfjJgVlXJ3oF+ROkFYP+i+WxkOuxawzN7KWF8ikerCtPcbXEnCEbbzHEJ/O3nt
XQJx0c8B7VDd1TmGzgLln8WQlXtbZIunEvPFj5sD05jB22AdBzlVToMQBXVzAXj7
NYxId2Lnit0exZHBkLqr3kK8GgSwxhW1CUkBtbtI++niEiSvroYsJ2NpObDC3nbM
KWmVerKolCzdtU+VAIaB0CcpNQkNPtLYlEaUQUTehX+EjXdVvm25whSy15B6zYh1
8hgNuxETqkqd6pXJIkt+MHwSbfBZRip6G9j9DYdywg+wzQwfKAkpwtLfdcQwqh+n
r+RUS+nSerJlt7HenFuUZ0HkPgUrv4Gu5u7Cq4NT/Q3BDP8lY387VJJer5RLNe/h
GnSjPmwSjZPdykd7vIbPKTmww/yE47t0mmXRrfzDEJfybyQqhlnRlj4Tj4kl/x0h
WOOQkVz1xzHt1R8cB59ZRpOxPgXetvfFB5kOU5751l81Z14BPhGHP3kVG7D9Nj6e
pcmqwHxoqkvvP3QisX22+IHQHgrn8uUPUlKRdfg3e+AYWE5crKUlqIRGN8WJ3vcT
LnkVFqbtsqcp6CES/DSgNgamkZSEmRV3h3UBj6Oe/8LaxkYov2dsNFtm4HL8a+AB
hrVh7pDDgx5gtC2Kbf8XM42/ZHqLA/tLPyHwmCbCpGgQjjSg81ZI0M30BebTule9
8u+/rrajvpaz9BkzG1Fq4zRQnUqQGOwH1WnxbdRsoJ7U6CFWQZegNZV25A+FMimF
4EmDG5/DTM6jUB30d1BchCMFQZggAsDERihc8UfUyO3l14RB94hupNkrugO15iNI
yZsoECGhz3UD0TAwb7IaPqYtij0v0ASAi8CiTnt1QT/V6873pCuPc+6pTVLQzBdM
qVsr3ZSeSCwNDIg3DQoMENxIUxOgFBCjzRQQe2Afkh0KO9NYcXeW5RVpYzgcSmOa
DACJ4ZRcVYrhKSdmVX1JNB2Dc+c8H4RxzLRNsKwwbOKA69pAmHC4LsNImCd8KrDj
T6ZTPbDlToPyOZVXl+rxZBXzp5ynQ6NA++suV6HDdALeYJ7lnkdOW8TFs0QNk8zi
X+pGPsSj7feu3MW3L/qtUdKcw0cTaNBLpMZHX4YClt3HuxpYtOMi/Bd2XUAoaROf
IAHQZzmDogFUy/tbqzJCbC3jUkXPvFPgqdDZXOt/aNRu7WyQJya28Hjze4giDvo+
qSPPCdUGTLSIEWVe0VLbCnme20ODmMWidJK3Lwj+ok+ah1laksOnR4lJKpKeZ2Ox
EdEBMIvrcjRuwC3p+jVD8/FFxs8yQLFahPDwq6rZUeauZFNYG8w6Ou1hiljp4s/Q
HOR5lKc7dz6ZEApgWlCxioz03K9B+PFhPFc7gmqHPt/6HPipdmNDhIB+/Ro9/Pbi
hHXvwBLPp0pjxQJvirWRJTfVvaEA7HmR3pAgGMAHHRnRC4qWoTH+q4FW0ajyPRxE
NiyICsBL8KG9RaVuN7w+8i0aBQmX1HhIUukfVi7lGdA9Qg/9YbXumRonuAvl3jLf
MwMmrcF/8jTbmjABtFIivYX4276PU9QYi5mgCC0RoeFzDMvXMba6Hjyi0nm4iIDO
ZMhflUuShROH6NeMWNTEToi7e/jtNqdRIeeYTLXfESRbKbhER/nN+vV35Wq1quYl
8cqZVXWaRUVuAI4IXvBxz8v5JAe+agHaw8upaweFUS9XclWsRAA/WzMPKBxC5g/C
w9AZIlevY8QJ3vVA17xa4+xzlRNTBd62JPAZUz69ElkdlnFIxFZ7HY0QMk5OmpC1
jA69ynQyEsGaq7cCOPQwaT22Ww/GuwkVY8Vy0LUgS+ynsuhTKQxUrcv+bn7EZzxp
QD9sOxaWMXDkBbApcUKMp6qPUmCJlVofgUAYtynFFyHkHqjT5bpV7MweViPxycfk
bPx6tZocKvsUPGLDJMW9mK+1dupA6YhuHjBmChYzKHvBHd93s3ug1+/gFjOw9u+o
O04h2/nOU/0QImhlygY4CwWJOiFSWm7kZd+QLdP9fkfjXTgneGHcRZj8fKFj7B/R
xNYnvYm4gEzfX4L1uIhqtlIk5UiFKzSND2a/q2VyMM+CVP4sCe3ALRaBTcuXmPGu
/tbcUK97Qu+ros4YMLgA0bryzhxH1oj1dAE1aN7IdwVtLdE6sFwE9796ikD16BWS
cU3BpKMpdq9VGk2MkoZ8HpMdACExwczxHBDbgxZZ1Ul4aoeZaMrBOjHGlmxZqvb7
9ZCRnCmSZWIObLMbKqxhdprfbwSoBDI6q+QyXrYl+OlLS+4PRkbuCfyndk2RMoIF
SDr9Z900J0WfVMhsv+SQxz047nmS4ek/qBTnY9tr08PFWBTpaxIrO6CzW59P/9GD
wLN97+o0GG00AXigHyIClTQ5FdEXoLrv7X3sP0cUY6ZApEHTiygkDFh7xhM7c34V
P5ypKzKkcs6HbRJ0GH/3ba1vfxJ3W+3vIqfW5u/r9Yljmu9fvWzgatpNURDHbjeC
pppmXC7gb1iC7VZDVD7bn+6nEXFPY3JqlJyoX+gZ2BPcwEiJq7oorSxaePR274Ly
s+IK8VmxMvFsnO3m8TmDZw+sBf1dlGwfNharJoBUKN+vLgBvdsLkib+BXw5u526L
+UocTP7/xpT0a+0E6sFjel1GktvOTj2fAuDwPDoT2UKi7TWqgnezbqZUIQLbupZk
0OgtyOws37aKCd1PCKXgiaBddX4XrkTwLXRTzdxOUlqkdcUZ0R7osLc7DV7G9EXb
SOtGAPLmKYWZXHXqT27Rcs867DHzJrx2WLC5u8/UnpP0dqWOF2AnBt42uQvNvK6/
ynYOtZ8Olt3D6BbTSjkkn6zRiSMahfl/BbqQ3FMdOxMu5NjKIwrdp9zG9NF90GDf
kmQdsCeRVPwEyTqfizdNcmvmB2a4E9GkETOZ29WFQ0KiPRs0ZHAaCZiumzlwFwro
zOjAwdt35BfdfzAmRn0fbrrfGIrDK2v6gwIhWSt8vB/z4Cw7CntKbY87KCrhtNXd
XAO+l9D+7Bg1aClCa5NZ6UqpTH06Qh2Mo9ppV+gU+ZbwslD0pVcgD5uQVarAMOBO
IgD7gUaXYpm25XqzK4woUJw3A1Yf43bCC6K7bU3cfqZ87RfVll+21ioCPjLveZ6D
m8/cdurszdLTgewckWTtybu9GYXqLeH5229UyyhSwP2nkZgwgCORRv9Opd+PVnQh
uwBqpSBPn0PwnYlVM1l5KOuQW79rhwYc0gvHPlgEjREtcYc8yfP19W/vAuH2FsYs
YNgbW1Tx3VJi/IU6RnRMgBxp6SO4xP8qYCZQrxHPRnU2A6yoiDH9+B4ecvmGt4KO
SN2ow1THaJoIdFdelsHBOcTJgKnwx7S/26THAdYvlnw8o6efNO6crQ+ohI+Xkliq
hhqI+NlF+oBDk1Ubb2JSeFfwVAva1J71aL9ZgTFUbYgAHIDfRcUWzHOGKzlD+MEq
AbiKHrwiTJZOO0zGQ6lrBZUzfXQeZXIM/HN8R9wwZGrjH2ojEjlRChCNU3R4g6E5
B9hJE3jwG3TXmDdDfg8xtLcCfoUvk2Xpy1QnlfTV+IQ/a53WjVrKbWnRwigo+3nX
si2YBdNFjZbKn39DqgXZxUXRPaONnuiSK1HajVArDSPwbctWJkcS2d4ZydaHjmUU
4a8sgIKfsY19T9ltweUeAfb5/mCKs6QFeIhTdYLH0sk5iQv3kA6lSffL9g/LGpxz
/6n+/cYL1ljdsf9nAsZD7iKvGccVpgm/tCTqzENyfi2ah+GzQhBZT3E05nKmqBr/
nBXuIZDp2006eK1020kuaczH+jrqip7p4Tj5CwfNrrXKWuG4mY/dII5Jr8jXr8cp
6imqcBNVkNL7mtQ6Js2Zs/Eqz1EDFomT4/hR41ZRzpUvOtve1cb/gpkOt2fvdY6O
X/GwO+N/rjXaLMoSb71j7lHRN9aFGaVm0pz3jE13sUBTFLIAxb08vRC+ITGfpvSy
LOdhVhflF0M3DPn2SbV4Dzt9QHS/Or28nYiu53sg7SgIzqKFoHPRlgd3yRM1o1NB
iPe2HbEd2aA2bNHPZvYp3u1yh6sDjXZI3uDhHecNXfHyIM3nGbJOuoWKAq/HSaX7
6si+sJxAbLxwaLG4p5jbxT4Hjz/bJZY0SEh49YXg5QGY5c/uEM3Eu3awIJAaGxU1
TsoNpqHFpEzR9LDzT266Ro3C2ItOuKJQam7iLFqnYkF12YkvX9gataU2oYsgJxtO
GmMEFViSdnqdH3E3M+DQ1/37rYx6GToWrTMztiNUhoG9Ke5CkQwumCxzR7h7AXAB
AaxRpCnwL/01gK4hwrvwe6X5JhtelxuLXC3WHH246gX5AJCVaFeZT4AtQYpDcyAw
SagM60pIGPEt8k5NRqf1hbCIfgEJn4jPvOApKo1eG8nN3/u+ZBJ4CSRYdqSIU6pn
hda4995yWNwvHW5aVrmkb0e+Ydfl5uBtCtzk0Xk042Nsc+eMHSAjdHSi3BlJ3TIn
9Ph4QKvTugiJilK1Ez9xq9mMr56RWBQ8tnOIPirKrlsVarduXQ1D41kQCbriC23o
UlCLNgvRVYCzizsDt/36su9EdMZ/crZIsmhd2zvrJK9a9jwI5Pa8QygpxopfGpsL
uGKuqNemZJWCVI5iEOCLZ5FFfGyVzIou/QXr/J62EZsusgvhNb2340wGqmCuXSPP
QV5MdM3Im3D6mmlgPFOgP7mmmfoRMHP07sFnAU9LgbohzY7d4aRz6XMiVfHnXvhs
uzZ9n4kUbbayQb9chd66B7h6CxVgC3DqYx4/Txi2Wv9wI3JXHchbPieB5XgKRHF4
8zyahT1SyO9DvPvnFZ/RMxTzNlvejAT8B2wYtRlUP5dmET8F1Uw/SF+1SoHWtSXk
Es3rWKbaR0wrDWgi1pRi9TMPlN99frFspLSCiq12ypQDv1vbs76YSAWmk2o3kME7
dlYLJZ4TIxB6lsg+LEcBFWlHqdlZXXLldDMVfoTqvtXWHdheAp28pnXRiOulgNN6
MmPl0p/ewGnWXzYg0Eb38u25BfwpUz2OVlCgtj/8si8k49X+O/kQaFiXcMCLkDhI
LA0vKIz5reSI5XTNvL47lOmLFXmGCJAbvufBCuhQxFuL0E8zVZFcvzToXiSeIkWq
lRGNXWjEX9QKi1zk7AeaJee6/s6qcjTnyBdVDAwQmIizrolPVEIW1NEyFrbKujBE
6AW6rI/lpT9ct12nt5Ddac62eKyIgRVEssuUZGdoUn87QaPUaQLzQCKDF52nWFUy
QUI62e8Es/hU1c09H29BboWpoTgvWGgB3tA95EIaOVix1N+bEhHlzdlfw47+vdve
lv2Cp8dAji/Ttxs2lAkF8Vf4Npzn/M6pvwIIGxhtesdOv+1IJhz6XnjNpK/7cuIL
/XZBkWuAQmSVIDhU9YfJZjuqbLSak9AiPuYctIY/qPzGN2HuSA6WCzFsJr2X3Z3T
UzoEN/9VCg4CJ2RCGRXzwFYfDykA4YxrNpsqPxRPfIoEMO7ErVD9oxUKU/1xEdh6
8aRJCwzJsdn+v8ka6MpUagSW7rDKFoVpM/p7ohdmlfJcUf0PvRcx9xUvTynsV78B
fZU+2NMQyLISYpRT52tqLvdzs4BB/SnW3LHnrTzTJpJl4owk+WsS+pryXydRtXCI
4mIvMnxrYwp6K3x0y5EurqYOMtfRiWDMr87Sowmw75VSc7Oee/RPrlbnGlB7BRDq
fN1wnOAe8DBcuiJLpIO4tmOFHs6x8c25ClImoRPl132+s4Rz1TclKL+DDvSNWrOp
Q01SgLJGRjPZaxEkEvTPPa+nzROVGdo8EJdykps0ncUB1Al7GWI6md0Kv81wKLF2
WyQpKH5AwWa2xUKgM3TUO8Sal2AcQ/bhFn2bvzwiax5Q8nFrC3a/0+MvjBYbLmLL
W45hB2mHn+UxRGsRhOzXe4je5W70VUyW4qAUQdRI2LHVaV48FE7Fu1vqhY7v6Xdv
V+EKOGVcN6xPhZvsUFfz9VcJnkHd6RlfN6WM270YFjNSFOzAMGNz0uHiYdVrTp3C
AVZjt93kCZhiMwff+4bBYKVBDVKyP5KWdgTgTpCTfR6p1yS8Et1I3SMoMidX5yV3
BleY445wCdFZSuYFQmUiwKqjNzuCTNFjdVuVCRl/tZrPu9zY07GYuEMC70xWmVkp
Y/mcfJQILEKXBvROn3ZGZ74qsEfwUVJ/2jxLgMM4V10QqBy4xHTv32A3EC+4BSN1
z6/BF53xRQl/HPGDKeIhr7OJ46yGq3um7PnIEPfJBVpkI7+yzwhKNTSoriFMhY7A
2AAqzdBagJ5IJSn34+exBZJPklf8IP2JjdGlVU7R3WFO+BrT4P3HRF55+TXo3bVV
kxF2AT7Rr2Bx8u6TS73MexHk7sTx6AI3mf0ZogNwef6b//I1rk3cUeMJDMTKmZJ7
Y4b6PY+yqrn/lKeXXutbxNyiRbq3Ltoi/zcaZpqpIP19SUPy0HNZfE7zx19sKy4L
lvqz2OAbpkz5W7Suf6r1U5dHWnEkExh8eEam2FuC5igQfbgfoRMtq1jmNS+Bx99K
E38Zi7v7t2XVt42YlHaY7Bw0opD9rBS59l2nEDml0zk4PVgI2WXExG98Ioqzyz+W
RocFuAJUyzw7EcojLDUGoaJlxegOL8ax1IBiQ9fbUXxQTmOQNYg4gwOrCVTNujHU
GNF2oAeh0oMcbKBuNFqHS584ocb3e6AruwSG5+mJjJKhOIPvFIdBpybEWzBlmI5u
fJdmMnQv6WLkQ3MH8kZ8L4MxqZCczxP+h4T9+MRrJCHgtenmy5TBxhQRCmSLGWD3
cplTJLcivza/nT6R4s7SM11mG7Mm9KEn673n0sxyMxpY9pz9Px1oB0Py0xBWMhho
THPOH+BueP3utITXfaU0jOR24Zq86dvaCmCpBQu2TimprCyigvcirqzIwVRrRFD4
/AEhpPVF0qHr/TH2PSUakalLguog1PK8+Fh9w5R5DR8G678M+7p6g989RrjSw6R8
XLKww70KSabtQytYs5npYvnF/y42zDOjg/BERBU1L/eF85MZbdaJzfXdVLYpjHsx
5Zmrr0Fu5d6oTLI14deVncWib08HqZmjHGEgyoQ6eZdrIi+v8NtTAWjMHP4l1E7T
mqYTqCpVs7PP602GUleA34ON1MAcSRaVpHZqAzgPuHE0qQlS0a7LefG0dE6EiSWk
r/XTkiftPy/bJj1D7rugcvmEPvS8IIkO4RcnA93numn+C78cuHnw8/nXdRz7VAAj
fDjhx3x+RQK8MJUyDTLO/llS9AHlaYEz/iwRaGhmCIdg/YSMGNb3w1Ifhxaj8a0r
ZL1wuZjfEd3GA5PGjzauwYes8SWzq5+jfDMkeoI/f56RxCg8IsOrogSPMxPa5bSs
Y2JULnVmQ/d0LJf2ZB+Qt+hMZy+j9ZNG1x856Ukdm5Esly+BwIewvWXdgujOVxaS
vEthF+1xuU68OxuzjXJrwcbUMJBaMRMjQbPFOENHicTjOBCSeGYjjcqyOiz1M1Lx
NnKGT42jxsoIBjnmRSpdQhhHQcgm6IMCeoZC0ZMnrfX6sIcIGJuyOec0GjUfCnf6
C6KTTWFBN86qayADAnf57quOk93NtK8m8EUvtLRc38NWLzrre5JeYN5AK2vSmyyH
hoP1sSB/+RwiEIvnbDOBZ4UbdmwOGreytoxzgGhmzmUVAS593I6XXe91L1KZ2F+o
DUavwYLytOwZBRorqLgO/rMk3a2U0HndmP91Uzs4dcr9LndpUnXE3A9xJB3TsWiL
IS+xl8OX/G7o/vdXZA52Xn+llL1g9p6mv7KQqwTzJJ7o+kEwa+emz5u014phH7pW
Su6vQUUE46Zms4Gcd9iqD0zs+/O0WIAJeiaKjwwI2EoFfxYDGC76J2pwxTAJGKte
ocnDJk/zY8NHJ+t8YJoTT9ZLe4ReO4Ey0IAYFkrLwx4cXODSmPhF2w6QPJRE7WYh
PJonmBbdqYBWxW9CLS30wvzxJ9/8arB1Rcq2u58xKkjjUvJE7pTJHlukxlRhfo5v
HTcFijcC/y9UCyxFesm2bHF/NqGk48v/LzX8kVRV6Zx2S/7Nd+bwCaosfKcNyLd4
u8G4isgm3lF6qdv/wD1ArqBA62kyOWxC+cX+VjTVWtMP3/m7VllfiuQmjYyDi6WF
AUMt+I3fta555FmIn+7Cne/L7F2auQUTFgQNqEmcDtC4eBlyEQNuXojFPtCjAgaI
fSZaBDKHkXP8PRpZRi+AaaeaMla07kH4VY98OATazpKA+vc+L0XntZ7cch+lNoRo
GmMI0sTqSWjPsGFqTvJbCaQbHtd5grEri2Z0RJHfmLHAzJUqSpcBTPbVyCEbT1iN
wyCJEsyUQziFnc8RiIBXxW210twThMlRF4RG554wZnXAnUK3FrQdVZxWga96CO8z
ToHAr/Cz9Z/lLdSJUBOyktk+ijMMNDYbX4Hm5KDd5jEjOWYmYWERygzuHk9voHZH
QHyEqJU9mne7cucY2tsKWfjJX+ktZsAIoQfUtOl2wDsGYLVwquFtymhAY921/Av7
X6KM016zPBmGEsYVaxRmzJSHHfxXLMJiVRcrDtSztxQGmmV+qp3VjYMHSKza6qKV
Hvj68RQJBF1qHD73s0CNHxSKuTCZ7Ua/X0kncUdgdM6ryef2vxQtlzJBY7V+IgPx
WdUBLd8UZljhr1cty4kZPagvcKK0h51QSaUP4FSp9RV0dk+8m0Ty4Nh2T6ABtyHc
7CyGaRrQJ4PHrSWn1/7Fo7c8r2G7C8/B3bmNAAHAhZ/aa3WrILh6jYdFc9S43mQy
7vPZvRPe/Cg5oDojIEJNF7bvDABj+w6osH2I3tPdGHpsH7DC40+O7dvQSTbXLtS5
RjWmQUgd+mlmbhNZZ2apEfGcJ6l8F51+lLljrawnXNiw2DP03E+2o0LY4methalN
k5vFs77u2+H0PPN+d82hkrnVhf+EHiwoU3Wq0Ax8EAYCWaS8kNCUA0KCdXs0/Khg
WdMNwM/F7ER99ts7LM0UBgtWFsemYwPTCmpp6w3dwEP8GQBibbXyL1hWaJ6S4lwd
NIipOAFexTitOrAAFTvxemIG8OhKigjX+qYMS+s7foHkD4AZILNTmRqYt7Vf62mx
ZHXPCWEyaFMtWu5M0VlFLlWhd0FxFyOWXpjSz53vkWjh3ISfBsi+LCYqJp82T0JY
VoYEk7Ui7A7FicToUVxkVjNDFaa+4Bp96jRfkeY2j3sLxf+4041ZLvGtztBJAIx0
B9ThI3y4eD8UmIETI6yy2roELJb+lwJujnWKlRzT8TEPPnryyP+0VpcpS1PtwCSb
46xuklnayrKwacbI/I+YHuaI71Tk/WvrCQ58g4f61VQP/yf7hcsM9UiSnJC9kHa7
fZt/xmex2VoFYm2xvijzC/k7cq/dOnR7yYK3k6FAQs+dCW3aiu6gU7LmBRNhyZ6O
koDSZRLoRw5jz0IneGLrEvODbePxQ6snL1iLkXdc5zQ3NsfRApoC/VaRd+HL0lJk
Ud1vti8H/UFlREvIeSmattSlXXWfZtclEb2O0+3BwBP/c7QP787uGYeWQzWZVmxn
wNLrCkBEqCSblSRAKljDg7VLYB6k4FRD+rPFcuUlHmqV4OQWaOrnZmiV0dg32QJ2
eKii9cSpIgbzkR2Sf6K87bC3SO3kHc8TojhpVhyDpe7s28i/D3N06tJsyYMuNXEB
9KwpA+mg8AyifWhfL9Yd32PGiQxP9hQBDicqKf+Fmy85pwa+DyoNo04i4zlpQ9W3
agWfC9XwBiRp43hQBWonfhX5acYIKAP/kFgUf+khnFx/6QP7ZVEUYoYMkgzYHjMK
mS/A464BWrl1GhDcY8dpzqgVW9ARVl9Yn7fnYRl6JEJ+qc3HPqpXZ2hD3xwNAijA
pokxvF1xKJipIvhEhcbHdNEhBc3j3w6vlVABZ4+Jo62IxvnNlzimeUfitVwj2vTm
vgjWqDNwbHRd/11lsYVRKljmdRtfyVwoa7bk0jgHBSFrikXO5z1qqcpIeGOzo0N8
UmGI5J+vBcY0uUOkXvquFXFAHnJU7QgNcmc+pxe/JYtnts4jSPlmvHQWoL+GMB1d
Y64PzlvQogmttWZL3kRBqyUONw/1/LfHGL+SFp2T4lwzRcyHEeggHm+a9VeESMtz
rKPoVbPn92K8X9P9NdnfYWYibOmxPEqeZUp6Rg7yHpR1oByYdfF81MR8fvDSllzR
Qav6uqiP7QvK6wyJPKCj/VcO9gVmDnBG+t1vf4YBblt9UCIwUKmJb7awtvomlQcp
w5hqmKTqqBniSpCggZtCs78ut+Iwd9M02U00++g2MwCNWxXc09sYGYlJ/wwA4LsV
ssLcKAQl9FFMAUPTkMTRicHJsIQvozNqi2vweojRCOuE58eddQN9kmQSP4yn9oLB
yIZNdjcarhJnMunrAFSVLX1aGAesP3KMJhMubIoRWbfLDwJcbnMlIrwHOXLYTBKd
V47nQzjLbdSxaRlXeMdCiJiOMKwUtWblPsJZtuQv2o92h+vSWEkvVLOn9d5mWTF5
Mrj59lShLta+DUJ5eb6NPtd1kyPf0fOgsxWyR/rcKdFC3hXNjRpcqKVBQ0jD0m7Z
e0g3hGZS3cKcm4tJbmoJ4vxcA56uZ/YwlvroP2YN27OIF5NodgsXAH4SO2Zr5FsT
MJpjmbIakB3BRU6AwNG4PKdhExAd5nAAQWmDbd/JibOOVZxW2VtrD0bHr96DDB+E
OY6XQuWVwgrw0DaMgNva1Ro/7klbPGOB6ytpSkahzjieod6cDtGhIsdiCJI0RrRy
iZYsIvCirvDpl3CaVIXUP3dZLtfPsi3pFWm2DLSZ4P2ywIZAs/fDyxo+nxVkHs+F
ip5U9ZS2M5dAQ0jFsYEmKgsA4xbYvhqdRVPkJTmwD2rljgorgByZ0dxD5xnULdYw
VvIZiv9AG6VD5CJUQUSba5L1iJL3KdhdzmH+CjOUsgE6pXKZgmzWtGMtlqFkte4l
o0XJdHd1QmAJ+5KmHiFNzSGsO4wHAo43m4n4xH5LSQvbIAorniplCGSigxezVANW
0D26bSh5WGcI93OJZGnd020OFnLU++fBRBbzByxVPzPWveYqzrbZaQnhs9NAXRby
z1CYjCfxQbPudhFOeIy6ngXYxL6vdMGcrNegcLvMAggME8vl8rRS/GczB4l0XMgy
EdnJ2o1kVOlRS2XRbflrH4SsTpCDkx0LKo95wV5JJ1t0I7JqPB94CvbcZsnzvxYD
lWdMQBe2Y++hWGzuYdDLYa+8JRmDU7sou1Bxzlu4r4QZJxu693zarrEsW7MMOfik
S+imqv7i87U/OaMHVqXBdNv339dupKLx+F5Pshx8GKKuF0GKAjm3+C0JLekcYs3j
8x8EGPOUBp+jT1e/b1Tqfb+aHnTc/NOPSivC7VoEPQqe0gj7OCda6ioznGArdIz0
dg7So28LlMGmtyFqrHSvjFPmh4JCaKj+XaRMKZND1uNloSnwALwgjVMqOdVn318t
2z0w7XVahaMEoU8ee1DkdnR9MT9LTmKoNPJNJ1XhZt3HoEx0MyLdN13V/W/UKkzn
JDXH2Y9ieFQ/MUR9Zc8mRjnuMo86nuCn6SUYdTXfYonRF9OHP/OR/m3fmoTZ9iUc
eRNLFGj7CSLaZ21+ZY43XdggtJYDFSSHD4LP+IZDokOCaz8vwbkx4XAKjbIQdW7l
IhL9voz3kbobk0IdEzZDjYY8NG3+NVUCC1HQh6AONjBxqheBO0/mjktzaA1rlXOc
S+FtM1YfiPNayiBZ8q2P4qVQSC86TeLnqg/LtpdJ9Ez7M7FoU4uPyVlwvA35nIEq
07zQyQdR/dRUsrQYkeu6/u+BX0t0e3yfofkYFSpYimmYimjRRa/QmccxHcARRbTF
PZQQ5iBiF2hJK2ZGnSLZIC3oFdtXZ3R2P2q8Rf0908RnAao7SCM0vMO3yCPYBtCg
Gl+sicxuMYn48+KxscgG3KBPk+4nr95ptf/TAbgkEpEO7nm/vSnMAsXYK2UAGDA0
NOzKEfs+NeDPxMAovb8xyRnV3CZZ4083L3+DbbyDVZA8hmUPdsnOK69+cmZKec92
2qYcb7lu2pdADqdocXziZNq054ERPbWWAOLzpGF5LGND6QJn5DqxnfyoavZUu8LD
Ez2uiKPnZE0OvOIcs2whuiVOvAHyXopf9jMOhx9BrCXmRqAt3mJmzSgPmvkPHAPM
0Qc13h1yula0PV3NfbKACPGBHM5uKADck8SUBNkDdNvfvRpv+JXcYzhDsE2duZrM
g1q+6Il/iI+nkf9QKtULZ2BuG5v/GKtXXjSZeYxD1WR2v6WtGPH0xtcSUWNP23ii
Xgpg7Z35eBQS5Jcg3wCW8XaDdGXNlQbVaBSE/cAKtG3Y7Na2Iy7zSDPABXkEHH5z
Z5K34N18XR3UU3eBftRkdVN7BkD7vHKXrr9U2doxtn0m/fhvDtSV9Q7NClfZwsYw
rVLMKX5NWKbSDesiXgqngYR2/8w3RgJuxlLyAYZZn6/KAYzsJxHyRowrNULnd+GP
x2LQXFhg9HBXI7zk+sQbVm6QWPgY4gi7+smBPz4iF/ttr7IVw3Buo4zIWc2RLmu5
FW6nASlzXP92u/iOOKQOrXUVZ62PoOgVg3AslKcChUf19q8OHxc2CVwbNHJVW9B/
E8+/B0lNbPym6NkIV7HWUPw+2UAC4y9GDWd8yhNSPBnm+5vH/Mnh1B7xOHa0Ka5O
RBeJWbPm7VU6/3sxG+5pGBQTytk4qWOqwIHGe2jZLgdKnKn7zsoTQkmMcgGk03kH
Ot6KZ8ZjXCk1lG8mm5DBg4eim1798rdE5UIVgaTdd6JmykKDz5RYP/VoK4oYXteT
w7uS6yA0DI05nv6OjV0HudSGXyisYXhCrnnTWpynJZ+Gd3ezWLgX+U0Au7r2SF4L
wW98eW+SQ30xnxReozTi8zcpRFSZvEGq8l/kq1DC6mD7iDUJuZdRyu2n7DUxT8DX
XERKVZM/O9qlz4uuDu5V5KuGnG68JmDtoodFS6Vt5ihF8APtqRbCRpPeMdwWemio
3FZ7CWHWVb08LrrAyHDxownpxQ25XjiMFNuuUR+eC+qMPfm7iRmsjI27nOTD3/yK
FEITqvDkV20CjqRAb266o2yfl9ZLfrLGuDLK4MHOoVhCAkxQa31EGKdOUrt8/sgx
tTZ4Y8PMunfwZjwSINokqN45KBsoNRWm/MXS91WtfJgHaZ7S2Tp1p+sHNjys+8F3
xQvNQt5XyWmE1xpFlSlP2MfzD2wVIFryCD7KFFCehhLjfAHB4Tvb4tZP/gdDoUDE
vniVU1bWIL0m6t0LVtWTDOqMdscuqp68OwPBt/4JT7h4hUFr/b6z93EXgODAHc9H
VHhINxB0PUWTD3cBFpXUWwS9yues2jQAGp7Db5dJUHi6ocvF+/+o0ahWTNQS0JMI
djnqc/aavmgqcj8ed3Xbag7iqbPKRxXr/olauzSX/070TvxnVH+fd7Fkzwkd2CSH
3E7FYfQENJSwdUJ6vH0pzwiuxPKBEyvDtB2o1TcYn5Ze1B1jkACSw1PVD6WP3ZWy
xf1oDvqNQ4/Rek7oqe89yzqa3GPs7XPxnQ++ma8jzZkmtUIUhRmxDkLX/ZxWxKsz
I/rq91Ug02O0fzydF73PMwnmhtoo0FJrWXwunfZHAHQrL6bo14n5lRU6xysY3iL8
VTNvq5R0OeLCKLVZh5J/yM1TfC96FPagVxs9PWvRjwUH12JFTPfa88mLgYWqCPqd
w3CbqnAquyyCvQwvIDQ7FemhnO3oF3mdovKzR/EVWiQMLCYjgCvD1gQRAhrH2320
tESr8uHaqMnD1k6a4M9QJlKxehRG+Nn2plEbpcsOl/fk1Y3CfIkZBu3Il123uYRt
05VfYNQ1K6IOV17h41ZsujgxU6my99q5Klocorxx1gOXsfbHC/GZLac2jxJpm/cl
bT4SoaJ9HxH5vfKYrBri/0Mc2S2ZRoTqDczNoU1JkPvO2JrNVN58SxRS84uhLLtR
78cSDgBKA9JhuiM8Rd/o+W4tPRXezn+41wMDgsc1SrcMEegZkhv3MWRERDV69QSv
ymZCp7BRviOL/jaiM+DK/58FsqSZ3H1IDITBtp8sPFoT4Mh32AfwRQdPHS3saV9c
wC5pxAt8Zxqat87UCBLtWmvhQUi6sPFbaiNTp9Szff15rQm2pOOIEGVJ9URZzWJZ
0Eo62YHsZ/pjBUGlEVcHRUEv7QO2vaeG0s74ePxvPQDE/fSf14Dji2Xp+BxIcVyN
UyYUgklCDtIsN3JjxRJXKdTt/3vDH+ZpozeyJZG++ZBkeJXJq4c1ZO0RrIwUlNF1
WK13an6QGzJT9wTeFVgZeWcj5zoWF5mD0Fci95sC+9IJqch83ivsAmoLlnqgbEt+
MK1J5S+KIAQz/Dzvi06I0R8A2kCfwxDhyFWZxgHOxERmJ44R8K5wPgBq9Vr+VwJI
2OPupfU2jfBTf4/RDp4MXbub+cGtVOpx/UeLOVhOAsyUJXQ+DD49eal4Fr4aAgIN
xmy0xrJJai7L72LV0M0QcZL1HG6dnB0vu0BLbdQaon5ngd+UbekQGcYW0xkQoWSJ
xymXi67oeYlYY2KiAEzm2KtmrvKn3aLLU4gllPPdgujFqLrQTWlHcjYsH9apDW4d
rjsIP7zt290q/ZOYafE+Fel5h2GmC5+fOHejQrz4XKiQJDpC1SsE+rL6RtI4TpE6
tjq4ayxcq8B2UPp5+nl5eCtkWLhwRrx8bG4z5Q5b+hG8CITRrzeYHG+Zljc5ZnUv
ZO5hzTYsrvHacNTZXKot2dnJnUXDAKjdHe2u2a+XBLSuol8CfqaY7c53++amGO8c
wheC1cTRgqu1+BavXjEDahreb9tsNEwLXLrhEgHYavE1aDTmkgIS0AeBD9+/nJbx
hMN4P8VntYdD1rpeAT6uVDlFlpzXg2FssRDH2SP1vBGw1O3guYRphRrzooiXmF2o
KN+KFzfpQBe3dYAl+O3UX3RtkcjgWpbq0fCl7rgv+jJflpa75TiVLVzSEpOlTibW
0mj9Sa/lSb2nNy123qfcdzWy6r7DFSGZPCDJfkv+BHSMABgfcn0wCQCmtXYgxZkB
27u8HG9kIDHgP8woVRGdm9Mwk3blGpOLVmfLytK4+0f70wBiYBqMEhRcA6GDvOe6
UD+UMcq6tZrK97vuD6VAr2jcW5i5o3GbYPWbKAaZlE3FqoLOcNls7y4TLhwuKg2+
TXBIw3lb0ftB9PqlATv7rqbN7ykpNfaf1ZQXKM3fKGYhYeUHPOwNkMGzdWShzP/w
MyhIgGK9R5jhT/Zrnn+lGAy3EVJ7SHWMlqUDfF4II/f8MPxvG9pNad+WUBbyZMJe
7u65DKTGgRwZOlfB3hcIr9L/LpYe6n00aFY8/kQRfzyJLR7J1EieC31Jg/iWAo5x
oYCwufIyWAajKL+JqCJB9fiqqqzyGO4BJzXhVOsZJsLUnr10st/TzGlutsPFr5w/
J4hlWRi2Wp6NbiztKT+smvjUC8p4PRqEQc+Um8ox2qRVtYWBmXNkUcdc1WsuMiuk
vlUfsp0RJFKriYUaDc07YnlG7bAz8ONVSfq27iBzQmAgG0cS8MRmicP4WsowgMNv
k6llCpV0wLiWgWh7n/eEJwklqdxAThmvl8AfWxTL240ZYfmdY+ySR6onE+Pr1myS
C0QAigwM2q7azgFnszZboMWRumRO+kSHt2jGW3taBrpL42+QmBWNmmkPXEFxXNAv
Pn3nIcsoHy3G7hiBZuedOWf/Lo4S/Ej7cXiCrDHNT471AcUZig0UR1o1War74yT0
h/GkHYZ7CmUOR/C1f13lNvdYygwQPDmnUQK1fmQiehP+RifuMNd/n+Xi1/oRfLAf
1T0y6QaxWXOKqfyLukdbO1i6T+YyxSN93GWt747cRIlgbo05clk92ct0HO64RXcM
gJn8pvVBBD2bzESox34URGNVAby9zLmPI/JlUDcvvGmmslOQgx2lspLwyymWnOXW
Z6d6Bu8ybcmgEBMEJTAlFDIfoh28AI331CdCq0pOUfDFV2iRwnvhDMsKIx0TwtPz
Z8k2KMTNrsYsXM9HEQ7XJ6gi/dZw4mc0fU7aPea3CGGb0JViOgsUkJeK+RvCxVff
JZpCHI82gkaqSmVqoXcmE+hb9ASfYOzcQI5ESJICtyQ2JI345Z8jim3rqgGrhkrz
XUnnIylUer8AUcvkMJd2RPSp7Z6HdBPEG6fxgaH8hdkIqToDhscaD04ONyCAy4/U
qrBpd2aBzN9tyLYNz+Cj5E6I0P8YlqjfH0ASDKInNSSo/wiq2CUnXWR1+L6ajqhQ
fLtc8gSaW+d8To5p7vIKR/r41lA/jtoTObARWM4tTJfbTFiNQq5r1CTfvm8hWY/L
i8lYZwyiTvt9A/No8RMhyV/QzGFzazo/uHteQhwSUClOOqDqCvCrJIsnMAnH56Id
igguCRVdg7WJvtGBDtRsnC0h7DTv6dHiXRjaOZ/C8R7a9r3eOXCE0CpRx+ZAosFx
Dn3qPOdkzKx+ZTeC5/JgDUz7zCc4JSlgXp3PkIwAtHV8O3Wnts71NQNGwimxF23D
ViJMvdCFf2c6Bs+n2R6SqZrgpwTn4tJywPIVi0h53T+1VJR//bsD9QJRlkohRoSA
9p8vRTfqNN9AX0Z/aYKlsFdIuhwlbFPwj+wTsOSNg4Qse1YIiBvxSXbGZ4NQpGjC
cikcG5zfQaiQWloZQ26278w5hg8vCMpiihymzGVq6K3f+5Ra8veJ60vlsLLZBPM0
cQsZUVLdI1R1zsDxvPr06vitFOUwdpbOLCsiGlfeLLDlnpkFNo9thdkR95MwM1Vz
pZYCcQUsiDqZVeeXfIDLyCTwboh+USEXy8Yb95vEmiAmeAi5wrM+EvcnrWAT123o
iNuScJISI3FuO0gmLjf+tjSdQFxEmbf5ekY8I1Ey4qdN3o6oFlXcV4E9fAsm6fQu
TdS6NJB6T5zybvAlGrqNVFV3L2UWr45ZfX2uHq7hhPQfogwxo7lTOgLQtN9wPvY5
5reosldTocP1tj2qoiIubDScqZVc7Ou/aMDBhA5uVbylEQHauTFpNy/B8Z61Y2Rs
3i8dCyn/xNDWR6O2VE0a0qBtzWTuAqzY2ASzkD6i5sjoN1heV+SrWRej8t0xw1q5
3ItuDnHVMWyAPPjuatc4tIIAitBXvbnqLNUrjSuHUgIxKQnIvCTWYOmu1HrpJRK/
KAhxS1sfrkxEkU5vXaYwhjepwtoItAtaiglD3Fw4oeuzweZ7MjoUBxqjVwqnnST/
wrPbFtljeHxqAxICuvMHQWYhZQPhzig7LBLrSYYXUQRnnXyAHohF8DbXmHu3xZXN
J4+jtzcOMxei+gUOIUmSCHf+R2UFo6OvW28CPIya/DIzGZXPFMBrpXd6Uuk6UQ8M
6x684eQsoq5FSRKI1wuqT89AOLKeAF/1MgHyw8uUG+tnFesSp/MyiSjVH7z4zpLy
NQZBHfEUe109uX6NI985+Hx49/JZVFoUJvY1DyfX+aohVcaZHYkKkRnKZ2S1d37Y
4B7w6pg0fPr1sH3dUvd+z6sdXeULIJBfu2MBP+Uo6b497u/5x8Ce+lOzvOnk301f
dpBihqU76Y/958Y/L8WXwBlDsJ/cWhgP0EhEWctcsEusQOEJ3gAEVZT1BPEAKIYm
jEqxz66wBJzQoNHCo8A+oAN6YfSRL0VkJIYkhGvMa8II1mQX7qyyEB9KkP081Z6x
74nK2p4PXW7HSyA/XU6zqJyue6YBD7yk3hvZfAT6P7kwjT7VeMzlwzQAbrMWcbpb
0Kf8M7g44IHNEK4NTZBTalujahFqkroZ7+h6/Pg3/mdFyCaUe54fJ/8zWqJ6S0TB
r9q+v46PeKEvVvU+4YE35kOKgGawG2X+14tUFGs0WMxrHsRIvXBdpomPI2SIs71k
FGGpDF+aR7yBc66YrWRIt0dAuV6nX6Bxwe9EcP8M1Zoxq98k4nbqz3hPRk+1tWMH
1pcQ3zDPnXszCe+BEgsdHpxb/xK6q2Y8qS6iB98FIIlo2qnEgKshTCeBYR6aBP5w
72C6p8Yxll08/R8s6+pR2T2VfYbbKo9Mc6aGBTByrPbIPJg8j0ErfjABaGe8KfA/
FoEoU//Xdy+zLYbU3g7xrGYhY5k9uR28yGnLtLu1uaPceVs+BFS+7BdlhDDmaH1i
VJfGfhJ6CnFTvNQ5icLG+5099DSl9/NWQlcN0wehoOmUFvQZ5wDaOQUeg4ejKJ84
vqAj/Jf+/4eK1qFkqnlj8AHq0xbpVnyoWZBGHpRZwiS3cHyFFsUXDj3okr/CSFja
aoaCIIpdWP/mZYrd9Z1KqL5CMzpF4GaNe/ApJwXxLlp3E9opgDZ6Nda64SS4gSmm
C3txQkg6haxSPzULmLLLizNosZ2kMu74JcDRPAEjLOmcbcXx/uW/WRzDxuR2tIr2
gB/et12d3WVt62bJOmAomUMdusXT8ScZtf6cwmKgGvS1J3FUXwVbbc82J0JaaoNN
8oTaAXfCtDmME0BYB+J3Z18N5URgfbS7Uv+iIBqH40i6GQdFzYgEcnqgpNdeGZn7
V8DELDncXQ14fSf452YOm3TQwdVC3UoHVSvIt3wyRDTGEpaidZW9DboHz473DfQQ
rfKDeKDadZifJbpn6ktMFzPD3chiPsoglpXRkMSmixNviwNMULERAXKygVI+TBK3
mgXpNvQ2sND5iRxgMBZ4qrKwPSVdhGWUaq3m5+acpFUvEga+X6Zf3JTSlvKDysHw
0xF1DGb+5Wa0wKlWEiz/TKTsIQ4D4kuJku+QhfA6zNgd2yfdqbt/VlBJtS5wLoRd
4GXjtvDnLuCUvxv2U/PfZk2GVU81vsR9GKNGRaMRUfUS4rf+CjgmYknlXYBpQ4oz
oDnENUVGHc7JaShqjwTLAnfhPj7Bs2tdFpswXxVml+eTo6f7nGVeng1+dQh5bw4+
/Eo+0Jf7XgOFRcn5YoKIaMrcmtGj7nU8A7QSs5jOWLOAsq0NI8OCFlcLqnewA2TS
zwiC9iIrBKIe4ALXJ/PZtSxxoHa0fAfr0BIpyv2VV2pPxKWGHp07thDRbUqIHCOr
6eojsBbivdwahZ+HJMJQtMwVzuTBJVEy9yuYLNXn2mHaIfn0Gto8VFQ0ZmVXLmxS
VlDpVerfxFxz10ygN3jdk9T5QhmgFnZxLj3jelulR4XOas1iLc1EESL8O+OvPIIM
dbhgsDC5lF1dH0fmR6+zikCYk/moVgAwECLL+OpS4S6Ifzd0UBilamzVddBwRBBI
Yzee/yo+SrqM0ECFK5Xr1AlgA4D8I4Et0YHG5Obd/ecPyX6zw4DsAKWcmgCxJEl5
RO4gRe50Y9msL7eGnHtZHXdnFqHpqzOQ8k0KAqTV40Eo+kg9W74MD2h4mz6IaIOn
gmx87zBuGg1AAM/+mhN0wHf8LfYHSzHojKo0B6ZymFZ9dzEw/ZkotulcSrTvVzhB
CjD1IKoCbBIKaiWdVwECfGg9zLE1ULdl0B4g5mmPsSFOAjhvELOJW0dvWemRgNI4
kiAR3A6uhkRpuVSKX+v32pzdmPnwfswDniJZAwe0/H2vclzGPLcN2OsHLcRjcQ/K
JcYAzxchi2COWiZoULjvW1tg/WTj84VfHqieqbm8k26/d9jYFCp1dLlUR8qdsYPY
UH/VyGPE0J22GnYVuODdEZ06pZtF+8OM/+95P2WX1oABxY3Sugch1WCuXW02hbgP
k7/qfCo0xGs5Lz3qYkklCtBcxsexVHPJt0IzerBJjMp7sDBCR7OnpHo932a4G2rw
93hXkNOIXXdpHhHkwiWH5suo8QgaunvqjANstaGTenzqjHTIUGlGoi3+4rkdA5uo
3htcxZrkb9wZceFn35t6RaB9OIrW588dw8G78SYMH07x3433SgKXBQN1pCBo/yBE
DuUACXhut/pWaTYIZTehrL/zdtRELo+6mZaZgJuuIrNhuovLUJh+g2yVO/hS54Bi
XtVaB6v9t2Gk9oIhg5rGJdoT/HCim5TZYg5Ik1hfV1FKMahq9YyN3I/0oYlV2LYs
6sWw5BKA9EjLRRvuTpy7XOS3H3BsMOjZDaNrXYI6Ddf6iTRTD71svsuReQIAxesd
B2rFT3gSKj028cJqSRXDKnTxIHdldOhbUxeBnz162000zEuvNMf3dNx9GRuL4xts
7B8P0y/Zly/Z76jLeCyZjDG+Zs2xGIzscXlcxLRycEuYcoW775b12qExp4Z+g6OA
AlxvWlds6ogutmyeGr/3K8sxoQ8DWeJj9rVoixq68jg8GD9xTc5UNq/Nr2ari6Ok
wni3siTTCPQQG0lwiiUEB1Jm9h+HeQCh1bnW+BldIvK4yxm59ut2xSYgYGxOaSXb
mJ2nsHTbIBxyzGSf7OHxeMDIkAEdwisbOr5jUukegdFEwk7IPfVEPAgbk0MLr3Bv
srDAm59UnxHL+KFbFOeHnY6xCGvKGMErG4mQOdWM6aVB4dZEB9QT6abdAIoift/7
QlvUqT4MPHp5uEIOI5noNx28YkHs9CtbxR5RqEHRvk79x9v8+d9A7LCLdohKeo0Q
uCYrVXkV1QYYt96ppK0Z1azfrdnlIG2/yf55JqAwJMJ2IG8jaapCsslFHENL8n/3
LqmJDkuZtBKnHhohSzaRPsdUfwshyjdDMHhX4rhFudNNapNMa+DU+fTZiLU4sc72
39tdnx/B6JaIv6KOJIEk03PEpTVUOvNo6oFzddrnoi03VaR/aZWKUo6nQNnq+u+4
S/R2l/gOF2tohLQe+5qOcyt6ZZAewzsY6eTuhQ2D9rXC9OIIeFkkgbWeoI+1LnXb
WnT+eWV3rVZh3MTt0u5Dbad32Uz4+hUi6g/bTAzRIC6Vp/7STqe+gEk+QQ8LzrSY
d4xZVTyVhpbJTw5f4IA5d1PysdELN/RF9rVObxpB1RtRXhkRuqpi8iZbiEyL5DLj
dxBSu9Ibc8hMuakZ4PBDwoi0Xry+nOhkMRswnuh00zimEZ2xz8AZ5hnl1RqrvD8n
8rlV9CYhGxE3Tn2AAjfDKfSQlJcYgxpl5ynTlX/ZxkYsdbhEQDTZKzu1lkM9Va4O
cKuAqTbt2KEKMQgZOK1eeDrwbQGXYxUXz0Y/T3fh5b1i2Ozb827lNDI+WZoovaE6
yaZ/Gq/8XAkYreAVmub193NZ3nkIraCxLvP8+xb5axx5yIzBJ3ULUH07MmKPhMCJ
XiHsKGgELG3pdHpf6w0XNK5W/8nifjGWPH2oyXvLp6tIMwBYVheemmMu93Ikn3R8
dT+2eThR6kSK1StLtJ8w3kf9Iav+j6Fe0bcsqAOcioQr3jzDFEBhLcLW0jWMW8g+
oQ5Kkyg1lbotgK2Z2eMf+DzAhMBn32RYrdKQxazHSNLkOR8BMrL7aWBI/tNacQMU
bx4jQIAH0SWXZ+lE2dt8zGiGv1193oyjuNRqx+Vcc9zykvmWVUQoCY4HINaKz6hh
TB+l8rKx3gd2U5qpTF7EwaSCZjaNnqdk6O5b3KPrKJiNFlQuEwx3g3VL9OUEvkUh
5jeKH+ydQcmnyscEV/Hj5JJlzrKTIzGmTOPuNvaPCfNkOpnLZ+aseaGOEEgHJrb9
J0KNYqRb2qXSlXzjywBNeOJZOq3F46EhkvLDCjKvaiCExmeLxP2JeRu5cAMcPG3h
+fEs3KE2sbLwvi3Y8NCtaD8RZ2d4tmgE61YWnF8/JqthiASwMDWKeM6rfWoM4oZf
GV5mzIT/M+8JUvbL7CzE/Y1sImbxBDgNXbuFVLlfJpY08WQq+JiZiFV6wC4HrYV2
5AL/awNazKJoNWzactP7LJvVrWV+nPJkxQIQrCfop8aTacfkF7oZKUCrrCFxXCHQ
sZ0vymOIN8Xyp4jhaW6Rj50kejIjp0rjU88kVYJmWHoumr7c0HTb/uQnnvwJLVox
MTrAtYj9R9ePSiyMRH2US0n1bXw+ZKKJpLi5rb0vtYKzAySdqeGoytbWL3ZKruEq
IYYiNeCBsNjXNkpAeq9nYGyYqjRkGViAM9qfLYwhPyf2jKiUbNRyQVSzX8zj+idP
2B/y2CL+7MGEOac4KO3C5rgH9WadefnRiPkqijRf6dDdkThTwnARrxDimN0tuH9i
dZb2xco0Q/AYr2LcjvyDKfSmghYpOALu6dMOmxUBOxiJbBRiPC8cbsbWH2xr2fVO
/J+b1TMnsGBYp30IhCSFqAPKFfKOfLv8lkvro/7DS2Yd2OjvLdc120UnXIaz3nHt
JU2jaRd8noqs21DzqmcLj9Vvm+7H6gUV8QMRY9D3Fw8FAzYLvAU7M6tv1j+wfUv1
jWQGjgNp4Wuv322RDYWSCwYnKK93wMF/ownJbuNzoVL6fdNp3DjjAEdxyFFlqKS3
Or2lcaXjRksRbVMUVcxnG2KB088w51lL+5pL9eW1JGcr7R0UHgqu8t539PbPvj4s
J50zw/1362C61Z2XafqD/tsT8LRdvQ1klCAweSs5V5hj0G1WkEvYnz5qdVenkt7+
XQ5K+9XE3XocpWLaS2A93hOCqQE7JKJaDXRYxlh7M8wL/rLUVLhEW8vdJVapknsl
XIcKk7Wg/HC8nHDuXTqNeFJcqMADJHtMO/vbQRU8rI5xeudJaCSL5Boor3tvBV4B
f8vY7n/1YjhlUq4zx+3Eldw/IXaNsHztNNpf2z7D4sebD6MvnOKWBRAIVdAnDQN4
zwMagOPLLu/iO5Y1LOgJzcFHl1/zHZi4yJ3HBwCM1ZoeVofwZEkJv1xQPCFT+2NO
yfI6WSAHEnhsXvPqOylZpLEELA6nm5fGyv29q6C3MVVq7zdetwzGvfwemGoKnzL3
RPq8BBDUvCpuI1fsLwCQH4iX3qLVPRoUUTHykJKLw0E7jJ6tBnApNYELoL9lmDKF
+wBf4FYNx9im4ZIUrf9N4IX2YxnfJyfPR7aIXtcPO2aTQi8qHS7whOomNmRKrPwM
6/UR80AkMhkOCsi7EOJYDF8f8yQ4UvzDgyjCUyh7StzAgIuUs0eTbXPx3aVVwYw7
oGXPsI+dA8kS40IrQ2eBdhY0ZUq/pIYaBdwWxqLvZZUFsbSgAF/eknm6+BVNbn4J
JK8Y0Z/cwKOVoR4yfem5LjOUUunBJBotQ6sZMkJ27wX2AK7MeINY9coYds0i63lj
BR4gP9rg/2IXCHZJUGu9he8DWByFb2Mu6swPZ8KdQAKgskYusxOLla+Ter0Lf2j2
rX0hvSGa5ewgPlwEYPcTGUg+NYTYAukpiKaqeibzIph5mhg2CRTJoGo4LDz0s6Sw
jFtoPnJgi7i2/DmrseVRx/6hWcFYZ0jExKWmxrP0XyD+e58hJnzkv9QWruVWR0gL
AjK6oJz0e3xLqNJCL/fGBqW+b50sW+KtS0qXfYdNRfyqTIpqKlhisYNgAZ4/Zq3K
VjPGlrAODfM1A+bTTSqCoC5cQDSiLof6mgS80w9+Vp7GxQOA9o3VdoAjHTXxSiMa
ijS+IDl4TpMHElspH1HQEG9RwYTBz0TNr2CkicxLGT4sKkAek5yAEVqiYz+yE4V7
Xk+JlMsNaVct0wIz8eNYV5cOmcAciOz2vWTnRWVJ/tJTVaFJyJ0tDd+t+br25JLZ
AQp5zAVPjbP0kXnlqNoRjF6UWxIeZh5kKMR19GwRuDVgjhrnl4G7AKkX5vPrn0iU
SmtJYtuAQFT4r6LhHMl634+Dlf7SmnFwqkz/OQMWMWpr+EBGjYrC78OCAZpKhe28
/477G8qtEZ/0yRETCd3f4CQuy66lBJxp1f/GGjPlJGNmc0/28PShZ5tNtH9y11ds
+GPm15fGwvsUFZ2cR5Le7lbwXkEc6Zo13skzSCEdzxZklvYYEHBjlS0CXoE4VQhl
4GmSZBPs5WbBfSkDyHV7nYXghDtWFkdnVg7xpbUSiiWJ5TRZUE73xY6g5cxz3Dim
LWxMu0cA1wSbm4z7Tw1/UvKtdqKYXgOASavByMstFiMfl7aRRoEs/D5Uxy/ecoE4
+D/GZfohrGAzGIEIHu8N/dRW/517XUhI4OalR/SWsxy4XyIN1eR9b274xrp6nB7E
XDOdxj1Fw8DWI8LuDR3JtNcMw29PQHsN0ucPilidcxyRhzjtoaqEKFmvaN4/NfYc
27pKlhEO25j64xEL15pSYl6zZnXhHCiIWYUNROoPoRsN2fYvNqdIyQcBKSXblDDh
IHEOalzsC98QsAbVH6wv/ya8xfWAFqBDT8S0GPxXXYKMz0iYFU/QGTc//TF/8T9w
87Vp4uEUZWPIuvlm6vzAQTBFbqH/3MQkzqfjj5JHYL7oDePupnLXegnKSYn/AyLA
TIdlcyq4VgYZUzWXmqQnsav0zO3vmtTk39j9I5PIVKFBH1tWprjmQcrKLPaLOKG7
/rM5FEHT+RhgR6UI+7z2ODZbYSQ5XFBgN24hgAcwFQ8SM7xGAfVfEWPtz6tjxoTa
ce043dp+0RdtitNU5itZi8GnuncMwUJXfMwxIb/tpLFgf/7wAOgXiF3ALCKW4+Ny
y7n+Zb3ZjpgOLjrj0L32GkKG3CFhE0YLaR0kQ6QJZu5vJU3MxBdoonJIDr17+z+q
yTckJBfG1YIL0qqGAzi2AdFqWyikj/Bkgtn5GKxwJknoRbmNuB/1k4WaabZUUwF5
oE15pS6Rfc2uQB9nCV6uaHUHkIGDXuE8EfOp3mNN23te0TObtpzoqIg0eMSRRBMo
Rre+EjPEN4QQ64PuBjwvetULExkMPy8cdryGKywsyPZDt4SyeX2gLwdaM2DdAaBc
7ZZFb5179tdCje1HGW74FzdlR4aGBG/E2Jn2oMrDIt7AA/IMMiUcTXNExyuq2TQX
nv1tmehIuPtVjdfCmxlvbnxDWiG4ZuPBjnxHTGJo2CeIirulEHDheJOaO3ZbKceD
5JCd5zTwiB+6jjC98sm0ZVWaAR66NPBF552fhvNaJXDS5lubMslMiiesjeW6X8PP
wZQD6q0oA8ulEIcPahsF9cev5/99RMeiRtPyUdwUanbw12xs2qZi8YHaramoT0Jm
+ipdHXagHfUYPQu9zKntlyZ1KZCvslP1psXPp7hj9SpUiy7Wd82grc973DFxemHl
9U9SRa8ejkOrswmYQNh/5MBPy1t9uWM3QODLI31yun41EJIJmZ8xGavxaGKDMNyR
4Vsfc5tSSuFOO3C0OU3Ucy1WiJJmuf4j4LZaRBLE+PBM9B4z80v93da/W0pBpMv5
+ipIQNOcQYwlk/BodsOLImjDIG2c0PzTLRs87FAaFQKFqcuZdBe/tpZDUwdbcisG
btNO0xMNfs+c5jFWmFkfYJ3DkkVMAF1opvLIjwdn0J36QZJAZjkQNt9eQzdGYOty
7wr7+8cLuwOp2xar1ydNGRP3VthgvFdymyI64KJguHHQEqCG4NtC4YqRv2KFwz0j
zcvUtrDlLh2Ra0eCJpDApJ/v5Qu4x/BwEzWJroCu9cMALkkbEa/gfO/qGVX5Uc7F
hGSV9GGdT7BUtkZsoXsMLiMFiiF0/As0vMRvMR+q+uh1CBZxYbkmciy6Dk7QJ6KR
kmITjxiAo3rhybCT1P0Bqo9BN0swLhmJfE2VSf31HDPAUreIb8sNhZmcpzNTH1Hs
XLzMeMyVM0cIUs/IjSBUZFLW1gEIArHs4XFSbaQviAb6yG1x/bF7HwvOD39WIUso
U3bcDvKIL7kfnleZhgVTZkAcrLV7YQs/IzZsAwO5dENI5gAN94NJaAVczP8pcKAK
5lrOxnK3MvdxbcRcqV7lyONzvwaQMvUBHu0E454BuE6dGwPuJZgw1tE3urt/PE/c
n7KNAc0yhYyH8xPSBMq3Q7zcFBjNmKFXj2t2f16MX7TiA3JcNC1EfmEdKaop6b3N
KlDjR8632B1ySGPiO1hUvNlxmG2YRN9EpyqjewF+n2bWv6F7TA67CevCSmu20BUp
HI6DMnzlvuWn3H62gVxbuf8ovP6/jChFZDu24xINF1MsxTdRd6B9mNuRwpyIY5Jx
y8EVw/NNMFiS9PhTSeoUthknePAcNA47zNsssQhMZEBklphPmcokzXDla1SPwLBy
yn48b/xpWonftVALGkY/MVUBxZcJMw+NijOhthmcNWhlNY8sryR1X03q3Rxd3Loa
q94GEw/V9sVVoA5DZYO2a9ETeLGFWnOAO/ksKttWNMesZaDJ0ZPi1IRvEMaQvoOE
RKgDhmq0IqR+KSvl5B8OjItC3HERx8DIIbWQ9aVMkv9Re0Yllr9tQT7r4VCAit3e
2EFI9SgEWZYyc9czKuV/rLTUpFlyTRpAi9abHRrZLWvUKJpnzWm0fWEBAxSG0b1y
OBT0/vopz+kjXJ3arUgfxfomQXoOPCQIYf7HJck6rukpcCSBnYF3m1BLJUtemdRs
u2EdjcnPvWKGbn5Lejoqn4aadnkw7T0OkAeyPhE6fi1cELEWQd7BnfWBGUI8g7N8
DCS3UwDPKKZb4I/zDW58sK2j72mHR4GyM6MKnbJaeUv62ADbTDFKYn6jqfwpgHO3
6we1uF2dLLRX64MgDfVdkwxd4cI4gUHZ12wVqU9pbysuEzN64O5OPW0qhXLAIEA5
3FW3Vn5GDCUCcMEfT4sB2NiTZ/OXODis4yXeiKzDckphV5QpwsNpBNgQx4TP/CRS
gGacYECvgJvt08ZMKFBddD55oOAeiT0rv3rX91hB57ISldRHIO3CyOGreXE+AGGP
Oj/Xb7vTRcaQKSdk7goN84GcUl4qj24VvdUYRIsj9fX0EK5yIDg//GNna3jCyK7p
gB0GlpBct01tss5/MuJLhOrN2OtdE/iJhxd0dJij+4vcRt7hE1b0NExJ4zfhVZOK
uP1Hw6Zz+TkPjtDC1DXoBX+SPizabw6weJGqDxfx9a8CZ7qvING2kxXypQ1+6PLA
EFSZOWMc7+qs8Cm+VtCQZertLIHlsXifqSDLrcl9xr8fsjhaw+mZ7+Fl3PNSvaA1
PJW7wxOTpOpYfOqp9a/z9KMpWwK0coQioE0w5Gzii7DAHyjdqob6A+CRicaK4sog
s3pUx/G/bDJTsvsMmcNmnpZJ3M3JIZADKGIGnMtRqxKrYno4o/MWF1Lb2TXhWp8r
OrNKKlD/UYkLMMPVCl7RbqERoHmb1FAMZbWiu6HYJ8UhHHaplk7yBUmP13bcbR4T
VmV0kemp9Uub/p8ZILHXMTZRhlLz/V/p6hAakUsiRzU9m9x+0Ty5H9EKG9JDlzRx
KEEiSO2s13SIdjtc4HwatmpZezqW8W65i8AZB33bm7yzuSry2mBwgmva+qft5RXp
kVbCDvdpnMcxDAanE1iJzc1KIobVbT7oJZ9yaAvk8SkekYxKA1kW4NlNwVFwJ/9F
AqrsCToKTX0mircTydfDVAXe54r4mNejkaVTiVfng6iVhajXwl4P1xxfuQIETi+8
82NdFIZfSpLOv+7uLYN0bJY/79bIZlOOWRyOiqzErhAggnnBpgCfTBq01yd+YFgW
3sVK6SkfMpYhnwXRNe/lzn3DOzoPeIAxC01fpTE8L1ZXUc9iNF/eVBNkNADz6FOB
vEQnAG0HQX02tYdkLHp935yPWuICPHPyWl3x1s6FW9iP1Me2LoqPzOfCxWdqzQ/M
SA6QLKNVHpAiByZrC8YXw1io47A5CIfUG15OHHY7cSkLQnSL9MN67WeTO/nphG9c
P/iz6LpXqJAdxmn7AIqor+Yqzr/1aOB0yPkyzsqfup1x0c3dF8ta3sZTL9teO4ij
oKAn4mBgQ6qxcDldXEbAS4wba4LJXNuWiB7bQbgT6Oj2sujMZqIYLfyq3v/wIDSp
Zl9fxFBY/aALrThbgYubUgMyRfvw2YRF4N4/XYdQkjJMji9Np0tJVcJH5nUzGiD5
wn/lgBAXiTyupkSWLfBIsApLd9I994XqwnwA0VnL2RKUil4nkyZE+e7XHLNoFd9e
9sVjSgfGsW/t4BpStQ4FDExFfhDH57PvTqWIOyAFNTJtLT9Yqjjc84CkE4uEFnqA
J0Yef+DEI/TKALNS6aVZFiVP+m7aPburZJUXe8mY+fpTs3/Up7clYsZO9MNL/vOI
wCbWuQ2d+xDHSCLwMfPeIN5RMBBg0rgUlzY9dfK6yue69FL63v7e8rA63Oe2/qkF
m86Du3+WbzQvJD0ymvWmWokwxjdWTdFBy00zAo1sdKDYoJbfWdGmR868IXXhTFXx
tOz8wd969J34Vf9DeOOXK0PTZ5EW2zVPH9HOJPIH6fKDcvUVhAHabvs12UUpRcCk
sDgOjoicJETXyg1lWfMgBoBh1E/EiH4TbLtJ8I3DhyKC+1b8KkZhDLpUALSo2+MV
KlIlODyFhVs1upM7VBhVjFsHsNjbDL4ufY+ypEJyJb37HRjVbFXfKNcUKwrYBeXX
n0CNsrLkEL3tPafnpiJ3ko7Jhk0hNhoEn9JtIZomYB+fjJ3Crc85lcPPZrKribLq
8XiRIbLY8fyrq2m5AebXPe3KPghHI0Ud8i/oK5YS+IkfmuuQoTmNbguDuSXEiw0+
L2XPaV/2th0RWaHuhoCB5tFM+N0oY8OJPWXr4DlyqrH/sZj4b0dseHmOUvAYoVd1
vzs0C4KYgecNrEeBr3kRrldNdrB3DY0mYr/EUyZHOd21mlyXE1hXiJuaCMOh8P2t
vrw9Mrg8tSK2m+1MJ7lU7HKNNLmcZVkUNsrfpuSzyKyYn2xqyg6ZfqsPY3NwdtBR
WmqTo5uRdScTAKlaW7q7DOg5gDX0+unkSns2jxM09NnenpmChq0AriU4yp71T1+2
oVytk/K742Wf4X74NdoYkFRDsUmOYvH7DP9RP+PYadlKXxraGYToAu5h4eUh+V6d
S9+S3fIGgdLNWbEZ99VUwf2TMb0hgff/ZUI04u77ULWron9e2movsZyh4AggFk1+
RxvQgF4w5DhorG4xG4grxBu2m+kGIQtOHlMALcJ0zb+9oDQ+ha5EGVPV64+Hz0E5
O1t+lT8VwT/RTfyWf0ViUdbVBRFUDGVMtByBXa0hR/i/dMSPmNgz+p0XNguV0dr1
C2O+SFFCAdFmFPHFhopI5j8/ZtzwLiLeQD9/4Bqy6KBZeruLRsrZ7W8GmpDOwxw8
K/r/2vmb/1um0HppIdQjoTQxE+nuWEP59sG9i6yGXzw9iLInX68DqCJrFAhb5PPi
QAFgiYQn6sNSxleMjskoNI8S9Dnp9YtFEWE4ptcUMdKnPMJUksYlMNAsrObW1Uk+
n1IAhontHD1ALXN9HsV1r9BIwHX/lU1TZRXZMQEL5NpBLnnB82lrvLnQIYNeF1j7
iMkKbQLhF/sZqTHPoT6v/xW9GU+rGMJ8+7E/EKnN81ftIZbJPncZrrTlTAlQFYqn
jmz5UnUJlAi7uKMrHRm/x2xfxFBQKrjqn5NO7msK2668tDu8C1bNjX1lYg2Lwwy8
wuvbUa3ljVKqeWRx/ydWy7GHHyFWJcN0XwX0HkrcU5aWhFio/CUWdNxDr5RGKw2d
WU1xDi4Vn+cO07QxC4lMFtEXdEf54mZXDd2heiKZWHb5lq2I7iLEL5nzaRi2ldfe
llX+mMiuhLcBAhsSCOpoY1DRwYLAKPXX8mfyk6MhmdHPL1wFn/CIE96Pr8IEYit4
oncJt9mRZ+N6rdcT2zUt/BeArgAB7UOopiQFBXnO4gA/DZ2AThsiyoXFw6woRwic
PIFKGC2Wh53+toTHgtYTXRDT11/ZH767vDhAAdJJhwSKnHHyVRd1J3nKRj8EtYyO
Zda4jBygsWjzJNVr7xxr99tJ4uBX0QN557gfp3pMcpEJqtZ6EQHOBP6BPhWp79pi
lBX0ZWeQvuDE8nG5Kh+KxjLN8xGFVNwaPimTFuzMPezD5NPeA5/jGXGPy96GPI6T
cc0ijmX2VdvBp4pK4Quk/aqjOVMHwfG5C3Pm2VQJJXfT7CLxa6gjyKJYYVrlpNmG
Z/3ieIj3tQ9xXF+QXswe4U+JndoV5beqv30v+oLq7pa71JMHCzQ7FWi/+ReLWkmf
OFUIlBYf5/iLPw0Z0txZ306YsRNZ/esq+aGgcCeQMSlF7l5VKJ1gSuzY9EsQAxjl
t2DzyC9UVltQbtdA2E7Icf4YyJirCXWaeomPQf2mmTqq2FHPaW1CHBAIuctRNOXq
Fn2zfVUnBmKS76ucZ0CGZUBeqd0T4CwvcEAWZewZlbHDNZrK9WPG245bRhv8bKUD
PuVud3lZN4f0bkoTq4ZjrBLSD5ppgkEmIFTAM2yLZ8X9he085MpV7nWRMovRUZL4
ikZ9DWPNTGeBXCTHM7LOYW2AANOclEpRpLD3w4jx/33s2CTSH9mey0IBVBJrmsra
JYQLqErOqdsf32poVFb7eC7slfuK/5mqrJIUtFcgOG7EBUrrdwGzjzuwetMLQpIF
h2EVYOgpVZjewIG+jRs1srgJvlcROEVcYSm9dmO++c+pdKR+6cCh4PL9bFJ+fJNr
PVgQyRL2CF3/HBzCVGX6nOeaqDTZp0asF87HxvMibAFbbEw/AQQx6+2feK7uMvYY
gRsU4B1XBXItIIeq0DaBOxn3DuUdARtUaK+Fzpsgtkh/anIW9CfX+H34xyubqi/s
DOqXF0pP5xmo3+4uZHsuuaflYT/tizxRuUtaPYkcQDUVDGXdt5vDe81fhD7hsPbm
BNDCQuGn/HQGq+pUHq7GZUOmNfvzJW562iLgTMUA+t/l0arJ4sR0Uz2GoK+UD8MT
87/7WDKKMMT7S0AkgjL7QksgyuV3D38Vu3LH/2zBZ2pfuBPuqZjS4xCWdwzE0yAG
SMAVHMuJAaBJVpjfozTlk+92jt7pRYwYkMRrJi9EHLDdmiNwss6Td/QzndWu5+7W
lfQs9zZ2wehF7xN3KtlJsl12uhRkNadsT4FKRVn+0y3PsZueW3kparLqQ6GmbqID
+uEompOqm0hqrB0eBrKqWGDW9o/iwC3nk6kSjqqWRBQ381Cxj7sZdXWcHIpCzU46
P0olBlEB32C1ocKs2YqBfz2Oz8t8QmmlR6HzkcJuA12TSwtYZN4iwtjwbiNn9bLB
J9h+gydmA254yAxuf34IFA+rFccuoclhKU1EM3IFK7BckrVxzlwuOak806btr1BK
nnWHrZ3wS6vVG1SXRSo3x8NddGFt+Fv6CIvrwSL9mRyw6CPQEzyUQL+GobwZpkkR
k8aJAk6h4rOeJ4W1dDkx1svN9Teo5EJz2SVrcel32nvRE2XZH7fGfVqcrWNzFaqk
zTUfsXWLbIyLfrftsDlg9THBlfciZKlqiWOExnSQgVG2/NjwoUNjK8AyHfjCTg6O
21atDionVNbBwAVvdP0j1Po/W1/3cwZZWxYe2QpRthVUHdTS2psckss+fHXFdMgS
xqtkxvj/oDWho/xB/sr1eYvVuUqxJuHHy7S+ebdVC4xQ4+W3ROaxIzAnZrbILlgO
3WVeDpeltLpH9P6g/XPUjhu6KFQnLf/SeXb0y4ywtTITKo5aVS8GtzytVsTrtFIB
I80yC71HtZTzZLdB1iq0zVja4m/I/zk5dzKjz2CBDjE2hejv8Hfd/5ynzLEdH7a2
TRDHEJtCjfg0ANUF5Zi7yQbB1+t1fvv48HDRAvOPDbPiLmCwleHHg/VRA82bZpcr
eOTQ/q5yZCQoZmc5HKKl3789mWqaveLvbqg6txCT9uiwy+3eNOVA98t7Qu8qLJ7G
qzGjBhRi2WPDkVjl5lI9WjHLsK78S/VrQ2eEJ8H1f3Oyw5mhZUOueUsLGNnzofG9
eC1eU7R7ufXIKbn+Yn3jOyjXugPXSsJUT5ROALCFWnJSJaUyOL23P7S2t2Xy50sZ
4y4ooWoYVcPmkub2YoCpfDRWTlEfoxe2F7s0BZU151dBl/wDBqT3cjFzqZM7yQ90
+LnWr0zFuFmHtRNxC55jyKK3jlzp3IkcRrqN5hVwbWcmcQKhpDHAAW9uNwOKyPNK
rY+dkJOu9BMcMl29IlKQayq+yQPc1Ruoca8NIyZf8JebZICzK/eX3P+Ci4kH63SE
2gYh5AF8szIh3P98ytQHLlGwM/lBq7u32Y5mEM6AcswsAWOn9WLrUg6jrNGhlZa9
ezOLeZ5KSRAqKPS8tatpuAErilL+7et/MNLorPzzsJw4txXVhvZL8l6N5Umo89tt
q0bqo3MAixoC8iI1fUP8sC0pwVVQs7Ev/v+acaJDuGZ00OV6UFM6gvkPdS7yKQFw
6ySHiNl+eFwUwcroF1LJaJJQYLYXPd/qynKjIrkuBnnT4Bg5G3DBw4lsqx8loVTA
6cDsRSLHXRN2WCxtNXGVk8x9KKgBC2612yEh495UBor+J38GD3evd6cX7XZHy1XQ
d8Z+61PogmBD8sXZbXtLSo5wNLbgb6XA4p+FPkwRNLVoi8FW1aNSIcIHu4RIlKul
n3a7ymadwruIOSEb0CSEuWDknhIjVyLLmaJjrAraO+sICWNGHnIcwjVld+oB0NNo
32jDp4JL3AvUAcR+EYnNOSn3sFEiNU3cmnS03NpiSnw2kKg5zrYV5M58UYi74V31
mruxkUEYzLZ65f/oE7ytFKANYXyY6j0IrWBD7xMJvs7vs/Q3idQhi3Sht+lOO5DQ
lqSHcg7NfmB9fXULH8SUnaKQImIXbSNoXtJ3B/bQEWQo3O0rfK6fQPcBQyVmngSA
fWI3+xzh79+QSN0IA9lpUVkzl3FMJ1UVQXXIsoJQ5Kn38pn6AP4lBGe3vZ8AuZPF
wQtibVg5tpZeS2wq+RiA/yqZbM0izomG8QCDMZE/qi+Fj5XCmCX8x/8l8qSergsZ
XRgv7F4bCxUYofV/RIIg55/UbxbGG2K3PdxoY8kZhE5rAFjVI+J77b+ApCUZsTc1
inOE08Mdi5P9JZXuGHDMiCkzbVmIcgtfVSb3cJVvir4wtEMf4FxMnxsgZ4vIPU/q
nBiwBRQdVUvpODiVw2BPFg9N64R4RStdckHX91PPM2z75v+3cQThTHh20MYj2ZfB
c2kPaNYRMkBwMuPT4DUDaK3N+J/OJGcHkZd4GJQRMCgWsXGEW7sBqkrqQLV74fAR
o0Sj1IcgJwTFS34C8ko84n35JfY+xZe2ed/f9U1+GUz9zT3rbuo9Y4JsR/bL8Kyy
eeKTdm98MzNHW60774+K888CXYDFcUYPZF0qTYbKI6vqpuUEl/2FX3hy6559zco0
yfVpSZN1y3/nnUdHG6GWsj+rCAXxfTHBp1cYJYWLNJYDhtqD5xrXISQJa32g/x10
qmeqoI/7Vjx9t6F7tNr2dVPx8zYpPY1p5imiOr51/Otmi9h630AoxtprWaRrbN1g
xQ8b8S5OcDfi6uVcxSMwE0glvbgLzJzHlB5MULjn0WvQASvlrDRCXjXuJMSMfHrR
k+AfKAsrqDfnNsYr8WjYultXORRMg5YqKXZO+lyih+WfnCDxOcJu3ByPO8WQDdIu
xOA+1kBqYGZvX3/yM1iP0I9O7zG86OVh+tLSxLzXkp2nrkVXWvKwPNa4QxzlHP+n
Fm+wN4c2X1DMHbOdB371dgX7vkRqVei0GWHigl3LsxhEQyIt1rLzjyQVI38+Fj9x
o52mPfMs+kLMfngK2+l7+xCyAK0bUQjMciCUrmsdQxZNhtH35PKft+trWDqO1gIz
9ekVUKtSdoTpIyvauYccwO+ZV1j4p5QVfSu19lb/2Q9V7tzdGiCSjGSZ40E6wgxM
+VYQSGAsKOvpSketjjnl5ZChERRtO26oCkPGNynrOegZ2BjjVRxwVdozRt6WmR91
1nGdz/mZ23BZfN/oign50yT/MHJOyevrTvMWMvI1AOpUYCTrtHbMDSiHl0bCAi7/
ZgjLbxi8upcKhMntBP00+o/seXyyPN6yoMApVb1HGlYx8nlRz1dvit4fU9MzFK5Q
vB5DVmop/rYKW0cik0+FhrvutGqrg1WtTm4/af7MZD/Pkkj1dsU9l9ULjiS9nMNK
MuHEzdeu0Mqk9EGpYuPzECgh5E2FcGePcJU654FYtRXE32SkTfsOERlZ9HLCO1ks
033GMVJJDA/dv1muGW/MGqSRoJUnCZS82UEvd/5FvFTOh6aLgyYo/JQTvIFe9ci0
wi7ORR4HQMT560Kyem2IpnKgpyU7tZ6fbEFhLufAPWJSlwP6n+l+IfsQ74jMXseM
ZxsrnAsCJqi0WI0WepJs9SiRPr6azg0iWMsSCMZZ1rxNjpXg7EpgXJfOO26q/XCS
rAshJYlT1b0qTltzOQg07nxvHYPkfWT3q1yvOc5dT+hNH7w9mif9huL38NmGJHrP
0CmW0D97/bKj+dceEmt2kY/qI3DzOV3d/Oxn73+c9V7oZEXyfOsZDL9E3jdqN9mY
eFi3no704cXLkk4Dm9QCnPDbW86hFOy8y1pulLtw55eo0FBP8pcFREnev4dXDB3a
JpXRzvIzJyLwCuxRUMkK2v9zXQrFglDdd2yl7O/6Xp8FvioQfpc34jGyFjO6d4lp
qOI63yWw1mTHPmJ6oLyZGl4QfdZypTJhJCwmXS9Ir6qaH8juBQVh+T1psBKSJiwt
XJbHTYIzLk+lOhmHCliIAPmn3VaPnHMooyZvpsiyvnJz/lFXt8M8WrkP2ei/coS5
5TBe5w+CrnifyJcU2Y39jskrhaUpOZAHLJCVlOPIsCcWPCh6WhsdPrHjvtIwW6rx
XtQBN8+HBZhb1MbW21Gb55DSAe/7LeiZEYqWp4YH/I/R10UF9+k/MJU6EksYFVy/
n7K/tZmpx9kC+pP/9PdJrRsL4hu0muTluPL2iRe2vNNpqXlG+oDaWw5PgeqzPZPO
up/L6+qpBijL3n4WCe+Gx0U09Bp6TLce60SvB+t98qDQfDXUo9cy/y/ucupHAfBT
lY6R9sNC5NDRkhfi0luTh8e1MxQ7CgqNtzrJnXu3wJBLeRpLf8DH2aG6CvDrwOUA
ZTvTC8db/tDgVsJKwAvX7qInoxVuLBMsud0HZvZfEh4g5lwqRIqT1L86OK64pw87
fVa6Ab12DF+3IC3NVYLUWUEZQmdsBOZT0eWJb4MCzLPyC19F6DfWohF/aWU6eHJ7
dW+smJpaIQR7lHRtZMkTQSR4hdzK+BZqv53xZAPYao2sgBlCzTxRdildZ2J8tavS
2ZTkvwe33ZU2cp/bUalt+MXHhMaTzcQgdMFeLO0V9cHF0IRHU1MkPkyubbJxFAHI
5AZcELVKRFi0Ekc3ABhouG7GVL5akGq3Lnlt3SVxQ8WPzHpPYtfru1xdUg71dmeq
W/uUQyh2Dc5bRIqY1JvGtqp3nqkqTvYP9AXWHyp9uaM7ePgoQfGc6edlFz5c2uTE
1JVUz3uvQTfmdSwnozWj2q4WW/fm1s63jc9vtFd+HebR1LJr8ktQefwiV9ducSyp
GYEDHSWUE1YTrM5fUPqmU284OvDlH5cggcpdKU5JdseiUFxoqCX7rlGhJHN7/ySX
LzsaZnXd0feEfnKRRS9rK/qjW6jAPf2rXkrtxS1+H40EDiSGJCNuWADbviNXS643
clwer38KyzNJgdQEK73ZiUR3BXHlTddxTztfLGtH0M3bjMdNCHJoo+fNHwJ8WEQK
VUoH03Uo41b3WTQh4cchjDdmzfTdPeIGP6EpMF8tq5ir9FXUEJZlVqF7AkjzfDSq
7oUa1MU03qxsxZaGmr9LU447LXOmBfdniL25b9gCZPtCq91zq3a6ELIZgZYgzCoB
mdOsNqJ2wf8klVJmgsXOlnGKLKLGg8Ni0EETSsdIwv7lq2YWmoOH/chOclqmssaa
qUMG2xHw5xqSwtei+q0BQIqexwY3tIiwFZpviX/KlWhh7lnCYJQlR2X3acHMfXNG
rnNbfRURsj22xWGZSAyhwvsTTnjP83xYlKRuoTMgmV1L2vbhX2cNoTl9Tkzjcvtd
8Q7WeAzt+VLT7skh+oQ2EIOo+hL9gasy2QIP7f8JleHZugVP6oSjxsI0VfA6J2iZ
qabXwp4ilxnUD8wP1tWyfcXrzeBjNAS1Q+kp0HfG6TborGVCHpjBG0r0CEtb0nlk
A3gW7QcL6Ifertoe9wUNp/h1N83JoH0ezdBOeX6xna7tOLxeqGgkf5CuOXON5GTE
kpc7VTLGaD7A1AehiUOJX6sobYKmQRciyBesLklh6s4uPxP3nSrbgQYOsYnxDkXl
G/j2eVZXJzZRu16BlWR4FkaJoppFq2LtMPuX9INGbBRb/PW1tNCwenl17PplQcZ5
nuCfAdLFbhtm8Qwq49qcPhZkQyx+80MtAu3UMF4yv0S6rHQVlBHYCTsBhRE3Ebue
r6KOSUmN41PcEEJ52FrOxB22L23ZnKH/6nMcIlHpiUMh8634U9vys2nflZsh8dHJ
Ma9Wa/QZzr7sY3MYnmegZ8YhaLye64LMXtUv27sU/QRTjuctH0mFc/ISU7Oi26/D
SB0NsxSemnOyIvTnTPvrVaxNluFwbgmwCDsd31UHYLNVws9SNy9DSHDVW6UtszGT
ry9xK0j4+k4CCHG7PIZk/KJ8eIm5S5HfhaIHk2i2uqSmKhOE8jgB4cB55wmKNeMQ
Iodk+qAQMve8V7I5BbXieow6UxgIvEGKBdqRvNhpSgBfqwIWkSrlhpmmSng8SLPr
OMwfucOEmvporpy0gmDV4BiotEXQeH1ZySweXhmfOomBxd/SaALhHnUPYOOwwN3W
u29dgK96+LfdTSmnbqJFzRfYdT0iKiWMwFD8vUL040sH9XJkQje4BSZLUFaVNkHX
3apQghUoYqg7DoL3aBunmlHVAUqjkE4IQp3abc3cFwX6ykHfz1wvxcr3VpGnyJ9L
MT2ApMX9CrMxFeHO4XYMxDhD8I6h2HvCAYrmp/wdxYk+8D+geARqud1xOrln74p0
RoB/2cX9uaYGBUfux3Zk8mYLyCn/bD13PNZFBCEeYJaSyvgYULoBfwhSoCmt3TWr
e+/8q63Q7Wj5368Va+ZuKC0MPwQ/iT6UxJL7dOVjJiSZDqE2MQF/CC+MYsmTe/2p
rXk4LIoIc+46IK5G1TqlXHDis+MEPlpBbghoZUhLGrYGVgTOaO+zn0EEeWtFurmC
gQ+MPNPuk+ZT9M8YUNcU25ERE8eH/UJNr+TrEinVP/txeYMsHIu51TSs03ga6JNk
8GNlWhB2oG5q17u938Qnb6Wr0d2derYra3PwSSQNxCY0SBXXOoFrbk07Txgk4byZ
XmmSNONqgeNiKPFfnWoPwjJx1ljt+fQp5mjx831a6qxtzt6if7M6oHaSn4nNVGn4
8Pa33tnqoryv3BJ9pfBWNXBw5MahVwQ8F0h7e7cDD9G5gSD1yScNZlPtXgnWdyDu
1BvPavqhKUdde2mDXs2L66QHGbM7RNF6tvEChObbtvfMZN0vq4ScNU5WTjJySJdM
zU2WbItiKmQnd24mlBzoDnYDXV9XHwveC4XMxGmNvL0YrVHGFNryIfijlgAiOuWN
z0mbvTZ/FmxuqBHm1HDa4uDhxmACzRpwRHmRHI73HegGiPLKnnrXeCyKaKq8n3HP
emMt0UGZZtWrtnaHMO2PZdHjWBOdUJtfoMb78KOSh2/ty94XU7rYDTTDqn4NJ+tF
tgDLSaQU2ch+JZokay2YkjBKGICmo9m+aIu/kKM8cdjVT6ttAh9poRdeK3B/sS3q
bUwX0CwyzZ3lXwh7L5BIRaMbT6r/mpu35QzdtLjuguHuhvZrWs/WArJDZxX7U0vM
uwn3Zw5gfxl1FUmF76dakY6Ega67dya9uX7EkTeFvHXoGTbDKHdRCVJTMG2Wf8RX
BODGaq1IKwVe9SjBPPfgEgUq6HdJsNBH4xfRwi37700fxL9xUhe8x+knneYK4MUK
B5xmno8+T1MjTRQ1QlQLwfGbHI3OlycGf1Nl4TVaD13zeY9u29MzhSHjAvGgjVUz
ojV77irPp6mzuQPNn00vKMBfwlBcoyMOdtSn61EzOonffK67skn90eKagq6aBb1L
PR9Qb+ILVaxAX1X6RWx2gTdWPXJxkCC03V9++BSO5ZS/V2EK1YcsGFOVgpStGkK9
6Hmhw+rinl/C6oORo7q4nAPPoL5XUW5SY2gyBMcVEwbvwtNfOnl9AcJyHANrZg2/
3ZR+ps97TpO8AHbIsOIdnf372+nUFQz9QFcPLrRLHSSjAU1+ZdhVdPhwcwpa2S5O
TxC6HAI1Vx4kTrzSDLU9GOQzNwE+g/6fPileT2ryg/KkqWlgSKnYIGybScIirMAS
b2zY1mk85hwGf72P3TDlIhtei+G8O3gHu0a0sklq2mBFzCIviIlsBJuiF//OZwVg
9cXqku0A4E9EowA5eoZPlTNN7Q3+ap8avUtD42U6EVZxvwISXPg0ksMNnbIDMXt4
zGYGjR4T5hbdrkP9TKSYjvN+eNVHPAeLYXC00wdY+/l8mrR3WFjAL/tuhze4UHm+
1hY60tTKPAvDc8my1XRyKsfyt35/MOgpr3IQ32jK+CIqetwJk6WYs1QASaGEkLZl
xwMw8L+/j6e8ADCxCMpOzXj+Y0hT3joMtgR3iU1gIre23zCdaojUD3P1JCEaNzr4
jv8Z2EkTcAKehEW3kqf/mgaD6JhQXhyWpCQNfB50z3XIYBGFgoV8MEzKvl3rejrA
tbQMlx0Ld65RJd8hNNp5j2zYCb+vLddfpJRd661UKCZ8jwZNxRgDr6cCd2/w3QlL
srceIfLSVGTnHyb6vqrGHRV5TNk3RsUvOwgmlNiL+ukYFEtOXE3lcvqpd0B26gER
mlK59TvUdQUIt5wjkh7GJ/G75kk5mIdhUuH8dFJg8/OyTJphp5EU9pYPefWSU/0c
HVr5zVjx4uhRHk26Y4B4j/tARtbPajs7KICg6Lr6UuEr3usvfsYbPtvdH1OH0fE+
+rz+yx1k9KGAX3MQMcZeXE5KNipNNlKXzpYEk0pVfV2ni08ym9swBRNBNkOeUy4j
cIH0rd+GHtPLYv6LcwCQGEiQP56J8BUXcS7fP15jyBN0TFw474teG7YbRBuEE+vg
ae2ZDnRskvDoHP1cZkTFzuYYhqeNOQqUfNCVUzSK3GCABDaEfhdwIhOpc3W3gnxA
tSkhLylqVbsRsnj0AB3YcUMjAkaBZB5PGs1sod8G1ZzxS7Y719XRdXbxAQgRWEX5
Ec3/iiE+GaCDR80IqEpt1m0s49BPXSzanxxdmLphakgKl1SoZo7Fku0gQiC92znL
JUIorcxOnJkHOi8tHj/hsJ3gbFBc5uQ+Es7c7B47Le8nd94/nqEh2qx8DgrRrWEc
zjRm0IWMi09O4Xt/5TvfW2g7dbrvc0w8AOH5iG2HCmUWKDAk3jyFmwHcLtDEonKX
dX8mR8AtJ5kIEDHzrstAryIkZ8q6xJRatvWN3RYrPgCPHXf5NxC9pOFtR4Lvi3z+
pWXAUZBFdgxkf+xec7kSeThc5jkSc11LkCj4u9nKqbONE0x43SxwEFCDN45WNnKr
UBXa/4ZIpMJRBpnLLPY1U01GxlHLD5umdT5l0M1VYvK1kKJum7/vgRcp+uEws5qq
8GGnEZb8Nqs5Hn+pVzaZJIm0qVzqwHqU0X05qyKupTfYCOmf46R4LjSNK44Rwt+5
JPEL7l4PKX5UGxCOtnmxHqIihE2ORAFbWtNkTdE0b4mkeFvaNz8gYs4rP47Hp0bW
IyWW7gIa5/t/Hz+aiqVqLj3Ui4ZU7hcIq2OABa1BMT8vbz8wg0s2rkAOIFFMmBtW
q7nfM2bN6wkyyT8xnvsZlgILALQV0gBUVvCaj7HgDd7yzxtYiAd/yWmSwCdQAoBE
Fe+PvWfxjoWs0YN63F7uS4xDnxoVZa68zPFNsFR5f+IUhVfva2XgHk7SYXY1FBYE
93kqI5mfGYoxgOlp8FfPs1hnQwgqNO1rtdrlZi/jHCI9Z0WDGbDmiQRNgfr2G0jd
mlmYentcpjQPcBE5h04Lz3MF3CN4gvlWBnzuELF5dauC1cRVzzpuKx7Soz3SLChj
DsXRvhgnsJb5ob4XMOkuyMETSVA2syX3bsNSMtuJBcPtbH0KS036/dhQl63kx+Bu
vsxSArZB+8tbqY96uoSGzvcu71HCYw/etjDZq+KhqbP8L3z/nrk476eU2e3pNQ2s
nnk3CCY9noLCD3MhXM/GVkV1EB7jyBykZb72VMFsL3UiWh+LkYN00HI/m8p+er+q
E0ZED3A0BJY1jE2txai6RfGbDPCa0aHi6prbkKs8pL34h+tQWfBnnG/MvAVzEBjB
SxKJxF9xRcaVjR0PP4z/eMQdrJ9kPqN1hLU5jew1HraPfDGdktmhikQCUgO5bQoz
IVjxtrHCtUoJwERXgzA9ZH/jHeIiCh9PJWI05f+Ih2cNI/o9ijMFngAyIylwRfjk
ImU/6aiRHJAyUOZ8GvM9omyq6Hijak6jL4RbN20lMN/nsledGLwfWwbqj7ip3tI3
WwfjL3ciJTUQe55Fm0+u14jOp8nIiqEFTEbiEVN2RMaGDYVitW+NODmCa7IJtB5e
5BBkyMDDCnrBPT1l8lv1LJoq36zmeMalSUx6n4GTMuTLj31oxDDFbLOtmv/eUGQj
VHUDKUlx0leMizfamnYN0HJxnozsFL2u6yIoL3N6ym9hZ3jeCVjLrtE+SSvPL0Mo
tOh0gEYgsGG3eFdpbc5NgaOzOr0b7QlthEUY5JLKP8qx0C5A8lCHMw4nQkv2V24D
P2HLZSW9gEW9CcsQLz7eG9a2qw9x58MZZMx+cXIAJ4l3v+f/DmxlI6p4zeIj3uXA
6CAFHxBJaA6Cimc6IPh9di4mW/c7IyxGrCqCBpEl5esqj8awpk/AMCbtC/wJ7JO9
mr7u4NNlJTCXearHp2RY4c1zdxsTSW0WDS7r3O+szdwo8/qef7uEc/46pTEVG8di
otB0H0eVt5+UJKpuGA7493qrPe6sbbfy8p5dyzedqaFLPaEnA2SBd8cMpEvJ5kF1
qMbm7MJSBJ6iotIB5Eu6K+R/d4pbgqWjf2THDIBF21Dyc81zhxtnVHsAaHNOnKUh
YUpDLXBNXbRbtOAspg/fJLVfE/l244sNTXxEOep4Mev9anv71geZrmgGIBo3jRJp
RcdlRvDsGq64EtJ9mVHi9e6TiMsPNYtFZm0Gjqh4Xa2TY9CKdO7zEMgQezZ7x5s6
+F98ne34s7CDReFQ89+AXRSF1X1SP5agTXJue4l/NqdsBF6SJE+z90uGaDUCmtmU
shvcgTFjKxvECFBCwRYSU/vqeo4wG6BjsjpTSV9t1tnXk89jwBqOockknAceGmos
E4Sx/Kuxox4OjGA2wDAC/+VoAl2g0cb/TodmmdkW9PTY0mcp4vrK4BtjXT82UdMg
hG0AY0yJVBFebiZ3nayg6CfpYzCOnjfOC7/Wpx8YosySxrV+Rm46wE+KDRzeI+9b
QWey+6V2ekHj5FArNm4VCAQl0AVJqUUw5RymfLmggyHjJWKb854BInXhvK0Jwp4C
PK4guhTIws7Rkaf27kREf03Ict49z8scXzNUWRbKS4LLrsJOs3KWBZxHicCs9eJY
Aa8kUSc19O1oW8+VvIY5VUkHnFFVPvO10GjNmx6IB1w24mY9E4btw9O8MSSAcfQi
F/EW3kM2+w8hkHYMmQr1JlaM+BV41ubXWapd8F+p4xeSBOowHaTYxb8jpDnVwcCC
c1l4ai5W3fkzaxjAs+F/tcbeUy21Ji0qHokkGYqNkn99Ntrt+IQMLuRj/v6okqCO
cLxRkq/Lz+vpjtMTrpEtKhZD8Ee/ko002jpm6lOw3fCw0+k2RVxy70YGF1b/yYPT
43NbC5fUrcGINDPv4XbIhLtEkhlvVPy87dh4yA1vX02LrkoIMZgJeC0yWUDeopXN
lL/WNiA4lr7AxoPhKLoWl7eeS+u+LGPoKeoPlnv76PSp5byxG9sU55PLipRMBfiX
GNtLPM3z/8klIVt4/V02GrS4hLpp2NO+8L+b3Rbuc9PYdS8oeb1oxijelQphXDgX
3L3LMPajmh66Cc2nRaGCaaIjbbJBjMC9r/0VjKqVngMzPtghdzHNB4RElNiu+oNB
SF5ujhi1VeqvjYxi8YL2uKvoPy8fb68SZKteK7jgQqW6nEPSO/NMYDvmPdds4GGz
VX1Pp8qr4xmyZQun8HejavHnQB2IMOn67pFJtnNlTWafwDEebBzuWuGmyZvZ/1Yb
knGHq3oCpf9lkMtJwz83cJQRRYfLV3s1g+9svlCKQqVsFvBDrTM/QjXrnWZq6ti4
C5oHp4TKyBIJEk0Tw8xdBxhGmYRXagY6/LJhLRLHFYqJ8BcexPwJ1zRIzk8mWqsi
ylppT8ZV46Hueh5cphk57N0IX4JR69mz3X48HwKwcJs9WZwk/2q7vUXVKP2CK7gW
Um4W3+JVtwsbZgLWjvROXm4lESZQtVTNbhqj5fSPDDb9RARf28ZxFENVLZ7HPMoj
4/1MMmbYVHbYdHnrXxIDc36jq6/68Ow6KimHJnc7x+93i7itEil5l9P94JtLRHVx
mm4ndc6p+ia1OUbiobhcY+GeTlwzUAbGTvVO/MbQMpqaXnqPilGwlQ7i9Us7dAlG
4L/h4T5NWqUTJrOf2Q1YNkb4nJM+1qt/ufR4AwrMQgsNb51QURLgvqQgCO4IZBlp
HbGb7FYTd610ZoI8zvnEkjOX7mUqKxCXJuAKAHaJnTCM4fzUF0Z1kTxnzShkPQKc
bCmoV2Cy9rpEIYctugs9sT1fKenORORfkhMMayRfusjI2Wja/rNRZnaanxCbuLJP
CLvpklID4FrLOXvkhij8spGuScyAtp8uCKEQbcKCcC525YStNwBksFVGikrhcW3Q
mAONEEWOWWHYPemG5NNuofiI9thAhAUXPZ0LcJ0cGIzqSXlVB6vPfNXFiZ0vVooS
d9XE3qte8988Pxk8Bx1I9BuvYv6RTHVUHIbLcYK6dC3yXIamPywoBbPNQw8ewMh+
umIYOTpGZqzv7AWvtVfPqKWu+o66ouAf4cF4iFjaPOyVGbXynXFBdqhLEi2svsV3
xDNfIHb0yjL55n6PhQSukDY6+tFXqgt42UuT+/WBcne4w+9a1LMOQFAD2rrWM5Wt
HuYb5SmYhfxmdQXKyXzG5g0e1GYHGNGgYSBEY0W3KkQ++RxL6MZaI7pzEzIpFc0F
hUHsvenPnEDjTdvc6ft7rdVaA3Zv2Kw3qLIUkBJjpPs5dug2Rg+H/hUd8Dee8pmW
0hpqGD15tw7UP9g+hM2C+mZKhKb2Bq2da0iOImHMLN+CIVjFp4UgmG9TSmHwCnUE
udppaxVVMF15QSTwn3NRVScZYWhVp20Uvc/e/cW5pMzzuNSIEJf8VkW26kCxcb5q
yw6PXcgyd/aiGuYk22gnm/RIJieRRPQClbcQI4IdHcs6hwRuzTyiSwD/bl3+GSah
ptJ4kjPxd2GGhJuH/y55kB3gXc1J/VrZq9JYnrGh0UNCX5WIXow4yH4V43hIcIvp
FMI68gzMNzyr4Jc1gXerIrhU5mlFigJBoHsOgLbnqQtnB6HsU/GGWismv6ZUmn5h
fyIXaiiwmzCSzqXrCbF87+Ke3FzZY044S+swX56qB0CVo+OCZ9MQnP0+CDHSj++1
kQCwJ/jc2kbeo4EvuIdEez2yQMb+o/qJfkSaqLuT/YuVIlePdgOLU//ZBz9m3tuq
Qm/rx7C3sHEp5Wv6ioSxM389TC2adhHuMOIl3rzrGPHQo8J/CSLBJYdL0AzoTVrM
rYoFPwLg/aDyq6i4ftcekHS1GYL/Rd1Gu7TvWUv2Er5xImG90i/irc9K2vG9kwdp
Q+GbGEIXHeoxEIsxdO5kOBnpsB41aWIZCFJcfUJEdWtjqkX4PAwrsgk3X45wW0We
2h+18ctNjQq/8mQZTTIYEN20sXN3maf4402rG9Ih/gFcM59gXTDARdRYxtfQO6Gv
Lb5LAuSwkWlPTThJWjyt40JEuuqSylG04ZSvRti07q2lYXkiNaO8lFyHD8kA5bh9
9pdLRsNMLl9dCxQ5Wy5td8H4eImfaGhwuRmYz0YaOc1iG169Ml3La20nPJ6Vo6G+
pkqyJIkAQ0bShf+KQfQbTNRgOcey2zCi4MrtQhxCtr3+UFiFzRXUUnpMMhgMhc+N
dpy9uZGm53tiUxlUWBv5VXDogFRiHDpygn72bKPrQvvBJM2wAWex7QnSzkvW6One
/LpLm7TAuTOPXilqDGDhYX3sV4RaSvhx488YaR9UGIZzKNDvgLyrENp4BMtB+hNv
RuWWGDi3x721ZxGVyRPpBQ0nnDjNCyq7e9R28NOP8k4N9HENe8W9qy4VT6EzchrD
ZTtXOKu4votrqj9s/w5MfwPlX49JR9HJ3rrYZ0zWsGUBejVRlgjbpZHrA3SWJ0Ty
4Jd1MlvUUa7iGVbTxqlhMciRYeKWW13tVVPjJObzIVm31JcF6ktvTmArvI8ZEVvm
8LpkU1nkbHr2gTnCUkyYQW69o4G3wwB28LlKh0PqbB1bXePR5xjL8w9iq+pcpWrj
qmo0FrYJVGUT04r84Ao9hpmzZz589JNvG2Dy8PCNdEIgS3D2RoEFsHhkefzl9bZs
r+3+o6Ro2vZtRxD7Ug6ZA8Hk2FjQaUFmZP5HolIWGza5mh4Uu44OUOY+uOYzL+oo
bV8mQCf3z1BO6bXOmwhC2fRCbsK0vN5iI+L7QXpkINO8P0zgJY3EenIizYn06Z7W
bNf9buIat+pfiGPFxozb2wUHmgDPhHN/c700/1CVvX6KBX6vunf04lz95XYRetEe
RCYwYZtI010ah+mskARMMutHWnpfiquz1kO7yS8g0E/uZiFCGFztGVwpOqmbaO3V
omtcl+aYkHHQUd13Zo2QiiG57hKFxTm3x4gv+rz0TsvLT2y2YcQzeBwHvAEBAkI/
ZcRT5yA3LIfkDWrqPj80XaWDBEX9QDa1drc+wTIF9Q7RmpHAvPrHR7hlG4pi9Maw
FUW+v6ieMiHmJyTSbfHcJjvQimCp1xg+YIPpkBKQEtTqcyze5pRpLqZY2B00LciY
7FhD1HdWlBBLjTcadB01MDvBb6xb0n2A4cekK5807VaEDi8YGF33NoCgO/Ymliid
/3O7mBwt5CDxiBQqXt2LXA12Jm69/z/vks7XMUPrSCFBtDIBBvxBpHJAxCqFonAj
6X3wcST8UtQXyeKA26bI/bTwmQ3rAejrEGHfUMTSlSlBjGxvk6DkqKnF/Ny7we1U
YeEgmHXgZl+z+B39R17F41goS6jgw4A8j2NKyIhpUJRlIC2bW+C77jlMogS1HxMT
oTDgmoyXe9/O/PMqEZ3EViwU94ouB2TqLUHWVt7Cg3vsUecmy0uQOPMGPijC2pKn
QuWmXTQhL2XVLebYyGeub7Xqx7E8DZkI3jM1suqKsnjzadW4+HFIdD82uT5stqKv
CDQgRsMz2lJQPA9uggGI4DX6gACnuhEmBzEdI0BlgzGgYeXGEcAvHBdWkI10HiBH
yDJTknmZnA/408LJTsEd4m/TlT+b/9ngHlyrUIhEIVZETktDQ1ax3DgjLRsSkk/9
BCDKK9tQPRJVrOp7BwCABZXpTNudVenM8mockwZto1tbNVO/mcm818jIjBnSz6+u
XdyibFH8c8FNWXFizG3dT5gNYQc0uD8TNR14UCRsDa5nA+bUw3uNTSdJIGzpvxrk
WrlYRwEbzFE05cYxCasV7HydXXx9sAdBEEcoyXykisaaSoid9jNx561lDznTls4T
ASIfJAkv47oJSW0g1CbWjaCZWHUwgTFohFBlZQhxuJXjmLfDiA22AzkLhXfGF8CE
1PtMJBIyli44LT6X2IYnF18rcOwhfz6nZULCmtUdM1wl3hQMHlrrTLDBK4n3psEX
mJ/xi0FXrnWokbZj+r8ogbtbL6fKtoA57S/SA+Kq2uyLj2b6vlxn+PqHZTFjhUCk
HA4gABA8+lIhRIqzo6/BvP/zRV85llcTBU6tLt3Vq3tHRcAF3j3oP/S5ES7VsxVX
9cLvDTY65WY8MYT2hxKnh+PPJiJ92WpBrGkzrqvqZa6IWyHsyBZfzg5L2LUxvLCU
k0dt2gNNsM0OHc1WrzDtpuo3Xovt+PdVZK+zu2PiRitRezG6P2oK6HZp1tEbMn/T
/i0D3aSAHQ/h2SEiOIcFjAzx+UnYgKGkxWE+vK8CVQ9hRV5fk+XOGBtJez+E3Dxm
J11fv2vyu261xGfKNvdrNKv7YNt3K0g/UAUhYnf7sUT1FeyyXRlx4FSLRSZYVtC5
JVN8P4TKmBrTEilOK2I4drVbh6pRpW5kyUPomQ53AlWx6pE0VpWC912frPWDRYXA
8ZCnPw7S3/26YO511RE524c5vsWo/p3CU0zznbqx0gf8niMgwWUohkn+RyQwY+rm
JSkHeiyY+bYZZWRPKkXDO3uWBLMgGA3QYqOVb+cbtccaniOVi7kdLIxynA6f9V67
rVN3wcF+pJXIJhfIpTwtw51ZHMQTHCcdg55r0GMxtEkEJVW34P+E8UcZDzh28TDS
eLOCipWwczeX8OKD8ffAaeeAqgn6gWTmamdtn6tgWmfzfu1r3geV8U4mwYHKc2kr
FZ+ZUZdq0NGccCKJjis2YJ+gygjMIBHcptV4c1J4Zg19c5bKkyCRMyjlVLXAZjwT
beDv2xhRxYLOvZGeYZaKUS48bdmMjQGWVkDGp+i3oaRNZ+oTOjSLmTlq2p4OCaCC
hX9crgUaVfioVdB3PvIK+wg/isYTws31GKIp5hva3S0Kn8i0SS+p63h8s+XpOaef
kOdPUA3XEev8q1wXO/CvbvOfENmFEqiV7aiVRM3kILjY5FphX6al9mOCiSDWbk/y
to4pKCp6dyo58Z7MqxKJkXPcpZMJr48rawjgRdIRUu4IlY9Ve8xoPr2Wutb6yGhf
k+4wRI9huH5u/xyu1HCvE6UynLBnhuOvRAe4qv/7gBlTjooEy9alsAzbVTY3usX/
nmobSUl9+Dp9WhEJAUGFPpbIZPBXewsXuqM3ExcOfKviB72dOfgHbKbgJWewkXR9
fSjDu6oAanexu8SwMdAgjG4EyrpBVat96ffefb+lDV6b2sYgan0LbBqKUrqA9xR1
na8ZsRnBc39OgzSrJ9qVW4fck+IUUdutyM7b0uQeZwcB0vkpTOEDWeY+pyfraYs/
iERHs/ZjfX1EEkDEXRM7HrUTw4N1VDeYXP3bMi+j5JxkXoJ5lZoS4qnVW0icz5sz
xl6iunqxTEq4Ur8PNJ+lynu6g/WtzGRCgr4NyY79j+x1ljUojvGMspefy39sJl47
nzwg0Pz1SuGDWK3SLAaDS4TDV5ZIr8f8n2GmAcdTczaaNdO7LmOam942up0Q85y6
KgzG0359q75H0UQnxB0ImAxr8tNEkIfeImQfFVg+YOKbPxpRLf7LWE4RVJgQwPGN
+afrC0ve7CFc1QpGB2D+omqGdl+f6J8WOvKfGQvSB1+yipYdZ7dmmCsM4NUe1Zul
nD/PQFWb3XS7Aus7a1ah4TDALNsK/E9QGLVZ632bGOnmGI1GK+NBSxDf37mZU8xs
hLX4HDknznq1mCQ5oHrQD82rFqIUbMKFcQUf6Vdt9d7y0bqJt15SHUOBtaclA7hQ
bl3akBhXm82oI+T69ay22ViYlx4rzOjiJFxcvPmPjIGd/P+9kKH3/BuirVi8m8w7
OdR5l0S9Ys3eYnIVA3vVe89gBHOX3QTq2aUixG+OZBHlL/w+lF4CMCu7H86uUmjh
DeHbIWhFP/0vDLNwmoe1ObqtRMGLXMgAZzaVuEXZuprbhrJblC/jEESdF9qCX+9s
FacjUcKC/iyZW7Znuy5LFTI/JJULNaT7dtidCgq4cR89mFBGjIjKdacKbKaDPI71
qXRp+03/NZciGYa8Qkj+qmT6PBQltJ+cOJTiB12F4c5U8eqAcGnHLMX3KwWwNldg
VnDgpSnmBgFx0XkrRD079vNSY/1AOQV/Bdh+y4+mSbTlqxmr2wPq7xDNZsJM4XGy
RV1IrCohcnTDVSCSBq0z/TJO6ZjfqagsFFKzht6nRdDO4D0xYpucqRAL7jdgdxYj
Kbe3qcesfqcxAm385tX0IZLvAF+LAH62UG9PnTI9wLGFMI4cq+S1DggtRKEViqmZ
SP/DnMUxx4mbnZQHWUJ52CgcpG/1GJzL1RfmtPVak/GpKLIM/q5Iz3haAME0EeGf
R9Z806NpysEpOI7Qco0P5yk2+OOZps1mabShj9vHgnNOgXdb+HfTmm/dtnYz0uM8
CGAGZQWQIcOn1zJV2kW4eq9sG4PxSQ3ubjabej05iQYOGq85PNzeXsf72miEgdyV
vgVYpk2Y4ZF0ipcXbQWdQ8A+JnavLebI8XrRAuqwpervTa3vB2fr4AfmMLd01sIb
Y1EjGu4zddsld/PVNvhydJ3joj4IM+OFDYvuWCshgBHVVjn2Yotwrfl7QaV1Ubal
TMC4oYfJ1MjrzI72p3VQYLQEMHTWr/PqABpRBlIjvG7UaU5N9aFAbiF9F43mDmEO
yAJwpY6d4QgehfbE6EoQ29qLdrotI5HaK60bTZzIvUGQ7c1ig21q9ZASzZZ+3/wu
VJHbkEDTb+BUAKjLcnV5sJmeAhAD+tOdWhyfhkl2XpnhUoSkkmAwA/1H9UliAMhH
mSf5gGBUNPMUkonXhUrnqA6/Sbkvvvh8Zm/JKgo3Fcx6WyRL7lHnFoSrw2PYyVFt
k2CfIMonpOMHL22jKW0g6cKHgaG1z0QVdWeFEZspx1AGAH95xZCRYINHAB/qLS5T
nVcbCVvBVQdrptpMG0Dmc/TA8Hz7omurG7a5BSm0fgWo5RR8Kc8q/Oqb3/2D8ZO+
pdKEwlCAwL9kuuAx09Kd/mAS6P6m+v3GFS++2DkUk9OuoXK62glnjMdRHF/nQqN+
4eCX2RVcGVJSYBmTwDFuUKBb+n7XQVH1dC5DI3fzpSbMCkTLcswBmdKOAyEwR0CV
tTp27pWTZllR6Wl7RpU/9IV8YNElT/lUJiwXNnxIgDnMf1Yja7dRT+xSX/MTRnV9
93hkPwPUnbNOiWSwSAJSFFW65InKO4Z8vzzmXTnOFoOCcEqQXQqGPJF7+hHTqzlw
JS2R9gULfM9lQtmRVIFpuwYZoaxJx3kNW1j9A5Lm/xCDG+qQQIXdbP/kJioueTeL
cL3+0rK2/8w8U0nxDf1MKibBaWEHE5sfaPcTkRYVtOheBG6RlPf6i0Rm1F/v2VQ0
9aJh5zEF8U1g9t+TKqQ3gu2+fdfwAEzNnOQDY+rITxUmDoNraMvegfkNcwdrM1ks
EP1Y4O/iuwar7pbq9aa9+TDfLnwJlOj2Lu30/gZCGfJ4ymhk1HZLmrRQqAcSbCM2
QFzvjrErlfRaSVSwANfV9pSpbmMTKJlOBDc4aQR2TwtLwbVoB/ZYOf/c76bUMQHT
f7XMTydljSDmCVcSXRDzg8uNlagYgRtW2XyfNVgY5V50z5gDInNpPZHqR6WozO4D
Ae2iyCsKOyZNZb/v4iw63CM1rcuFiDzBjQ39MoETQtCILTETFYLsIsmmI5XkUOta
xIytg3C3v6yHnleM0yV+fI/DQLkK1/k22P2DdBi/Jiw5uAKkJ2CNK9dNE4CMk+Aa
Jfd+ErH5AyL/ex6Lm84XFHO6rfRYAJX0FYrPJfHhL5KnB9un4hl0sLEVlrFXvyL+
nUsqTVKeoswFFLQuGA2qk9mAcZkXETlHGjbeQHjn5eHQNCQYJXDeCeJTY75wsiIf
H21MOJAfNqcRv6twQLg9fuJZ9uEIXBnPCTOb6Kcg8f4OY5l7ctOMwZvo9vrEIcoK
OoLcQnsXAVhqPMD+PzyP+yVkvkXQi3ps30xb0Lyg875eBliGvKx1C6TKYI7eLKaJ
kyZbR1T35oIpsPjJiMGXGcPPrQ6m4Akw+zn8XiVsRx+VpcJjbQDRofpk0139zgG3
TjnZhCnD5QbdyO7UpXdcEicyuLZPMkSV7Jw1tSzAVFrcZMtG820wAwUWFniJillD
Xy3LmsL5w0XEp7rXvVuBREiTcYjHmbQh+tk5/lajsntyqBNYgPkmihNf4wFP/cSC
H5svAVw1/QuCAm1i97pfoaosQaC9vuYTgbo//dnLKCiy+DBjQB1ABe9ZyH3xwuex
umnrLtQOsWlF/lSzT/o7xr1FK20HZtonQPRDIeybVtSHmhgIHmWeGxBZvVQotUCy
wJB0Cb4yPeU1I27rx/0/zJLozUqq+EbpMUmczfCe3YPbI1/u5MW0jPwc3qoDLsso
wZhjH10lY9smJQXKk6AacjmerH+uZ2NOYcBTXix0EQ77CJsNsFaPhP3k4QhmHQoo
aQkqRt9YVXXCKguwuLqpkFcJMSiqXZhYToyRHsjFBPuKnBn2rrLIdQuHEffl/AyU
yNcoygV5YDgis5UzGl5a5uLue8tFcGpj8j6+05H7ebniY9oIN3y2wLS9lomoEJBl
MGAJBrmVCk4qzzgOuG2PumBUjhFZmle/wtfRiUEZESOZV8PqQ+3/VuW7OxuKInbI
VPA8cc5hNETEpU4OLAqu8zR0rnhtxA156imNLv4TA8rknyjlz8xaaabyMZqlgaq9
OR/WVwcHJtWa2w/YkC5oImHMO8tqoQV+6K5sleDH9O5LJByJttKihdvkHfaT377E
s5CUAItMBH1HHHBC088q4NFsiknDAllnBzKnbUKNtk0x9Wgml0dsVjM71CJ3rI6I
F3CoWbT51iIAOK7sEAQ8bRAWNDrki+VMKHkdmxtWBJC0apjvYU9Bq1toLdm6EM7N
tnQ9PGg4Wg3NJafXgHmlnnSwl3HdAxWm4G2Zn1g01KfHy9E351rt5Ouk8ZpocPsT
ozYIorAAf+JXUV6bn6dmi5pUwwTdPYXaiRr1Zl9jA9SZOe5kWOKJK0iRiIGUr8Oo
Kq7nzf2ihte+5bUoDqFb6prY6nD2DYNemlUDwADMMKjCWyTB1OTE26pxqJeoMkVY
qH+UXwRBhfD6wO2PeO+2/nl0Ufc7GW1+WbJ1sjYkGcV4N5uMGvrVujXKJi6VnT9f
L5oAFSkMY4pVoB6E4uHwmcT1NEFMqB69IUOklyVjzbcwOR7WlwNIqOgSmQVHK+yp
qKl5y0mrb2NB8p7J2BJ+EeXpJXThRcmFfe9vnoL397F5slP+/M11OxlGQz6xE7/u
5C7/M0sqnsEWVTA2ZxCLBsNLiWnWx4amkG0Z+Vt8jE8YtGIX+5gv1JePDrks6rPM
FZ1KPNpsTSU7rOiqn+scIrmDWi/VXG1sAYEVSRTX+IVBlNAMX4SBpSb5v50n+TNT
aPI3kgP3RHx3mGztxmg2LfGOpGHpJrXex6WpQ/xd0V6J68RwOiLTPTH1sY8bBpNJ
ldYKTxtb78OdyKL6DwqAdBrvzynfh/zmCEyu1BJke/9I0nX3dzsWUmV6N1rkQptj
Dhp9C0RnH6YLOj5XjifOT8gYhjUQWzmmTD4Cxe3gLFMQdaaWu7srv/Q7IW2rEZcB
nhh2v9wawdQ5L0pbPw/zoG8U3kiqEycI3m7DYshoHx7GVjU2kxPKtVytJe8Y1sPn
hBk63GOMBkILoTT7LYkufYEvnjc6gVlZoCiS6NyWPQ3jdlfFdSqVaj/C9G+Ox/rt
Bm/f7PV5GxYAKTVXB+7Aohl//DlQ8M4R5W0AUpsus2sQNUN270/zgv+88z0EH4gX
CVxBf+kP3lAeaS+ojAvWNMFqsaMOZ6k3XwR7JqjtzlY5Mwzle72xWSy663idQo4i
5lcf0qkMIWkbWrSqMbd8Dd7cIIewM6M7CZyT200aGGZ5H7oiMKbjdm5RNUi+iq3D
KwrOJ1PI1skZDir7iOqjPA7R7QbJCDUb3K+wk2I3ztpM7Fiph+ItKp0SHxn4c8+o
OydElFVpxiUGvIXvQPkWUCR4aZeWVQMLgErzcicRnAsAabxF1288a3NFUjat0Djx
1NldTwwnfkC5L4rgraARjMjoYLx7ct4y2ljFWJhbIC6b/QmBBjoaJBCSnl8T1WHt
5tGC/9ztgFmnSlYPV/L9r+uDITJXU6kvx9jWLDZHBOa094YMy4gsHgqPrHYRofIL
tiGDIqLFkboL2UREgL/H1bcg1Wy8/rdB3va9ORj4epi51ToMATLsv3eiXZUjK1x7
CfLaLdLxEqOcfK0qRNbKlkY7BAy+xjcl72n+ZB2Euy1yP9jf/ypajqXNqkUjqRnS
ygMalFUXmUaPhX7hUIrG+iyk90213BvWk/xxgcqhDXT5ampkXHU33BNwklMaunBD
rwRV1C91igTpmwaLYdFowGtcYPCTIVNVLvC2YxrCYA0DEUeTBMKy9h6bNUaFQY7Z
vbFIylFTDsEQ7KWuUdf4LTUiSypwflMpfn2Fk4OSO5ypY/ibh7TblOl/Sca03TXO
7FWHxh3N53DayaTSqVMS+v9sXgrw+Ea9QR5guq7aaf5hsXQTGnB89rIY7JCs2wo6
TXBEHmnRhWt5z7e92TErsvOYP9VLW9yNJ54RzwUK1mRKYw8pH0HEj5OzNP6ASRJm
OYe4axBWErqgwkGzAtj1P+94XjDUcr/gTfC6SB2i04fXYpll0JVbCho7TRzcx9ju
rBP5TUJXyyHUcwqEbkRoAIE4bQrwxv5/d/8dBGqPUS6ZDMoDXTOFLKnRMvqA0NhN
lOGrQHKzo7iuHbxHqLMUuJrxVkeH16HtYRnQxU/Oq4cZdFyQIRrqDev14c/uG1OX
sWFSOs60Uuzn2GsXkr44HRL2MzRu96RQ3GYDpds1ITsmWjwgCY3/sqDUKGzJ1CxX
6emN6F579hfu9+mGNb4OqwiEnT+heVNF4DFSMOU7Vvri04szZ1ObUmRnrXqwE/V9
MG11F7dXPyH0BpZvBpJKnZ1xd5mm+EzBfQutYgu/bwtvLWleinF7yqAaxTfT0e+d
RTaCy1C303fxVoMNf2+rOnez0n8FdjZkpJcz3l0qUL1+2pGhSpPGdfPsi1oZ6axh
sFdJLWi65Q+4kR7kL+nAZBRtdprD/C8749cMk3N3FI41ssCGjwS+XaKAhIGv3nts
0MJO1fBco6cHETC2sRo7SYAl10lz+K3HTb+GW7Go8aLY9NiYbHENOmMUrH2xh5qR
G++cPuKnOJM8xnz/bhFfNLjZPCbuFJgaj1reM3N6NqSZ/VqPyr7GhyCjTZa1/H1d
v/gOh1aeY70EVw1GaOi6NRAFxVHJ7BKkhdCSnwdgFRIM/ws4YZOZnWxTAhZiW8OQ
ZOoSuNWZab+CvRXjjxoB0xE8e7ztQlVQiSWvhcvXOhWbXJVsk1JQ5bjFF2Z9npFT
+KBuXfCyd8mAafldtTGBqtizZJ1UftVlztnM33RmpRAn1dslz8A80GYTA5tN7VWO
OYZFkaimH8X0J0YQ8Ck5XZxwlhNCSmsalwwNoZISh6YLDP6ABKLzr9iyNj1SWs3H
qGK9zqyr8o/dqJolffSwHJeIpQ1b7lZbXrgC0qvxu5oVEYkNYN9vLS8LQgX3FhoQ
0ZZ9u7XJhj+Bjlxbjap4mBEH3jLCfvbHy0g4oiRm64gOuxWl19vUuZcW1LoymUcq
qh1Sa1QhjUSPcaELS8Y4b9+csCggGyhR+JNXfTJg/16FZepqpbjUj8BNzZOTixM+
g501RHZp53hXcG8KZElZih5DJHi93t7Mq4whCfKafr+k2noYrcwQ1EKa8xdO10JS
Lc3Uf0QbJORnXH3cRXO0Hv9Mst29aEIVDtHpMfR+9WOCVHM0/JDN2p/VEbclraWB
DljRC+U236mDPm/HFRfG5zoq0K8PNSvNGu6BHX+3HHJ2kCiUINABEaTTEqcOoBfs
LqqiGRQut0zjcK5P+OW8IaUaafxwV64yLSAH8CLUulvVOMRHQbUotfAqsx7OTrW9
4zHNvJL0/JkPT4RNWNge1d6wAwGYQS4oPd63DwVQMfQM9Y/iD1QL9b45f3forWyw
jafjczgJHSiNkRsGJp85JayFuW/qMLkQBCYop51fORVmkNqmgCEoWs6r54cZ/xzK
xOT1gjdTw6HIMnMdXnSTj1zhjawF7kjYrDhWlltUiokI8p1IR+8C/7bgEUwN1vuQ
Hl07/p7F//P1rwI9zj/ya7pnbD+dqF9mBFAQo5WKfmBq+0+fQNoRxp0usaVfIWac
iaNo4gHCVso7oIR3WhuwMaYmKgU42cCjDjMWVvepcuaRRLJ8R6I2WWpyp9f0MA3U
1TfxQbts+Uqa1rJKQeEro8MUrL6NCMD50uhO+pBvGgqzfHmJJ5w1dJ1dZsivf6iB
q0qFRZBjzZbR8ei7Dx5iPDrpQi18rFWdilMqJJPuPeP6NkYGr/IdsunH50z46RHJ
44FtDQUUYc1OnYggSIihe31wLYWGBVJUHWwJda4q8GhaI6hNscjUSrNQ8ac8cavc
UkVoxLPNibuKDHqZ4o7QmkKoBDcbUB9bsfpHcyInAaMu3jELFeKly1u3pLm81YCY
0x0lZva9lzvk8L4y8QMn7QFxiUcLBcS6Us+1DicP/kOeEKgdteEHdzg2mSpjLCb9
kEe0JEKBI1QRmpyIPIKzgX/YXeQ/4iOEMuaqyZWLMHJPM4TxBVvrSNgkc2dbZxc6
KePclYvPjlmLRj8eq47HFeHupX3XGIMDE2atscl7mt8pV1OFM5qPc6M74fwYhlZo
u74UPQWCKfBjXQjnmB1D2QmvpxEDOZlWNTN1gM/UDH5YGxJ7K/2Sb7nxhunecZYG
UJGxE6kugJNkwDglOGFCvzy8y2mwE+9u/0snRe5VeIgad0PF/cEYd1CIddNJn621
T5rv8FbDLSpNGILOFywn402EP/LxQvQBO9iIFlYDHDZh7dy0jRwUGi2x7lsqFNPt
DFgGJ4rLIo1AtGnGETkc1ChlhsVMJyYZSTeumNfOj3z90JRC3Bep3EDAsoWZAFmt
y8If9S1aT976vMkSqPqSDIehf9ZUXcS2eDnxXhaJMokn3ND2BfPX1dMfnLAsi5b2
LjEXMXK/mFxnmgVLKxg+3Rvsp82QT3fbDwb/rUBo4caDe3emoiORxveQ1Wfo9EYN
f3DLJNRSbZQNb9XoY9qJYwqbwrzt3tLwKdZQf6PjZ8ej6xeFxkB0vjG8BwGfv1Vj
slYGRIy3j3pq7cmGqOBDAgUmKDsPElj/+6TISZTwf1V3eCo/7dwQbKm5erie7IXC
+1X8btfQPVZKw2H8fslStTKgNigGwBE8wtrD49VyIBzGl+Rve1B0D50vKqqA8cfh
xWH/xz4wwZ6fU1NjAqNUlUnuVuENz2ZYL9H5YlIJpay1qfY9qjzdntrMTEoc8JML
XQ+QOxtpukCyJvj0lsBV/pp7FkNIcw9J+uiCXMZM1B8uhfTj+1fXgLi/gLkWua5h
qm0NtdKdSNsmj4etB8xfsPx5IFC70L/OXwI/7oAmLqcCfxqMWw0xgRgMI8vMZZDh
0ms2DDw8n7uYhxLMFPZ3J8SJ58z5qemS/VgN0LlY4+lKs+kAEVyqc7GzGQBUO/A2
I1KAEafjsCWs1NExv5IX2xUgPWe2YqWxf2tstZsLJMfIvJ7jZXCxOC93vfj6YrUj
xv+g7QI4PPZ/cnqF/StUyOC6/93/TXDIm1bVA9LwzFc7+1NKWU3RHrc2nlHC0IfK
CBZpc+B23Ep/lkY8PL1mRjW77mOzV3HOhL0A8AJu24fSzNbIL9MpBJk5sKAxCH9w
kV9Sg2NMV9g20APgTRkRyaO5gbuo02gGmTBc9BoePiSAfZ1bR2PH9aXj2MLmME2h
l7u7CXjhxDVmMoYRmpGMK9Qv964YRUD3yEXPuoR3Irufdc6AMaPS2HMH2LfHW9YE
Q7zKsOTES28qLYdNGYqKpJZE0jwOrfE/wyEOrQwo/yUI6knE5MnLSmqHZndiAgkm
VK0l8t+/HZcNW9sJm/Qemr7twdO64ulPO/8kUG8SDiVtHyHGkukZJKanFBgpHfWa
60KOJ3g0wD4EvjOqCUK2i1CHhvEe3jXAMySh2yLWsj7GEh95xgNAY+7+7MFrGVjT
5kw3bEZ3WdjqSuTwX96xBCzfrDQCmfW13vN7Ot07Z+AJJy7xo7ylU8EO+1SEUmZK
Mz6vL5AalqLFZvcWXejShjV3J9gzh6EDVrgT/7dx9nqC/rJ2QpW6bykHlDG+j3aG
yUl27V5MIx4+QXHu4YLsmc9MJ09jpRDKeOUSwDcVgka+K/0maVRYdU7p/QpZj1wS
4dCYi2fIItFKP8x66r0q2E3akVbidWMlG06i58L2950OwSog7EUMaXiJZS1BRWn9
MyQhR3HceT1jPS5onV4NmYKYDNlXRL0LZymba2StpdCefOepWp0ifzdnqJ6K65BP
wxTTCzsW4wT1Op0oXqsGpiwwNAqGPXSVQcbD3z5XrylQkkpBEY5bJPuOm1+5cWze
ApdtF/KpAlyHu8WCFy8jpepPEj0mstHFYq+mbTE9+pIpd0IeKpGGp+mhxoMHpxzD
HqE6YS7IJvE5XgyWpgACWE23WDcyvjLfMNj4XlhfGk+nQ0bQR079DH06e26ZLly8
TN+kmvWB1GVlRp3dzy1GURyV152cLzSUBy1P6aZpkLTHdXkfQKzH7oa7HoSqxdwj
1hCcCx/k4iPwV7zzWgXF9dA/3V27lMRqMIw1T1KgY1SQ94rURJWQeLHkAhXdkPPS
XjzTJDhWWDBpXbU7zaG+3iZH/SoNYvs2xa8smfx6hHgtn5oL+40BvXugqVOTueGI
pzHYQ87qFQaM/wB8fKX4lbOipqjerUDAoYM5PeaNsFHxc2aP1EdVkO8RWUlth5l8
9N0evBkvM+QPBEJXHGtfdpK1ioskBiUB1fkRRgQpCuDWdBe7YemmJRek773olP06
35Zpxqq4vk/mXxJirMuwShCN7MuJon9rDT/hZUxmJ0o/GyIT3vzDUe+qy0WDn5Hs
bKsWv1HYjW5rFV90lKWaksstEq0/7enmrIC9lkYVtSgezdsvIC/VeyDvaDegp7KE
MNdiTXjyJlUjBxCiscSljxAY8pWioF72W5LE9QWORD8cqwVfnWCYOUoJnffuArz8
byPfb05TD+leFp0tZCnkmEs1dsdHY1qdAYez2c2Kd7sYWj9dMySJA/oBPG4LWY/0
wXyFTCZfaoo2WpjnlN8k+W1qz27D4ykLTMmYy88j02zAbRE+NWmZ+0t8F0TqL538
JYNDPfboOdY4Gn1el3JTmWE2Xez2lyygEUwJH+yh2ZMx/64wMOgHGwks/1GnyB6U
fXOqiI4TcQCZJQGv20awUGQAk39eMVJQxEmVzfqJLuUg1CBRV2Pcb4U7mHSow30f
tytcJ5YsCfyztwP0Z+5ErcE+RAaraeyCs4bc4rErhwLnl9WmKcmWQpw1hLSiA+Jf
r5Uk7L4H507ioKZfd0qdb7390VqbhZh92b44jq1deIkwQAcRY8qDTdsxh/vNPAyP
JkAWi1UdKd5jefjo1JoYV1ddGs4QEGdXtYQgPBIxVygInouLrCybFxc1OGuChQBc
LKUESZZucEnJ0tgHouobaTnF+LeLzbvj9gk+SYHM1IuA1WGLF0yvJHMmaKHLX6s9
MtUmCaCpzVvwXus0c4Vm6835e+Fx36sPjKw4MTOLkoZmHNbdvffEC2WVfgmq4pa7
zhhLvXRF5Ld3daNFzkQH1XW/OHoVnyNF6d2Otd1x2GhxlX5f+6/rAjv962xwfci4
Z4Lxj6uqRgN3acjRYo2645/GWICCjEyaj6KewjHQ1T4A2IPKwYThE+gUR3A5O0Cq
2PLoJRkwyPO+UxN0BHUUnPIntt5gAwxrM+VAsoWieTmrRvvGfOoKA40RNynH25Y+
lr3pWCMpi5mGpvUSojgsK5cavdmRzEl7ouoWU7f1JZC76/U/TywosuQAXNmAXCcQ
twYJJPCD57cLrM7HqEMxY/o1Of6mVUsVsjkj/H/G8LLLn/w9YNxfGHH5aDAIX+TM
kodv/lz+QpBve/M0cvUBawiUiulEXVd8KkbdiRnjKJnuXhlcYPjDoL00AnYPfSSu
aiag6PDeHbwDEszgmK69b598AHm4xyhgzOLExUeuyFtF3O7ybFe3Ol23uvkrhKHg
aNGotZ68W4Q49vHYaeIuBvHVh/BN9BXBZhJOhsl3Wxrz8sXkpLeoDbq7Yrd0TpTe
fDCroWp8qIv4Ln8Me6K/j7m6t+xoJY1xaYTCUebSWst48Xmeb6xTKYwwo+fb+bQ9
FkP3i5QO1a3N7mvn0Un/Y3Qig2ZE1MY9xRSroHGFTl2ozvlocvA0OtcKnyscTBRh
ezFGhL12tWTnht3a1cS6OzOisdipdb726G5/d0xsgseQZKClXnqCLP6g6k8NNb02
hQnvZ7GmWgNHYrwZFTHTc1K9MAUQ9GG4HAThDpStW0qsw5idi96Q8DT1aYaOte/W
yOTuEcJ0++9VxqWLPSv4d8IQKwgAIvhJmbg30MfTL4A30aRbYRpfSkBTlQphOI3Q
fy5KFN/hXwLeNjiYU2VarfsUvqY2gBh09nIY7DET0WjWsgNbLK70ccNrLlHg9hKf
bljTurt3SS/urdMEeA2C6NzbieRWr5rZgaQSPcLjbvlK4t8F7ocsir6YNjRmLSRI
oekxX6KX7M2cpq4PmugAay9NKRC4SQn8jlsW+dTEvzJAvPg0QpHCjrQ2YP+xzE4K
H6yQWZMIL8W18FppExF9KhoAskcvrrgsGF3y8UpyPQM2Mgw0SpjT6qCH0JrP2iOZ
JIJ1EtdkroZ1NEvIF9xlnW5svc7G6CAHlDpcVlS367uqMbyfmdbwqSnffTGpg2/L
813DPAFkauYylVZmRVMDcV5gXgpz5+VKDUhS3IZwTAkoP0zEFuhnnjZms4XAQl1n
FZDSBwi6kopag8F3tFdtK5Xf2eUfMs71nKZjbSW6COKOlVah5SINN2/XnEP9ivYB
DxbySlYMC4iHrpI09XQicUx65smO5YeZqOvuFg3M8V2uzf3OxbEVgwcl6lZqaA2+
Pas/zkSxggJIhJXixt4i/svCKYJSr75/pLWQ+xI4doQ8f5L+LSFm4PNLIHnxA+1a
xEk5URIsAhtLyMrNATwPqGPIpiZIwiRiZNksaqsQlwQ3kTC/OUTWF90W1v3YNQrk
B1Zf++aRSySiAvmN9eGkpPHs8e/nNi046os/LEDgdpyCI6lwmECTf/m2Lhv13yAx
+AkdLzr3xXfzu4ggDfFDENlFHhAz6C7YP2+mw9SJqNQ564Vv9OTJp8jPcXtNuoU8
G9LhfZKEA/6eldXoV0OoT0zr2sZ8XopLt1FBcMODUNuEqACVbjQqEtsKjoNcUtto
3e+LmFPBjReEWuGMJNUrHswe143WjX9SXqGUMmpx1E/lmYGeg62/f4CwvXiySmyV
RN+ytili1kXUFMERtE0Q7e1YyYCFj337JbIIpR9agk0zoi+fu9Oze5JWq+3uGoCw
AEmOJnnGQpscNDztLyv2VUigr6VVL7UuO4Hvh9GXy8hh6Us3sZ5f510l5vWwBZme
ENiJQgpW1f5BSMP/xxHh06BR/RVPVoS+LtPmHa0D/jhc89PmHIUPXr4sDE8dsedq
MeArE2oTPD6SXik+t0v2bljxMek3z6Y2tleNKHSn1hbFEM5Ic7JsLVy4MSo2Kq3g
OZngSx2Xkyhy2A8eqWIxVB9o4ZOqYE7ZxpU3eZrpVzWoBLCtnyCIsllFOVD0ZzXz
oKdFRz11tnqz9sTrDqT+PxG8sBeje3756js1RKcgeEO1haXpnZchVZN7kfFH3jag
5TDFokzNraZu1YlqfiPq94n7rqMkAPGY38YIyKRiNLCoy6uw+WMcDOqbXskCfJjl
Y9DFYey3VegX2lGAbtK8LfOg1XD9k9E2PVXFF3rU/NDN1yMzk4Q/t1cu+ZazYjjn
8spRQ6TZ0gYo7Rdmj7JQrGev6c3kM4lMvSa5dAo83lS3BGkCbr4jJR2vtWIdbYcI
Rl8OJ+E1s57L9RnrKmxR5jdtLGBQqGlRu1vhbZ+RZQ6/oYpzSYZb3SuhnN2G3NrB
TMoO0x7MyFPZ9YS2HJBOnkisuYn3w46skPAep7vhLccYsOGRO2KCsecWfYuLfq1G
6nZ4150F/GV91sQ8BPO+rKLF36u3JDFhn8DHnR3i7m/ZvL/ea/e3xn3WZw0Uvg0s
VVOgsgHhaTncLh6OREiyayAf+RoZyRWIxkQPR0RNo10ycllsdzO8YtSFY6M75Xbm
Bpd6YODY1MrKpbUjz6AGa2LMImpp+0MRXmrnnW0W3ZFohftJ6wJrUa4ya03Lb8jW
pjKMALn0v8AaEiJlknOfypOYlAsVXi//sbwBedz8wUslVpwtTQt0bBQkanq4VfPD
XHaDYZCAdfmbrbmysLYsONlVDH1/tbIZhqGstNXwXsHnADfAxqp6S/NjlrrCUIJ7
xx4bD8zE14RcrH1+AUbtN6Rc86tPr9piDAXmL/zh6bZVrFxOVxogmqiq4Hnfxqr6
NUW7mqPP7DOrQfE4P1toHsBD4+6XSK5DMu8xZMmLPGpnb41ZS9ZT5VfKoWDsDZlZ
ISN2mH2vQLxqNID6yjRUsss+a4XQdkSJG6NwqRD3yvc3SdLA8hdw6WPMMdTmqEL5
mrl7tSu+gLBRP3a/9vMfam5IuQb5Q5xQHS8WmymFln93qp7F6FdGb7NM49ndl88O
OSS/1B++z44HMuwSASeZv2X8w7qSvkx8mbkwc0l/Y3FxwiJ8QCRk6u64T6hIv7LU
N573XB2LRjhdzxt/5LcA/7OrlyHrgkDrmyMNwFSbGQbVbx7FM+mKvAh1KTsO5Op4
SjrB3+2bkThIy16M6ujvGaoSyltCWV5NukN4JKhxr0C8hr/GISQB88jkhCHz1tro
Q0vs8r3IhkhhEj39n+nQsK0mzColiAIfDDtihqIpRbxoNrMaPDI8ADY2kHuOLKf1
WUpuU1HGewkA+UYm0C/d82BbC/g6EXNzg3DPZnWNgy27xajl35Vn6k3dtasQa2Ki
DmCcZWRjFLIcizvX3ikO25m4X4q+Ttq3cdusEamAp6StRj6ddZWp6Tle2hTduJeB
oI/FI8wFNzmzKcuMfLBqYvjg9bncCiXefSbAn/Bjxfl+lCk9lc60rOqBGWzDLpNs
2oYWbcivty4WRQJLFCtMbS+RSFC/LH0apXCwom6y4u0SZ9N+y/lVUNx/tcYMYfam
GB9H6+QkgluOacZqesFb74+aXjNd7ziYLMXHT/thY5jqxBPjdU81uKaEISdyxLy5
0HIEGtgboni37LZBMoJlygehphVmMfxi1j6doGd5hHz6QAhZ+bEuU3MrPbZ0+Q3v
yBuTbETx0fctSwBxqR/gSIhjhKCE4E4d1Ynyc3ynzk2QfpjFnNe+3UBh9llagXv5
QiMw3bHKlM9VV9mfniA7CPa23NABHbE3X/aWEz2qfOX2OViSxvD33rwu83brvP61
7RU5BZBKt4UNpZLA4AP2c19aGdoxQ5wvIGnO4PZ51JUvUmq9fwnpOlBfK0Z4os7O
bRe2IiUwgZudWJpy+xVW3ijDpvWTYETD2IaB/FejHn+Ra8qljMjVzF+k0NyyT7D/
/k4Fe6cKGacLVThBVpR0Iz0J8TDJewo6wffDGrS9dP882qvDFcXYerLwwmT182Sn
6t3z6gwcDJbjzu5awCqGlUDbSGlYzHdRg36DCgmwOekagkBZBh4FZ7o+TyYNCll6
mOlLaINYaG2dogY67xPbQwDmRHVGy8VhwyLNNA7zebNQDDE5o/reZ0HgqCUyHWlD
bluGdQ6uAsBO6Gjlt7crGPqffRbcsgF3o0WklW1IAMOkJX0ei1WrCXUXXxq28Se7
I3n2pzSkwOGnqu2D+pHkzjUsaNndnCtz7fr7++U9uOSDd0+oW6FulNNwYRZxd7gl
9LNmRrXKRKir5FZN0KfyfgpptY81hqFbBzClF+50NyBqurtWDYudawS4ISzxIEd1
DqdUhKBqLTeeRtllRkC/I61VWl8bx5fq/vgUaJhsXS+NtyXqtJMYBIlwa091SGLV
xLISZf2pTJt6uWlVGvdfG2v4y9RDxEZRUEAii6mnlwZ0goIntU6BQWLKd/KV5Wuj
VNkJP7H9bGxvbN0wsyUgH2cSC3kmPYy1ET99fxrwuuy8mUddMkDdzttD4BYhlwcX
sCRKW1AeePP3Oz+/6dlMtYZCFUbf71xap6cuMyvq4fNrfRx+DvvHZvFDJ+SimQUc
QnndmSV+WMNvrcYzPPhqmV0qxWDTgrenPQ3DDISZDq0PmgK4VFtSYyd/V1JDUF7V
VihwyEluClTLeq1RBJm8fos1ujh6InqXG0pBsLSofX+MyYZ9vznD61rvesvV9SzA
Jlq7kpPGozYyI2qk58UPyvOmlBX6VKRVFf4AYKT/mbUx5iB8Mmg+pW+dVHGEcDkd
G0lKu202zld5ZKr8btawU5fl/FFE19NIDHzNvKj3pKA57zeGReqQqNYGUglLTlb1
DUgEKcA1vApUdU+LWSATi5nZ8NUVN2k2UeMDslnAA2YXzp1wjaCWyZZv0/ek5+9w
fGtPsQJ+HuBWn2Z7dUM419A4rj1b3JHIWZ8xpTUOJeOr1BkQ/29IaSEOWvH7jFxi
p4J2u9SO0sctoQrgOJi/Zhb011uTFjTXYtb46ADNoyDvOVDH9GvRcLhAEEm5aCya
dmXgaryDSgULwkcil1x6FIhbl31+eRyK8nz45YZrlH3X5x9idyN4VZ49/IpM4icr
88CtD2H9Ha5W1AvQZhPyFq9hzN06yuDV+xIhRs8ixwsbqsznn393FT5ekcRo3Gss
OBSXR12HPTvU+gq41gQRi3L9vTtObfXSxZcGGq8WfKUdX9Jm6J/812PQb6jGdNvX
7ylA7clUZWVeuQQMV1fSBMOG1mAW8R0CIBbZJG4gridUSkJ38dwp4CSnkL8PedkR
XcGIxWDt9O3uYR6wruJdGrTieV1qbP5x2+c3qdmascdBeaH5vmHKZhWwl51Yd/Og
1zM5pVwCeHR1diefi+OjVKLOkgCYpv0L/g3X2xiyVKKGVENGiIUktEPJ+wTR6Fcs
v9rTOY82vwWjQwmVSKxojHkrMYztpnMTF6cbyJbx0hpPHupmvPKvGDknfLM38ImB
ycx5OZJRNiuumr9iFfn/SRwlsVJ1f6LOEM5PWpTXBw7CXWX3fqPj1bv0vEw9DZti
jT4h1jf7BNg6Bat4Xzl+z2dnPcsh3ZVSCvWY4rzic9YppJozLzcqZtKd/rlPxT9K
7O4H6Pg30umkuxpnil05lY+/nfsiYEsR2tz+Jgu04bjNf78PkxmP3VnIc/rgN3lL
iGEW2OEmZYtrAiULnOKD3ZaxhS4rC8FJEEkSswW66Tcyd27UNzwquMlI6cutv3BW
5hiHLVe5jEIl2CQ5PtEy3a6isffCm4C8pIBFbtmxjKOdA/jO14xLtVmIF7AP+K3t
BpvyWKfhnXBZz5xJCfwOqun525OTZ3qbpqbEd0/P6tnL/PIm7FjvGDtAF4rLjTCT
m53Ifmawte6mOQiq9oEQnVvcMXCPSTLkzc8bdQOzGZqgBr2cS6yt2VIN6+HB0Bk4
T4UrrW3JEV5ZyL0n7KpqEo1DAnlqHfEb4K/UA3i6Ae5MMLxibh5/N07FWiRlSxHy
JHiR7tt7cQioSPLA8NZo0WQQhmiPP7CamVEQqknau7kkaYxvL5tVDiw9GA9Jv6Up
JgGwnzH3lKrJHCyewtjZ37g3SXEWJxmDlfvIa5FDGIpkQJHbBQJGLkKvC0z8lJB1
JDC6E2Ah0pYXa57DZPHlvsmVcRikMxpVqbcrG6rd5YtWc1QvnVs0opte4oQmwwlm
e8oa2nDnD8GBolr2Ja3zGzZvsqHr8Mb/sPqORuNHBz22Z+u/IgXEGoCkKLQPy3OI
R7P2006FkN65MA5+WgCOqXssCbFYvnVh/S+fvsKYV00mxNmJE9mJdSFcVnnrcM9b
grSvxwcQFSEH5fI7s4a8wZHnw6WzQAX7tQVhnvTUF3nc5h27crExZXyzTHx/kKY9
dYUAeZZFZkTGrd205dPLmOZ/sQkbmTJCtBe0j0+I4tW2Yxd3ddqqTjWrx12eklet
aIS3pjoDnhu0XcE8HyRMrA8bHZr8IdPp7gaE50haGzhkV+CT935CMHN3jX6tqQc7
WvtUzftsQ8KYM8Yo3z3IKu6+7zNi1BsUTuV9Qtj1ZjMXst6h5kK8yL3Uipo5J7C/
NrHk7j1Smnb9Ok9lolxnmKvb6CsUpy3hkiRI+sO2YMdhCL/lbA5yGC6jJOcC/P2y
chkju3i9VZ2lumoBCg4v2g==
--pragma protect end_data_block
--pragma protect digest_block
hOnr9ggRfZZ5GIAI7XB4eY8Z3pE=
--pragma protect end_digest_block
--pragma protect end_protected
