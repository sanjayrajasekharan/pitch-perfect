-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
cwCTMOUjW5NuXzGFrFQN/Ijaw1/ljX1ZUztpMn24rfAzbYpMj/IccCrNvPiOBRIE
7Iv3tV05d1bCK5gcCy310lcqQ0PBwfL8g0F/tTzjwlrMNRySS5u28LIJp7BmmD0J
NuQh5SgsWQEoytaFPjQCat0CzWwHNaDbtPFtU1afOAU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6080)
`protect data_block
Tu/9iOOvtRz4Wxt5ItTuO0GPJRpRMKULD5hl+AvETsTAzbAOcbsbfooKlKU9sRCw
Yw5jZOIcwgzMP6aMSihofH1JR4Qs4OEq+0MdtnGSH0agoeE/npAg4gl/g7YhIh0Q
kc/v45swptA+yoLZUkEPgC7ZWH9IZo/qe4VUcVTUYcc+YQanEDKSWho5tWLUikDS
XvUMDFgatKJSPySGN1JmegNuoVoWK6BI/l48NVr5pkGs/i3m3eNGRlsdxAM5sKFN
G7NNph0cZSD4RbXbrBinENXmrbj+5zq5BevYfi+iJ/n9UUFN+gX6Mcu0+WROoyhQ
ipUTfEZNM9MIoG9obU/FyKG66/DtMPI3Aa5DAI1rZLGbiH+gdI+Qad1732m8PCr1
99pGfAgQ2aMgjJcT9nxH18pBaxRyTP5Y9M4Tsah3KcmTN4dDe49G/fcX7MlyoNAR
M35euQLhHv3pShUKbwY6kpZg8TuNe9sV1tef/m0z8L2+N6qMCsyrjKwJPnjZaeqq
Kdy3NWA0qW9OMpKOelk5QqdVs79kVMhsez3X9aggMrt0UcJ97ggo8ZK0faIJxt1g
eligtwqIsQMPEiGq0ogZrbNsmZYOun+PGTEjMqkFfOMgWHSdyJFh2vCNlaVJwS88
aSN6Y3jKXhfCSZjOCAUmUABlye1ZUHuV+Sahmas/Ob8Wa8bp8yeLy/QupVh9ujh2
MCh7CmD4y1Nj+0fc2pdkOFeJmM/Ph2DqsijQ7K/8Yyx+sF5tluo76AWI1baVOgFq
CyT43j0VBQMnI0tvpyKYLhddOpAb9UE84J1f1feVCyus/LKdqNKTD+kSHisfdCYY
amQOMeM7xmvYnLvXZPKglYPLzqAODuuwdR2iLWBr1FMSYgcNCHW04Azh4/6FKw71
gNg35SgNBpyDYGnWCE8w50YzZvmyjB01KhjwjZRwCusrLzChFYrIcS8NX+wM604p
gCIEl8mAQTydwtGUkAO4VSWdjST4MSmS3vpPilTrAE3r3hKek7xBTBkJCVFdU+d+
QghXPpFsQ97sktG6DMYLuV7suMxkd/HjaalXx7ddmSX6LckNoxKnA1UQZwMnCEh4
JF7T0td81/gG9Q5mI6AroAIh3ABmZF1inyfhM4y2JptdtRGmKAw5XcLqchfFTZPK
5Ia3+eDXmJmP9XEvVrzgkIZTBXk+RgLz+EuCUso4Atxqhc+aocdRY8++OY1h9GV9
JdEEehAgHU4tybJHaIR5c5PFZNqlpGOBFTna/6QFEmGiR7hODSjzZCwNQHYsaxKi
KzoGOf0CHdRs+Daqb6la4H8gJ1Ol+aVeo/r47+2pQSCaSgPjatgFnvYrmHR/NX6t
wUbiKoyyr5MnHQig12O1dpQM+jJ+DeO7ucqj7rDhm1fgsC/gCbNdQB6udr6Gm8QB
v0bhEyp2uzOAIJrVNg8fXcJvnKpt1raeaXz0e3+sM6vcQ7Rtu2wda7G0G5I5axv1
OAmgxNNRSOSJcdSVPt4nOwFU8Xk/ZL7aKMk3no5bn9hMHb1p89eVUVRQhCWWEG+v
Y/6dttlT5B3pQnVCl+dEIc2m06cqSULIgvHugIc/gueCoT498wWeJ3tySMLoI3zc
Fyjz4grR6D2CeBBiiecuM3HVymCwgHuHdCNqTF6SsM+vCZHqz22d1oCmtSqfY2yC
cHTuj4zNiP7g07uPrIrnDJl1/boX/k2krPYg7uoTh2+JkCPuTlVovRtt+QX1oMNl
vyHqQtuju7JxoaKxr8ywLdcxRi7MqrqGsaZ6+oHC6cnIvFTQwyCZ70WNm6wkEz8S
09Nct7vgLqlwSJZOa8Gq2QqXBZStQY0p+SlOfojcBHa+1EynR9CYMqT0HURvWT0C
zumyYykko+TGTzmd3qH4QcxHiZkC0ajS/JFaRNvoBQGWyBXG7DREnz8+YVp55kE9
+R+S2FP0tw/uPo2Ji5a/vQ2OeDvWQbfC028vBMfXaKJrf3/XzXg3D7Mrjw12IFu0
HcaA2rUfpzKG04VAEcqIuQM5FMOD4wLEsKo3vXiEPe0TTtBBX1S6D29/mhVWIy23
eos1eNPo9Dk4E/ijlsuVn0U4alIO1Xk5PMsibDh+54Vmux/p6Ohp//uSUgVIjXFb
Cf1xHxjOZkhskH6Yqw2K9H9kStS/cCtxmKQbZnqgjznmqZyd3ectxSKzxCWteUzc
7p/v56o/4nqnK/6L+CCIxlJZQH7gC1trXZrdzV0doEfWVrnEk/QXXqd2LAoRFy9y
KuDJ2+hdEX+kNoVj550Od3L0fwD15KXSfowk2419+JzzsXo6xl6ZGkVgRXG7HVoI
9IfuJdnbEXSMdzs8TexRIDJLy31CatUg8K5V35aTtD6PNbhk74cVN3AzepB0YnkR
TmloMKv8seEPSk1ZCZH5kmWzsCWNwfq8qXszQ214RRP5ebUZw3Hzdk1kYdrceFwt
sAOSTjmVZW9Zn44NVtlk3v001pndbRg+U+wfuGP5WhRaziSzLzNNtjo+xYGTDT90
WrJYboc1JGnzjUm9wIK+cghYmG+8y8AjqxG+Nj4f0Wfrm4MQFDSBASa2A+S2wdcY
rZnbY4Tcr52DlWY2sKj4dd9PEWew/r1lhDY+wNUDksQZIHXlynLhQlWMZ8EYoO0y
4d7VlLgOmOJ9MM7jZPBGuZAfFKfQWeOpzfxv/TSfkrBiFg9xuug84Ja++Wi72Of9
dkdj9E3m1Y2H8JQMMDmdGCeTYvyb2w321u9th1+IuaQJxPdaf0fNYvC5PAR52h1T
R+/G9Uk4rRy6Y8TrTaUUX9KaFSiDzUl282dOFaaWa4g2oDLBAnu6ir+7ZuiSW2nf
7bWkqu4Gj63xxvrDR8UcxHTR8SNe+tcN5zXTz4ZUJkb9DLh7lRHkE/A0y/WtSbqL
vytNsq9cMvOiZYYW+sE3OCpnCEJc840jdJvLE5reddmd+YsgjFMMMsiQ1N3hu2tI
pW1LzfCWoU8IKdfdDVtMnFBJm310/Bq66+9REx4K91UZdrOSGDuX3ZTkx2J0JAnn
KOL0w+YzBlmiSoo4B7PEJeEPCUy+i8iLbDbjfpVzywgsp0K2mAZvm/4TWEnxZiVJ
td3GS8Umu8Z++SV6AkLKzI8LiRQm8ELgktV1E911v8DPvfR9OOpfa9xUmWk3C8mP
hP4sGywHkVBPQz7ONi1T/tDY0W4TgR9p7acOUc2hnNlEfRuzwBczuKJ5xiunuuRC
apVl0NN9cirO0YtQcKyHpj7ItOpc8AWRXIQ1QaKA2G7vOmM9VWl0n+E1k4Xv28jN
hqT3nxAL0cyci2rn7oToitjk3/cZEZNBExg4xFairn9eEwlrakftOtrbbnL02EhQ
pOrbAJn0Ow+pKNmOwfPyIYWWe8nx30QsYkuCDV40f3K/BxmLHUJa/a21zyrZcLWx
jsazOQHi4NePpqLamDpYcUtdh1Td/Kq0AypfgGxm1O/T9nHO8PhP6unzxwlJ2t5v
8ges3SR0Ou+9bmhu7+k++gnbtuBnSg1JOTJOJLrdxz7hxpx4vf7t3xxGuk9PchjG
jOm0ol5rklroCrU/hCqSMvy64Uy36MCF2srWkK4+EoLBIp92vRrXUGMdYGL2GOcq
1NdVpplhAwOWPCYKsBcuAlRcDsr5wXDwh+hjl984pJuAoY9mrHLl1Gch37rupU8V
qjyiUFAkMf3mfAYkoVE8SaKAKXkBLQpkNZJbSPdOiYuUlrPs0v0vYvgtbx8Y1/mm
x9O737RsAX6jzUW7nGNNnU3rL1fTkH7X4q9RMGQKXPl2KfAZuugbwR2A5ylnesOW
aI3J4OrXJtCPwz2VnZeQEAzgw/rLOsVGtv+YtPDgNR4aqfmVb3B70ZZh8kqXHrna
wEQKMqb0L/9NYayb2DZAPkDmbr2nmwNsBA1Ct7RFGaO4J1LMvJNM2LuPiXb2/RKy
evhfQmywC6Yw3Ua2jqsNN7DFGeETxAYdIE0927keIMzEFYLq0EtFE3myoHLvl/fz
00Xi5e4n21Rp7PE6mSzv+AyXz5G/OkhUZYcRnRh9c4CnTsMXLdBZ+bWvAi9bKGUU
r+MjbOC4s/mvrmG54QHx1eQkAav5DgpSwT8nYSbLhPrbDEsvWXjoKFiO2YFdsyPV
M08p5DWuBamItwjWRHvL2NxYyrNkfm7BnVb7ZKGYENhyYEvAFqWmJFW7qETZAAUq
ElUFa0vgj+HugQyVFUqE0Nbt4EhI1lQi18q78X0b/A4yV2E1Im/M/TVlLZ5lCBxg
zJiw6gpFVD0rOA6m8/NKkp9vNK1FVKuA0mILZq/t+OakJTRo6dtReNi4RNkaA/Gb
aEY3ncSryOO1rg/ByX2zpHjCNesxouEs3GE9fgjjjd3+L6y5NEVIuE8D/CUlIYxd
iNapltXX/xLblXQfs6/wcIHMQfDtB8ED6uLJUdTgtJlX24VMmgwGWcaTO6r0kure
5PKVFVnWqb4y9PAR7BFoQG8k4pORl9pb/uiNqradQmi56Lh/KCGtU6N02ngNc1FQ
RJHnX9qLmnH+czkRPbArX/6KW3qwNQPHkB22rat37hiRuo7lxehvv+9YB1jSBUg3
RQxrHXJZApgr5w6+do7/aGGiTn9qcz40FtuY44CEyzlT6nySZOEwtnLjNVVTHsxm
NGvgcHUw7Kvz+z0hJ/+XoyaAz4rNuFz/hwwMJjN/zYbTSFxxrzFWwKs4V+dI2BdC
IdJy0KWjAmE81NqV5aBK0RUnKMDGUS6Qo0/Bmm+EwNwsM8KeSi2YHJV5IapOTWi7
32rlyaBofhs0FiGtsEux9l17my4ctlnoCBQ7m/hEN4Lg9QM8qizlF0zVAgk2/IOm
8cVBGjKU68MB+5Ftirpl5qFjEURCW6tCZSnbdc5dXOvPsSF+0Qib6wbzKfSMGDJ2
iNaQAFvUjhlG4CrvmiGRUV8UqbqFow/s7I5PvnbVWCrMtv/Dd6K+bxWFWReeYY4n
7k0NivWTkvWAqaZkvaltAFL0VByB/rTa8ld12SdW/nQRCwfOoRktXx5r//Nf4JEi
Jb1MdLDXQdxYtzyEhjlT7epQMhH9r+77mKFNMS5khag9IrztsU4s+xWlR9QATmZ7
TIbWrBVCXnRVQK1rbO+ayGFH6zpOQDWw+lrbdwhL5xtz0MuJ2cQvq/TD+iNaX/Kg
7g29+5UNhbNnmddYQQTHQ3KSTAWVRoaCSZIW6tymZ4EU1i4Dt5KkoIg6lNV9Ven0
gqEt0zmUL2d3fqInR2gZJ7ZACHDIYJknqgjCKPc90q5MfC4MEnF8kNfH9LLou3SH
/VqKIkROap45+cZ27REsC2ewLnDhqaUrGu/CAu72Z0eqJX0uDA+RpD8RU271wm+t
nWhgr/BW3nT7O8KrTXrvsxVjkW6dxwkNSVLCGLkt5ZqO6+9sargGJx9B+y90HlNG
tFpMlEff7Nd/S2DC+ZVnl54DEEfJM3FcfzyNrYjejXgYZ1quORbZgKwIpBoSswHy
zkv07zZ1QInldA0VhGzOprK3gmQ+eNhk9OdCfwZ67ojehh3+bq5eG7mt5iXsQY6O
k6GBk9HyScQQZoCSNtlxSnmwG2v1KpZ6fK1TpSCA1dbd6eQ0DFVEphxQsX0fWD2P
LdixLnbmgg0k3Hx/xctdhntSLWym3vb3k5GrrAQa/az4CmUxnUOWMHW3sv/vuKqb
TuJ/gvH5/U7K6vEJtRwXbW3MmYR4jkhnyt0xtSNf7b1TEbR1Qe6Oso5Wb6iRAONA
A85An6iN/lMcjcUyUCvuCeSZG+/jyr4qcUXJ1smCYUid/vNP+o2O0xvOUFJ93+nw
C4hi5KccSqTt8y9FGCqRyH34c6Dl0TDKXxUxcefIv3QIqQbi7or+yJ+RNL4LrDMS
ph+pQtcVOFpKYZinSAc60kTb42hiS3fPvCsDm3rrymvaaewEyDxMP5n7TYZMoSKP
0XMpSTLcNPgDRYJchaDIIw6XiN9kRo6AGs/n780OWXepwmPdvSOMzFliu49QyDCl
6YQq5rhU8mcDMVShc+msdlHVlcBAlfTTh8gOZgkmJh4OFoljs7nOk+iADuYmBA1m
3m7m6/X3owKK8idJlq+ghCFg8FZaRDj62/v6zQeUzAlFBNQ9/yjdn7ccJDy97z4i
S5hK5byM6PBo00/CZHJd5BTmPYUyNVytRQi7AwF4UND6CWuZOycVezCZhFyRJsyl
68IR9vwf2kDafXDbbaGMcMQOE3Ev9O3JcBPyLwOUiRuNK43ZX6vQYWetqI70fbaF
DJ3L6GIuVB9QAC+yvT3nu0S20muDufdy1Q1YoNCQg63+jbWlQzodtAOToyz2eDTu
Ia8Ib17ExczDhroa9JVngEqUE4/LxKtYqVeZOVCCocREfvksAlXLsUK2cZVHNBHU
IZpquj0GjSnjBKE8/P0LY7xJxl4/ceHY95pbpyO0o6rpLl26VWx/f5Rxj0Jt9BR5
Xdj8NQkQqUSkDURwYBJsJe1OtGGzuQRNbJHCtHDRoeWTODqMwizDgsnlWcl7PlQW
34r5Z8859iatae84aOfzlbaNJj2XshvVmghHmgPER9p7drB9r0NrdywZlb0XW3mC
50muzJfal4XDIPSHrFQyz4AdUM1VuMhNZF2F9Mijur+9kJ6G78w6cb+vP2wrY0ut
fYaC7YhdF/Q5IXgHPM0B7kGq9fiKcrYjGFFJyueSLl3/ZaDE3AzUsOjCJlJEiACk
onbnu8JprJ4z6YEM7AHW/fxOuY0NGcxTTceLTO7XUzmZiVLK+IJCn50TaEnSMol0
Wgsq1HaX9tcj1crcMFQYwxHG2cY2O6xVD0ApVe6QH/At5H4SSl6zfpLtFCcmILdE
stA8bOCu0zQgdfMclCWBzNTqy7Pr533L6ZkMVoCvK+l16PA22Mg79snc8U3fi65y
AhOsXq2jlBHpALFCmRo4yttII9qNz1Om8ZKmN+HwIu2dnGQUkDnzBwAWRMHROuUG
V40nKGBbCxiLLaMmZWyU+POj51REQ8ljvbN3TI2r5lAcYN63r6UNja52sO/SCwkv
dORF0iudkp0FzwQ9IYma2vwtxE0taIdcTDeIeHsB9IGOVNiJ0Xf4UeHeCvX2eXF1
tXHE9RNewVg4gGiE6nWQV3UDgU3v0oDPtusFrBxWENzEaI29UF1IK/fP04JMzBmG
JS4ajJ+/YJc+cZK5xFqiGRty2aMpygXVK1YoeuMdzZ+gpk9nAS3rtArLimCfRqDo
U7jCM+LVdvpyiTAD/riAMiHTPqoM48Zd1UuhAlYPoSbIgVKldDrsHj00wSxhIr4a
JvI2a6qtNt9cKq4dNbIg2NBl1tf1n38k0ycjoO3UkB6KHNhBtsmrWrrbcGDl0Prk
WB714hwNZ4n/s/JZU7h6ZbC2Q7IxAcq3rg9lHOnCv4lY3XX5dmZCy/u7JbJpiu2v
AlbTFd1PVZt698qoyWUa8FizadYt28PY6bKCStLb+qcL/OpzIUznAgWELSqUbEd2
aYkLkxuH7u5P3rBIFAM7HOW9eZOX37w9qvgILOtfJiXJjGfPZ3kO3CjU4bk7/PaP
+RIwd8eZ+CQMurdaAz8kpC11k4+Jfk2APGQ3qjteOlFrqlQNwbF50SNlN2tn0Tnq
qM9QDyVPiOHmBPsZvYYXo2NloursRNzTVAoRo2k2nLqCkltrlv/on+II8r5NEfDN
PH6KaSvmXu0QLj8m9aLFdrvm5Qbq6DCXXx8pWJND+ouBy7wmQAJw3L9rb72UNHzg
VZ2S7+1VBfSLdKiFxZ9yLNCU2sRhw0EgKlPvvlZ9MORWmP6cbOIRafDEChYBdlSG
Q9St01GNtX2hFadl5+idY+XZaxV22r4v8YUv2vtArEV8nwtgWSn6tbQ2Fym0WpWX
zB32Oq6m1jF3WPfUAXsf1mbuGESt/02w+FjcNp95xkyH7BwfgNngwcEBWzelYMBU
iAXA7LUqhLuYhv7DH6Yf8qT38y5/3fcizye7qTPj7FWQAQm2iiZzsuHsDPP1j9yf
VFbOQMA/9MK6f0nC5yFbS2y3rzlrxdZXXBfjE25HYOIOF3ab5ashddhTIN3iX7P9
1Omyin33JfBUhGJTbQn+KpH1j34IR+jUzw2R6PFyC/z0a7CpUNLv6L/tpKC9yvsr
/uJR/Plf4UOysL5fu8y7CVJ2194KyaaBWHtZ6fElm6M=
`protect end_protected
