��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki�N�z�-���̦ܙ�C4�'8<�%��u�z�T�/���K)��u������_@�<����6����Hfq��e�/ s ��s��L�����7�ܨF�]�V��Ϣ��gT��$�d��uO_{]� �Q#�����m�l,�f�J4�P!�== ���p~������
������Nl -�k��Ѥ�j3\@0���,�{Aڽ<krZ���l�e�m(��(0�4�>9�\(^+��GC��N������?���`��� � B~���c�?,6+VO1J�>vNjG{���˵jF��A��k�N���p�,W�N�Ր�/��Ũ�y����*�����,�L?\���m�68��F�!�&�c;�ҏs���3���r|�8^��4{ۀ�$h��4ӋK0��Џ`��8�hH킩�� ��f��>l*%� �M�Y�\1���IC��C$� ����xMqb�W�g�е��θM.�����C�������<|����N��s�m�̑���1]6|��h
��>���>;�.G0����:��&��Ǡ-kc�_��`B{1	����9I�`"�#��cӳ�P�ُ�'�S��vsؒ����n�J��Pr���'�W��4/1�x�|0M���y��E|�J%Q���^�r,�4Z.��lf����`�B��_B��i��l⣕*o��J�=�����~,�!+���/4!�a��ӓo���OYO�r!�	�]��(�=���%��3�M�Q�o\IOָ��I���\3J�2��=�H����x�{$�F7�t�g��<ކ����
;�b�c���K����(�:�Ө�'�ѕ����ϙ�sT����9S��,�W��T,M����"�m�I45C�6�����
Q(<F��̯���Q�B��x���s�
<��'U��F�4�>�D"�3�S8Q*��*0�g��;ILT�:<6x���#:��� ����;���L]�(��I0���8��&{��quPݞbt�L��E��>E�:o(���r%4R�1p��G�cc���p�� 6$�8>d���l�3�:���Fx�(C`����+|�4�*|L���//�^ve4��_Ǒj�VM�"Ra�u	�P�ʧ�Y���nl;Ň�[)Q�|���l�V���k�N�m��R������%]��Fu¿��)�U�]���%�+Ro�$�5�G�C��j�+B���m���k���g��Z	�$��@��+\y�Q���t�/
>��$	!?�|/�2��S�J��L��I'dE��T3��_�B��}�˩�!z���WCD��
/��d�-��-wd�b��Y�~����i��2e�x3��u9o#1~��!�z��l��9����^~��oX�C���.ց�N�$`�%΃��C��?g�/B�Q����c��-u��mۥ�0����l�	 ^�cj��=���Vj�ܼ<��N8 ��OI1��	b��t����Jw�P��x�Z���9���H%L[0��u�/1)hO����*e:uUό㕫'�e���eYK�G�;w��_@Y�|O�At1Dۘ�����.�r��lU熵U�'ܨ�lC���F���^�5�/��+���{�锽��e)U|�R��}��W[�5�����ejx�>��������f��ڛ����ie���xdS�F�xwŏ`��,t��hl�2o�9QʬN}(_��#1�:��<>NQ���n7�օ�V���J �mI2� \����yL�������+�P�h!��W2/œLZQbX���<�c�"C�kB�|��W�j���\j� y35�,��!���Q���g,���f�u_aA0��x�\CB{�E��MB�M��xP�O��AR��.,�͏�iV�Ko�)Te�d���/���b���� ��?N*,�H���!��4�guz{����P�HBM
�G:ז�tu����`�4k�8PI������H�
CxO9�Q<�S&U>'^<�vZ֭޺37l�"0�羬�F	V�%E��g��_v�\ �׆�@��Z�ϴ�������L�Ɩ.��TkWN�r幽p5,���}�����Vޔ��@�ߪ���ɕ˔�%v�G�`M�3�k�����%1C0���E>g�����9����GpȢ8��sZ�K���=��Ȉ�5��U����[c��B��"�M;i!jd����d�N���N�..�9�{ם�	����	I���>��M���?��5]_�~�y��y���>ɑ�;>jAf�>�7�)�؊��x	�2�k��'�#X�;�ޯe�Y ���]y ����n��
���sS���L�F��7D�{G#��3�~+�C��QK�g��%etV�bn�{UIhm��;:���(��-fvCj�[����~����H�m���`���Ȃ�^\4K�XQ!�����YI�b����l�.�g�h����_~��n��rF����Z�O0��$��r��� /Qz�|ީ��~V+�@[I>rT�=���Ue�x��!��5�A�c��Xw��#��A�����e*�(Hj��x��ӫ\i�E/�%�;:۬��6(�H�6 PXz���ۋ�_��=�}~����c�����Bt�Yq�]��ԭd뫄��W$�e��4(���t�c������#U�d��{��'���s�@���jQa����0��Y#��HdO��d9�����wf�ld�)�Z�.���t<E�y6%#���nc΄��m��%�n�D"4�9"g��|�M���%���k��k�`��Nث��8�:&#�K;�ݹTP�
}�lp$��;���Z:�pҰՙ��
�h0�3ڪ}�z����~C�q�YE ��Z&�N��¦f3G�緀�ҧ�.>���s�rm�_�X�m�N-�#�:�'�8�YC�Q��|�&R3v��V�y1�Z?LH���DE(S�4�������{��yI�~��[d�-s�W�:�{��@���n�gߣ ./���)���h䧌:�WgGǋԴ�x��$��*�h���R���}�ma
��<�s�U�o1)���OV�y�-,�6��]
�=y�IZKۖ�ZQ�Am0Sҁ�H���)	��Z�K��;8A�$M���1A:	u��n�~���3�G_�+n("ə�)_`j��*�h<� G8XY����E���W!�*�'���Y���$��I?M	�.	O���*i�	
�#'�Qq�5���
ٵ�����lH�,�F�Mgo޿O�3����#B<b�6�d}H�iq��Oː��[/B0����k{C�<��฽��ɠ��C������9u��֧9b@1�j���%l���
�_�g�$��^y�=TNB�M���|{���0���l;zlX��=~�_a#���	�Dnn�<��;C*�*]k�`g��iF�[��&@�q��`(M��ϑҾ��z\�@��]��V��+:@?��Y�]��\6�3GӮ����u������d�o*'n9N�c ��n��6�W����d��+�d�n����n=�A�����W3�M�D��{P���4���Y�>A���4x>˾&F��;�y����&��;C�擹�sV��N�RQxNz2r1�cՉ�$��T�������zh=����1|;{���g�D��2p��nn\��m�O5!@b�gSo�mhk�D�"��$�wT*�j�/���o�c|���>�<2�S���)Cw0������I�sZ���F2�MvaE�.YE�5����m%��j��X�È=�k۫D���*7k_sѶN�U0���t�ng��f��5?�#U�=$�N�ʣ�[�kP����>���C��z	�q�m$��1�K��.������&����j������49h5>D�\�KB�{���*�j��A�+$��b�M+�X�Ъ�bD��浟"M�G�4�a������b��D!36i�0Dn�a!�����i�˰��{1��F�����-�J�Hp�0'�fbH�p�|�#�����6�v,Th�9�Tn/�q��;~��4e�����w0_Qb��ȳE<���'�y��Pr��̘�Uڻ����&����5$&qbƔ"�(�0r�p��Ց��]�c���S��{�TډΎ�:�w�h0ş��ŭ�����f����^+蟚��f��,f̬H����`՛���6�A���lY�LT�yK��?~{�C����E�s�58��\�-��!��¯������9s�~ s���6��T�k�r�al:�r~U󨥷⩆MdԈ����]�s�F$��@�v�.����IT:�^�s
�M���p�\�D�b�}��"�$�Tt����^_�Y���ǐ=��\,�T���V�VIv���v�7���驧����U���ԫՅ�Qsw岩]�t�i��7I���`�o�[hO*9jܡZ«��u�q�z��[��+��m0�FK�7B��DFD~��������
j�䴆!c���h�9�k�S��hr�(����ꚤ�+�0���0�p��r�YM�|_䈹M�ZM�@`�"��:;�YQ;�Gv���rt�s;�(�
kv���ʘ��d��e�#d�j���5��y�U��,Qlvȫ5G� ���a��:�<VT0�_�p[��!Þ^�K7/'{J�
,�H8�i�����j����I ��؂��O��J� <2D�j	�>D،�F��U�a����A?���aW�p�ȥԽ�M�5��*������Ɗ��`[�k=��}�U�}���U��]v���\+zq<��
w�)Ake�8@��G@& �4�������9c��PV9Ȁ6�kXV�EĬ#'c��/�3�5с��KP�ސ�a"61򇧽�����l}��Řs��'-��&ɫ�W���e&Q��
�1�)K<3����	��Z���F��ŕ
�����m�����ՏY��ye�I��jb[�`#�~2�з��a<��&�`�,OV���~�����#��3�6W��<2N�*T�g�mC��/�j\H~@c!kX�y,Os��=��R��PAp݆�sޟ��~y�S(��1�F�~������j��*S���cj��Ɲ�!�,�0ë�q�" ���
���)=)g��E�$L�n��b?2������� 2�����A�����NT�w�dIh��Jk�"�k��S��yd�޾�ɼ�ň����:�;������y�2Rx�>u��O%��	����#(%����jW0��&IRIq%S����X5�JXؾA��P�����D�� x�h[���@��UdY+v#�xL4�J+ބYƺ0��r"tO�~,�y�ې5�q�;�g�m�ߪ�lP��g#�ӻ}��1���k�����(w�O�W��?*���m��Loʿ�~|3�_K����o55vBc���A3l���(�|7)�
T�?@,��F6����a�ϚJ\I5�Ս�!�P�հ��g�Vu����Շ2Th�����uQ��)U}]�֣�p�K���8$g�qR~y�*=\���1�H[Q���4<l����R7�^\
� |� �N̏L|-��
� �F$���`��k,�5�Iݔ�oC�W�g�R��i�s�hĳ��O�^ľ���1���;�&G�{��Ă��æU<�uqT�)��)�X|�	�ՙ:C�2�ἅa�Q(Х��PF"��Xq8!F��?("&����E�_[�����lʯ�������ͽUW!#	>T�e���!�62�������r])��q�Q���x4�J;�����&M������6?vQN�إB��F��&�=G��)$?%Rfj�Q��8g��&=� ��D�S�"��ѥv��K�v+�Qi�Q7UdF�V�J�Ť��3��=�pQ+��x�Z��us�{�r��-�U�^7S#�,Ͻ��ɘ<��Á�`e�v-_+�I���8���8)w��?�ޜ�TPu`����,2��H8�t=l7㜔R�_t�Mgt�
0wT���$s��O!��Z������``Zc��� k�⹴VA %�`�;�7]wC�!�+Q4PxgS�yw!�V���r!b�ހ,�|��}���bNx���'gT�����1O���i���c�}�(�o�9'\�:��$-��'���A ����@K]P�~9c������r12y��I#L�5����>��R��"��yEGt9։� ��U��
>h���V�cf	��b34x�'��.�Y�rk��*/���F���X��I�DB���������ՌJ�z$7���N�O��C�GI-�0ٶ�c��#Y`c&���8'��!�@C�C:��@n���'�lJޗi�@��C��Մ
��pw9��M�$ԐZ����y�c�=^����R��H���y��1�/�zΒ2����=�yx�N�_ �O1�`��	�u��;g*?��bB*㉽^K?'cwju��!$Ձ9Ļ�k��87~���.�����fl�  ���]Ck���Y���1�[��/��Qd<�d�E���)J�{��}8�n-@M����!����u�`P�5K�T��ͷ5�$� _$�E�=�ty���	�  ��PG�(V�-%Ҹ�O��U�l"���F�����=3"��Q�AL�x�'�	�P�b��0���4���;������y��[�����eC{v���3s��b�~��_4�F�I���yI������p�Q㌈�U�^���CkAY&ǝ���J��y G�T�tܖA�{��cχ�T)9W|P�&��c�����H#�Qר�B�?J�cf�e��y�]MW�&B
鎞����C�k%����>J�g���h�P��r)���T=4�Od�|$qu�$�0�f�s�)�}�73Ң�ư���|?�#�J4�g}�LPh�Q�d�)�g�6v�5�WV��m�����{罋�R�V���$�>�0i>{d�i��2iSE�����a��k.h�naX������g��� �h)�ٌ��_�	�ܚ�o�RQ�抒��9�gdM��+���o���m�)j$���x�z��i{ Rz�q�ĺ@�%��H���4w�=N`�Ė��t�RB`5J	E�e:'��&Mc��(��;�խ'�#nHM�FkF":�w�vH��Ƅ��+Bg�4���i��mY�:��}�=s�Ԁۜ������V<�Ͽ|��лEA�H�v��P�w���h068�S��D�;��v�p��Mڻq[nc�Re�c�|E�;'}��DsT��۷�s\�Q�@U�:��VUu��[:Sh`�OL�;���I��}��R�%����M��Y�To�#��������v�nM�.�X��恺h���;Z~�I��i�c��}����T�P���ʅ�~�"�_$��L�'��'�5��� P�E��"�a�J�.^��(X��?�C�Ti(ɮ9��UV�T�̬�����;���ɛH�͵��i��>++X���pڔ�K�nS[�1@K�"bJg��wu'��͕m��?�w<1�[1���'���]���e��䊿Xԑ�%��w�Y�M㩽���b//z�?���=q;,�\�Q\#vdA,�g���/=�l��}ұpS@ަ)�(B���y�S��<3�G��ض-�"�]p�����n{��a�gNVTJ�jո�Ǔ��:u����%�8����'et�����4&k��ԡ L}�,�����s.MpT:PF�4|o����X�T�Ӱ��ӮfF��6r?�6��]6����̝��9p69j�JC8v˓Slܽ+s�֒�����������B����cz{,��Y�a.�?b��z�(=��*�
�n�8O�
�
Oj��quX����!�!)�tCt��цX� �b��F���&b������)U�7LU�_�I�d&xC�R��r�R���1M�	� ����d�7]��_"��h�)<�9��:Ґ,~B�٩ު(�J��E�U��b 1�T!��{��`�TՊV���7���?�^Q�y��[�(-���m3�=����%�:��tl�}@SA��%W�e���GY=w��ɥ�>v){��}`4
����P�/�q���:q����}���\���b諉��}u��Da��a	�Gצ�J"����abUa���S?��O��>������>j����-���`�p_�d|��U�T�x�x8S0�&M�I3�H���ΖE���'1��ԥ
�����H���������[е���~\p"�+dT�iQ�������C�T�^6��^O�P��:�	�z�d��7xT�PO=
��|����fC5w���Q��u�����9vn��$�ր�j�[�GϦ
�>���0>X�s*� ��{!{~ıx$��?���Pq}oj��=�Zr��_X�����Ɯ?�g#I!+�n�C�X�c7}��YqbW���CR�p �u�D͗�!+Ӆ���0���Lӽx7�?����U�+�\&BF�,�::0� ���n�q/�m���w;�9Y<!uq�!Bf���P��HR{��i���-y�/�@��!�qۧ����_�ƪwK�0�DU{j��m�R�Nb�N�
q����]��&����E�y�mN)���2��	#d�V�Kx�~�=�Sb��pDJ�Q��9��7��R�ev����%���_G���{az��$�E�M�:��e$�"#��
�K�	��m�:��HQU�@Z.����k��pId)��eZ|�\޽��a�a�H���o�5l~W��,�ï>��V:��\�qn0�_.�ߦؚ���wx20���#s<Y�����Z���g�}��[Kur����L@4Z��BWԅ&D?s��ڻ:<�Π�er���a��7�L�X	P�����?��(�Ent]]�}�-����9�l����J�~��HsK��D~��Ԅ9��a����@� ��ފ�J1 ^��$$̈́�g�� �Ζ�R��*�E���]D� ��c�1����A�\�%^֛)�e�3�'F���D�4pXP��3����	�&*:Z�~{���(���سr.�t���|���ӈLn%���+M �>ֻ���Q˸ �6x�Z���RbU�ֲ
'�E�6i��Xz��&P��6��p���3,����"5˝X�꿜�Cܦ�߼���9��)�ǰ)$ �C��`��-�0H���#х�5�v�Y���N��Z[Y����X�ȕ�%ݘ�iaq�L}���R���D�o<��a2F��2���d�jj^h�O$v��������
]Eƹh"�M���+,p��{D$��aaW$1N|��X�a�{T�ϴ���wPvYD@g(::�A,��D���U�r��r��FX%�W����ԓ�H]�d��Vu8q�,0��Ů��8����yD7\���B����CN�O{ic*s(��\��8)W7H:Q���GN�e8UzP}?!C�t�<i���çU� ��Z `�^�TF~�7o(G�Z�m�PCB�%��W��v�bC7�bS%�,蹔%���l���_�M��L�>��Gz�'ڠ.e�������6�lL��^� ��h0B�)E2~o�k�H�:ʸ�*�8 /�����Tτn2����j�"f��,�{FU�a�X+�{���.J����W�p��9����$�Z!�u�i*-|gZEm�d����Y5��ܠ�i�z�Y�TiÔ�?]5 ~�+�XP�~%���V'7,�
��;`�Q�bI�t:N�r�,c,���J��ٲ�1�pC�D,�Vnit�I«�����_'2d�KE�p�ʙ�����k���	w7����{��fip�$̰pw2� ��/i���#jԒ����ց��:��#T����ח����>S��#	�:�e�;�X�ֵ��jV��o���v�����ܞ&�a��~=��2_�0����7��_k/e�)k?�3������5:(y4'g7�`1Y���"�U�LOWc:Q
<X�x�a��3��]�":�͢���ןw*[��Hfӳ'��� ܽ4��ׄ�`�����s�+>h�	��<���=g�4�FT,�	J��~UR��UP��o^����~a9��]8���wKnM�p[ ��F}�2�(,k�9xl��4��6��N=G6P
��'����q��޺��ů����t�t�/���3�,ȟ�?T�_�� Q̓�H!O��Z����(�J�H��6��V�P����2�yh��K�i����XA�q?W\�5���(�b��1��K�<o�q�Ie֏�Ҵ#-{}jK����~pVW�R���O4�y�QJ��`���>0�m.�]���t��?�<�����.3�t��8�kl�Y��9�[XJ�����5�C7��/5{�«lkNc���H�-Ƶ#%Y��.F�*��,��WV�oL����rI�U̼�w�y�S���d�\�n�@仄���%f�9B����֣���H�0���,�[��^(	���8�5!6�}��J��,+9G��-�1�&{���J��WS�3��y�C��%��_N^���0P�������o�\~: mm���f�2��G���#B�z'&V���7 }�%N��/�I蓾��V��
k(d�{�!�TY\�����b�*�Y�$W��G牺 �=7#%7|J0�cڐ�)i}��d����^CR�&��,��~]�ki��	���Ge� c��!��c\,:���Vo�����6�}�՛���+4�"��0�Xw��<Y6Y4u���JQ$��s�)⭊@�들�a���ǩ�����@8��a�o��:�Q��7�ǚ?W�Rw~��D}�:���w��{>�O9�#z��CPm+ˤ�a�h�S��'Y^���(�%�bG�M\jC�����$A��,Ҵ�S�+W�&ۄ�ۣ��bb�������du4E��p�c@���w��3T�m�c��B��i�������Y��<` ���v�`���E�`���T-��ƨ{��p���0z�\S�$��G��iEg�r�N �яB���[i��U�e�4�υ�1�r��M�]0a߯��5	vv�J��K��V�u�@{L�T�PNz�5��u��l�M�g\�?�'��nQ��I/���� U��������z�E��As�e}*j9ՙsƘ�������3KCaַ��L�J�p@���P�颼�k��̠�)��XifҨ���}�#s�;��l��M�(Sm��3E����F����+����O�t�H�G�+5Ԍ��iB8^����>%�M��^t��@R_D.n!v�3N���C�v��� �rW��	�4���o����H�#o#K�<`��[��U���P�U$�n�3��r��� W)4��q���f���L��'`�"�^�� ���EN^"%�i��9����>�ޟ�hg��K��B��,U�9ܫ <L�d&�Y�����ޗZ?`���{,bC���	$��.5�=mZɬ��4Ŧ5���k6_����-�?/
~����}�wb?c�
��k.vA�ߘ�Wd�*�D�A��0~�BO�Z�k�Q'>�<%å�?�cD`~F)��\h�U��4�~!�� v*+|c�6<O7 :�4��L�3��������ފ�8�+������q'��Q�W�h����@�ǂ�5�m�k�R$r��~������U�Ad+쉑��D�f��1��5�M��p-<��7�jů���N!g4G��FbF,L�rMg�ĝOaSd�l�3�M��������������"�K]ZʠmԢ2��iUMn�=)#�D��$n��A���.�7�C�����ڃ�w�ǻ�����ꇻ�3�uh��a;�
SXay���/0|���~ ��0/ι��ݿ�f#�gz.�������U�!Lx ��C_n���ˉo��,�E�gBF���$!ƙ��z�[-�N7�]*˙A��|��"~�:q��//XB�`9ml=|M�����;���c���I�Ė����Gl��adD���kD�b�m�5\�?�D�e9�}A�n����J�F|����PA̡� �l�D*x����â5FP�7H1�p~��7:�t|�B#˕}I3���kd�����ܹkn	U�a�ں���{�+�2%��Y5���<?l��>�	cԌc����"��Z�p{���?�'� ���q�e���V�k���\��>���G�������V(蓝Y��C#�li�������ym������գ�~,��w!q��ӱ�$�=�L7�D��tj'i��E���d�kM|$���=8��<���`lA��)6�=|F�P�ו���n��"!�w�չ���2ٚ0��<�1
�� :=�T�`X���h^gּ+���ʟnV `D8V��y�ȁ�I��Y���E�$�g��dJ����5�	�{�LB�WA�G�q�n�Өe%_$w��{��o���k����ȱ"���?9�|%�u�"��]{�J���_ݑv�o�����i[��}0�P�,\=�XfӇ�Oz�A_��1Kw�4�2y奁�*=���߳>-+R��k��AN�q�L�k�VI SL�y��{�2�[Wޅ�$��a�1�%ϼV��:g���p�Cv�f7�|EP��@!�3l�ueX]ێ�w�7�o�����4�1�SLp����C����B �ٻ������H�Qu@�/0�3�E3�� j<�L��I�FQ����$^����}��f`�<����M_�A�q�]R��59����F�&%k�c6v���������#��+c���ն�	\�n���������*�Z�,�oi��~WW �蠰
��O6��C��Mbq�!Z^���|�����0T��87kuˎٗ��wѡLP�I�A
5����o}S��i���� ��.;x�b\0��uĎ�3�;�
�8l���/^�s�B͍u�Vj��vvvM�9�)"ˑ�o�h������Y��iH��_�I}��7&|c 7\�'M�g��c��Ȝ���cA�/-��'��!���nl�T�K� Ρ]�m^x�D�ē����X�o�����u����;�'�)�ė$�vQ��޿$��&��j˗�C5[2�C`�$E}���]������{�����������/v��e�D�S։4�o�I��&"&`ƺ2 �S��<u3���]3���2�Q��t'��LX.R�u�L4�s�2{ԥ.�8�95ș �
6{%zV�M�73�y7��9p���S��}�'Ŧ@D��7�	 �D�9������~�0�wC�_;\����&~(�ͤf�d2��%E���_����?I	��m��ٕ����d	Dz_������y���%��o�{�' bA���S5zO50��u<���qW�e�!�B�x�.S~��[k�(XjA�����1����;��La�nw+������"D�HZ���k���:z���:-t��!���Ӆ���5��t��/ɳP"��v�q��(+ŕ��Wt�i�T#6�i��Y:A�k�h���s2��#3�
���Itc�eDӉ�銙L,q}���q�T�CN�M{8�Nk�yX���^G�V����T�#D�4��e����@��}=W��%��w���LDg6�v��� k4z�������t!͗";4�TY4|%\�1̀�?ل�@w�Kl�(yPfYW\�R�R�;v�u�}�;�afx�����k��w�j;�=lB���C���m�z��-���~
�h���*=g��@ڳ�؅h7�H�w#lU?Ǧ>���L$�;SO�ƈ��q8�[-��T��g�b�z��KS���AJZf������9���><,�Er
�L�@�����6�*�
g+����{��������ST_4�D���阢,v�R��D;XK�_�\������A�z�����jRl�}&iVq	Weq�P��1d�����j3�ᵃ
����v"����~�:��8}D�e��}3�Y�̸q��L�6:[���#�f��m��o�pgT:��`P���F��_�'^1�,Я��\);ƍJB�5���d�́�,��s��HXf����g�w�"��:���&���+�xJ]�pk��
�{|L�Ӗ!���a*���w��S��p*�;R=5/8��&�cp�_�Y�s�r�Qī�<SA?S}a�`��(dh��P�����]����(m�m[^���C�����樺��_��� �f��)�X��R>Y�w;k4#!)�~PY������	�x �f��GAy�)����Jc���@�a�.��C�4XD��q��ʛ�ث�W	6�����!���(Bc���-#��L/��d� �?ŉ����*�T\��>Bp�Q80�N��A�����-s��h7|NUt_��Bm���r9�UbuU���i(1WsZm��:�-����`�et]����/�p ��h�6cq+?��T��:nf�Reh`�fݴ/�/��شʘ��L���i���h�p�����hhF�����Ě�%Db~���E� �N�Ĳ+����z��s{��'���2 �������m��z"��gsj4�
ۓ����+�0cj��.����~�	�t��K�=+$n�5�������]2�iFDҐ(�i��Ĺز��ۇ��#Đ�?z�w:{�ȭ%�r��4g4�!�/!����[6�$�[5�ʹ)7��:�
�(ʧO ��� "�v.η0���d-����� (�x�"bОzԷ\;�.-i�(tQ�����<��o'��!��/X�����c�΄��MZ�S,��~��`0R�Q?Y[(�֐��C�-�-A"M� 5�'�b�f��dh
�-&4ڊ����$�v��:�/[�Սʫ�!	��f�YV�1Qa��̠�D�C1�0����y��}xN�DFR�OQIsF?����J����伫f;��*2�â�]���UD3ֳ-��P��lDh⤿���=8���x])�;sf)B�#�)�_�V���o������+F��0����ys2�ɬ:����-U�^'_��8ۯk9���a^Ht�0�p*�3o葲�L}J`A�)�1Y�9޴j*Ac�د�P�,k�1����oqI��"~�=�B�Ih�v�Q���LD~���P ����������0���`,�z�xޱh+G߆�i�a���7켛t�Z�>���x�o0�o<��LAC��w��ߨ��Z�E�ԍ��и!��j(%	W�ǝ�-V�� �v�c�&0k�??4�D�3�(1��ZЬ�7A��n�j~��������L�,`�reЯIp6֐��랕[��{M��t����\�?nw��&�TޢQ�[*�6��K���.W6�8ŀ�߀����E�n!w˭�r�u-�w��)��V��V�L[�AJ���/j�e����߈�^P^���O��;`�jLc"iRK�2/��C2K�oҭ�	4�@i	�v;B.,�:� ��،b�x�ҟ����$��kۄB�IB?���:��'���YGf�b����Q9�:�|���8O��@�:��Ǎv����^d�[�"NJ��_*�c���J�Y�9��!N�?�c��7�B��^�?+\P�l{���w�a �6R9�����z�j�E�~'3��#����>�r�r�2W}����^04E7��������"����e+���߀��t��Z�8���f$���`mC'��#�؟]��U(ǀ����G��ɳ�Eic� 8,�H���54j���X����ݠGL�U�nS5_O0�
g��ʈnKf��S�ՕG���!�47	��9LR��aMo��{��k��l�����kx��v��1��r9��_��ǿ?���Ut%o�߹,��F���D�Ai��mYPc�l����D@�P8擴2?i��(��9�V�����Eg���4b�S)"�=�㻠�<��{�0{�<���O�C����[$6ŉ�9�j7_���$��[`cr�
MD2#^���O"A��AS@�5�)�V��r2�^��+3B][�C/N�ۢ�J.̣/�K�"�b٦`�/�5٤���՜g:Ƞ)U��)�'22��:�يo�x%�������]`]�cր��d�\BT�l���ri��!����[�t�0�^.�6�E�X�����Mh��绲���@5�D	�J����%rg|H騬�)����M���x����E�I1��H�f?���deOu�������ɂ����݂eyXF����a�Ő�\3��𥰘�s��f�{� �D\^v��7ה�7	ߝ1tq.~��E ����w�a
1cX��(�)'���|�O�0��s坮ț=3����N�h/�Q��R��{ƕ��۸A������
/ E��ba�s���f��>���,	C�R��/�*��;Ȳ���Tg���>u�N�(~�_��E�;ϒ��O*<�]���5j̔W|��PO���"W���?$tm�pk�bQ��D�I�i�1��N���t(����-A��lu��4� F�������6EY����[M%Y�ס0G��|�O��I��7��B؄���#���E3� gc�� =��+p͙����#�ͥ�T,��'�GÝW�ۏq>��Ⱦ#�T�G�� ��߹K,{ �P:pr�{�tR��&2�6T�EK��zXg �a�hut4I\�&)�?�� �qoߊz?C�tHTan��\3r�����qF����`�q=}(۟�$�@�Afr�o<��f!��p�y&7�4�Yf���p; �*�?w�Y�X���i� �|��x߫��	�t�WVLj�NS@]Oa7����6(�����db1[�����V��.�����$+<[��S�ځhN�����;��W�<~0��J���M�G�ڶ���Y<�������T*�RI�T�q$��]�0�xˇ�ii/ӎ�AB��&E�|�� y�7�n���goF�:�����;3� ��$���d0v�?OZ3@Z8�1����)�lӚ>Z<}U2�!˅#l�V�؃7�Sdv<k��D�f�F�*'8{��Q�s7�|��'F�%`�ţ��:��C3��5�c�^|�È�b��6D1�Q�AB	O�Ľ��T�vS��N���a���b�C����bn���� �A��O��-Vf�-`��i�5�c�ya�4!?���*�@Ӣ��И]�����ض�3W̻�۾����8!X E�����A��x��r�#��?� g��̓��u�dQ(���T�`
��26�fݦ~����5�� ��{2ҍSE51+��y���ߨ�76����8�:�!�
T��j����>B_k_	��]��z����Ϧԉ��x�I���*h����"0��}�NQ&ܩP��\��9c��"��`��V^h����`b� �$�]1�.���j���'��j�E����~� �?�<g�t�>�E��]��C�N�WuZ��1CEFl0�Р��j���?���9��/�B�k�b��NOv�"�401�aT׏�j���x�Û�����9��n��g��5&��@���&���64+�1�c��j"DC��Wku��:���#"D!Ӻ���$z����i�1�� ��>m��iߛ쨋�`u׬]�+�wu��&���Pr����>�a-���I-4�g����N3A3�췙W��H@7+�.R����r �-�Z���ur�!����|i�p�iyƩKi�!ϕx�t<����/$��
ũn@A�j)�z��I��E��׼��9��1�ƕ�l#��� ���7�1�|r+�S�=�/�
��$7�h���3�K�� �HZ���������҃�S^�ÈK��G�{��Q�t5�p�z}�$�\�_>Ux咂,{TJ�Ay�["�x��܂��B�/u�3=��ɥ#��-[V R���Np�&8����*�U�^�mhy���-�w|���׷�~���eGn|�=�-׾��Q<QK���d�����
�����r�o�pG]�k�Y�������!����G\���އAYϿH߬;�rI�4�lH�J1- �SmAQV���~yw��~C������"����u�&�8�o���nJ���0�Β08��K5o��J���O�]7��K�4�����2g�����LQH���(����V�d%W�V�^AT��T �H5�I��һ��-[@/����)���w���0m����_c���g��� �y~�SS����CG���l� ��� (bv�P��"����6�u?>EB��M`�#0���aj������6*�hk��	�����!OA�g�Tg%�I?��"1��q�3�����(E��57{:�����0h&Ҹ�.�Qv)��h.��0)�+���j�Y�������\�Z7����G���<�vN	Z�qӾ�F�%:���&}�����N�}g�H��2b�(���.,c��z �t�'�+p|cm_@=�(Go١7�"[�D�B�tj3Ѧ�x���-~�Z2��(���EҲ���s���'}M3A�lsSn�xz�Z�����D����W@Yz�n��n�˪�рc4J��mU�4�{�֐�1�^�r���^����̆="
,/��U?�9ڢH5�VVY
�ᮨDB+�Qz���y�`�y��?=_h,�Ь)c�D�~U�����L���V�S܆�-mnZ�TZ�2�5�`�؅���d4i_B 3��I�,�7w�]&Jˊ��!P�]0�٪C!J�t���	w5��,�]:��j��Y��؞q0϶2M+�}\����{�R��2w�I=��zi^dz_�y�]p_��z8��R�s����|< ;�baf�� � �Acfw0��	-���ȀL�����,�f|LTف븯�\�A-�F����4���s��M{bl�4hd�O$�Q�
+u���FJ��w�U��YuMiA�aBf��q�M�ޕPH�l���7�V:����y�I�`��l��	�=�U|B;݁�!�(p�P],D2���!��T$���������e}N��X�y��nk��̣FLd�G��+���Ğ*(�A�蛿�k�*RdK�p�k4|�We�{�<PЛSk�\5׺(��dצ(K�R�[P����_�G��[%a��`�N�b�;bf�TT(���zD�4˃	����3?��0�{��6��4b��O�~O&s��8[#˼>��cQ�`V�+�R��[�0�������V|��&u��x���3ٲ�ٓA���M'N�xa�5�>I��lpH��o9��(AGK=P �db(���䵿����JC�9��>>a%���!=p��v��)患���U!7�$���Vև��NY���#9P�h�0��K���ci�zN��<��8YH`T/�Y�H�{w�}��C���Pa�X����*Y�.g��Vl���/����µ�w�fb4�7]C۵G�c��WYS�f=7=��8��⏩'�Kf�"c�?X9�/)^���^�b�a��'�!ˠ�f�@Q��rz���H?7_�x%�ϟu��ϳ�� �A�!'�u��E�k'�"�/�Dq?���铚5U�+��}s���=i�[���J���-�	���rN��@����o;i�uaO}��,J2�&���i�4�_�p^�z��d��<~��P(�+IWe�T��0��=�:�M��#U�WU�n��w�y�Ұ�~��n|����?ݦ�/����	_�p6�&i�x ������gD
�wFa�&�c>�G���Z�9�mz�wBZ�;�B��y'�xEde�����Մ�э�P�1��精cH��SD���B$���_�fa1y����Wᒵ�g+�]V3�F]'J�!{cq�Ϡ!)��m'�$�w�C��/�ܴ:��=W!���T?!K*tU4#	�O]�^���L "�_l�l�z��]D�����^!#�EW-z�>q���/�0s�R�_[*<� '�T�m���'k�_s� f����qP�o��-��P��d �3a$���2K#��#Km��m1u�_���w�����_�f��`E�`�|T���| �����D���No*��C�c�?U�O������׿I��[��I�hy�r�Qq�BX\�°���yO��Y�1&o�v�du�y@)"#Eipl2<P&���ћ��聅�6�/ͣ��)3'w� �V�k�Q���J���I��V�O�X�V�؁Q���O�l`����C.h���+g �E۲/�p8�jl�qd�A �X����0|�6�([���SR���`�K��_�K8n�U0g����I��"`v*����cn}�i��hQ�\�ގܧE����Tt�6kY��A�G9j�� O-6k�{U*��&q*g�~{���۟��7ﴔ7H�9�h �IՔ����a��Guk�{eS�����!��,��~��ԝ�(5G!����h����x_�����]z�l�����ڄRN����!);P�a{�R�w�����Pť�?("hQ.�6{eW#����W�ʪ�1;8�2Ͽ2����cJ�t ��y\���,\-�g�E҇�Q��1��&�S��ʿGm��ڐx+c����!S���ǒt.��p�B��=�^�g�BJu�V��(�q�ev��?!�ډ�{=i� &?R�K�khDD��q-,�-ԗ�@F�O=!�\�s���&�ź�)���*P���H�R<~n�b�;���)�c8̛t̕v���%܋���K4�y�+Ô��4��M�Qv�_T�5߲�`��:tC���!�����Qb��e�y���7c�
��$�W�`��+G�N��Y�8�ϐ�W�ɰ��x�/��E��l����q��K���\��+��1N�Qe����8Ǳ�OZGL�Ni�T�������E�\Ge�o��,.t���&�ߌ#��`���Ճu����3e���L��@�~Qf	B=�.�|l���E,s�XO�
���@p7#>�72�&/����݊r��p��MN�G�M{8�3����-Q�AR�?bӊ�rר����o0	H?�a��y�m�uPP�*=�dì�'w�B��ȃ�[�Q�[��gNt�o8\��i1GK�j�*�U�%�- `nH抲^�L�Oy-rػ��� Q��,�Il�S�b_�0����Ǝn�ʉ�/��s���9����yȶ�6W��gN�db������u���U]���n�0c�ģ,\�ؕA9��Z�N�w|���d�@ӞOL�e�[���T�����3���nG`$��"� �U�a`+;�	4LA܂��DLYf����'����q�9�F-N �`���B�",:[#�6�.�t�SQ�f��_��~����e�&^>���B��uE�R
�<6����c�"�<B;��ed�ۜK�~ͺ���*݊� �ϭ��W���k����%�XB�MJ��w�C�%M@�QrD6�G[_"�uȳ���4dd�pna��P��*���K��e�C�����y��Y����*Z�ڙwYx�����a�E�0��:�V@����w���UBlE���ݑ�+��ֽ?�߭�Q</��1��(��۬W�x�}�مf?�Am�e����,��çf���av��W�oP5���cꙠz�%g��7M��0��]��1�&�(g��i�@��"��ƚ-n��ܙ2���8�`{8��;�&�8Є/����J��c�
|6���^)R��J��a\SڥU�.Y�7ﲁ�d ؃z(s��2C%��X7�|�)`�L���s¢���|df�,�xG9��
�w���C��T�x#l�0��i9��7�e�d��JueԼ��l��t�S~�R��6ȠG̵?ůV	*j{�^�y�O5�l���G��v���#q�;2�E��E�JM���)��8�4l�0�!#���m(8{�����֙�(�Y��u:�0v,=��{n��麥��T��D��D�y	K���; ���Ɉ砉Sl*l�Q��_����-_p�f.�?�x=LN~	�rU/������>����Dr�=�$��Qp���tꭚ���
�O��¡6��s��lB��e��%l-���%d�J�N
��������P+�23/=�H�Z�t��p'�B����ԃ��~&%�N��wD��ǂq-FjĬ�(ƭwKQr" �S��A�y���W��Uh����"��}��Q����㙅��uJ����笤%������6�7q�ȢE@TV�I{�$InD�v�j�����/���f�b�%�B��gݷ���OɶѸZ,�99<lq8�����_��ה̓51hE &����z����%Y�6�з�M�8EI���qp�T�7}c����cIyO[۷㿖�*�p��:$��#�E_�탳	��c7$��u����a�U��W�[���7��UIOje�P��	A��SL`��$\���C��v���SIŴ����(o�Z�1M]xj[Z.�f1���Lx���7"�	��� a��>\s���n�֫�\N��v�"?��G��]����8�ʗt[���$|�Dr�q���c��a����^ǰ/�������e�d�-L�B��_=󖡦wk������ cve6��Ĉ^4�����V���	�/XA|S�|�i��wnú&��}2Pꖔ�%{��_%8�7s�[Q��~1͆���g�� ,�P�~�3g�q��=�t��鰁׺?���K���������-G�+�Fn�ۆ����Ω����