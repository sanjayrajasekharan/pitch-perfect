-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QJIDENv0ihFkPDTmssQBkxjS6VwUfC6SbPR1L/EgMzV6hm5dCmgID1yQyOCm+bNM
f4FM0TP/NOe8+DRmJVy72IIjEK2T17bNkGb76YYdD9ahlgK6IZ8taAyzHg1uSN/C
MNedfrqz8JJpLFOBtM0/A6obMOmeR9JJ1aFi4PX6xqY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8003)

`protect DATA_BLOCK
ZrzZUAKVb/PNnh2ExzyUtGwYZlZMXAG0GxUEH1hU8au8nT+GmqbIXLaaCz70+IJH
ED7lbvNd+267gOKETxWrA0b+dM002nzu5ieqJBIPU2+I9uP1tGy8EnVolS/XAMOB
f6pDQGgt/4gSf/dv4mE6Ml5OhiuRBt947w6sDVHZ+deAMzLyVj7m1nQ8FV+0rghW
VIXigdEXojvyfzFvGoLtP1DI9itBBEQkH77a/r8DPC31xeSKPLG4POEIC4vjes4O
DpJSjgD84Rg6TTvbf0fL4Tbr8FENd3Nz/3zvzzonif7cm29n4UkjZ4/jEjCR/wSk
LCXf+0EiE2mtVSY03Q/g3IS5rvn/tQoOVLmElmxnNrZZJUVJclWq3ySeEKOoPOov
GHct5hqddykieqMrMrjXo6qDj5gc8JRWm62OtvwmAJ4KX8vtFkAuAdhyl+HyD1RY
g55IwH1XMPlbo54k1NYGua4LCPNNLts7jXDyvJPQdEqKV0l65b9dbqy9Ps85sFJP
30TGJE0sklUfdVOGUEHeaRUCqeTyPeW3ujJkMbThCDDzP35c9bvehO0FLhV8+dXX
qjAM2QzI0vtg1v23jrWHWk1ut6MLH68DJMr6mL8g0UcdChXMVhOc8IwqdkNuKw4O
iuaICGZEA0VIZLJgZz1AzCTP2aDusAbDvQvrvSLzCy7Ibcy41E/+025sRac3GSCM
R124NmI4gzSnmpgjMiQX4parL37f70mifRzt0WHycp6F7JOcntyXYwsh8oCb/3ol
r9ZF2vbR8Glszi4FCyjbVzGgR+EzLb1Ea5fMlq3k7IT34Tje2i/eFc8Gi2AkP/+M
p7WXgGGlZasu31FgKqRGN+kGC7yENPIkZmFFiMjAnrn2Zk6lGe8XcFY+IGjwHaTF
lQ6AFZ+WF1ZS5j1uXYZ7BVx1KurxLEjzYm+THdfh0PYUzPARTtSR3JlIhVG8Ktmp
0sjH2GfIR0w8DwoEJGLQ9BOAoMCSfzKyyP271I/O6rxs0QXqhg5ylXDt+50yQWeV
xoBdV58N3tfPpcRWI2MdAjOpNuDnJG9BNnJMv3kdO+Ff3QPDCPk/pUXO3Zn/gg2c
jZ4rprhJtx2xo5VxWz4hCCPq9sBBxM9vKSaqWvYARHF4J1nP0Ck7+SVco3afEUL2
4p65X+vymm/hu4D/71B7/S6CMOp3YlPX51q+yrtaPnksNvUtphND3Qdp+S5nSHo+
Y90IOYH4fsXX6VximHEQ7Yv8rGGVZ3SEMZ/luesgBslJ4OWRQOD7C2ysVr5jX1dJ
rXfw0y99zH0YQEUVnKJmXLIhYEUYft8MQOhaCq9JIbbC3ph60FKA+85AcffDknuM
6fJBwrjQjU4m3uDi3xk4yICQCwMH3t9JS3WIyx9sfZxhufEOzFlLQ4bBMY7zEk+9
uJPDtJQIdsod9NghiWVYx1mJwX94bb8yO/Oy5xzrrD15+Iu2JUYt/dnLjlezteuR
Y520+2VN4jw5UgTLWsQZsGgjlkd1+KMtkczGUqqcZkvzwnjUkxoma4yUd2+fhVid
NF0A990+PsO0I5SHx9g77XpVYIhdVItLaQD8IyRAJB0JDcb/FJZRhFGFUwaikhL8
f4vOwl8RUZp41N9aE60oaCV3eSxyR58dZR0of1Ssle4xgu5a5h8DkFdW3BOvbONP
xNeTjT+3IMCMt/CNwwLuJ2va0OuEWPog3tsETjcvF+skAAjtVxaTaqEIzu/m6UZd
S5Di4BWiIswDAlnIjSwdjk8DfNLKR7K5Qjq6D6ZUqOkfWu0Iu/yCwgBbrIu20ubl
42hCsl9jtKHSAGKkAmYhzPiHNTlEgieYCl1ITNWZWNPkEwOQ9S5YqZZuR6nxBzq9
yYbDKaAImOrvXL9qTSaKH1xTatMjXqZBjIkiBsMhCBlizhfFXY1RE3w6xWpW0Qtm
oX7bsHuMDuADmU2SyJr7VF4PylmuiDupJp0hkS5JHnW/KKT1PFgVe8ydH70H+dvN
GweFFjvczd0J8+QcDXNX1wDnv45s+8mhRTuJ4X8MppKWJ3S3qJ4GcXKZw9+EaQvA
vuWTe8hS/nebg+xWc7T5babJ6zQMLdsJNXugzNxNuQLVkqiIufRnnHGHA6y/M2fu
7VwyW8+3H3XwENAMVu+i8L23LUOu/s/RBELwtmgM7S+I+Iivb9ma/nEm0RUlKMwl
zMDZluiMbp1jMPNYZGgWkFepuldAHf8p6juXfWCjN8i76lacoQM3s/Gis8x9ozSx
9diVRi3wjmFVp/rxGC5CbOHiw5DSprtiBjyDW0zeS9Ct8beO7RgM7Nln7HQJes1k
H4WAi29QJqU7ZsNTW9iQGiwHxNFopDowHst5xa6A+WPYTJDRbt8UmfgohyISi4B4
u6pfGOyu96uRVmulWndS4RCRmo5ar6se6XVCqnwWJWCHSGvYHUnEmKq1a1aWvdup
TCL1zbok4wSUY9lARgsJ23WZYTRu0PnBabgEtACYmUYN8IlZnRazBeJ9gVw/m0tS
pNMqiwbW+ZmxwlvLRrlfrpCcmtbK/DmETk8iHkgKJjPwqsTNX/CRoLYneeTVw8gZ
TWbEFVMoK5b1nP8H4cmOK3uffmAmdNHxjpM7pMkv3QA/vv12QNjAogJ3c8XrOeJb
b60Va51bPum78NYuTIaoOqC8YzTI7vuzrn1MrHOQpL6FXkC+9W6iSwVEMMv3EB2Q
2+JMuVirm7He9dMPgGnM3c2PMvpmLq+hY6aEVfCWx1CKiP6m+0r4QNNdQ8Qt4cbt
lfu3gkF188u1okcuEJfJIskp7o7SDZWFTt1yRolUhcradozmqNK612vq7q8Jz1XI
iyNYJMC9eYNBk6r4bpQ5M0rp/mG6sumjAiTdeOCPNOWRHsuNe9AhK73czfthybIm
nz92Vj52UHMbV+AKmrnHlkp6kYv/kpIh6Hb6XxwEsPq36npGYORNHP/4AqiV/TNI
f9a80jhriX8WF6wnRs+JuG269gd+tRxUVLAcCYTdEy7cAeTpInBKy7hzOhuQ68cQ
QfPoShxMZk4C0j/przPdts9m2NAGCB0afraHt7Zc4uok0jVVFFy9Oduq8BIAoL65
FUGQ6UKIkiKoEDnUPMYBCR2gHebRHiRVeJcq8+FUIl3KAFUdD+FoJ4txe9zFcv0n
Fte/WM7Pli1OPMHYdX1tLdZL6DuSaIFJ+muMvnWXooPJ3LYTRk60Ea5+oDNQnwOo
o8sIO658sm7ph1sNSEqUcDuaTO4pUFWM8drZxTJ4UXey0AZpYaHZcA8StIYE+/pA
ovkHoC5jEVewCEbGXUMLNyrltoWCslt+IQw8Rd2ELEllY7SBnktk0EifVSLlX+a6
8tdnKcEv1gFJxlNyzodF4GqZ89C3izlbAhncJD+xkTEjnuQdURilRatLRM8tb4uk
BtwNDePt0luXdf6/lv8e2lFI93ygFadCrOwq/1Kd/8N9muYmjpauoV6RamblH35g
mGY4GpVlehktPJ/p0kjiu8mhdk1BBqJ5W+mXnmFADZD97H95jW5B/Sfh3cnc6G1L
UGVm2TX4/2fu5dnyLFYCo+P20SHVck4JaAC+IzKNImr6ohGrKM1YDg3liuzkpcA/
L5icR0BXVL7x1UCfcftZ5etLBlks0V4T3PC2+SHOHKQl7YM3rd+fQm08HFSRfOUp
uS78xa8WIyGMFJ9NPTS5DUItwKxSEkHwGIYhcIa43NiLYom9gaDrTKhR4daus97u
D/NkojqYbIzPqhbuADx+ZODYC15bNIg2th5bF+mhesF30pDYyu1phmXJST18JSmJ
jOGDodq8Dam9+8c/4Ng0D/+5t9ugnUZ6ZJ5dLdNfHM5JgSFby2rSuKDeEEupCNFH
Gd9HB19LdPRoCvS3wNf4P7yISAqVhFpDvYzvTJZadHtU7D64nMAhJDL717ImREv8
Pvjx2iJWwc1FiwGJab+sWq3mjWKnrsnP3yOmz4/UgHlB54nEkahEQUS5luGkAhkG
3USSfWH7i6dVNT8LYEzeZ8lahFwzmmglBriDvZl2K7scDidWLc7yi7ia+rvw06pC
Lo1oP38bVHWLYQ+u/35eFeCAlmM8y8b73D8sN4KSCmMl8/0rX9X9m8GrHPtcn52V
IbOgWWEDjfk3bZj8q6RMMYkWy98FC4tfEF66mM/YGXNO0O8h5s71z/U2D20vGlMK
CTy4hvmp1W5oWXE7HCZWOH+99Z9tKTaWoePbsTsodJ4M3umuI3lhcZJXFNEkY70h
dvl8OZhoGmrsT3sMZmm6YWOH/s7KkEeK6kobyr8n9xdGTITNKfduRTKUrckl1070
2NAvcGD0GNdSgS1sZsJgq22crG3cpnx9oc2ka0ptd3vC8IT+kkznXfEJUTQjIMow
Al6V0Enq64/2f9hWbDnDBSVm4V96Jo/AlVb765VT68QPdWDhEe8ZRnzY7HEENyrM
8mO3uBOZF/DEXE6xkqLooJoyp1d0UuDjX32D64wu/eK/Zkp9JmM2fq5oh455uX5+
pMefKnfsxWf4K9pXkzVH2XTqLggTqvNEx/PkIZOO4WsBqtbmBVMe4zZFafoY/cv9
YqIzJNjZX6cexOn9H1uRIEQ0Shbdq1ia413HpJSn192TF3eVU5Sg/l9vS+Trq1Jd
OraMVyiYwdSzf/VHrVmNmcWTh6efr/IMh3CjRAcNL4xEky/fuRxvcM8qxakS4OuJ
ix5E45MjEEE3RZsBX49QU7C5YRpiwcRPcaDwDHX2hCjiunhFRxW5jZSrmRBILCDY
s/V/OrPUtz0F4/EFXr4LtQrcI6y6V2n/pYH+iCmTapqtcAlLOKK0WIjS8ZwAfyMr
UpGaaLi7nFOBsrwxjX/quyL6NZD0lGyHIfgn9HHDzfK5KrxHpEENOCNz/CG3Wy7e
UJGta7GWf/YFCD/a6Cp/scukbnqIZ7wZpoO3PUG/OaoJTksEJ5+Xci3vZVUMIpxV
+XlhOLYoR6uBVPcdnHQ4iLJeovPGA/L3HOBYGacqkY6A+GntF11AXKyFhnBcu9Ss
w4ZYlHGhoFgL90Z1dT1R59tKzGhFc26qkLh7WyjC5bcKGSw99aK0c38PLGAYpBzu
ZCgs4C/ReqBmYf4prOyvvtkp2Pee4WU0VwVDrCp0MsqoyJU8rQ+w/UGbdxCbl2sl
66K/mVgdW5hMAD4btMQGvnDOFbAggFOADi5YkbjPt151tlEd4e5GEhDDzBX5BJw5
SoB+EFEmTkz/+5rXdRR9jG2yRy4c0ereKbFgF3duSZAm9v6PZiZuGnEm+ljYKY19
gpc8GJXDtodMQ0r9Jh0+u2ExKD/jivfjy28gTQNLBIfPB8SwGoEYkw8yVeZiN0eH
ygY0dKx+/JZSWXZb5QrQK1JM/TqLodhGv6U5A5YYKF74RTi0HovcEPoDiWYCXlqH
d9ceJMSToCSW1v+EIUKrJqZG+yOKNGA68E46qQ3cp+JEFi2AXSSgGmywhK62ovCd
QsIvzKTscqC0MHLoiZDIU9PMSc//jFVW79y/9yFOJJdpyXvPzjE5cGNYYUPfoYnh
+ZMdHWrMUD6lr7wdWQp//us4a+grCzA+TAIXNQR63XXohsOmPRtgGC1pd/P8NJgA
KYR4PACSopvdChThv2N4gCzt4n5Ci7Q6RGoilaUpNY6UPUsMqkkwolYq+WvcTbWE
pZ9IyMG7uP1zqTJ4DM8p0qjogpguj+otJU8feBFrPR9y7rA7t/vRBLAt32NC1WvZ
Tsg7LiO+VdtdRzj/kB5/XaAqCmZaYDhcAJpEepQLUQjvIfRw5VZn2Bgpex+1Z/OV
o3HxQgysZY/9+dP4V2DcgnxwMJz4LZjx1ZcyosRhhCa0R69c1afd3lskpkLc8Mse
Ik0kOF1dVPWjWGcvAntNjGqbTHYO2+LQgT274SUiUAnBOMlE1ZJ3TFltEkozDZU/
hHYodlx9ZzK7N3WqMVlE/162ORWHq1GFuek5Jw6OAqCmq3jZp5xY6XxGzhkC6/2F
XJvMUDeh/gKigPmDYUyDF6x1i+Jyz8Kfhya0pYMM67/SwW07byJCTMcb5O3C0niY
SE9dGyMeAXNNOXZ+Hnz9XSQZk3dAmas8heWIIxPPGmM7S4PHiyOjHQUkKgluAhov
zk+/7OOl+7Em7Ny8WU/NzU7o5dXulMA85DMnax0U8pDkvDrmdRDJ5LFwQOaD87Bf
n6dkH+8UPjabi71htUIk1Itc5KBqSahH2FoUmeP15ORmjUAFV5rFIe13ybODFQyQ
W6C5PllTeVkBnloplW4tsekgbHih20pOYLk01XCgf1+DHqRLm5LoRXS9jp62AWbY
+jExJ1oKgdnWTFq++m6rbDa0PSAMxhAmQ2YP1AoRXncX3Wu9MuycNbQ8E03WEiS8
wbF5HO1KLPl9ScmVuaFYmkVMiFleEwNTJMUbrWxx/92VhvTeU2BWF/k39KjbKSEZ
hC30d0r5ntC0LKPfrkH6Jn3iI2CTgpu+RmklVGeJTgI1c3DG+kWn3lJUOfaPaabP
IvlYRotK+/UO3T8olmiF7KqGJdHLW/28rFCmIRFYN//Tal93Wi48A8isUk4G9cJP
9re+7UTWR069JB/R17HtGdOTqcG5xA883E3r48h0P9o4Spw8kTCzlLNd2Gc6rD9i
Vtr0btpkhxGvue2ntQGKVLJX+U156m+sDyAHUwmmLMtzj3z6wAzp1l/gK6Svp+th
NGbGVU0CovBzX6jDYnXmtOWB9zSppsy9sW8kcKw+PyviTVDUpmVsbrtN0hGjqjVB
n3LZm5+L2eioxM2FQs9BRzPKulltT5HX+S0HpytQqcfgEnX0OlYmtZbzGk/Rnyju
UeHWgqZMxTWgKoz3DG8TG6whPWPlBs0uz5h8NyFScpCgmHpGWBoZTeTKjnzvFe1e
KYUQp3vRos9E9TohlRCao2c19gojBAeNU5wR34gNmtGic1OYwNmO2rdO3YTzMKIx
+tFzIoAFk4MImu3IWZqts/gaRouEsec4t8D5bozEhcT4JvPsgUg1ZWEeabnxxDNL
cMRfJt8OHNuzCBr7gSlkVBJORoGiDh+9x/tYrUkLJ+/7/fDURnW9NGfGTrIgMxRz
Hk2BizKYzF3pKvQdvpLV0eEFyT474CfJW0RUjo0fEMPuLP6IvWFuQzARTwEa58ii
mqVMKRzMkZ8/qDGQzYbp3WOnS4sfSMNUSydRaEkVsxytbktNKVn0KrYuJGI0IRYr
HhhsBOjGf9R9c5hVzoMsZ6pGyDMDODqxm2Y8zo5roCHM7yfwa4HcicgyZ14Zdqu/
HS1RdVi3gzjWuq6t0WSdyAc7dGXlM+Ra7qJN+sAbtzRt4rv9aw8etEFsnvHDZvjh
xldDaUkW8EOCekt6f9K8WSRBIp4nhfX+NhgBZUwZ7ifCXVoU07LCKTU6wmJBXQPq
2m+vbC6gyy/e2es601ZccoRz899dhb+vhUltDBLzDFdWBydA9z2cunRQF0LyiawK
Sd+Rc3x3ggsYP25QUrQWRx+qOqC+51QtaLbws/MBpJ8a88QWvoRL4iIY3buqeSn3
CNC63QZN0SaqE+hET/hPvDJZkhv1DEw4AAUXvRlooCPdLH4klo91laaLax9AjwwC
aElD82gzyVazHCx39NAgrXsi9sXD/+c4dxlkM422Up4Mw+Gk9n+Wg/ehqQK7Lz9f
ir6yFJ0WLRBfVI+vVSR6TqB5m6TFM2SAkKcgEsVHnBdI5b37tq0A2k6AFwFBKIxH
ou7COlJErOR0lFTDNS0XXaHmmLzt+F85qHVuBR5TU7EzuO+Aq1kDIdJspM/hQVev
xpa5bJBk8ktejRtCJuF6YDJhtV7kgNo6q52DH+GDpTdJN+rc1qxJqiqiQ7vjX1j8
NLY0gVk9MNgIvX3kszX7t7ij5VjlJRh7Yy+PID1NoRSARPbivbtp8IxaY6xzOU+4
eE4T1SYGzmNtYAQzJ2+BMcuzRCt/fSkaXszTYCfkjhQkPw/QC/x9RwYv3eDHqW0Y
gwFTA3HfChX62cQ6awMVkoWV8jsOgQk87w8PFuznsuUkZVL/dHwP8kDEhX71e64+
bpPQyEM36ZCS6Rrn16qRhXO72jl3z2gxwZ5Gg7VIRFI4chfD+W9+cKoOdtT5aLUW
iKLo6ooCEg2aaGSXLsry2CNhHOpdnz3hDfALQHmmmzphar+Ua6qUz8zvePX4A2gc
y5s8+urUHN7mKSoR46KmnxJDoarsiU8B8hQxoEK1uRVOARTIYf5L6UPutiRZTyJr
+Gqaal+d58rYWRGFjcQgDegUDA4rYthgSxqOIDoWFEkIbbrrpqiKVqhy1pLnPE0M
18UCIlbURKPJXc9OiMG6CM8OZ93KUCloOMEILFJvXG5qr7iXC1SpkZ8crdTmejS1
X+VpNFWKyiXASVUv8k26G6n6xj/XptzvSP0+1k6Ayv39wxPYrFNy70jWZu2WnE+O
eJeIQE2ht+01I1Z78tSg3mtMQN/ed7lpOch9nki2XYe+V0+psSMwXN/h93RE5lko
Wkf8xJMp9Jd+Bce2ZOp2mr4q1Kg0AiERreJXiVBV14lXAcTZyj2Bfv8RAVNpbl3Z
Tt4u1w6JF4hwIYqT5SePpsUJOWj4uFDld6b6UGKIeIrfG17r5PlE/ck0p0s2Nk9F
rZ7/7tv42eT+g4K5BrYC6h5b02qjwCcjm+E4QKrS42DxFPh+WJmehrsxrik8QgMg
Yd/fqGKYLvmCMP9RsjPWPABJJX1RvPVdQJNxlGNhLc7Su3UeSkWlR871Lw+61nGX
IMTFxtsiWFNIasxew/w1brw2fBz4EWn4AV030vQDgm1Qpw8nLqKBmPY6Xbs5IJnZ
XCu20s2IWthr7PJZQkV4NMb2CjE0o9kV7O2n3jFLyyv0lJKvmRP8JowQ/FnfceU3
gBx+PZFFwmBEoOoWM1U7STWrgYwyp7vB6ydX/qhQshjTC88EdmO7dIZsuPPQsoST
RHf02s8+CiHR2i0sfqlNDbOEpPghSwoxR7KoDkM5V4eehJ77puhgMF23qgPuNp48
JIUqNmlBZHIhQ2oZJZVDulhQ4OqKuRp5g/USAnLC3DI0vgyUmmCYLm4VblrEh014
tYiAEmQGa0/eBzktpmHNoiwpqvs+BS5UnGYLPtfZ+FfGx1pHus/eOrQE2ryjTz6R
kd2F1o7QJg2gcuCsFP0TlwkPBlQ+Gz7clqUilZ2aZy9tpUyVffomt7aa05Dag92a
O5sIXX22cPxNpjckLR/3FrP7xC/swTnebEXGFEJ4eVT30O047ZHxv4nyQBauaOax
gM0HS47zhzvOO4Fi+10J+aLtlwzIxhBHCkpLdUWJRMe5rk78T3GEVN9Es4+mfw7X
zrCmNyal8WPjCPNdpUbUWctKbjYON6YdqNMDN8XSvmTBmotWFIzcHk46CqFwEtCy
QLN5l/R5W6ziwmjjRTq1LfFTOyhe36FZag9zYCfrIWVc7Kd3EPCQ9tT/qMLVjGjS
sn9w+r2pp/z9pVuniMTnbm+4cNTXdJltyuraOY+zXO193Q3x66B6pKgAxit6cBRC
QouiaFQHz5Qnp42VR0WTEiSKCo7Scw+kYsYWzzM9GCqyQIMb8allbfsefI1cjNAc
oU5U8V5BwQBPV5eGLJgT7aSc4oBkCxHRSug3zmZS35uibEiOzDfbYhyfcZu/gZ25
SZVhEeeemAntRhk7EenyHPQFytDr+Ma6rJAPmg4XgKGH9RJGeUZ6M48+Hs2srym9
PZa2U0DDu6g76/Ze8125dAtbHbm1qTyyOj0E4WDJLUu2eT3kB/+ETcl9qOeMV8qI
scHUZPEanhAe0IE26R7+kZ5SfyXiubvDsMkWGeQpI2hmDvdadEmxHVbVJD6R/90x
LdfM3qn4JpsAw1kOohMI9dB82TaTUY8DtQPWT1/jINA7a2KaI9bHQXnm2Yxq/9+9
gvly4MBfm8LBvrELmIJYomipniofVxghIDgWWuRxXiv6gyp7j/d5th+kzl4qi9m6
sJpJq9ElxOYTxLam/O3+w4WsUqskr9XLye743S4Upj/G9ANQTSnqXQ1Xmk3A2XNF
i0cJD0p7CNu84if09n/1T0eSgWKWmlwOPA4+z/Zy7j8zJcmdx8QkuBDM7BThrjTg
FetIRlpXER1+SucASI/xCMB5FKJszR4ko3vHksV0hebMj05L3Ae7G3qKA9eCPidD
O+uJharDVdbCVSjvoVMB7M8iVh1HgbpYOSLXOpdcr6oE0CAp6U1/bp3HvzqJjX+W
BiMVqDhLKfVO9d+c8MqPWlb1Fodv5cooz0b/MOmFcJ6pECf1aT002i1hVtPSWP2p
rJSb827o26h+CXvX9BAQdNkRo4OEHSba1L1nIuw8UPnjbGxoOb1S1+majIzSHzLl
NWp6uuT5d4roFbU0ZukVaku+eywd2ZvKYCWHqcA47RGXFt4LqhNNljQt0LUEu8xZ
mud/oX+wSBRyzDNkW4L8ijEZSW/vBXDDtsVyYqi7jcMkT479AVGApfsgcHZDnMdG
o4RRBSj0YIjpy+xEbtAuoDYCmd7IlfKZqlM9tEIqKPgSUC5Zh6/OEr6PoO6LphwU
2PqWVUWSv3IGsTlm5/U1djY2KFIyE0BVPDQJ1NLJTLX69UE8dIDfLqJTlqyYIfPr
x7ZhQEUY7NTP5f1jy/z/mw/33MO6K1Sh5xfK7zlWHx8FM6tHuCa3Zy+I2oD6qiwK
iJVQRskLjQ1mINCwGc6OPn8lYtDqGKUoXyBJ/e8WqHISuvmZOhpOVOhhNBTLuzoT
pNBfJ2Me2xy9MJjUNVYrHQ==
`protect END_PROTECTED