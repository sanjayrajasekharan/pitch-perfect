-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
P+LM4HoQ9tALvgd2yHMg7ggknoGbnxr1ub93ITl3tZANbDrjFEd3swcaBJf57yzb
oe0JNhnAxKUl6u83YQckL2L/z345U63v13AQ3OtLsLt5nGZjYQvKAN31cp8+dJnQ
Ojc1oJSyvmmG9YNtEZ5+0G930SNgZ/hsV8fJSeZ7Pd52Xp1x8f4MXQ==
--pragma protect end_key_block
--pragma protect digest_block
xiivBonXfXiAFTkugX4OHRudCyo=
--pragma protect end_digest_block
--pragma protect data_block
+wMhx6pOpecY3bjkHvIGwPqu8WS+13L7swaG/EwxWTDxkx+olWg3f7piZzUDx4US
upKgtn6DwUwZTPwS+FEM89WbCQH05Pi/L0Df597silh7nlqIyyGFyxxVO3BbRY3/
Fbz0L2Nn0JuvChAFW7HHwnlxfUb722umiUGuO17sa/ls2nFBxVXUwCyuXU1ZPk/Y
zS9yUfo8LGsKNHL/EpvepTaZ5MhZLmd1qXxIcjOFV1jj8IVGscFTWpkydVw1FQkd
KRWInOEyq3FrVGjwmosjv8qSyam264JUA6OPbVpMHXZ6u3a62S1MjCS0vyyFWaoV
dAbSYkrC8IMcFA7+nvrZm6fdjwuBoDn77WHQ/EQmpiLuZvGTa09N+aT6S4xhyov4
UlIhTEf4GHgKJLHBMSAc6FgVORvkOdUckG4n8tc0O6nf152fnSmobI8tg2pbcgjx
p5zdl6lPJ8gg+wTq/ktW/6WZub0/G8DJsNfxAeAQDfrBKZhjJMvz+qOzxmAsO0LL
KrNcjvDmCkB8Xf0yboClKw96JqQe1t7UufYrktr6o0JgRObH5aQS9JF80fD2syKw
UoIe72Tu3NVPwdNBL0Xeehk8Ya+HkvUVY090fnW1yMri0bun/flbKFseqaUT4tzh
Q7D321OOPPjoLrXWL6EKeNoy2yM/KSKVXOiF7l0u+re1g6qs+60aedV91gjJPEC6
UikAiUfmxUwa4KmUwrHvWhiGmgfQs5hNIigB8DDMYV81VViauofQd12baZJQ8fSX
CDzglbA0h49Xy+wpN+T/t2847yvylK/kYTJACt0Lcwk/ZBAcbix1WmqsHtYtafY7
9uRpG/GkY+LTqAz12dqZ71yrPxe63/4UBFIhEBtcslarm8j6lhHwQMJLgYI2vjmw
AneRvDj8tjF6XwYXU9k/ig6yZhQjDD1/J7Tcpv2TBHEw8GLUBsVVcGMOuqDeNqeF
g0RSKxDDuC1aw/lekpBLNulAGal0L/376b27/Uf52sFoqDokpta8jDErjtmz/k04
ZAOK7on0E3yC7jVkR1X8+KjJPa8y80rljZ8V/sFZJEN8AsQFo42nielO4/72X14H
FwDTXzw6Bmu60f67QkjH+r0/g5fSAoq8vyary+Saw5tuxyl7S2UhOiasBA+zUjdh
MorIy6Z5pJrVaTa24e8Paz+CEfp9r6i4bTEkzfJDBwo86oJe6kbZMKkj6eHkyQR9
QG8oRApgHoY1n7SrDjOJrg8ZbSSXrOQete5DT+bxivaZmiFQaUTq2S80rKMxeu36
HVRoRumciUwGPuzAu8xBjQsX3ux5irQ6tgNTn5DmylD6YzcnCUB221Cj4AtROi4W
cQmENjUKPrZZ2sSUbc5+O4cDAU6DZ7xfzP4iM4OPA6SZlTQcE97mce6dWYheeB7x
aRGXKQ/8iKXZRD5Eo1syQh73Nv/AEWttFl0Idr0LYJCxue/4FPuIQPR1FhzXeUk3
HeQdeGgo+sLb3yjlhcDtJbVNRUHtCnCclq1TPmvdESSP9tr/CUch1Uq7XoU9HjjH
gGDYfPjolYAxDrcIwhjQZQsXjtwMxXHMW8axfWnUD4P41A4LgsVtVcY513285FAK
cwBixjTM641LdzQTesLf5ReO1nmj5MlFguRGsyxIFY3SRk+pUXXToXfvUNQOv1km
RsRRpg6ePev/MhfmUY53Skf+wB8cHNJ7i6bNO9vLyo25KE1OdKnCP6hsu3ZTul0u
HpPAp+XfytmuwukLpZ8rJD35JeUxb/I8zYoooo9+7xDaUSBYXkLaw5HiEnYbzLh8
vOJNcrAgFdXPOP3mtHlB0PjsBDoiNwprz134GJxIppMFebiv9i0UMebEuqKyL9rU
qFNsCJCzWEwD8M0QuUggnZWD9Mg8TYPfczgzoOQRhRf7754R9DVU16vuaNCExW6s
Zdg3SvgAKA8TpvAyhCGAYchdKsTZpUtu39sGGK0YsS5qM+ZE0w0R88QeVJtFAd8+
f1fOIHo7Smv763O/pNzZztGlhU9+oKjAhS2rtXQdVSJDYMw2Smw8SX9CkG/Cf3We
fexoCwTYzQOqYvgUICcXDBB6dO6c7Qi+HGaNDY+KF1aH75whLBShw6UfsPR08pkU
rDNbB0aL/ceojvVK/CbhL1PK8qnzb19bbnXhTsicKHnpOaS/MxDIvG/DXfF9XG0X
gysT0Deqyh21gGZ81gCoUEi5/7ea/yei5Gu5OTolunv+339E2njWgJdGCuqCXMNE
psi5yylvIVkysVWqFtqq9smEf3lEnmYcMMEw9wf/DmC/UYwI8xGQNi6O2kOXk8Md
gcnZjoEi+td8l4gFBxbpiPXatFl+hY2JGnMOz6lfJpbY5ij91JtjD+LZQL4Y5p1b
5IsXPeGYicegfw3sG+BgQzVmmtXsUxpAndhH1SGTLi/fTLrd0/niCmGOHxkNgGYF
F3vGxkyHsuXukfCmG2VBPvZqRegvUg0p/6R8T6ZqnKLbvq7HD5A/3asHIEo2LSg8
X6BxXA7P0ee/saBlyjhzhcxFLlvbP6L96Vc454D6PRbSGi0EVjZESuNjLvlMNtMe
B2c3Fi02hwx6YGhKxz0i9ivT17GsAQujCcTxXNbOhcvnGqqMpcHVTjZ8lQ+t+xyx
qE+9lDxkPV3Bb5PeJKYRivOP1qBzoxxxw0MvgiM3a4A4gClHFcV4rbCkVP9xc+kF
KphWubOeN256gUv/t0qyJ56ydUZHm1JR1WQwsfWj4sHHfCOE/r6pcMDFMmQLR3r2
UuQHMirD3+NHJX4C/12RWItMpgwItpS5g+SDc1gu8xpE4LUbbgK6C0cgaRbY+6Ym
e4Eftj8TfMP/6VYGSjd0zhvZhOxJLTl4ESXP6xuuSQWTfl6s5HzCFsLwWAlELFP4
74cnoaqjmD3HCu6k/asUIyd1rQuW8lOZhs2t3WkMoBwFZy7a0Qt3F6n/MfZXngYQ
i0eDF+TKVW/gyDbhDHCke9A1cI2a78Z5oWpv9r08QWxn47ErfjH1sf8j7n6sCbEO
+NxeDwyAj1UFjH+2d1KQK5qfe/IOqZGdnqGEciL6jSFRuWeNzBNpBwXF66DojMlM
fsLZPzDYSUgViEplemEXAPmKIPcDXzWqZ/BOa0yGnI7zTTxS28w6Rt3mop7pZoBN
KNzuZHlLI0xKPeYJseMLeGvFQqBOhVYxYPapgnthhLIHH67MuNG/f3jzN4XL8VmO
5qJ3mtHqZFdH8NmAd0NumvNnWr8JeZmj4yj94YAd8Ig7xI3a8mtWLxUpitdB9Oun
IH3FVqlTqKjm+7pBNn2Bu0pbVHbPmA2BQvGDzYjOxBXYYobkzeImbcWZU+lSc5Gh
V71bpEPolNETJK3A6DDISNyhprxMtQPkZXdCYxDPUTommND4tvzLjP+TObdB6iHr
+fsc9LGvNCDhwoPJC/h4twpXNauOepNHsecm09hEPTXxlF5PNGK8gMXXonEvUGQn
bjAlXM3Cu4Yv1FgkzH8DbjtSOeSKQjiZv4yA1T840DtEjsnsjGcqVW2rvhD3y3QH
zBHv3abvRX8MymqjZXQgBHTTsedQkq3ozDEsWESLZAPyypSKJKCGoFNB7bf4DJZK
ZWDxRbTEf3B//qHAeFYA3HULJwBDAbhErzyTrX6Oy0th1UUvSzpxmvnBntLTFUWz
ckDu9q2aDHm3IjupDLZgQ7YdSG1DWmMs5vhr720K4zZOq4qogBBBzVr/4JlaYYgy
mRG4QxgXGPej6uN1pAYBn5TfM2dUtMtGzY24xIaeEGLMwmCg4fCwE5jReBAWkGJk
F5sqdiHFTDS5zLq0NGsToN/TwC8Pk0hy1YfKO0RKmCtbyQMo2EeHa6MbBmt1mTY4
FoGwp+W+W0PXcuSDcW576u82xOrRKfnniklNNIDSWcMEy/dp4LpFoAGXLYBgg9UH
OrF+xCG1Mj1GrhRmSYJhHv+N3amDZ5OZr5C+oUF0zXWYfew0S+ZMdL/Vq7Ypr81v
Df4AiA8S0vZBfjVfPK9bJrHVaZI7YTk+IrUWLikzIOelNueUW/jAQHK1u8Iqq1Ap
YQRD2uuMB1TL7uLm/lULAJO2xWHIc9LHlSMzpw+pHXEk93CJ1VW8RS9OEczngT1J
II6Van1I1RJ3bTNfc2Sx4eifCL/5i+KwE1WIIxNwLOky6bw6ig+huJ4JANqCYhTI
wPQ2gdOX9ee/ZtBkScGHRHFC6B0Zdoo8mIl7MyITQO0vgobSPqYONwLW0mbhTnnz
HIwk17mEywZ0hviwrNPxeJyBYqj2EiwwJTaJBMWvd2TJHnmrKDn7Nz8AlOgKKSAj
3/NuO8MdNnminehIbvAfFR1a6J0sz5dIGcpySPCmtSjvJwg7CqwOXTjTcHwWR8q9
UZ8R//k3g4zPpiG268Vn3hlxU964NgdSmv2IeTTF6SPhCJ88dkpFtUMWRTauLNGc
AqpvqZ1+L1SBC5FSf9QBYbrzIvIWE8zFvCpsC9pQEYdj3nzbnD6gvowaQzPUcRYj
ibkv5Zlwhhd1dLgvxr1lJKwkCVOMhE80cWEYINqnFBVUN3iBlILeexZkAYAEevyn
E3zWxaoWA8PrQzMN1ddZUFsOBea7KDuhuML7ePKylxOTeYJhgBs7BuScc0Z6wwWr
mqorvfDs3npXAhbjTgmZXdyVodmmx2ppK62dgXfYDkG/utsAUNtSIsdeCluJIBkb
Ul/bkj+xgSRw6XgorQMHB8vthAc4wHU31/I5VV6Qmj8+NHvR+F1SNXYU/LzC32zF
FRUuOgxCRakopbPPWbhB42FsqqWz/HftAZWQ0Fy2nwlIwq6kyCxDGk1UK00yAccI
8YrgZ2qHfEI49Sjoj4ur0GV6bb5YFMYnvKD6rTiYmgWs1PpBuG2e84qzMKYLCKz2
9blXHILVWabfQjvqB4hR9EKBVhQjwnrMAnYltDiqsHOnY+9JjuWkf7F8dFuoxNuv
k3jdfR3iajhXb+F9p0p/vxVUJWaxi3qDXMLzXUEja9vGJYQ9qaJYKbcUzP+xXsX+
7imDOrdaSLVA1nS1cTQdPWYjZip0uUP9NpbsLUsAzG5Ox7n/InscOznP5xZGBluZ
/ic8yvaX7XoF8KvVhgVeZqecjMF83MZn4DYNxJ9i/YsfrMlQ5lOO2Zet3ecYf8HT
VReGUrEC3ejYgBHvUdA81+vZBllgq9bQTUzsEYXuG/2HIBo4iFLF9HGxYnzAiGMb
3HBu0/Ou+IzLgZFqi8b5lp76VwjWIy3x7OBJTR6sLgZXIVSiqH6ZRJJQfhB2yWic
lAQLznt+owYhVxCBx57BBN/o3CJrl+ZwliJWnD5dVSxFUZivGZvRkLrdPnxiXwyt
i6jIcY4HaI2ChxbH6zVsMJNc9MDUGkF6uwgOIioKeJE+dmM3SQqz0wWp5Ch3vppJ
sYdZEeGzkP9d9JL0LdL4ntb3p7C+SnXQU5GTiqwzApBAD17CFsycMUytbnMEGpll
mqLQZbLVHdhDpZ/GTX52qdouE0bufseXuH8KoG2VFcjWeLzvbSuktDcg+vSC5fnm
092YGINqJK8p9jS7dNh8+AHyetGLTL5fX2UI/k3Mv+1/BxtsmNuyX8xH9X9UcvHV
3jhxRIWzq2Okr6xTVBKScyMdTXkG9YOsQsi8M86V9moGfSdyuSmKlzrTdnrWS+vF
X8wRAii772vgE+Xy6B5dSzgbnxQvUUGIJKS8b7uZvNX5VoARIJOjjMyWA5jtdlpa
z7xJ2otnBFWTZt/2GzTCdyYdnuckki5TdHDlgFytRdOXfM3UUq/8aKeaWxLa9EtP
2XqjtoXHvIpTQ4yJu5vAgv67aZouevQ5Jyf9Ev7WcPOQHsXv9ZubQ1ndKzMbIZLA
CVtGblCdIlAcP+Sr8zi/GWfNjkFABKHidfXYLvSad7CHv1hDZzq8C8v4cyI6hMlQ
ihCsI9HICYQQjuignWNn2y81C9ufbLigGO70B3zlA3wVP69iUqC3991oe3IeegCT
+UFoEUA1CoDo0c7an4y+XOBOh1Z0zoBTsVCEBFDrINTytBVnPaaM+KOqK0HA8ELj
xcfXa/KEPd8QzWOIZoq6KJSBAu9HYWf3XOc232cpZWTRKvS8AS35514izn/n218O
vR8VEdktwCkV2tj/P9uei3Q0yCFBlQrWp/a9sfoMBY/V6XoYrL27I9nTkBAbus+P
9zgkLkcdTBNtdTCHFVkkj14okAwhkFzHUEs28DeO53hMjmpTdgO0Q96fvAStelun
a4auWl2GA1SAnbdAI+EgDdtdmrO23l3Glt66E2wZr00qWS7UYgsDK53/tNIsI9yl
HrrZGUuzcdRWRRDMofW89IOxwqG5qOABfjYkd9f4VBQiPUakXDisU8XX1kdkwTuJ
XVic/aMpsraxoYShuMP3N7amuBV7lMlLH0Bwz0bUEL2BZmXYmjNoe0xWcdXHCoEf
vE4726n0AVlEggsVJC+J/lLRdZ8lO0qltFYF78nC5oTlFCCyp/Jvy7cLFm7mt12n
fPwzXDb343QXFPVW3Q2pjuQNU4KX5LdsI30+9DtpN9mRNt+9Gdd2uQG1/Q9/dJ+u
drt4e0qXSY3VeSG4VjgkHqBQvlNmphZI+dFNGfkWDU2atXOoOOWC/Xn2xUxBh0wm
XExyL0jj/pkAdwzyO7GCLxIDNffkBBzCAqhUogYZ9UqseRsmKWOtdJOAlqNL8n6Y
fBt1PRVhrDBzVhqKc6dlnoHcPS8NvuLI67wyaRRcCeS+bxFX8IdLnEgmAME/C3Ap
/AvP0TFtz/24Xa8qfapuyiIftvo+uGtQYTdnKsXFAhmXtdQWu8pimvUFWRuUWfQx
gTtnE1V3yoXODjAxxuVwXIG8v5jLK3wa14R+WlB4pobTgNaobgymJT4qKYaDQaDe
fj6XDwzQaT3diKf5wSDHrpI7ZRHtscwIp3b5MWC6/Rb4TEKLwXL5bYm7EntD76WI
dW5iQkQsMUUFLTpzgxYgJm6VTcIUOPmOJNbOusVmWms+mYylRfFL1yyD8kGtfuil
4t+/yuHKmLObeapvnPSbLrLIcX8TKF+ZHpOGxV4tL8r/IEIdvw34XRls/26yebNP
3/dYVhl5KIMjkzeswDcQJTBsImQoZr0P27vpnaIDjAGyBSjgavXCIbHfQwWVKlwp
hrztZBydMiRgIYEw6PMK4WDbeAbudX4ldgPVL75cTAmuUbGpCmrRhM/ACDgkM+0Y
eqqmbvFtuJ6r9dZP10JZaMjbe9GG+TiDnE7dgoM171si7UO5yKeDxpAs179yDoan
jtZSCJg04up1Eswk7ol3YkJXafPWbmMJTS0Kpog+qd5qnUGbzQcUqCXJiQ23xxal
NGmkeG8VeJaz0VV4mzAN9X8lgDaes10PBMhmTgzKRKRN3FLY4cSZTX2KJErKyqiu
0RiXJOuO/6DDK034IBeDLvpqx/b7FPWfuBxG29Ib/DdV3ET3Bun6Xhlx+bcUtHLZ
gzFOyQV/E3VflXp/2FbaBXpSOLtti5p1tITLs1LzUCHjozipxHZCbyOvIVeAMwIc
QHO4hDEp76EkkKx4zR6WRi1wDPrKyEvpWsVrcMoIj4JFjPB/QBNHoZcoa2skohWv
LP1SclIuYKv4iF1TVT+bWGut47Nfht5F3kv5u9z4F9ScQNhSyijBg8uKyV9a35ne
bbNVAHwqu5k2bzsXIlPNSKKhwRxpTSeOpZSdHxZXlwfOMD40O1HIdDDE19U0bGg1
waDqBxU7NlEKhMosc8LxER5jVFQpvQ/IEcYvwGpSwzRnPHS9hp2uDLYwwpP6VqaM
H+Upn4XGBvv24lPKWZbkyM45DajV+jqEXVLvJ0z1SAgJfGVJuYDvWFeeCOVzxj7H
QfnYrEvMNWXjnM3ZjHAZWFKBriN3qIzlfqfDA9Kl2Xr6ckCnaDrCo20aWzwZ66df
FsMJQTLi3dICG4o+5p4vrNHApp0Sif2p6zjY7Rc15vjJ4UypNCSKFVIOWLF/sIH8
S2yUnX+CZgnuWO4FurYCQr+Ks5PDuHyy8FiBCoG8Q+rhJFBwnuB0dgIKXROBDA1x
EV9f7ZVStiRyKxNX6hZlzcvLCgNNWpM1WlcWP0s75rvb8q50Ous2MnhXDFDVMyr+
krVl6253BgOm4ymhe6T99w/hddAEYkAuBmHFt8vKETwwgRIsg6bohuSreqFNZy3z
+Vu8wqbyvHuCG9tKiCb1ARX/JqWh5rzPGom1fVypUi2fAoZ2U7UFJMKhESCOzbJq
CTXF1HN15JO33I6Y6+fZLf0xY9p9MVPM+SODbvsn870WBu9lF2j54FR5/NdQLHeE
Y03hRPfA493y648G3yfadADKamChoQJkdZc2M6xm3kYIjh9PdazcGqi+DJbLWBmT
jmR54PFDMxtdMmuLKHpYEDnDrIZsAnJ6kk4QmdbsLWsai6JBPd5pcu6FRzHLuRtg
ysIaziZZEutrUs9bRLhdyiA569n+fnAI8Z3iREhNrsy5wEtYnGN7j1WpkvmGBbxC
AcgjEdF06lpe1Dl4IaDoWJmuBSybWvNtktzivb2y6vPMxUYyXiQTV1fBpsi51Mbx
4IlRjPxnAmCbdfOZ6Uc/4mN5giThWly0rxjy9DmpvPFRz/azKQuJ3RbylFjjsksL
G/tLPhMR9PjxnmYhdVl3aYAXjDTpY317Tn6kHlj6A4fWQm83Vuzg5oQc3peYs1xv
LP6n25ICwzr0NXescq2s7ObSO2MwB0uU7PTGMJzKSsJBY5UVXwrwz6VjPg7SnPsp
6dQz0OT38bgS7P7pESWfWpw2Haatx4PQ2G0wSmpDu5uEEHeb3LCZkPWd5aCjduwP
6QThqSoRAInZXoUTujzw5VD597uF6dpBL/Tkegr+SEqcTmIlPIS8UQpfp4U8nwoR
paY4bfNfkIDzz5UNru1SlnQq1N379m2bS8VUU/kq5bxGn3vR42n0TcNtJqd1iqYU
/XPfK0NWydWK1Dl52hLFxD+E3C/FkrlsJoWTC/zibUZHVCt5ppdDKco7sYnyZ/pb
B9ZyXKpx5sagF0LSHVyeZm2XlYk0sINnkhzgRhddS/iTaOxnp6oUzY8m2gMIhxx6
CyvMdvoDIQGHHFcMjb8e5sOxivqTGf0YiMz+X73qKO/xZdLAHzsKJNmQd46joBrO
fW+irlNqccI3J9KITNDsHB+9slJcd1GnawgIe8IA690KEAVy65dVBEpAN81vwjgP
e80Hwzs7V09/ksZr9oi2xSlwz7q3sMKWDO+FJr20CpIY52/Lgln0i5N+ulB2+tHg
YCdkUU8dvbyqMD5CKGMQxPdFlvNLTPf5+5TpNEDy7nbhDdSlr/+cvxcO7/JBZYf0
kxhQ8CmVsn5e6LhUc5fjGT2QTzuD1WtlMhap5ufDV+P019bH93JHH1lbTbpdOlQ5
lowfyNytlJ/RVIyVjQDJnEEwuRD6tFexpg7Xd3F+Ib+AItJnswxkNr5EfqSieMOc
+e64pWfeY7iIzakPdAKYaLidIM0sMeoan/k13YTfUUVm/gfBBTb4C/QQimaiCww1
FNAoh92J20ft79oNlgyd4lytnpz2RJx4HyZz+wv0ttDvETD3QgP7ng4m/rSXKLe4
7zlRbgKyrPFi0VW3Uy0FyYF968yJV2z7HI2yFNAy/6uteGrdRzbKjz0VNGSsloCW
LUXPAtYl1zAioArWD1TjwPHN7A/F4e0NbiOK37kxZcuuGwEG76f00k1Zctgpbtpf
gH0OKt1Fqtk/ZBkTvq6b/Dmf1k8iPwKDg7mIWNE+YCxsWZFTFXo6OD/AcYLKpUPu
w6JZtPWdptuLmLWXG6nBJ5fb+Pbirl7rqV44iarSUas0rFR+XW/KoT3qxbafBkTX
npdLfUzd+La47b4eeKcfIROAGxYsAaHfI+wwvtxerUcTexSBC+uq4VSLlGjDyZjH
9B3D35CtgS7mcw+715OKG5WbyeggWhhacHr59vvdSD0usxUZVJrl7c7riEDWeSpE
d9itEFCNGfntvpLvIR8WmeH+jcFFy1bUjR0QsuK2LGuz6gOS1nQ7A3h6AqKlcxpz
VVZLE0EX+kVo+6oQMaJpMtM9k6QZWzi6fiAaEvRATPYjwLJ7SUz85UUHBJdbdcLX
AvY9V0usNeokb1xowihbOovVpaidI9/Cwr20t1zvKsYoXPlZ+Kkh2ve0MNa6fS1c
GQ3+/ZoFDv1hpu16vEKwvMN0Swl3YVpmGK/n8Fnu/PsfoUiu/1Xxo8qb77kkhqWe
PDRc6ElQZynE1VgEIUuCDGb0ZXgBSnY9lFDMB+Xil2ezGYKrFOAdYUPzZVDS1WAc
YCLwMJKeUP2EtByOuERoPknPEEqXhCvJ/W4jPmkAaIGyOPdwIyTUbQpVbPnZGDEn
p67Fa/k04m5n0fd2GKUvEHTXHN2UaF/zhE6RmsLXsb3ieJ2moKOUCC2RvAi/BwAV
G0DAOfLZDGAhqk91hyxx5CyM66+L7q+6I52G9ntTQ51qFEmuhiCV5YdpTOVh4pSJ
r0HJ37+fzy6r/3U/F3wI16InZ/3rryobZajDh1VLLT4UimCgbZTBtGRX7c05AOMM
pkoyGxD+py8AVhHgKjIOfRcUJ+yP6UEya+Ywg5Emd9DZH/VM2nLil9HCAEsCxYou
5OjDmXoLBQ7s5IEeztU+bxllqiv6YqD6gw1Chk43yVQzVQEPDmBDs404EqGS0h9d
VFeTRTAPg83+7UZP0AA/0JP+uc5EUJkoeL00sZaNe4H4wnpICdaahrb/IOjPkSr+
g/M0qP9DV7E0vAY73MUK8va70Z9CPFOBZLwy1xtlrAmkC0byim/6BE66/o4qvD+O
QGD/kPQQ+L7Mvr9QfnyEA3Dz6E6YTCgNvT/AvrOsv2qVL/9Owh2rcWf7CXlWt9Kx
zGb4JKztH4cwpT/wivzuIdvF0ELbEAe90IVP9xcjg4VXajPST/SjyYmZT/xKD5H0
jJXfbV0HlTSVp1hyuHn2DgunGhTi88n7Xmlv8B6sdYzEv3Lknsl+SmbjASHBl7R6
NPxHq2b6nYe343ayurgbNEWYtAdI39+9zthkbO65DxMJS4TcZLUBEfP67nnPJYYB
6AAJ8rupu82HuPORlo02iprUoNcLqGs0qfFNK71gmEcHHMznzte7b+qorOBsaA/5
L7Q2EP9m7mON2mljWE/6YdvSUKM0MFupM4H6ZP/IRxwKjSZsa8oKG1cms2VSZTDQ
AridkdKOB1GyAg4sNATvG7Ro+yJv/xJp5BN3bDPlxrQHQzPanJyNpjKdcWLDibpA
rJtYNTJPBE/ZtDZmwgKN7EAoquQnq/ERZMcY3u22VC/nI7Uakt38/xOOZZ4/erig
AD/u3zkfA+DHU4zk4nlx0lyVwbxfvW4DTbPlTCRZidn/HK+ypGWFF/4ryNrrdl6S
CgJxNS3OU/GC0HM8FgD5muXGQy1k8QcHEKk1HWhqhhnU4wxvZZvRdLIzCMMQ7tmb
vOC0w738TJ4nJD3R8+I6HM3QSkM6kxGBBeV3gxoR6/U5LaGbwMjStSTSzSMYs0MG
z8JTWT3UybdGq+hvcAUrPNzPT8rHhR9oR7YHHjNNBPfZ7FpkLfQG679BsQnjCWzS
YQPEDggaTAXu7sPoBeP1sEDL93y2tPgOAe3LKuDSsJkG6a64zoSSedgEG2hdvA5Z
1Pyh73yTYeAwNED3MmD+6fqPr33SIdIKsB5Ustx4RNtIeAJ7FU05YURrISzBFVXQ
yuelyWuPUBq6H/CClRJuJ51BTp2QWNaHmaGbnqGMYL+H9g73xSogtU1kC4bJtjIY
3n0kV9A1PY5P8SJoZvl/mP9SsQEJaqQ1eB0UXs/YTKRJurY2CKbPpTFjUtQpcQYO
sDqIBz8naRAkKe5ShI7cddJkVCtUHOjWHL27dR9CNU3AOCUCxX3/NCvdNtGLqEcM
8NDHv1cNkqI0JAfwEhE3WHIXknSdyq0fwUpVLmGC2hwx4PAx1qJxwKsRMvqAprsx
/AjNMc2fxmR0g+F1xPqy/csE0ENBfEFhF8pui6U1Uj3ldGnR9YSU75NVZIDgbeq5
boj/OUGLupHFUx+JNMQgnim3YEJ0IumfupHo38VQCu6VnH9TQW1/Td7nV3BG5xIM
FZLzNKoodXDK717KhHaEeF82gb2Y697VOset+uRoaggVgU8PSMPgVgF6jRMoPl1L
gnij89xpRcQTPKYTTp9uUfnZAPf3PeA0hBpoXJv8OZ+O1q4CF6e5JOfRFEceL+u0
CrHPplFdcfscz+IJPqMoLoCihGswZXHbEq3cX66Zj8yoCrUUy8DhRLcBEUYAIIzG
KBqb7UtN+jAWUdaGwZFX1Y7hLg8cSmw40QrCQptLEgiwcVSdLKm2J2KcHt6aeHpO
/0tk5dQQ0Aly9BNHof/Ou96fZYX7/1FQFOgd5VhZEparzoZ7SQWsw6Q7TEncL+dD
c4WQsk13F5UI1ZUNv3X9Ct5ODKYvLGUEIsK1nCOW4ER3H9zLmDh3002NlaBOr19q
6YVWs7Pi/MeYcsYtSn3WPDO3Jsry/eKnoEI70DCiO1vkf+HYEZ/m3hhXfRD95fqM
cx06Hbw0Ix2GGGYBbjRf4W1szGsEedGB5ggdgpfWlZnAGTFvNi/HjaiEY1P+cCD6
YsI478DuSY2YNJ82r5iWvRYJ4XMYkYKV54Jp6GKmh+v/EjMBJHCQsXvAEVgo/eMT
6HDdDVirPj/RBq4rXK1Ogk23h/i+ARXac2F4Ih5mkx1jKzpyDDRCaxIcuEQqEm1t
R/EUObByT4iYlfmtm5LQS+/g93aCw+fp0dvzfAp6CYFeyzlMQz90ILwQSNgMWEas
aLZj+E+gR9zOxdoXGUk2NDQ2U4s502rreRfjwnx9eYSohsLcdTC/rgF4hpW4j7OM
RI1W6xyM7pjzFOebnrccUyx6TlH2jIlPTUf3XBAZxV6Pt2rZ/0xKE7e0Cb1tUeeq
PlfVnFGSUYcn8qGd3nM9mqXIxWafeATNrm2JeUKgFb3/VDFALXdu24KVQdoE/je5
9zd6FO1KdRu4NYIhApjXhhZFaT4TX8igcroNgY5RUXY9eiSxnql2pBQSixf0jvKj
mXzO6caRHfMrOIGomSOVodkQ8KFbQnVsbcvA+6ORYR4h3lCmi7qzlljJVHnQ8u0o
EY6RMMW/UDX9eGQfktYww+sQMthjCwJOIv7x5nz6KLODeq4280hvTk/TN6/RRmVr
imyJfZ1S7Yi96k74C9SmgNE5a5Cjf2rvmhc8pEPdociBQSXyLZ83eQe7yvmmpzBS
jV17Bpbkkd1SqdrNEV6/0RwKMgMhuY8LyvtPV9Ynj4GqC8yfTR50Qblffvhofg+e
lLW1zw9fuucFpBykZHxQL400tDFt3bGezjaezu2j/XM3XSImQYYQV571Y/CDnDK3
n5wlFonzptud+kaxOIryKUdwQLpBzBLuB2ckRYkqKuk9XHp79QqTuv3TQqNL9/pi
RsMXPiE1FZ73Yi0KbT3DZR7pIuGq+fP6VEplucG+82TdHTasJVusGeRPaaHN791P
gv3wyZ3WxckvY2U9rlvkVMANn4pTc9Z1V3a2rIB1Wr13MGlkjccX4aC5/ymxi+ZL
iIqdfuMkCgs5uN10NVHl6w0ubCGXR0qup+TW+ueIwqvCTGarc6mSe9lRUvyc6gXc
6cdXvzqK0BnoyWtCD2VQX8cU7AuhCgP+yuRilXXbte1LOh9S3yOo1BqzxLj3HUrO
bY6Ah1FbT5DxbyDG1NNMkAln68dO7+f7z7iBxVom6qbfc7kxPCJZX0qaqTkktPpa
X9hsUhWX7MZUUjjXAOa68rG6skk1L+6fU/gWjdJ2DJs8sw5Nj4rICxH2p/xptWoR
EZKi/5vEpmD0duOljwGpue/RvNlxPHAuFcZcEYIXl2ouXxbG9jkZb0I17SKvLhI5
3nev1JoDEZB3LBgA7jMH6h9insLomxh5xFMelI8YUxGcHOMr00377+FIK0v8udYv
e/LP9hMesauKE/M8UPnKdDTWplTc4zrGUSfWbulqyh7e5ldR2B7ReiYyhemr8a/m
S48Dbn7lGxajtQWJwOALGBN8S7q1Rs4dmgF/lQJ2qB+r0MJ2OLvQwaK7+ZZZ3MtO
VGMRAh3bgHbfwowuFidHrTwzFz+201i38BQsGv0x7AGkHBdyFBNOopxq+QM3x8VA
6bKpZ/DZTStsd5JJv6JHN9/EdMigZ6B6gEXtZnhZBJfb1rP7M1lQnBXSCrvIII+W
bpUgjcr2ymSy/84q5s5txldBCSpCfTIHF9TX5QNQB6yYXv8lffV22P7E0gMJrgsM
NbHFBFQzx8HxH71dP5/v3PoybEW+icuJu+z24FAbPEvR+Y4m11A+r4wrp8GUhJb8
VchmhkllFTx79JaNYg6YAOmvdRF0GCvNlZp/IqoGvP/SWHS5lxUbavktg3eskQto
86WKIlQ+/ULZcSpH6RtTs1j8hGpbvv7qSpzS0/z7LdaftJpiPulglQOF8D8dNq2P
mm2QEAbiAHO+5ja9NHuqUEm0w1c2M5gGq0yV+BvRVsZV8rLxv53DBhWUF7/IQXDV
VI70A2KKTv8ZQcYO5FQakgPddxZBvMtXNsq2+oEZOfXbD/DMEAhluICz+p2m/gFc
C4NRnlfxRAVf+R44MK/9oT7j3WFb+SEV8ozJ38OPPaH90Q09bJWx0FBA59ao+DrA
KbY8u+fGselremmHJ1tqCOrBWE/xTEPjYUWlyPS1A7vB4zy2gD8mvfsosB88jFlu
92AaZBLrEvtke+DSI7e3SCFQDKWJb1IpRGeDsqSF5W6C1/3K4CeWMl+nER/O+YZp
VGaZwrwDZXOrEs8GXZFcjpDOokwOteMsSm4rcMDDSm13yqnTykXtxA/yTgooP3JT
7ciW2YJ+nQkMj4Cqnb7DAqJgh4Of8D/GkYJSaO6xgGcVQ70QyqrGTOi7pqjF1ZEx
ZbMcpFmIFl6/od4u2LL7t1HMUDwkuMoFIhZ9sjczz9yZKcwER6aSPfp9DC9lXv/4
gRZnsz1t3X+bDJd+WpgKa+m1o53fGm+vjGh4AqDZ6qVYB28NA2/GSnLP/nM4on54
rQEA6KxE2K30L4sNtWbUyjSdS8LD8LIpGRVz7K1ZfpG3WlxzxbGg3sl1E8xiF1RD
zPn/uHsbtgzqTQd0p7ir7xKAvfujOBZ0rcDAl+E/N3OpfTxCYQoxmU3qMtw9Rx5m
yCPUt6JeJoQ6p/b1UIja8geuH8W+VkB6gO9zoJDDeIghI8EK7P+fRjnDntRkZdxZ
mO/uoEiDSqIkxeXmZMeFtYuJSLkE4KkXNqU7C3OmbIDUGZr8QjXZ2TleoeONfpBz
VeqkvRuerNXDEfR3O/v3FfPYuP0wT9onukOySACUKPGFYaBzqjhwKLMj0bOiFRee
7UmWO48BFAEwH9ZQmbOU2DHLgxMeVRFpYbdRMfEASAKM9Xqh1W+txJvWrWJr9wLT
S1kxM/chf75bJbe0dBVy4tZLI/YTSivRvUEZsYyOVbaJ7BdVizlMKc2aDfjg8IEa
bdJ4M1MRSZlPhj0VKsonY96V112Ew0JYFzfuz3orurGYHB55I4KxS6L9AzK+gfcT
HQ53HOtQoV+Z9qOQbsShtAmOwrnZSfdjUUn4CHIZ8WQRIgw9eukbwsBeKS6lwVXC
pNiDmxJjrcjmlt906qLGiDdUvKjFwrIOS2IHlMVKQivYOJe8Ag8ZiFtc8Bcav8N/
YASitO7rbYrsFGJ3e9t65HVWbnpP8hf5dSCXYUGfMBndTW6zqMosa9s0i8d5ldBn
xws06UeAJo1ww7r8cwoGdNZNePgO0LVCxlXIOL3bOIXO6QJuKgbwWNcfK+g0PQ1l
IY9XQUcsAXSCnB+HbKCJ7kTo14KWSjkyK2hfXT+vqc/7uXkh6jM03UOVulk2ECOj
+/PO8AubjV925ehqtAMPOArwOuA9zUQwKor0hdOgOVKq87fx3X02Z9jX+vEb09YM
HwHRw2cAW9r2SfdlWDDgseqY27WzzXx7dMTXg7PpMokzWqQ0LTiu5iYjtdJhM1mG
da9IrX1b7ewatLGVSQKSFmPEmx0iqAvdL+PdDFVtn7fSdFeCHN6a1yxNyWkVZUYg
X/Z6yNX5U/li8k7pmzzJI8SF/SrltRJ6Q2c0S31hWnIr1tNn6SHNBmMJflXhSbQR
wVC9J4M3aRCCyRhkWPxI2NNUH6lffpZLCb1weaNnx4BGqq8rii98vaBelwrm0L8D
nr7i/cvIAorRRKFkC2+JjCF7rLTDsjP47KWXBwSbK6gevpP7mb/r/eLzexAMW+rJ
pXhY0/odG+8l5fmNuMzFzAu+D3/teb2ld9lbGhHgACXaKAKOtquYynirF53eTSlr
OeZqiK/OEm6Kn3B/PZ1oAzJ/kPerauhVvMDgY3+Hkd8XS5LBLgE6pZ8uK1psS5PS
x5bwWrZl8MTbLxe2bM/1KkUjJevMI6iMW2rmBCdQ0dscOwUdTcts5thA1F3jvVgd
PjR/oQ52vXlGJf+itgIbnMBzz3j6nnO3x/3qGhhlC7i6FOo6tfRfHtmi4HCfKBoZ
h1qp/NTZS7fdwmgvRFzaKFjdkmY9JmYkXdfM4M3izdJKToUlt7QKZN/vWAUYeCP6
yF3fO5/VGGd7kfrhXJo77rBBeIeSVfFK8aAF8pUyWShjST/SA8EesK31ejS0qT9S
/RQhWvNqAQLlZmyK8PQlfxXv0OKDpp9yaLcEVB/xoDMLpUf1gUYIYoLql3Lrce++
oKJoCu7sP6i6AmX4472ymKSsa6qxfg00Bb1V5oY4f6ANawKDU9Ge/vUmfgkOW/qB
bAuxU/NvVZBWXHgHY9q9yJJVF7sNvmD6Gn4TCPwkUjqWxG1xizUrEZ27l3ppBqQD
JF0P7qCJnuGzZO5GkUuSBeer18MDhaPSJ8w1LJlb2MpIG6rg3rDnfh8QMNRx2VMp
GCjiz8z9DnAWF1V5yM4An2ve9utppQ7EDqqctqONVKc/TGNHEUKdBiAMpbBMP6Jo
t2yfNvSHjBom4gaSgTvgSEPO+VKg1txjYgb9xC5pDKTZcebRK35CqaT1hHeYDwGf
qtACNkyt6aSkB/rwXqgZr6K/y2kEq96+DzNmGI88fsrKdBNP3+KaViDz0dYh0qg9
GGbs6wB3evnXbHmsjYfQVlF39PyXMBr0nV1ePhcck+F1bEQ39mgBFZUYe3lCC4wL
tIELgvpTd3Ffz/AQSsVm9w73+rzolAzIBuQi+wuqTu25H195dgA5nkopX7CYxI3k
U4irU4jt3unskDVGF/TqcTrIypOnJ5XZkI5ocu79qlD5L+EcvO0u+lI0Lh50biTz
uWC/QkSSOggkkzohKYH/C4NeM7izpuuM5EubnVRtnPhdtnRLCjXZbhYAcsRVCfkv
PggSYz82qrLP+cM65nwdw6wrVa45/s6Av1Ln+VuWsW9VSl5K2Uav63W6AcbiGju9
v8cC0LKx0Y+MRJjEM3p/VL+sfhDLcS0ScFgIWTzgZhf5Whg32tboFhxwIgqdgSz1
1gPhsKKhkCiqu24IvCDZZgef4ZxT//j2ij7MIKs0FNbcuPd81Jj78v+7naENLSTn
aHxnlytSn5k7ruxQqYNTJ9wZuLrNdLXzQO5Z3LbnN/qWqe5skc2gOibFUsMe0TZX
jqFqLJjt73f3getttnInvGLUrFVBo/P7QlLAzc4yN6I9ZXGU6wAR5+uVPvV8Sunx
43eSX1NM0g1U15Dvl/oeNz45Grc3eMJFQZWzvzY/B6SF+Fme054LRx2+KTRsXwBz
Vto8DuiAVx95++kBQRsYGltVnfDd0/2nofgf0ek0f3AiS3b3XorwNIwe+dlk5vw6
gzolSKsOotIdnUZ2dJK8xjh54k+1cyjsaUhpdbKVQepUaFWRJmYyu0fJsrYhD82e
2CqLuWXTagiTRmqVrYCIoDQWu8B2CQl3FyMdCpSO5WTtKGTibdiJiqBI5IwJIAn9
ooOXOowwSUA6t7pTVQ7BkAwocIpqE82VfxXp+ujFkpVtOFGyJtZJ9WFEYG2LzW+i
rl0zMhLIwAm2ByxhbYLW2dr0UprQTUi2lZFs3GRznSh5QpyNrYdtqM22lGLAcNiL
LzQxRVcKwjKZUx19c7RJVgy0zcyx+v9/W7Y4vUYPYh/p/PXT5sohI4AlONiyYh43
WOAf7dMFM4wsSoYj+T6nMYP4pWsQCiyzX4MabzP5Kihd6O3SJ2bRqYLonGBmN+Xi
qIbYhmhQbrxwjZKl8zHHT1S7nI3fG4mJFyd0jnHtCB8SNSN+bOI5HYMWpsSPJg/S
PsSiPLt6q2gAFPS7OV9SIrS/8T+oMjhhI0HAiH9lMe+ixATwsEREvAyvdsglsSZV
KON1wGf9clDuQ4yUiOtUCGLYeWAu89bifgg3llUbceRWtvpiYWqClrTj/uZbNdQX
W9B4A3XHQhnlnas6/qRkH9HAWQv4qP5kVvCXKpV7e/dCTKUp1KdPaurvMotnuFQX
JdArCGa6UUvegDur1/jXUOqLj4RLBg7wWGwMzPwqPIRpfLw3noO7DB8Y7E5P6Sdr
5iQITUCdhF5fV+gjWOd46HPryu+PwMdxm/aITFgTGySzspXYz+9t/gsc5KzIqPK0
IMiLGnh2p/SV0vgjaByIN+1oDEPz7Uddx4XG3mFYe25ae2m46XmHEPKzHkJNU37m
x2jz/H4NXrVmAlvqVllyY/lftDHuhKF/WQfVBNjyOzT9lQs/b+/9UaU0tNT7QkOu
BKNI8lhIEAz4Wd+el2b18FYugerlPjydweZlc56Urq8Chk4DIMO1cAHkXGHDr/xM
R99NcCToetsviZn+U7fg/UgBeFxjs+XYRgDzJK1pk6O87LdddreDsM9ldsaK3D0x
n44Qf5vZvmC7imeHWDXkZAuPCpNUyvOLK6ZHk75BAb6ZBFEzuQ8cZ8e7ghQOonja
9rb/7ka7JMFi8dZJ9o8pU+AjV1+WKzXy4YutUWZNapaKUGMjGXD63rz4BtJIi5kE
pJn09+gdigZZDN6Cy7+5J6T57BALMW0gtFoJOEIS0pGPDdxrOWIci43K/xtbiuCP
9LuVPHIskglCO8lUtrRZeCQi1Hdu8KWBCmujdOYrno/8WGN+Gi/0IbCZj9d1ugkW
szzLRooK1QVJMIXfZq2DI+nqEcStQJ6WFPPhJQs9w8KLBK5u82XlQsnP3ExBrl4Y
FM9xJpK6s5V9fh4XpyoArKVCm5KoexdS5SOu8kBwL3xC2PJHqbcTeDXWdNTQ9F7d
66snHFBt19hIpylmMynrwdnXjoLLlO4zUs0FDjPMeAf+j9uEpwF/Sueq9m+rY6Mk
ogv8h0tChg0sX135ARBinHYz622q4zFWJ2G78SooQS98EJb3Tp9OGEILu3e7TK4Y
C2U0FC39zPLTJ+Hphj0wDH1Q36eyKA7aZd1AbBhDg2YG+MVA7DBA6oyeuyKV3bW6
1sEih4L8T2MxElYFSw0Ii77uQO/OVtR62RKgvXyeGqfnDNxMAnnzzX0kaOBuICG2
QsJfa80BOiTVBzNu3sxbdYfATpvyHI4S6QEnTBuevHmdX8b8IXzMFBFsZtcAK9pi
luY45fN0GmzTmBE33K5rCakyOp6onEh1xfPMtLl0WHCAQx+1I3sP6VZdWT2a/4H8
oqMtOk3F31f9POit3vvRVltQuQzYb/s7N+Je/xTK0T8m2LltPGw5f7rXfWj1JdIA
BgSG3eEW0YzYmapEV2HhemLaj7/HWiHAEwrKs8dHJUz4MHVLzp5aBeI20bzqisAl
Z22I6aeQwbNGXVznbJr+mW6hPcNlVq2wfJHfGrlKA3NrQuAveANUUJ6bRroAymFp
FV3D5Ybn+n6vgfcvcK2MXPd8VQ9QvtrsfQBYZ5OstVeruAvkBLZfBHXoFTpxtgfJ
w4bPbDhE6KnGiWXPTUNEh1vySpahYnN3BSkXAWAR3JwKAlice9PiXqL78/uDPwn4
cgdrCYaTb/qgFzRLWFTG8z43e7cSzIyx08XB9FAWc3cWeNjjA0IWRcpBso73nz4m
5MV23kKGiQALCsbpIAMZ7U5krclUwYFfDZrrudz4u1dbNi1A603g+NynDJOQZi6h
eEDpOKsYJMQf3187+OjButg/d5wpDEDgxLflbUbmlVtcgHKpH2oRi2iQto7CE1U/
KxsR273hTi5OZcI3+kP0ZxFtdRiX5NpifgzofSeNegGMumaxgDeW/jyTJdCwu0Sp
HtCo/bEnbigt8JG3VVyhdhJuwn00h5SS+jjahoTQieAtd66b3+Cjwu1DdrKP6kQL
/Jvblj7zP8tvUKfZu3TiIdwceokqLaC0r8lNHczfhrH0aieutA67I/8jqDRTauZj
UqWFHCDcOFOj3tAE6haRWAqJi9DIofot/bKol+Aex3Do8hqEoWO2EVaeRklOxyb5
FvPfok+zfgvJSjCkhFtCTtytNh3eugPZOf7iPcTxPPR+gXbtlKU8mZ07ykAwD92S
AldAgaeb4p4DKnCedp6V992xmxuDUhnS5JMKFbNIRbRs1cxCa+nCsLb9KjJEeDRb
rSXWz9OLtuubeH14AEXyOX9/ZaBkMafdk5kP4XTNt38sKrkhmpt9vH2yWemf/wdp
g9xxguf1uYVEQueVvr5p2YgoZt9H+ACUR2lCJKMBNYNJwM1khyOvCO1Z85q9EaVp
VWsH+P42JkEQC/eFegY9hHX1R4ZF1Vb7O8dhp3KooQ4YbzBuVjJh9srMTowyGJLT
VsHWcR4bVH20Ki1wOMu7kEUFSDSb0nxBE3aNN9qnBhGgMxGxeKxJPYRBOV32gauD
NUbFJ0vCTp7gee9mmPwC4gnb8H0R5Pj8JDGG7Wr+wshAVNEc4xHLC0fHXO/JkRpD
D0IdzOcV5+3c+l1f6vJPnHV3I2Xl84e3HBYh76OuL3bD3cSXWZ7Il5AecQfOP59n
dF04R4xXO3t7uAPHCZuKEPnPNx+C/JC1tNvcYEX8MSPiKMvK0vPzv59Rsp7cpZJs
00Po8ALjC2KnxdlyFQOXikfgh9b5mJWsha3tAokDipWyI5eHva2e64dYj+8U9/oS
E+yOQthnWvzc9Zt4t8IcD96UEkf05OUEBxjYbQ8J5nATEecw5GLl/+fRSSNlGBnS
1de4+pSHkcoJByVmGA0+PdKgv+7hbFiEDHuJD3rXPIl657glvBbpsrCr3ukSkLjx
nFnq4LZHTb/1H8HFVUpPO3vEl2WHHW8BVTSi+TUiWDdDvOOF0Q3Zp0SPHf2cylyl
Y088LBv1UFgQg4l2gE7zGS2hHC+U9lD803fnWFLxYatXfxtGUDJ5OVgEhRtFbYgk
0Qygu0ddzAzBD2LPGbIUiqdAEG6EYCm0ux/xKtXwncU2JPOYO8Xll7zBdaEUpCYM
pPJ3WJdNI4TRuuP6fEjd9lVjpnyzr+v9cGpmYBZcUSwXZGWUPm09rZ4+3kr061D1
q1Sq66RoSSbiR4ERrXD1f3J/axpL6Vo/Ovj97xe70fyocH8SLCm39RXSCui7RPVv
QASbu1YUcKhUM+aRhi/42SY5/D2Lf0V3iO4sQFBpj5DWUpU6BoFuvOxAhXaLAApg
u0DwzafYcKiiWk/o+t5G2yoOcvL7KIbZcHS2Cg0auQSQJf7twdeR+JWq6wwpp7Bx
rz4G1ZrCyvrVHsO671xNGzVs6qNqJFs/bA8S4l2nQvL/7Jx3KzdwslNt0jGUgSru
JpsUxnszq/5M/932XEzn+zd5JqMdPT/Zo2WW0p8GgCTZMqxub+zsJVz97uldESMr
ZPqJuYrHIS9jl3jb1ZICFXYb3FXNmdoDMwvPTS3zHjJsN3xohc/mUMi1syIrBx01
v4RLI/F6tVZjzdrnF6bRmi7PXA77Ueb/KNCEFs3tS8f3NTRCwtsu4dDhbBgiez0b
Lxq0Amlptc+g8N9UK7KSincRBHbCcOwz+FuShm1CtI3PsOdp4eleOVE1CNaNNE62
PpJ1NNcypHdogShRJ0+uQUOdLhEsU7KZSImKsL3yWKXusuvZjUvlnDnWHuWYSGqV
Ro0fL9ryW6pQhWreF5gVrCwYbpPNf2F03P+bMGyyh5pFS98GJZCNgJv14IBKNFc7
arX4JMWEOaQE0IlZih0rSm4F2ch/4rz8C+oDlCGDeFYGWdCobE5I+f4yCXsgWtXX
IbET8CQ6uhfV5Lt0Eedufg1eLapfg8CRs5fdcckgv8l/A+NXs4j14XqDlzhdPubw
5GVWU8N23/Z/QhpMT3YpX7wuosYPTiCD183Yy6WaY/bJHSudiqS1n5WgH8mIubmF
yac8SAEHbFLMUAx44jRYO/3K57dD074IUGncYbULUWe4q2HbNX0G+pUiz1S3YzLW
YKcXtrsrg2ooFnswxTSlmwakYDhDhzMe7zW7khj1Qc0jd7NiA4fL/p9cnLtIdwwO
KIa6zKV++ypbPx/AJkwI3sPMxc2yMJagjyEb69SZW0rnEXTI1Iylu/Hxf/abbA5X
2yf/psuzUJvz7hJpNAg/w7IDR12EPORWg6nJbcv53LvdZI3nxEIdXGfBu/W+dgH2
ZSS5R9g0klttCKU51sK5pIjqzqlVs46kVBnMnZnmXFoLSBn5JYKhI7ivmR56Ql4s
JNigJy1vI6NQI7xVGChyN8N+Ua4vAdGqu+I58c11qxpQ9wmrXvWXIuRA1Fc0TcIR
duC11fesFR2I3q5Al6aeh6BVp9L2ePsEBN0lOb89ymvqUVPqyRW8L0Hk/FxbY1kQ
DLwzglnlHX6dFN2qnACkTW23Jsq6S43pXgZnKhHySOczIbT45uXoDE04edxr9P0g
8mzlGuzP7B/bIJn6Lkf7NhAVTBvFl2IFa82nNRH8liR5+25gntMo0GAdP2JcF3fv
VSo8Y6VF4HAS30ccWiKoU7+VMcMcDxv7PHCqh8wugvpYFyuSFh0uWHyTjUESs7/q
hHpieFkWpwPSON5TRpzWLrmb0sRvKyIuA0JWlltHo7iiOEhX4ER9j9dDBQq9MUZD
pnnydRFih8LmDkdj2Y7sbumJ2HItMRc4QCNl7Ua0vPpfURtfafP9EVcDu/HshPSk
96K0Iow3DWvsCUOhxzScUN+LvO5rH4pq5YeJBJW+Rd4BXHnjwaOWXjNM0fyGjYwS
iasmyqmPAvzJO0U+w9XSMVzfPzmVNPR8A9t5DcMlQnMq0vKd3ChV9p0rsHNp04su
X+Cg2L7zzq6XdzOMG2mYk/b7zVelliIy96J1KUq2XJfMTNE3mbGHEt5kAGarLLiq
npQ0HxveSiKgecCv5QJ5UE+fuxZPALhYtWX1nHKJuVvRElU8IFgcvvxeTw33KtYk
oLv4x37yjFoVUA24hugQZiiHVdJi2NA7DIQKgpZQMilf+/RCr6hNffNNxQHZl0xJ
jHakNMbz7SqeC3HN+syrFTw3pFJvAUzNXkXXgCY3fnJYpXfIAG1jQ+71q0mnh+wx
XKQcKPgn2/tR9QqOiasEddp7wtosi6EyIbzgtey4DjLTM5G4IPIgKajw7Ddt0Zqz
FpG9wcAN0hqE3mb6DALdX1/zAcC7zXK265foxaIqdio4gWSwcHjwLPfmhYNzamjX
dy5GXszMO0sojgo5akBWM03Jsg0jwAtUuDpO4brq9AF6HjU7y/33N6S4zaxWUdaM
S3ytAdyzUAO9PJBkomi6Odh9hf38JWYQp/evTgLvnALZlFoNpzRtjqeIxDDs6Is5
ihJupK3rBZVfF4nNmJ9cY76Ax9TP3vt2mZVG5YC47dZtIrkhw47leyK1otkqldIa
xGof9rAXiO7YihOjGZj5+yLH8nNN9+fNAJd2DiUpFdvorWZ1AQ9Jx5XXOA0KVupt
fIVTkrC1MlgexObul2TPaJCiALQsZEc9rM0ho+JSXPmBRjcDedzy0EyKEQt7/X0d
I18ZiAdqmY/7HL/zE5P1c1D+qBt+nyHlwkwEhb1zVleNOuTIheOZkb9pvB1GUF5Z
6oOdXUD1vlUpxdzD9AjUN2M+19BjPSB9kmu0QRardnhNS0uXRXnlhKIGrSa4UPSu
hhkpca4MyVHDkGHxnQCcWcDbMICArgDrV6YyRdK1fjg1lQktqQOdpUuZDwQJ4Kie
hqPjP2ZLBtztjVAnF2+L97SicO+VjMypF8p3iwCRWprNAyJfzf15mdsRAwJHqsGr
vokkeWRLADuOU7xqLDz+Cy+dkYQ9Nkfr3CjuO0/OnV6kVxtihgHwuFyYiyng6aUz
eAycrQkVVDKw8uzPqfuaYFegQW9paKtWqYNteOTakOghQxHiwwkcTxFmw4JiZ0uV
oHWwOIE3STnBCFaxNkMGRrn3bMDkvdrm1OxYPSGOU6s/Dxk2m7CWAkMIAvI1uvfV
ofR+65pBQRppWsQjAPGi5OBJisN4zznkZ9SPBZgmoI14k4DHMr4YjN5mvYkqG+FY
YLdWeMBC/a0UG66qwrv8cqfB5u/iNEayQ9Y2lcQpSJNGtbvijz7PGVmJIRoAuv02
ckMyKl6WQ2cJaYOYUuvYkc2ynAdOi1M6/gcnYZAT4kGZ55ECfiqLnxRpZ3GYUa3t
6b11nBocAmO3Iayfcpyk3u+52er8BS/8RXmiNgDlF6UyeRdRPCfxVhMRGR0Zz/yy
5+IrC1nmlibHQ8Gyb8S9DcpFXh9YEpQ/eU52zJ8x2Q7ZD3VarDN9nhEVOupNyjoI
QXDzJUlBmkxaWdN2oNneMBy4VOgdCQhG5L0XNZdAKJopxjQCyWVxM1Av3Wl33c1U
x15jEl9bvCUQt8TBvc0glQ1/FfOTcipucFX8Rq/a96Vr9GRrubARmJWYE6V9of2E
FbUPoOKiyAI4wuQIgYuBI24YkudvTCijNdvFlN3T6z5Txdfidr4DnGsaWb+FDSfL
9TZmxm9C5j0akOq8S2LYBf2TFdKURzZ7UtMbnz0dHq59LgGxPw5q1Dxh3Me1bd9E
/4wUsZmgHIsJjWfVpz7vrjYgRamKKryuGRa89JYGjw71ayquZS5unHBx50dfVU8R
d5+QY4uOqei66Fw8vrt8m/WmPbs9IEqS2AJXaj7iZjKck4ggzYSZLFvxneJmk//O
XoRVlYZspn9RANthZ6KnipWMaW3n1AK+03U6Q7hEhxAk6oDnxChLhNAbhWA9KW32
n4V4TiwlNsN8BM9yY2bvaxrVc2fS77ENs/k30PoBhNnoSFNUY1e2wmOX0XvbV4lD
DAewLn+GOFiREUXY/+5vAI7gsulrPTKvFwFRF6yOn/yyVLf5DgfnAqofYZHE2xDV
Pqi3tWuk97pczDHE6DQ5mSXRMN7fkfiQxaBxUF8cSZbrS4VcKfFEvfsHrBVE0bQ3
q9XVWedqf6MXJ7iFSCLLS0vEEjfhd9cwpQV/LusB2SYTql+iXPLt6ZkeccDtpNTc
mFaW1nHCp1lPIWppJmmMXi39crdhm1D8vITv2wjxZ/TFoPrOGb0IKpfh1Att4tp7
VXu25Cqxo4E3fU7ah2IcjYbm1nnlKQDcDX8XsOnYURcXXrxbQLY0NTL14bfIXY/b
z2Iv6mFHhJ0Ng8x1t/RY4i9wucqofwL7KWC/IxmzSAPBCf+nBR//sKk4s1AYlAtL
MRt52Y5ZiUuXe1Y3Uy0azJvFMpTTsm6kgw8UKMm0u+jWcuR+6iwvQE1vAlFev6sw
ocry/9C0kK9DoENgAymeLyZNaRf/bCbTla8zVNljOVwWbEY+A1sti5ZLe0EzZkTT
aeX8I+36okQUVOMChOaB2VlmclV17ZjFAQH1y5nr5uu96Dzgs6QLvU+wkWg1jUYK
+VObF0Gy6Z8Ba9u/IUqnDy6YlExs31bH2+Z+S4jPj2TmmQXb+MvU0a20EOdV3Rnb
Eh9II/pTorDbnIqfrltP4ZHy8aFXXvPnMas9MRAObbnEwsQJXARZG/f+btf1uqS8
facvDiPHCAxV77rQ0qgGf5P8XfwNhmZyvqQDK1HvG9BBvQLKnFcebJwO9DS8oj9M
Ha8RtWUWDWZW1f/nZLmuDS0MGXrkQiuBJ/rkBZS6RI+kCtREcKBrpJ5gcl3HlYjW
bHL13WDDanI/iwFh6LtyJH0qZLeup2/WDHY2vhBspd2qTo3D6aoSgU+fCucG2Aa2
cC9r/BhW2YDg0+n7ZJtCYhw0gzsaEytPU4NuoUxNvvlX8GHGC8ayMeSXuGA3bar9
hwcpLCk9kCDoufJlPkldeXnuhv4Ar967jmhpIBDeG2M0tyMj/Ktz1Bjyw9CTyaJ8
xMw/2NYpJeUTXXIYQazJeCO5ZG8hL3KCnzBCrdcLL70wzWCVOaVN1kooyiOnws9l
Y4GtYqx7GxasCBSeOnJMMHPxLv0g9TVH8VqVPX0GM6CPkVOoUAvBhXYdwX0lk6cc
yct78DqLzkIc11Dz1t27H0Lftckqlj0qVryd3pYHicdhOi+CsmsyzaO4x0EHgGrw
7jPRAA6HRL8Lb3TuXJsg+v3W50uHWlAf0l9w33qmJmNfnNtd4VUC9tKtz+mf9N6B
9bsyPsnudCBqEYqcbb9KHZ4xh1cLYoJL3ZG2RfFbUsGiYJO+44X73YVksp0/ofG+
dcjRWue2qg7DOOu84blBByJIjNDsGJx0QRibMoRRqo8G5y8DUS7hBH+bGaX7DU0C
ktWiLDoarp+BgfqnD7MuHT59Odr3h6jMxLlmPDtadEbXstPeJvzG0YtOn7ojqC8v
ULbamQXke3WP++zJpJCoJXndEnR8AGkHj9/bERYK60uA7TU96ry5jnwwCGSm5ilv
GJazZdPuWuuUBdsGw7VFRVpxDF3hSIrmljrZa0qnXMnx7rTyt+ADF7fcCQuTHo0x
/j5/s4vinFNaQ3HXOhfqKqekOcp+A+IevfOdbAKJkGi6NTM0HiPeH3RXhBhLN1YA
HBholhG5HOKZY6CfKz7OWik1Lqb8Znk7kl7tMlOvjXgZnQDTVljMpIlMXOu/JqvE
TzRUbKHD6YlbSibFY8xyEIe+wPwiu68vakjRj0alx7vWo1cU4//AIzc++sHS2Qbw
XIf9vUNX37W8DuF1WlIW6lzexvdr9feYYnDq6w1U3esezzrfUOlpmZDUgJE+wiUT
HbnDI6DKaeplerJQqNshrGPfXwJ/T4RgbbqorcwftKlrnwh5yLX4Pv2Nuw0bKepJ
9bzx+V75OjQ9wl1mxCblI7DxX7ktBtZTyibJ3XZ/WXgL8jQdBusDidvM0v1VprzL
QYPi/45uz1U8tWyxqzP3bIb6OCusLWqbFq1TAbJRQEWBJxGMuuaSTGGg5ypHllyp
ivIEq+F6+ahgjiEf+K/2p+I4pPzn6RJVrSuqJG+bZUyKl3tSqBkEwhUKvjzOcJfC
kv8w4G4585K7jCSm41/17ThP1N011F9vcj7v1CBqmFxefqedFMp908vMzx3VIS5u
EBzy3WCmf5P5zEzMhxsnnijazjIIGYX5AWwn8ss70NM6vwWayBcEcAIXoMe+zvie
hrjthz9bNZEtEhrZWeN7H6KazC+cBefJcrLnP8GcPBSzQqsMdY71FCPisEYuRLOS
NpnDnuuO+rJt0L044IZFZXT4oWyMQclFYpraaHKnInjdoR2EXNaLbbdMzM1iHTjp
kb3iXhpMezF09uDI6tKv+lztuVIKkt34tAjMrpmuYvvJ430Hpl9KoWp1JguvCSUs
jeVwfIIOrb79LWkSJzg8c2GlbFXsn9tlu8vzW3cQTPz20lQbydL5+O8A43WyQ1AB
dVIkWIgryQ7X4cynZxUT3x0KzOo+Ow04dmmJeH++/5N82mY8DzspQt8SPx6yvQkN
/t3nkfWgLmzMjG0LDVVpBmdq62jNIZSWJN8kbaWWalzU2+6LWl56vi4rnZFDIpCs
mfk+5fzZvo1BxsLaw2W3oPUOin3X0CAksIJT6wEZqDKQFrpsT7VWn1NyIVlz0Ga/
btAurgT7Akuhh/OLx3ZnFUHWH953/10v7oRqq9DiMXbxL/GDAfpOM4FxOdjmfi38
UMoYmq6NdpQO565UXn3R6X91IPJ2BNUeGCTh9V1SfJLZ/cEkn92VvE9eklkkW23X
52pmnzPZXwMyo6Ta8aTYYyxtaJBXW3YXNqwDXbrgtvyJsFTPiDeZ10+DYr4on8OW
kwXfb8W9pQdM5JBL2TEBzd3oetcu4GJwzle7GVFmXyH623b2yAgmF/9lrLAjsOxT
m4xyuquthPuEOwvC/OLHyF6sfM1DReECZqe9Ws8mdAtw/PHsiVWciYosb64SdVZz
im5/XQfZbiPu4ouvXGIUtJwwW9GGLHG+8xM8ZmW8WoHXbhE8OkeornjYgpPieTs/
QANa7m1IlaHuECu5Kqv5j3YybwOkEC29zm0aEaIw/d2rW5UPUaKPVmVkUCTRlCqU
E2vZV9oMrXpCMMsJTTLxVH3quC0PUSoY0/TE12OXWqWYLGVULYGbS9hmP89JPu/y
WcT4TVpMfbjMATJoq6NxJO1B3En4J/0Hv7WbHnxPVdpbFutTTcaCTo2G1SKnsTV+
og/syuhZcibU8mpRnQdpM+/bpWd3k0XSocAhl8eUig4tmCR+9k1R8jTpqzHbcCpJ
9tTJotjboXBcScqA3Q7+54Z99O8PcPzsozqL2AJwZe4sexCWA4HbFOnPAGHTPz8w
4O+ue+dQ5/R6IVFawMJm8332NSHiywdUhTh1ZXwE9o7wqf5L7g2nu6IY1PcQXJPe
uyxVBVID96iVWKVQA+JhX2abrS3J4XYEoTo6N+sgNnO9UL/pcoe8JcktXhmmI6OK
nvXlIznqKHEJlHGPASi7CqkmuI4bOIGmcHwyCXGLKeHcWQvpKIYpaMLrUS8LV0R6
go6chpRmIN2tKLahn8rIwgpYUCvg1PGxlLwSqvTMq4ef/TJmiZJEPi6taxOymJ6s
R1chqPiHhmJy/9PaPx4Fq7i5ctq82K4m8Eav2OBWRlLeFtcGlQvGswseJf8sOUgy
oCROvPJ8Ypfuz0MSTKVdOEnGMeWo+qE7pPaDKLFji6HePEspftgpth3LxssbVxlA
s9Aq+q6snrk55U/mnlZ5Npk1ZXjfS+l6P+QFoLsxjD4D0MmxnSHYz/T6DQzEkktv
gtvtChVZhK/8geOH6t895AHT1EenM7fV8TU8cYqq/9bLtEFwdtxL69dx92ukjKKl
Aa1TiKm4f1c2UbquH6xnVqny4SSMRJiNFLuODe5jprosFKKyQoQGOTzhu0oQILWT
KRuH0ilw5TFXSzMRGypbB/KqLoD6PiZF9cRguy4lMspCpc9iqY7hqI7lddSl81Gq
Qacf4zPr+P3qL6XrMa/gK3wcd5+tzfXHHQOEGW++s+ubLWc9zcMMhdCl4u001i3s
sECjj6OT1lqhAmv2EDPIhAojzmAXw9phpWTASH7UY9DDDt1yHQU1hfjks8oPk9Lp
GCDlQdWN/hwmXdaH2cFw9c7xcLQFEjtBSfoWarSysV2XbPR6OVt8179rRhWessnl
nl9bWosyMebQCG7fE4RbbNeG1gqU1tP8GJziXgcoJMQzX24f/STDme4v2VhLYdF0
VN5NrooTizk8/KCFuNKXJ+Vtd+4D1j+2SYrCgmNPjrk2XcvjUOwEKYQM0l6awQBw
6l6WbVG6I0RFIXMSpGFt+VuuLES76KnaL6SA+YQg7r8bsQYUSsSc5cAQQJJR+/bO
g7ZQmABB4PtW9mtBkoJYeFrnqaScvACZi5G4yNkmm5AGxWGf7US5N0ohT5ZaEjpl
sqQa8e4TyV1XiWkuzwl6KrDe0B3Z1GdB1eA7a7MX8sSCW3LX3GyPNeu2mga2fSz9
D8RJAi8ZmD84uxF0QixgGchf41NGZi/X77AbLK26l155CFVYE//y+R0XQ5XE9rqD
ER94C/hKJ9EErWzevRwE0exECI34V7l/PpMYIaNh3dwgMmdGTwqnS9Noj6S8MmCx
i69nFGcTjxkvg9jCW/ffIgh2bA073r9PwcU11bzcv1WEwaczuVS/JYrwrZx8sqp5
QhsD3DNb8z5fSyO+Y9N4UI2YnPuzOwN4P2nrstpOnKneGr69Iq4JcXcsv1kD5wqO
oLrujrf48+O4G1XFKUwlVxGNtfU3sYHzEkuENYGWsVw6hfBNuDw/QmD88YG+dcx2
sIkKoE8jbD96J7j0YjUgoLnpCWWOKdYHhqpf94dUO9jGmic7u1E8Kwz9gDcFO1wj
b5eS+YrQHX8CoapvIqyh3Mb4PJnnmk/2jyhq8tQg7MZ+HqhOdn26D7P/wON3t+XV
AdGdV/X0G9B8CRpAJ59v8x1dw8ZQjnA1B+C83zRmFXrr03tmDO7i2+J9oSCnELeS
tf6puQLiGjTGGs9p8B1mrq4L9FCowidAO2XwVBawYKtoYdPsa5MbIw2q1aA2P/ty
FfPk76BAE5jCAvtnb+SX0QXrkzD50NGLfG1x01u4S/85rUMuI7qUylR+PEIfNJh/
WnGZSabBksyIXF9CO/knurb2sffwQO95cklVPkr/gdgqfi2zMbtSiGjgPDFas3Kd
MyHdp7ED9DzSz0levEV2bhrI2+syqsM4oaB2IktIY0psuWsL4hNPUcHhH0uAAInh
v6PAIpz3M3XWOVrX9m1X7wAW+pfbLIkV0UmZiaLKuoNPbsXINJDEG8jcaIelpA1z
KdhQoxQz9+xyub0nnuYe+hqkpkn7iYllDlpQuRXhsjeoi76+XaQh0ygoERVqw0tm
FEZez199y4IKKaXneIpwVABbkAV8ZEG7uI5bBpw75RMUSv4OszrpXlT5xGia91/P
eHtyRJ21ccl4+ygYLPsh6WwXzx0UMbn8ONJ2EcGBJ9zW0EdQGPYZC/OoTeV8O3+I
7HpgtMHPVZ87UlsutTj37uFRRnrBhGcHOVl9MGFx3MFolm+fKfANZCKOQ/cgTlhP
EdowR+QVfOYjNjdgSqhVYReXzNaWgCdCGTSQTyntgnr1F2EbF5SQTrofNEJVNFxM
PjyPruZVrDnB6WxyjL2b2zvnEm2p6m4QkauXcAYaHe1m1eHuQsEpcB1zi8kZShDl
lqPhMQnplDhWs7KWSqA1AnZ1ZDpwOpFxVhAy99Pnz853BQ4k2VwSk+RdN3+7cjJ9
/kICG2hPdUw9CRd9yZo4r4wtBsg7lEp+qO3JDDQlDTLvamFXv6o0yN+uxDjuoO7J
0NO5pmlEsI9Uxwmx0YLpVJoCspjhe9CoVOdNVmqJUr88Sn5+LLvBWfegY035xWKw
ps5rJ8pROuX5eR0+8XHBarDwE0NXYhSFJa/kyHqkRKEgf3f49+J+pbD/iTV8iNXn
buxYFiCU5AjPC6jP0U3jQOdc9YaetVAccTcbsQd010TJVSrkHMp3TmuTRdUpUcMk
GO1JDZT/pcBTo9BaB0t4A7eLLaOeYgKkBCFzHHQMwRfsrUq36wrYDplzTdY1LYCa
IMVclKZbn4APvHIgWsFVlGlIXEhAW1PXGcx+XXcuwQxtz2sbffs4cOJCdhsGuSpz
IZK/tUkEmZutxQHJVr0DxKSV3nkZYRKblrshikF0T7sm+m8jFkfz77ZhxEsv9bF4
4PAqD1q7wCdzRJAB8kU7e+HBlZwfZCPdQ4Y9BYCQB/ZRUAHOPMPcaDWqt7coa/2R
u4XFLgDBFGIQNSsfbj6uin/tGnKa+0bjEPqHvkVutL/WdDvD8MPmKmE3EkAcgJEl
8QzNargB0NKBJcHRZgxPz+LCAxKRrXT2ENIZP29cClG1bQhkIfaVA9iBruFay7j1
zziWBphYSwMtPPFcRmfoOKmLeUuiSDkfNR03G5QHDfO3FFxIv7FAYBuib6cB3ugQ
bpJkqM18pXHjYCz12aQqTyrVGKii9ECNRnBSoTV1ama31YLD/qBgyeDe1zF7L4aP
UUMI6U8xUFPSAa+tn4VNuGBW3f/okhP7NZqJzAn5PT4XatrDGQFd345cag1GIGYm
mpfFTYzl2diE5i92uRV5MV6ot8xXEJIGiFZ3CfzUtdwToTO5ML+AjjIWvzDIzQQd
7h3o+tkRggjn+Xv9VTjem5o2ORPT4d+QHzd+XvlYXFZiSr/scp9xuKdSQh27s5if
OsuHMXclMR55t3VDzLEZDAS2DCc3pd79zFZ/kz629sR8GkAlj/A9zsRpKfZKTlZh
iV7h7ac/pCNCMNo/SWI32d5wUpf8mINgLETfThM+ErQfaLlCz1nhO/ILzw7+7/Z7
23j/mWxDmdBnxON/qmTxORyQ/jdIZokJxe38ma/xnwpMMHxBPmrF/etiTarZAROH
uGRTgWgbh6IsWwDzeBt/yZ6Uu3ZXc6cPsrd696Ae0DLIksb+PbJzzhJPERofLmnt
9cAqsIAtVJBZqKEMAmbrVimfCpkzl3WDk3zhTTF+TsQmlUbvgBnc2odtSBEZTexm
UNiL8BFutDcStNHHBC6AQYiZlaQ5YQi2KWKW94BfECccx9gBHnrhcfIq1eR/z5AV
BzOHXNI6ToyM0WMb4rjJOUkIuL5HO+J0uN8whLMbLTWtNc4BKgARyO6XJVHqW4tC
1VEtbRAmsxHE0pAYE6QoGtHHiGsBjHvnVh6Yjmje1/6F/BwkbYPGzbwn4TXvv7pt
VQLoGe9ybzDSqpW/MFPGWNAOQUiXmIliwIRIJ/mI1TSbM+9Dro32CYhUijv7Tfs3
rNIAsL3JZBf5Wz2bfyvbQOJdoRI3T7C3mfxkHpC60Ed4piiNE9LkO5pjbBmloyx9
2B4MkASU+XDLxYDviRdICA==
--pragma protect end_data_block
--pragma protect digest_block
/DZE2C5cbuV7k/uL4XPY9P5DWYE=
--pragma protect end_digest_block
--pragma protect end_protected
