-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
D8KPB5hFrEpR0ttf6da2d8c+cQo1iETmWD8DZ+kSQJs848BOMaUwjtfTqrXqGTOF
Dhdis3Dw/tNOeqU2rBTDbiLHpLbPmZiMG5zhSnApSp0MDt4xxXb97FtH3BdYCw0E
zRhPWFZG+grl/TMsMThdGEOY8BkpIHGZXQRiayjNdHdrKqokNvvIvw==
--pragma protect end_key_block
--pragma protect digest_block
MwoKxxBe5X3qRJEU424J7diTYZY=
--pragma protect end_digest_block
--pragma protect data_block
1YipOb5X1xEL3m8uTMCxtwKLhiPYmD96CcecM4uMapJY8z3dGZ/9UXdV86/00QrC
Q/rabNSyIwXLd85yyC5VFzAXem6w8jvpMYL9Z1gNXtK4dji+VKYqjMAS5tWjVGLO
wUqKQhtqLGI8n6usQFDEP5IIINmpMS4wMyWd8CzBMaV7nGq3r0LlidGrd+EiBj7c
njniySFjkNo+yRCPpOMdlg9JbGkLJHW0U1i+Y9YjThN4vEk18LuMAVzylxyHsyc3
8eZaGYgc96Q7Fwgu5mYbXhccokbppNZPVOGHhW8s4WtH/9EBbC5DCvKZ9xLsyOmj
Va7uYm9oG6J3F55A0ug/YDMqfkADqIsiN8MdszRAhwtstdV7q9pVE+bNlxu0z/Zy
1GiLVuI3XJYlKG4QiZ2Bsc1SuE2W6uSwK6/L1/I1/J70I2p8Q9o3HsRhWdSmPOBA
XdGg+LZ2EBAXy9VkFYzKmBWSk7Nhg0vzByRhTGGagQcNoMo0KGyUlx9TAI0Lt5/z
sf/aB2SRTparLEwULjW1Bb134IopXXMHEUJoMNEPArD12UH29L975RbVHokZ4NcV
MXuGMXscNeCELGQZEPTFP8K4+ELOJb3r2VccFcqMsJAsq8FE+HN1FQyWFwpvWNmQ
9/cplwmdi09B/U3je2+cZK/LDB5v1daa1cqchaL7gMhhhA+T+khfa/KELs1YWVXh
YIaXeNPZvqhyTziaGSYPFM4uN9Wyim8iN7I98CLjmNllAD6KmusDdhyGT60YPxrL
I8nmqG0qI9t3YUzyso01bcvY7Nsa7mvzEDBzGUbnYUPsxjyfM4oS6siwyctj6CBh
+zGeDdIUKo3/WmJHzvohpuHJJS2QVA/CaYQMYH8ICvJkOMM5hgTkhsfLz6tNwoAC
SNOdBsoeFhC0WBlVxMGbCPbuKkf4dDvhXkVwHZq9gL5xf+1rV1kuDfcMp3CwTbKX
uAKDjWvXTspN/MWiCrCy9jPD5Ga5FIb4VUMlLsWhcn2qAqWg+nEjIoVycNPoQTEa
KdcKXDLtsZ6SOJd+IPNwI29/4+vTKD3VDV9kz1+EgXZ1GVQ7sOBLnpc8tYg3OjZX
pasGYwtZ8R6RKkRhvtx+ljxNS0F+8Ky2nsSclj5EVplS2oaGADdQmpHl5VMBHPrE
6EG7qF8PLa+aZpNXZckAcqdqFNMmu9yReiwepbN3I3o4r41mSsPNVrPa3+w+iy1L
af0qDn8LD+HYeddcgjQ4kZVKazFrSqZiuPCiuw7S5Iy+dWOKd4GBZ2CQVPomr4R+
jH78lCx6DGNTSQ22tYyaNMVgg17sefXn/XzNJ/N9JRNsCkPTjCPF1yXpPrPQZx1v
7qYLzjxVbfmvIWFCHdw19/fMAEh5VqnKzzVwBt5cBQD7PzdC/cTpilHpg8c+8EjC
WUsSt3ByYzPPgLdU0pTYEPfww8RElG8C3FcrBcgcoWfA+KznXBjzCsVyImz99h+z
0T24JXk8sWVCHlAOepUCuKgRCheE+FH2J31uVJYcwFLIkCk0i0EmJLmbE4/P6mDN
qA0TUJCybdjuQ/Pb+sSYTnru8xW7dZ6ZprSoXtr+rz1wAgC23p9PjTfvXWeo1phG
ABbF9A1lv8kZhPMTDJRvRAWSTCu3WKVOmAcDKL/7R8xjqhnesSLkOJcbKg4pZa2n
SWKSR9YDFO/h0G6oTwq1dKHK44Gq7Ti/vfCW8Jc27/qUbWMynVoKhNAcxlMhtINb
XGeMuR/jWm9K2Ht2Hb/EVz84f6nyqG2Vv0Uv8Zu6GCkWcsVOpEvCz0cRwBTEuSif
yVa1i1TMq7VijG82ykqSuHi4nSu9zCOkRhlaS3Yw4qOsmnTqq85rxCoomL2+2iZS
1OHL0hdS2nF4bMH1bmG0eqe9o//91oI8EHPYZrt0Iw+jZYrZat7J5X38Jyn+L/QC
maiPYwQ3BY3aU2PPcktHH8mLaK2HXWBDCIsmTzyNoSJgCOeuWOzCPsSR63MP2q5/
i8FF42LOefTt2HVTnJ+KrwXPTOnM3LX20XLkaVeUWub1Ag5YnaDtLdwQIToVD+Kv
TympW8UVbui2L7qDzgHTdZJ9khc+VaPuEdmJhGfFvpL2BY5iVaX+5pIpk0fAXcVp
nAy1fmOB1JKweuaNWmjs872ikd2ZCHuBMU+bwwSvq/JP+ybp4OYacDYwHWE1gdxj
BIj32XUjs7+2kE7rKX2X3O3WdvapKocgrSUcqt7PHovZ29ONWOH2i3cXHmq723wH
AShTLt7jQOgVxN6u0p2LHeyOrxWEbHYCgIMSmUKBtMh3NQ5ruwoVQhPgGSFY1/gM
xWobq1pjrcffhrv4tvW/PcUwzD7W6SkQhp4KrQhgvQ0xt1R4J6d+FxQLzBJXK65+
kMTbB47CbpFZYkPHa++xkT0IbQu/d8TlmlwiblvzIcAfpCLse9aww0Tvjq8izvN1
p8uN86noO+/9EN2kq46V1+sRrHnUcsgyOjy/k4DYTLiHeKCXWdF9jd3FOKeE/u3+
8/9Hu054s0PhJkxpxImn3nvE927NvC3Pwqsr2IWNo+k0O+1IOzXY8Ix6uBTLHAdK
/93bX1GWbjQt48cK4KF/5UbFpAiiKzkBo2/LOTcLK0fzD/1o8FoSvioWpPDsuO5/
6FVlYGy0+n8FlyqvU59t/Nd45HPIV3j5DQ1n2BM8GXLypKYRj7CtbIiHz1bh1EBC
ZMW6xRXzc7lfkWb1b/BGQUpCgfgeUyI7WYx4VWy9ITSMY7YyIxdBRNPR0a0ROIJu
y7JpR6iwJm0ZPCKYuQWcMdQ4Tijve7/XGg3nYJNXMMQ60STwrtHM2P4oV3d/8y+D
p15cOqfys8ThwpNC6JAUprUO/bI/lU69v6hnbw0Ye/ZHHAPZAlL7Ti2p4dPZDbkl
Jiefq5fMBt6+rKVhsfRzF3Oy8ITDZuvK++5laDLpyk3YZ09M1wL2J0clsitwoMzA
j3rgbADt2Pwy0rdsYDh5q8LclmO6R1mcoyHVjmNhWbYnxUfrbcpBMofnAhLpSGyX
4Hguf7lYSn0liXVQvcOteBp5OyBYF/9eF9ZxkhjTZkOChC3pn5f4GEzEDoIKM+1e
SdjEEXuqi6rz17m21Zgn1pRmzCN7/bCJ1lrk/1oLXdpxOyHyPx3flxVUAaVwJc1O
S2B/U9ir5g97tn9i63h9r13Kwkoym3xJhLIWdW8vX39yLKsycT8+MCN8rdIK5w6D
NFGUL/fAMqtLoNojFk1WKuU61McHxx8Vke+9Zpkoydqb6W0jUFUoF4QZB0vFf0U1
5zKm9cRs67f6NP06em8tmEsHzCUwZm3E9aGTFL7dhdRVrDHusbm7b9OjgS7ODH8n
Hoyz2RL/0OUDjzzXP4uP2PiTPzs9RqLY5o8wWL4vt1fmBSSO/H2Q3a4+61ffcLmP
JnClhcRViPjtE+u8HlBDweTOagy101LGoqnamS3M3DwN6Y+Nl6U4Uh1bemzt0oaG
R68TIqnEaRrbgrf8mBK5yxjKkAw0DQfpncHxGfmuH8El/72no14aC7tNO8kpUubJ
fQo1o9OyOKXUeCG2MPMkoma0DO9zhnB6yKwojTHqexTxcNLPPUqr6TU49XbfPZuT
BQ/8ad/QA29r2uOBDXUbQuqKCAAE3CPxBCgYHjTWx9JIVfsEM+4+7B11e/h4SrHn
V59RHY1CvuRgnQnoqkKO+4dPOl0mosrDhjEiIZGLdjp4k6UXPz1jBa9CY70AR+fz
4Q7o+VTTI8zucbktiqRkWJ0qaT34IA5NHmmKhruIk/YeapRV0olaywq8EoErPI+c
kOKkiTKbBj4UZIbWk9+4m1kJc90SJfCrGckG9TkJDb9w0sDEibF3kFZt3KM25bLJ
DOYax7zKPDSViSRRfe+I+HugbImZD/4rsJob4T7L733QZCzscFKBQdsWojYsC5vD
PShdaiT4sqTjXSWrhQlWAln1JMhLxorq6p+bxwWmNy6Oj2zRfmSMtgvO+BI/1MUk
zCI5D/8q+3yYsBDrMMqzvITGYIMkDo5icpJYmHdAeKf4cftr0ACZPSfuIQVQO9a6
B2pOibJMek4IyjeDPR5GDxd2bU9yIa+Ev0njYaULFq1DIsyygTUQW1WHpj9ybP/x
DQACCg7snj32HYXd9Hkv9m/Fijqyy+L/dMgQbh1i8I0sFCeI9rLC5MALGD3ez3Uy
nvQlsESYNeyD3C+LaMS3a9s1q6mOeH9PGMQYcrA1KTcW+/giUmgxD/EAezRgeBQF
l5WvizdKcd5zSd2iM1TeiLJn8CGwlpBymppckIHCCGl0bS5zLNHK+PeLmRoh3JHN
4Y0MyCiJKWGEPxBLBRSCp3dZnk4uuWpUnvlF7yK3kqQS382M+ourqfCBFrSY8Y0E
FjkW0U2OBIoOyL+KJUcQ1k+ipmfzYKFaNEOiNoZbYH9ziYZcEY2xs7PI1P9IZ39b
sPCOChbssJIJVa+TLRAvtRQKYPPpKbuJxa69u2IbBxEH5JXk+RLIXmdrxBbPwEAw
tytxrY4tiU/HaTKvspkVXFeHVSJ5Uo6ZXT9xGrrm8IXav5dg9afv7TXceBfuH94q
arcYp95pj+HLO2ghV4U8Y5H0xkDqqXeYh9fDYb26Y92JdRb/Nj1hIyguZQkiYL7c
k6FVnkWxr8i9cZzMVtwTEJ4n9dRqaps87QPfb3fWjSlyNaribdf4CEamoXlFhBIc
uq4UcUwEEQbzyBihI5vnU2HmhCSmPlv9tDfvAzGJx/AnRRdjhqKFBIukQp6ZuQTH
2Mkl4bC0lwl2FF//2hNf/HMi13GoovKalTIEn/yASfoH7Up8ulaRZDhfcOny5GN8
upkkatKRxIiJ2/98hdK9cYPrNYiHCV+K2k+giAMWjWDtxR30p2Am9SFYqfXUpzV2
I4hviBmc1vnTkb+gMzzXU4GTdjhCTahmzBlAB6bTxRSJhPdPLlpMPXnxVhkqn9vf
jL/y80ycC+UhVfHPmlLyEUXJRA8syT31TTIQjUcFfPB6s6Ce7+DLWFJlKpKUeUQq
C7aCmsscM1UakyoKn9oKPRmrWcoiPHsPsQd9HGr3/gH0hLHUidaBHkG/wj0OHqfW
DkxJbrtPMzYkHhTWddNBDl7LMsx8FE4koA8aHbgwK4aJJtzJ4QWmK5mOYRElERG3
BiTK4x1vDebfkGkzD/aDhQ3f0FXiAEhpd7KqyGQJWV295ZGHxkECC3dkIkRreBuF
HUTD0oXd0sEE9U/eDUHtvpvyb32D6gHLphAQb2VK8UgEQWC0a1uTN6pyj1u3cDtO
AMPOBEuDLKZzn9op33P1YJwOWA+TpRVQvSHowrJ/8E+SQyFaSYhlXJ1EZDA+UkEg
/ESlzAc+ReymWKoXSsX3zWaeGgOSZi/nqHPRY6/UkeQ1FAU3KHFt99jzR8exZorx
PPWzooikUiQN3zPJwQLN01n9uebvnpGfzL3rXlFpTxyIGnoMXghYHi23P1CLA2OH
VgCmDr8bxLWMPNpaBbUnAWtHVyk0/AfPt5D5IPqF+sfPoYkZ73fyEX1bN44Oha+5
WWPBJlK6ZeMfv5REA7o9WClQkgyVgzzD8UySwh73cL95sDJDueMO2dJQ5EmW3N/X
2DRbd3bTUqs5Z/HXM67N4+/O3TSiDUu39STvaPMVrqi0fHy57QaLy1Ouxre3ewA3
AAIfbKABX8cj7t7d3zQkLnBHPBPNz0WaOfnWLBka4Mbfv6kubJI5wirt+Xn9ATFa
4DVDeJQQDgCaty4oMwvbp3hcGDyJtbO/0cirGoKy/u2fKPKTjzIMydF8nEd2oaMK
TC3cqjg1bbR5sWJvxGYcArIBzwd28NE48lnKbh7SmYIMf9W37awvtPpf19U2uKzC
WHJs7rOAjfJU95EIL1bxdcdnpWU90CaANvF0fGkqFG6IiQ/70qzHOQFcsPDnmHEA
Uw+6nolGuWyUt0kzg60j5wMKMX5RoX49VJHGAH8ZLzLg7C3ThiGQ0YwgUSaUzAex
LDysY2uJOQhIAThsWTcbQZLaoQPFVdJJinMLczAXxGAZWpux/klfq1G2B/C5B/68
SRaWE6fVdlygTGTRmjii35R/vr4fmdNoH8wERBAAMrj9OZNYb4ElxB/ySvAnGGIt
0URhrTP4QXavHRJzvQ3LO4FFt8z13P+gzolHz6xgjXth22Dbo8QWisCsIaPZYmT+
pARHXsx82713BOCAMHlc3eko8b8GHaRv2QSSDaJmix8=
--pragma protect end_data_block
--pragma protect digest_block
8tT0ZGRNzGKGq8Oe6YCSPJouT4M=
--pragma protect end_digest_block
--pragma protect end_protected
