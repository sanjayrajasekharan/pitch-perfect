-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
v5UyAZ6GlHAUq04F9c7exokgOypURtpBV2UXTqadSQSchf+hn06+B7N8oH/DBNZc
ivqEfXjV/oRB9V50cVxAVORE7jV3/e09cqi3Q3n7y6F3JS+MY1FaDSjarsI3xKdY
57td00mVv7CaUZgNKJ3FPs/HcQLFbCqHGPA84NH1Buc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1680)
`protect data_block
R+teyHqU31ZnEfzLSvoKdftggzT181DRuSCQNvr5sHpaNIbY+flAS69Y09MbZ1XR
cTJt5HilU0xINCsRgiCgr+HTKbmx+blKsZCIOZQtVENh7PrfeZvjhIs3GRLSbq3O
MGaI2bpr2exnijOM7fhWY8BXhDVfgqbO2cgvqBnMNcte4hHSC3hfIexZ65siNYGP
zgCFWwqaQijQAgdv97Y8GrPgbqlNF5O6122Nbp2SqGR1zWTpn2BrU8f2qsf91vjT
Rbed+z0bU8S90sQn0XTi4MZpswEgeTd7TBXyECr6zZpuOK/iKxqGta6siAFgBjLh
d/o/lC14bUmFUkvnRtVhzCtaNO4H+9jwlwLt7gvFZuC7AKTZmsdJ8r8cMZu6evku
JSm6iFsy6z9lMqY/ITUTv2qN6r8iMNUFYoe5ZgN9O9kLx6CePeqHr89UI+JsyyHO
bKyFXrz9jxbirWvvBGq4vp7lMeqjpkcLJPEUhbFjtJE3EPMnJutS7JCPmxBkHWxn
U93A4BZrnl3I2zk6cZCypu98wJket8CbuUSdWuZDA/K/M4qKrJNTf4yY2EcMnEAH
sPQjoW4f3PeikiQyi8NvGTYlKtfdS2jqbT7Mzhe4lbzAd9NEkHX8+nKBQK5v+OyN
lR5QIV9kjifXCrxQRvBEqUttowZGithjw4ltfky00ZA/6z/S5H9sNYJomKa4qsmD
g4xygJvfRpMi3bLQclZU7Hh8PRLIdLybfuMt/bzenscfzFJcgkdt6u+Ao4h7ENhM
cYo7PlGvIeDTkqxTVxcz4fMUvIJHWCugpaFKtOL9oog4Hwue00jbObSTUtyKvwVD
OQrRB10abuyLzNXIAJIvZVmc9HAxDjN4PBj9cf84UxkXspm7WbdAziJl53D2J4F4
lckeKprP7rhtcoPmMp24CJHEJeZThVO+cq9FVMkg6JQRyYa2AHDAzcxfdnysEMQ+
IrL9GR4hyehdtGQbrkjo5CkgjuuGcV2cghA+0Gcf08dxHGV9vx5IUBQv3C2J0ki8
fu8cgByw8wm38uIXgbqqva5dNVDt2nl2E+AYNJe7rAXGkL+UKoC4vmuhupCxnN8D
txfx8zRturwLz1g+vAGyU/YAJQdK6ue+m0MRrIUIqk+XYoXnuY1UxFK+efoVQFmh
Pm2QYeAiXEC+uYV4t4g8nlkE416e69rZLg0uXVWX6LEZRjRr8ETEjjNX0xZtNYZd
JYwTiVb31tV7pnf2S98Iif5tRk6/a4OYiA+i30wHJd3QxMzvE/fhxyZTmLxv4wlm
FOTXJU9bh+JrObIwtpqZ2f2xzKab+11Dsc3XwCFx9e1pfXtVhbIu7D/Hinsp3u61
6VfLjh3DFthKaskOOGzcY+8naHF4J+4zouhajTO337izJjbkiFng3/V4Jm1KqW1M
WU2P6XBzeuzpmjPUr7AMrgUzn/7hjEAp2zk6TCbzWZke/cRDbabzuMvIXe5xbh6T
OZvjafWv+RON+Jp+sw+EBO+hTDTJiJdYrbuBJXFdAh8QU6kmoz8CWXUhrnHoJk6w
9PTZ/p2oY1WiOmdFCMpzxfun7bJ4rtFQ6L6rzbsFOy+JgYyJwmiupzmOHz2vIrE/
RcK105LMCgycbojxH7japDwzrODaYVDvbJ2bnuwZgQtNne1hPUYYBs77IuZSVT9e
n94YbfqFBTjHHcq/nCIadqoKZNUVhA4LBsa6gqmbAXq5N8mik45IvsPMSqj1ZawD
TTGpP7RuNnb6mEnhl8XrGoLKgUeim89u6oXCRImkDFw4rk/AsdMPsvCFudgusd09
JUGSjt1ipwXycqQCIb2i76+A3H2tNMAeGlcCsdrpgtgZwl1+zhy7vqxkFJerj+7/
xNVU8iwn6JGCtvGHzF/OWRqzmSzPZc/yL/+f2IsGJNWItj6wLm3BbNs5wC19EJZl
vSXSOxEDVi12Up4uhgnUPm86d2Cr1buZuHPdToBYzW2b0tZEFGHElo54qXCczqji
r7tLJYqzBqs4/51DlKjNtS4/MNohDGmvo+Qpbxd2O9wdZhzuxXpI80ASv6xrRD0L
RUh4kkhAaeWqX5ATPGz3xj92OE3wGTIX31vMBshbYwzOIOd0s7+N9yiKZuhKhxAj
IIqj3iQPkZx2TShynS+Mua7VokehXuJqITnKMF+En5f0W7X8wUQu3U8e8/UDiqh7
kbdnBhc5IcpEBDBTCzhSRd3FZSq7Q50q09gDnsTqwTAyL9Yj00oTuWMeme/BKg6e
`protect end_protected
