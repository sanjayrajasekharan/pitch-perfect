-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
brvCEzhy/cu7/Ql5YNmJUSYzHENc4qaqJR7emdvcgKoKCtsCX4krWnuaHNrmpyqy
kU1nNSlMZ3dJNHangg6FDagk6gqWxyFPYRgaYZS47v0JrSMJC9/DbRYQPfQYvAgk
jHsYXsa77PN2j+JzwYPHV9W6bjuscsNK/gsOleNjqBljw3kKQWqAlA==
--pragma protect end_key_block
--pragma protect digest_block
+Khj7drLTCg4t4HgqnKFBTZ0SZ0=
--pragma protect end_digest_block
--pragma protect data_block
uOce3ln5ZB/bHeIkjhnW3xd61f2q/glA9KOKxl40Cv62+eM1MDeGCMg2M3GlutPY
mN/X+oJKqBlmAe5ahTnXg/sMAkY1pBdoEuUIp2Jnln5B2TOcpaH7YjPxJqc5oDVd
p1YaZoTuUr0v/nCg3VpWx/hNailFoOu3FnO4DF0/OUqFXqyALnPcPUAzrWipjmEG
RAz1625N+wQ9vpYoQz8ZhZHBJ0Q+P3zgM8YQH6Yv0fB5+rcI0gXdxMu6SxFJrwoI
1l1Tf5T1uifGla74Auew7oR9BpAnBtpLYV/PD/vpbF1eKsah34Y2DcsFQAkiR4cE
C1mKqUDXhlxIFo2HH04ii3teiWik5vri7dXAMuXfcdYhqPWwbGc/gv5U72SKxhNt
joNyUspCfGOBuAcvytR/aoD67eXtKwZDPQs5StkdHdhj84/zFikOX+m8hLUvmwZv
xrxSC8h4AQ7BbMHFvww6wmvyY/+EENkzgUferkpzRTsxuVvO5xrbQdCINWaVAqTH
hSWL2zcISK3RBieeWxEk1KUatc1AQnFRG+IJQDFvwQ/jOi8RhCzA/BRwH+T9N7rs
gJE4E1Hp8R3Xq/WkzH9fGZX5ijdSN2lbPmgJ2Qrd0K53Hpw9/3knxspDzlw3hV5K
0AWwmMJRTPU4UrNdg3bXf8ZEzd9JHslN6lzrZlZhI+PLC3wXQj9ifHnqM65TBqyB
neHsV4VRhrfgJlwqIWZ6iircAdek6/rMUwbCl+SdWtr8oWHyRYwcizks/lYNIpBv
sygGJMgzWs0bEPqHfqLqW7Mp3vA32FWKLheNofdQq/P9C6SZ14B7bTw5tNHWtwmX
tL9VBKehSKvHrNELRTKzJzzJBer9JEgRXj2pqt/8uq3dXXchutlzZJ9CWS5MivYM
ygKeif2l2n12IfwM8iEMCHvKKnerl0+x1ijdvs7qHCaxJd3wZJ6sKDMxw3QRhXAF
wi0F+IwlNyzzibOTOm3itwO7n/hn7dcVQJShku5mUGPLSkT9XtCG+T2ZzSKJmz22
ns67rQ7ZW4UTHlb9uZ5raO7c17dLHI/XQ+I6cvpdDtsZUC2vaoTe7eDsd/KSnanH
dYWOaPG5adMF42cPBlY2tLc+ozrrD49Pm6E2AqTY7F2yEda0ixDTSbcTWP0fpFvk
SdLyx6p+Qpv9v5jPiRT9fNc90zESwCbqNihjjVB+ZJkRhRAuG/NzX0U4prBGGlIK
CpSoWAPm1cnM/CQRL7UBvU0LskQ8mb4z+nAk/fDJVbagR5nzKrrt1vQUE3eXjo+H
qfBhUoZ71jwReMymwDlIXQy95ce9jvC5Yjw56YxtbVfH8vcINDTeB0mGBcXqRaD/
pIGaUp96wPRaSAh68VuFZjIEvbs62PXJab0ZMctZJXJ4Ov9xB8XTXFY5n5Mke974
FfUP5Wd8ZeopsLIqU9k/onhbMgvWPQaw/zVAcN81hJ6cS3igh30MZlKJyi94GXOu
8WmOrkDkuxTz+qvbWE3DUO76FOs2/S/tPJZv6vz0r+saexkLyvI+iCRJ/IDWLtdg
PDOiZQZJBUcu1V6NuJDJDfWcFNuhCux7uOnEkC28M8otwAeCT0Wc7yDXpDGJpFRs
lMwtVjUBZt5JBegewN+MEPgRTD/z1Ocug+N2bwnMHl8iy86Fg+1x+29OR7VOUVKk
KhQXMWAflRmx/kzuPPlDzIx6qEZsYwLRXrh2yGC7wEC7h3E2HmGggLjM8fXQcJm+
KJLu0Y2kBVDDiNZFWsiUOCidK4bk/Ks7YEw2VqfE6CwPrl1rMtiEwNSXGkEO0SAh
5b14WxIS84ZBOZ7NUC0ujVgCp8bmc4FxE7KeugNIUwMXa+revEOamnu2IWAxRDyX
afAvtYspETRHSqtmRb89pD8mpjF9aCfDNSySlcm2qeQK5YmJbt+jQRITF2VVia/a
WGFTyEWvsKu9+w3DZjiqrFMocdJFDC7VuzmI5V0GBC9ii0nPpVxfIwq9V5Fmy+R/
8DIvNktqsYw+bpWpsn942F9B4cg2fFoxnSmAPJsP79UKD+PAEYtN9/nTX2WnHQ6+
2Lw2yOFwEjACvvjnOb+nJjSG/XpNPmVPAu+T1QKRCPH8FtRSWHwzLi9A3ZQXL25y
2jTVvgQVP01zj2l0oC2WwShzmyJWpUQj4AGtHAboklVQzq5Q54TXyWqc8dmk6oxt
iiwM17ef3y4XlwMdnLpD4WSJnQA8IW7uDomoGeJzBTZYv0Y5mbAAd9tq9pYvC51r
pWkUdywS3m7MSzy+Hq/0lOl5S63JUmSPRDM3JmfCTGPRJIa7AfGKDD/AezzezHk4
AVyZQWB+PWx2zyIqbh1g07KP6bWLLiaKF1i4eci4fhg7Jn1udv6kNq+YztFjjahj
QOrmoV4uG7mA/4XkOs3RY+ROt7M5zx3JSjA9d5Aq+K/WDIiigSlrxDGlNBx09Ua1
4iUM8BBRPtEt0HVdPLiOVAHvl1qULQL3lXqyid1HEqRlqzkqSfol/SGFQRamzpL4
hEC8Nl/XJIHKRKlBBrifHflOqgPKBEStekcy4AHf/wY+Hc6LUhx/Rs65542LXRX7
ONPhuE8plFsBorwRL6PNi7ogZHcrpq55I57RBYVk1+dl+7V4d84lo4gmpP8BSL5Q
u6MHNEtz1CEXWSakwwVMCUI2xWFRod9CvItoo7u9AOWZZHAGbUU+Sg5i82yDX6kb
78Z1xG+gyg3JyfxzyfrY/I81EPb0ilVroc0qGR508Ou0L4YUloQ4c8q8skI5wjM9
cIXvFywuWlgyRXbhrgycOgM0bxPtbStUMhF+nJID0GfkVuaCkcauSHGVE8Ahg0bM
KNjk9ciuj9cyGkFPVLFonSfKqylMyg0m0bWSj71fOQ9VLAMVLE4QL/sFZAa5kXMW
Um2al9kXbGo+ZKN6pbVL6pRFrGZvklNMM+l6FYufjbXjuQhoL2lYI5z+Fw6cwvkV
rQ5IxemjLugiG2pseFz3GOy5yN8fFCK427mZeMajKp8/k+cCEFBmYVJSusJ3x3KK
qxPSIZze1M2vWKBu8GTVtieTscR5O9lSiipe5j6NHiWWUL/lb4s29MYCkNPzziQH
jz57IhTwmHsuAg5Ae1jWaQt2SfsUhnwMR+iBjFbdEpaTO4wfV6OO0BnpmGeNKdyk
jZ9O7FhYSTl/3gzbAjHoYIqaQP166FZwMsIc6ZaP4k3CsW/OPW6UFGVu7di6j7B0
9RJoMMTIgaQxHwcnwXfW31k9oU5rBHROkN9dLMYvTYSPcNPclqS0N7TOnYrDGeV1
ICTKIWBZHdq6ZWFaUc82FhxIdAdSswwCtAJcwDfphu2P1ezyXI5C2Svi8hpH/ekV
wYAlRS43TQYS9wuPo7sLT090LRgWdnsXB0oHpahQkE3tapcgK+/rEG5txUKqUDgZ
q+Mg+v+Et/FGM/4FI1MkWjuVEQmfyEBLzL+wC2Esz9HSLNtZxbbLDIBVvMGB/RGM
vz3zMzqy3BwEd+AYYoYyh/M/qIpzatgcXfPxMNZCYOjwawmWV6+EWjgLod72BWya
rqsTjgClFvCrLE3hGAmCNBK7ffmX06h+Hcw3KZY2C0h68iZ0kOKOgXgHiLpOhC61
IvxZza04nu+k+USdPQPNm+t06YLmxrIADmtUgPeqU70Dzcb58xWrx38qkcJKmapw
8o0m3o3ACwRRjTqQ/yFAt5lVbDSmsYmUqU1vytmaO4NgsZ3YABgJRpMAFpv14SYU
5/0OgAh9grnFWhv/UzqWH4+Pp0XOUM5ymp8JhsCBx3dCvgkxZWP9tjdZxYXyMPD7
3ThE5nAAXhb8Ubqypk8NldcGBfDkEt62YhMJlUwsQ8XoXH2Ao3nV7yYWdpzqvwjs
gmgACnSr5pkN+ZEo17RZD3695co7WCoDZshx03ap33VFCuh8cshFkV7aJbQvNTFC
KMlgTH8gLzl6OscdT/5AFEb/CZ5oahcNFU7h6V8weSbTFe4ZFxV3kKBbDppbpDrX
4kOSPbZy7kRSMB7P/tyrfZrwqLpo+CxL0e5Q3dvgqoM2YFAYHvRIyy8/NO6MmL+e
MByaDL0zX2lDOX0hTyZ6eZZa7o3jw+evvpdMQfdCZCoaA+TVdK9TETi6gxHaSoMn
YuGEplCoGepqfgj6z2seE2od/7uW0fA0fpVNHF/f9qkQk1IeuLvrQELmxtIrfrLO
1Ra+4e4jCWUA6gKh+MhYnoL8xjEmp4fZrXPFa6CUj3dooAPc86w/sgqExrE0siWb
zb/p25VuJ0wdeiT0Ob7QV7/gIXbo9pzDPGDXpQzLFsvHQckuRTv+Reo4ZWiIy8/K
k4xviJtGDZWm6vmWu8Mk3AwhzmMI+Hveoy5X738Uw/AZHSfoPImPkhAJyjavFOLm
XzsOmne5KCkuJSjHTr0R4AHD9JHddJPfhpTJgNk7OZ1Js37F08WQhYV+82WHQoEl
OFXbJ+JLVGcSrSuc4QDrkAPdgcbJtv4cVo21qK9cTI6LMu+2gcIWy+XnaRP4aDCY
CwIDeqNqGkptl1nm36w6EUzqQz1d7XRKWhQKz6k/fUShMSMS6qq3CDEita6f8N0T
kH6g6cvqLLIZF1ZCGH37UX3xdMokXDUJ3fgnwr0rQJ45Tfq1dIHxkO97gjYmySr1
EGxUeT5WnYPnafcVayOfSmMC0PaJEOJI4c+SObbgE+/tMvML94nkKkUan4gHzXhZ
rHiN2RK1GgMCQgCKsBM2BQ0YhotURiGFLJcn7+chb3umRDc90IxYIryOn8EPgG5n
1DAQHH2iPBdrGoYb9vxxOGiPOwusGz6LlGTCmKu9l2mRJsl92Lk+L4BqkEFz2VJH
ygU6bCz0ktAGnnTBQ2/1Mncrtz1HgbJCq58IzJu3ZGfFziL4iy2776jtHTXGUzCl
8OTDY6pEsJkLE4M/AO2F/ZBj099vDNO2uuUrnDeKoPyMRsvGys4VKqU2gAnMEpH9
oxyGbMjokeHwlPZ7M8mTZOOzyyNtAVCEsO6GG44f9ju5db0nnhEXx7jx21wMhB+1
xRAWd9TI2Mh7r1XmZInE3VUw9qCDQEuTa4Qzb16A92lVAeYlOrR39/XhZt0HxfiZ
AT449/ISroMQrw4KvbDSdMwULx87WCtwfhQP4LfmcAh64AKbRBjCAqnZ/0I44UTz
0ePGpvU1LyPIr3dD4jlOSO5tpa8YGVe5DZDUgOsvwovg39LP23ABJGGMOD/ydMA4
9iecNZmJpj38mA6hNA32ZtrO92CivHKVeB4lQvaRLtIdodVx2k8WJGL0gGIC0j5L
I9q45rBu0qihptisIiyUQayB2VUh3BxvqhGTKoOX4aVcyMB/hD+2dqrowPs4t86R
gCLAhSSTTF0AbgbaW5+lboILKsS8tkE8L7S1/Gz+zLS+cUi8ybLOSDVXiVr1KEwH
7XKXObn1SDLAtHWy0C4OXqSrEpnimwl33FvuBiNvYzEWa73mpKE+SFYExpbneCYy
Vo6MuZS7vX94z/lsebnkTsdIDQTwBaiYY5NBT5DF8JSd/Nf20TVwzeEpiTIOx0pT
Qmwaw+yOL/9+ue5Enw7Xaj153LMzYy9q6vo0Wahr/L4Qrb+umOEEAcKc+V1q1z+z
FxfR3ixvZurNVFg6+UD8/hEjtZtz/eKTFu0O79gd2bQYwquGIK1agk5hMPVTISb1
ILvgQ9Ji2pmpHEQ049MZRlKLHMabIxW5NhDVaGBmZ/Rn2eAKLNYoh2VVsYpJL4BK
DBA6Vf0z/Bzdc7XTSBBG7ecPBX1bPTat+zXOvWwr8QJa3EP2DgcoKLB0Q81iD1JC
rU5u8PXNHRCt9nA0AwsyfwloK4CecpIFXpia0ch4vIKRuooWGTv7rx1hJFA+MMSr
rGd52cdV57HK5gMNzqkVjgqxC8vCIEn2mWarW3XS+JKtB9XpgIa2S1SsgWf7UYAM
acrniMo3EXhmkIRgX4HCGt4IBS4ssPHjsofY/jkf+DXy68IKG6nxG4eKwM8IVd2G
RyyRxRLEvEx7pGE8yuV5HukD6FV1UKlpgwGLMpEWTet58PoE0s8MRikg0Ag7hVvT
pAR+R+3YICgO43eO6MMFRl9F7XC1Xwroz8ipCE0Bga0WmB40fK8i65IIMwoP7b5W
QLWDkpWyJclRGHDh5lF5WqN1OFlGQo+6PGr6zXfsX5aDCl8zm2WztQ4Fov2OU55w
sXET+nK7U9OBpC5VaBdUBCJ1npdGn094UbEM3/QcIYYX2EhM3PPBfin58QsTukZq
2NP3o+F2TRBHlLqY6hTmiRotbRq8OTtku6q27Gqp+DlHCJm1/9I3uxEuhw6hM5bW
cpLKCVO2tmpXQvB5gl2nF/iM3OUceLZHwBpSjHAr8pUk2g4MP7OdcmBF7PsNb7Fk
GpGLsGdfU/KA+c0xgnV80ryBLM59Pg9XT5mZzTvO17cLjYoa+pxqNQ1D/k6BHri9
r5iADh8xhkQrdyX7jamb0bO8UqvMeBVRfzrsonliHFlf/eFyM9CKaQssHcz5LZ8G
R7dNKf78P9gQp/yVebDxaPUSY4KfVneIm43ZaHD8DzY6CW4UDYDiiWXR/sA1X3Gp
OlbD55U0WMjDe6a0l0CUXTppJGx5xqvZmSKz4m9wwnIKbBoYRWZr/qzIYhpdo6TC
QKp0gLMO6lPTCrZLZNEf8JYP1oLB47wqqsgFuU38nh8DsNGJpmjbPUZJry6RCg1D
uWKA8A8xnN9CDC5KFppg1xOZZJjtr7bjLK+VDh85EQkqMwO2zNdlMcjcOTiffxC1
vWtzzEEz/VntVE3Cx/AlgaY6qp0zKrqiJpoatuiNMWPrIVY+3JFYureBpta6fV0K
eycAh/s+XQNAS2RlDNB+d9NGXK4GPszjeBZpwr/k/rxas7wxtYf3ka6z7dMlMVXy
cXrlkYqFY1iZck5JFc+IB8G/D2PwoLgXAcUor03WwaA9Rycp9X+N7qdvvmFpOtqh
B0ixyFYWEjUO3WDiEO8g1aioMfh3EewlpkAxMriQoMTYMjTaLMSuw4nmaz5afAJU
Hblb9lBQGQCJWr2REjxPsmz03TNSDsovTawq7RIHyY6Qocyo1zTQWeBPK6oNTqYr
oe3IKHQL4191vJ9tVLIGNEGytafcCqlExL3G/1QRDlWQXwgHsfiulCBu99a6UXfJ
vwb1YhpG6pKG38ydmx6f8JEj5uWOL5Rhoalks1/crpycRdVBFkMeIseKE8uSv434
1IBtcrpzY+Riok+6waSNSkZ7FiK+rLI3kSkjy6SRSMucTdYRodFXr4ebmADnqrzg
CPbNBQyJAm6AlXHsl4YfIpwZEpA7rpQ5pt8BNEFwFF72nyTJ7seUheIvWixM9MmM
Nib9T2Vud6wJJF7m5Zh639CurDCLxMkn8u2458lFGrmhzZnDe+1uxXNImGSPlLGi
7sUpYZd/WJNMl4uQGjdhTDs1Cw99fNpmjFKqcCMyTuj+ri7tl+7d2vJwgICq73aR
AwMS1joVy7FQmn6RQXydtrz3UAa1gQ/b/j/UIm1+uAgse2VHcFY16U+Pfc0rH61w
FFLk3BIBhPF7DXN+OoIUhNB9TXCzAPKfnm32mKAmzAAMtq9o+jAVI+5S1ChmsgG9
+mCxWvOfEl3kxskjXsn2wKyK3CbEfpHOjwUd6q5ob1fSjKmk8inzhxo4KfcBgtxS
g/RRwqCwdFWHUi1P0OvkgRReWSL/FQuNcDmkUeGo9iWQebD8d+S0Q8b2Spiaqlh/
WbIsR1RLTnDnYRY3t733ID2HPtxZvrd3duenXnrEEALO1WgzSLUz6HsHg0CjifGx
kRvztAMKZGUx/MmLBx2lWRAjjSspbqpfOFFQCPnYAUkMLj6lqFN+ShU4PJJAnNue
4r1AJ5ck4QkJolb9D51wpHEnoGtqqKWzpbooJRV6Pysc+UTCCwuGFAd7vWUATaof
5d57JX1MpnBYooF4W6Y7i9ozo/Ht+7xgOcTTcy2jIyc4aTY9PBFW8lO4f8Q+n/lh
SLQZVjTX0sf9tQ+DhTn4mDW1bXAovn9efQsnDdwvfAK0H1NZ1rXLj7u09n9ChcoC
C15BB9T5TvDPnjJsqG2BPGgfKacBPJ6h4cVQmmezeL9Df64QNBDCKbWoqblwS4G7
tGq2Vlyn6ipXFKTZtn2t96/YfwaqEMsOICKKVg5j3VUCjEkypw8JCl1k3ZfyKP52
UnJ5brBjUvGHNNBQXzzS1dgKc1lKo4xAYMtpBZ0eID9o0W9Sosz2OxR1gOnNJJNF
wmPzdmPY2BXgboSJs1C75sMqCV/RIhMdlnXm/lXalbiI79FyT57En7JiTz/ceqNu
T5obzdlIk+zlcoDnurjrdxhFiKRFd4tawewS50nma2qsQenNkRY+68tQXe8SiHb+
eg8PgM6sMF0NcyYld4B3GJbkrgTH1U+Cy49ips2hXLMHebLbNSoP5zwfdZz/IeL4
iRMrD5n+JUYcITZ3YV0BMYfXORaazmIEK6AzfHkOVRF9CVgISl1NwcT9tMG29QlQ
axiY7ebA3o+28nvS2XNzg+S/IzCYxTumGSXUvIp9MIj1oQMH6y6kWB/XFnKsJNlU
RJxfN4jlJyssCR4yLxMHzgcPUPFDU7Zty//FMd1ahUZTm14H8SqNI3K7R1p+nH14
n7agkLq4bOr7URfgypyHwX5Hqd+4Kip14ortZ2bW2S2NTU3uJGTGmshHtYfeSbqF
OsPCUQi+dqT5ffpmiX31cBrAoAC9F9NAB1VUUy0psR2xqjjGOwCHVM9XHk4JVyet
nMqtIvzHccTRjS4QWBEahqLwb/fNrNcpz0CNpELnkFfavUq0dt5f2Vc3p2yl6qWH
vhiPnOTu/KJeOoWdN59eXZpuFWL7Q1hioVAvqMVNcyLxfV5V2AoL+57OlAl68GOr
QP2Ept6kIV2Sn/sEY5nlMfhyE829NXfN5jDdWxHE5534Bk0+Xp4+pj6+0wSqA8mh
sZ88LUniYObYC/RxWPi7Ym8kAQ9oIEm/FEZE6eXVjk68k38zysOpcrmb0IuTmXty
eFcnArC9W4MKwk+YYMJ+DSIjWhmkyx2xAiMXcIk8jyDF8cLfXdigq8QzTVZ4dMGa
1PkQHlcwN0LHphFZP+SqdWZY6wyhdF8t66r1GZ6oJutiF3YihAHBFjtS0A3L1jt1
AFamaHiOSpKo9PY8dDjpvCGcdq6j1gKWnVlBmVxdC39MTWl5+IE8+ijBIM+7fgJF
SMXNhy283ebWcUb+OdJ2IfxVY4Cb9F+duQVb2hoA9NdlLnCEJ7qkRPXKI8fJ+YzE
8jU8WclE0FDBvyGjy1pvxUci2bIrUtgjxFLWtX3uxPsdsRtDjS2uaUVoO6ubn9RY
4eAz5e0T6oeHNxfKPHzuBmRrEIWi+oNEMPG25lMjPtOEvPsLY399I3cUgNIm//mL
N998EBwchYXby65corNBDI/p4+PeE9E99eojXIhr7NOCDwXstjtSePX3/3uuKSiu
HApojQUHDCfkEZHY4wpPcddxbP1LxGIlO6G23IG2H2pUaZhAPflzzltnrIGcs4Zr
jp/P+fv4KfW77XoPybpG4NHg+bYKbbOFVUXOXd54h9EVYdScMTdyB1cmM5PBldE6
DJjLIuQTwxYBfkrstGd3zgFlh3skw+o7co/SAoRj2rDPNjwIBLSXHGjXvy5pKSNC
z/kyn3qFtt6GlV3FqXwAxLwRc3kGBSwk50vTsx63JIrHyirSqJFEA0v8rNYg8u2t
CO6wF87JpdnpzKxdvCw+s5PMaXG6GAs4LW1fJjJZogO0526/cRoi9yqmnw81JP/V
IJZCTVpxHJE5yHqlPVsTbjNBZp5BXI/4iUEuttaDvGyq31Ef+L0VWpzT9MemPYo0
Z4wrzPRYSlkNN0KP0GHqoSvp/AuGlaQMw/M5W8NnwbbmvFYG6lnd5oNKfRpCvqzv
DdITvizNv4yE+GCjQ6IoeFYwwFSvJo7z8aoI+GQjm5TnbEXePwgLlUabdq3vjvul
zsMOu7/Q+ZvyX53ycU0WkVZABKK+XNYrNBoU5mVc4WT1EvmAu0sGv/Tj6u+Baj4K
eXQ5lMpbf5UJ/NnFLcGvbX4DI7S1BL/Hi1W/T/eP2DGa1hH0TFgIE5S8AOkDiU3X
yM8s8GFWhciZSfdb4dLlV3qkArT0r8VyP1sqLmeXn+py5WyvYiOhYqogaxDJqPef
r5VWmsiPOQkxkfE+/HYOqBnGJgEWCVV+6iwo93/uxI7fWG6cobSz4C6UFsrPFInV
UC8g8LOZk4VF0D7epOUsyqfnCuSQVdC2YMZFteR/cr//jKCXew9CDn8lqgVtCaeE
Mx4vhBesgod4I9Vk1Cn7K7yGziAsXZNmgWM5pA7BqqKSxUBur9OdCgMKoCLeeJEY
2SYz99FwgXt40+0rNPrRMWXcoCl43zzhwulcFCBwtVjN7tmHI5NlkYczdMLficbB
xTB9h5mzQpEEbprXSoAWn8ZSnR6tgCOWvCOnvoxilFjwrdFCLaxLA9WAepiborOf
KEv/SwdFCkpABbfZgxRDV4HnFemYAuPl3U4eBM+cgj1r7igwSm3hEkZmtGIn5OD/
nG9xE5XuHVm9yETB/Km0+SIUDmMhLIWk0/4Ms2CIQYAv6MoL/T2U+93SDVEj85TI
02BsNOIH7z8sR2r9QQvoF5+l4c95T5eLmYxMliEgGw0YWe392ZkWrV65PFUXVPwa
gc65RaQez6tM2pZ4p/8mni1u3bOqO9XGDIQi+BzDnQ7ceaPmX3BWGLOZFUWHKSzD
l2NHPWWFdTm9AUeZYVDl87ul4j/Nd3qX6LMmRhvUfmh5+k4SkjhestnWI1QlTZmN
5OjdIep0WuycbCuignE0tcBNiy9o8ox+KAZxp8YxDUKQ03OOOyIb4F/aOJPjkk8+
jTT0PL2W1ZjDze4b8j74QdJB4BQrY3U5U4TyDIhSfKB11XCcs84k8HAm+djfiW8D
QWPHWlprg7C6MLaFEJa0zsXXXu78K+pBrDbC72S2EAlnsajw0kXFyCmywpn5tN3Q

--pragma protect end_data_block
--pragma protect digest_block
sw/uV/0eU5PCGo6F0VY+X/HBllk=
--pragma protect end_digest_block
--pragma protect end_protected
