-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YdlJjsNikgu6N50M70117hkHOLLFpxrV9fndk/OPaPXwMjZVTvjF14eh5jAtLU7HRaeI2/JjB2dd
bp04hZdtckFDGakb9KudGwjrrlqpE9RfM1PF/GLFOkZ4oqEM+thOCKivzKJAiqSqIWleT/tVZEZW
gGzxd2L+grAFTXewlbSVfMjHdI/5x+HVzT2jRZV+S1ZyfjMu/UFePiWNYIxcGlLNNfl+J27lRpdm
IqpyKKmKDQLSit3P3eHzSgvV1Lu7Lj4TGPcxmH22zjVaffFLg3FWcECuBXVKFH576M8MT/fjyas1
M38qp5ks5+zoQ2HWho+egY0mhONgw+9iFS47Ew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 44000)
`protect data_block
AIUIBPJS3ZnjSX14td0adX388a7gLXeYEYihpjBLXWHA+UVDJtOhf1s5z34PR1Tj5jLIW5r77rbN
2Wt2MI14zuTgUXgy/1MJ1JQq8YFxFdc3m15GF4ir+CJpIw5fE6v4uPM0Gqn+vHsSs7WP7ouCdMSA
lNCjV31KJS8PH0qmjwItanzOV/FOvrLuWOulAolkKHEiVL4w83ViSTT+hTQrpRTkxoO6SFtkUd3w
pPWjARDrfhgbjl3WV0GVb18iy195kh2xxYTv6eExQi8juKTcs1h3z5iLYOVM9Fne6FqYK5+u+LtW
D3Ol5bO0NFpJqOX7Moi3eDePgm7M/XwXORnhX39jZTORm0ZUxPLmAwJdtFgm2gzsDhYCjpCInvT4
wSeVESg5AOLZgjLfxNPfK7qcs+gLaEp2tOrhnz3GydWTIrqmJfYyMhf+tELIgBka4n0ZIpMG1323
oNXWPEmh7jYC4YlngKWYz757CPdF4/mACnqG8JcKiaTN9uZpFKVLnfEmGNPWV/Epqo1l68O2KrRG
/GUCBOlti6vo+bp0INRnTl59FXyZXVgmmGu1cKMwPscdO2TNcjKO4DHhU9rDrPVEX7YXNbb/jO2g
G0Om+F9We3mgqbqXYSQcldl9hxJVScuvOvPH382R1p5fs8LCZIOJpsCpVdzSF2SBvNQhsM1yenEb
fUB/ET1e5n2ccOfY4o0k2gRRwUcXwwsIlt8TcxeWbtCxegPEsodbRnyvh0ZNcj03ex6Mvpd1JBGK
IWQshEyk0gDZpmfjF4k9lbqOKzk0wxtYbiS9wpB48ZkZwWD247Il0stybLb4Y+tzwugwssfyAVFU
U8Vq2JvhNIRfjQnw2BVEAAeg4uJ3ZEuh3XeW578czj5hjIaD8zelm+row8u9dIeZMjVwpTIU2INB
SWFga/x/7rlHG6cS7+9Q4RCasjRkDjxt3qZPjsoijqocotYz8AOh9ar/uK8Fq1IhufRGXPw5mtpH
aRpppgfCEUyTRSheYve28pzcWL5MdZ6HZxYwlefyCwP1vPavqPZKKTkG5HYMvXvma1ojLNWuMtSm
EqF0lwYKuxwTIqVPVWH4liCiobda6kcjX5PQi04yi/UITxOkLA2IC+RBrIJZK5swLAsB7GMgrwiZ
rN7i2uRmF6tg9M1335dsER/+NBTtwpRkLP712VaVEgPDh1bp+hWPMJrjGp5N6BCKlZC8tZvBip75
rLJKx80b5OIxO9nMWb4N04q+iEhbjbuEpCbIZ+j8JxMwsDHteEuwcjgR7j/xmYVTwfV4bqUTJqJa
Mm9ufKdfzzd3XEljcCpclnSEggp5+wC+LqB0fIf/ikuoUtmeBraBEpUw1td/kndPbw3P7g5gM4C2
SrvYuMRHvotLT84mBBlvyOll0EVRzsP74XFwUGDfF7b6xV2UbX7Gy7Zlbw5qpDWnqGoFz43Ifn+M
TkghZyEqlmp45RRCqM3GNRTQIIzJLOSqWODVu6xnd2SYmyRkI0gaBVHcLO9mVfYZxj9hYol7RPOC
lMaZgjhiFeyMgsRpcoRcgUPXoq13TGDuf8IShfiIr6byUqnTE2VCpherfeHTKm1RILa50O2AHWQD
NQZ08BoneIKcjDeeK3I1bS5pC29cP3d79zN15Nzaz53TDANVEGborsA25Avwd//XwuHYHsuezAS1
JRsQencDhwPJnWnoD16UEFDqSgeGbSYTjW58y4JzPVWguNp4VYVUwHDjM7FxyA5/nux7GO/NNpC3
/z18cOYzmZJN6XxiQTL8V4gxVGCuNPc2uLL0SbBBsonZRUlD8Peage/zRzhDwdufbRgsyl6EmA9H
uYuS5U/A1ee6UsjBWKNkVfG9Mi5S/6/78GJpzulLTUIzqrCQ/ItpWg2GGk3q2KJdk9802f2Od6l9
hO2A3UmPADw52vBXaZpiyjrWGYX9psU6mGKuuUXQ+duNdF/VZxp7WCi3KrV5Rt8BSBOls+BNzvHW
HumalTmmcr5su0x3NYJnammpHMa1I+nXM+br2vIsV/TQUUn1WCAVcGfSQEaEp2Gs/Z/Yyz6ZFwVN
961+nY8oO6kE7yKMvBrdVHN3nzYXmTZ6RgcwTcPMeIy81hUHR59B6ZRuBQInKDKRO/D8NuyVhpwv
7f7gS0Hu/5qLITeHVh6+D0BnNN1UGVdZsohwZbiYEDGPIUwGYgZkhu/++i1XlZm5C+3SBMwrRvOg
CUQHxSr77cSmJzlVbIcDnIy9xxavYFCJLy2MmmrqNamg532HdFvB1R3uXgy9D4RQZT4Tw9wsqpCD
Qb+E+C26/ywEmRYOF2FDavPNe9MlAifg6hFJKAtI1g9vTnBVt/YU9ApQaboXM06nO+zonymtgQ9W
WRVSXXIZemwDf9+AzecDGE6djuJKdCnCIgmqo+14ipIjnkhyocLn0N1tmsRE8uJQ+GfP5Xn7vBVy
ZMsfP5tROpC+dlTWwk5+TRRa14BZzCI0s5PYmIiFZ79LzWxbdJIKj0dAfj81MMytBjjx9ZH2igpl
m1VtLcqA9HmoOJpTIt9ZsPk/0kfRel9pKaIUG+c9y66osmJJcFNdzm1UY1c1tqJYu7ff5WIOf7jE
PI5yUmR98nLwWKN8uK3QB+gring2saeVsoTxcogpXoW7O6hqwZN94UPD9PnD8XFajlG2+RvLVPz2
9BTsCJER0hMBLiqhw6kbDLcQHFWgZXlr0T60s78CZjXxowTIesLLj56NSN5v97eLuV28CbQre6mI
Zzyo25sr2mogIPzScQzGw+sw18jSW/XD5GsCIkWZ3MnL7QvMhidmIdfGa+bniVQR3M4WonRhE44l
zHXESSvgaJoYnkMTcGYP8UmW3GFkRpa7fvQoA+aymnADqw/siEwkuMkB9jupQOkaSftn2WVUVnqs
mRw9h0GW3yWydb/pE16VOfudZ1x6xfCjs0CZMZLxnWIfB8J7EAjN2x9AogT6761v23C4w3Q9F5Ip
jtH34JhB9S2ydrilRNahWVNQTdx2jNgapGmLZX2Nv8DA71MIPLHQ2AweSJcA6ZBckcTMZfIESBiB
4CdAngbydTl10+4OOYpdFfknzngu0quY0bQUlf4nawP+DcfmZAyEIZIuj3CkvAnbMr1iSrz85Xo6
CACXxKVBAeauczrS0EjRCZtQ78XL3aUjGkkOM4K/kWkiVed+Kp9085PK+P0xc1dVWiv/BAhuWYvB
yDVwdCNKrcmNQqfAofbk8qQfyz+aj8AgoWZjFoKV5qWATXUvquE4WQZmeP8uOwPnoG1/bNlMWDlo
HRnWHDm4Ps40Wu3EnmUU9oJwIWuPghMFJ3eD6bYzoyC0Y8Pul7TKX+Bt22erYylFzchjq20j04Bh
7ljf4De6glrp7ff0T3/ixbDri0ZHLsaGDB2Rfjlb6hZUgfoCduQYrSsMZnCb9ao1YO/ZC8nnaGdH
SWsds3ua1wdzTU4nlTq5Uqi322FRwIcHzLskBWht0SmqVv9WelZg7ynDzODjPolSXzehCtOUEQqV
J3fFMHTiYuLzasdw1G3YekRD0WmruS8NZLGsmgnLLVbOFusWB9zk4Evp6lm57ss1y76flilAc/e3
9Rc2PaQ3ti+QRYATWw18qHqNdlK73NMKozMdr49p1IMCQbcawFtLIJ1M8Umqgu/DnOJbYoVz+b8R
FfAoCr299kL3Xr51V2faQ1ZYdbl8xbIQdCCwKcDakiKlZL+p/fSQFWUfJxpyg1D1bFFfZm4Rut8D
451n7STjfGQ+ldz9yzcJsHR4CAsQ3WNEKCpuWXQ2Bxl3FRLmcflUpZj85YQlEx64ac3ErhbFYoRL
eWwjsjgc98sZDrjwyAzB5Bs2FZWa6C7sOXXucTilBHvRoR/22yTRpFSE3vHP7SF1z7H3ligF/42L
CQG2+D8COMwuRDjYp2elKMligKtbSiCBik+Bxdsb6v0zM8uuEQpqpdTTJGYSFqIS/ZBD37ZXo0sK
n1YLd46EhzVleQyd/vnOedCpBqwIUCxI/ueqFtgV7VARKcQVieu15wc1uiPfzjkV6FVFe7X36t4w
IHP4ZXcEHmPXvN130VuQNXh4Q51imkoxo/ZbPQEfUXEdW/n6SrC0aMJ5wntKKZLYzMMPM6aOxjmx
Fx1uLFF/Na6tas3Ma5rcwiiyfngDKaJELEv/Vku1djFiH0FCNVS12CXEx44aw/2roW3xftqdWeBT
UhKLbIQjp1SikBAYk3tS9SxWbph/8Lsr8D2hG0qSOhvcDmncjY95o39rXZBLogy1oFirZ6Zypm0A
Zq84v6s8ZHPRiNnXkdvso6z3ErnF8WwgI6cQeCiIc0O7LzC3NyWIWlVsORfMNg4Hfv6MLeXRJlX6
3by6Kxgb1QP4hp4A0sNX9CfEEPON1aNjOM+LsSphmje8XM8a66v+IG57JJ4QiMB4EWwsKzvz2FtY
UWyz+j1W/QDpol3sv5Ur2Cb0mH++TRsIUIzHbilIPgogjGLuWKaI3vjHTBQo3bXzHQ0U9ipLI8gh
EYc8Mgta4CimbbRsGagPQB4zWqogbitf8GjhNKg1T7ah58E3nlC8M6U0YDLninO+aKszWV3FukFU
5CAXGSIoSNO/rYFBLGEwtnVqF0QcWBhKwQmSen4YNDrMdb3uAMowle4W6/dMQKKAdEjr+DrVMW80
8CwoKznOewt8j74bRralPIOufRez+BCM7sSsemIiUqouk4TDaF5p1bi0koIRGYIAlti3yFWDZjfc
CiPKFWxgw9b61Pqbsifi+CqV4khHI2DzGGbPOfWUVTucm8JOWbIOn8UG+2cII9alE+PQfmOnAbGb
jVDaFfvOiA0MCBltC9PtCu4nx9+I08eibOVrZP91FNVJW14TXKJ4meUQ+zMg6SSiJ0Un2Ko33BcE
0k27eG5Cu8SQjcSIGD0SVdy1Rb3CmsYgRbvyUIh5ims63vV5L3fZfMsyqQ2USI/FOoWQPvkUo3cC
qdx6SHk8DjIJrBet5Dtla71VKnXiEXsiyHSULbYIHfn2mA8RLMZ2Jb7uiI1epcGc4J5ThQZVRuCs
CUxWzkEUyORYN7O8DYWX07AuulrHi3w8tjIPxEoPO+L20l6+lz+udC3jWzkFmzqfoWl1qdkpshrr
5dh26yAi7OrlWnP427DyUxsajTrAH3N20tqZYzzXCIK5jwdDC5XBFt9kEhgN1laEk9puM69uC67v
WDSxbsNKFotV3EzHygNJa6rK5IK+HZiVIg4LQIcvztTmRVBuOhMBpbXXEywiUdEJFGNdFHNtXz3u
ZO+G6x7l4RADF3IEXZ5GRucafngu9HrVB9fFRHnOAxzzL5946SPIyQhlhgYwNMXx9xDyXEoIAjmU
utHmRjEWGRyK8BazIiYqQo/b1FMhGQdupAoM3zjcwCyv/oLtaCk6Miy3DSksU0G3C58Mp/MGsb2e
dCS1Vt/V96EV1Usf2DXgvclyLf5koy7joEpdxuJGfO3EgRdWmceEeFQglUdEt4O0d5QA9FDKJ2e6
ZdwDVgvMlBOsT74sg1CI0OyYxz3jUcszVSUFAi+Bl68n88Tm68QGKxSjAGOWE3aV7J7ffZ9AIp3c
YQTqd9RryNiulpeHdiOzdOhx2Ff/zpd3DubnVGTKA04vNjJJ17chVzsCeO8o4gzoct5FLfsU0LO3
Z6Za6QoAl2O5/PUc3IPgC/tLYHlS1dH1Hy0HFY3CkLRL6VJi79OG+wWfiO382TvQbyElLKi1SHXf
Ifc5O9tHOgMrdzammemSjDMiPii5VCQkRPVQrnJDyDXvOxOMrqoldULpAUzsCC7yKyB9KgVpeBUt
YT1Kuady4fppluwZAiR2RdVJZ31x5T38hjMvWStxZFVCTR83aPbZx5me1pAgyPdlZXA/swmz8Gd1
72BE0blufUfqCgLXoNUPFHmkUUfcgjGnzBleY8nWyVFzPTSPH2ZIawLqR0FbtlZLxRZoM8Ls1PO2
FrpAEda7hV66ByWJc6vadRnHGAjsojipJ/o4COnQsy8wXrkIiJqvfi/BZNllXF7VJDerRSNGQ7rJ
X52/tYbFLY+U3yq1SoXPmB2ZnKvN1Wt8QHNzD4cKBXtTw3DyGdQvmf6qJi4o7tRevnAi/zX7pXce
xe//d5KjYHp2A88Mnw7c//5mk1duNl4LTOn2T+KKOlIHURAA1riAxnRzOZ7wtc/ud6leG2+7Jl1H
LZ3istE/+p/L3yiappN5W8cd+ugr47TmDquyUHJmbEvCOCb8J2l30b0DDqvmh00Ohcd+pVLjaHk8
koUJ3GrrztrSp3XD3Tj9CtKiGdNj3adDvn0C2Wy1bpBGwV7FDm9Gitrn0EVP21jSOYaiUQohBrMY
Td2/Rk/jwql8M9xUjta3HkBhPhCWkp0qjo78994JFjDuWY/Q3MaDmCcb2jdsa2v+91grj1LaGGPi
MMGuYe9omsJSmBsM564cQONKG342aFeHmDoi8JOxtyZ2rLaCa/PLVZcgRm/S/cf1rxGe7+a7izar
M2NzgbwOp4hgMbUShU8IiTQvD8TzcTuaww62Kwgd9C39y3YzZ5QOS8phQBAGk3QEbvj527NK+gpH
oREAlmNgRFhDIb7X35Wu0+g0qzH5qZ11fVkcJNJ/Gyqi7UFMHEDS5+SswxgXU7Ay5igtlVDu4hMi
uy06pPhYUDzDPFHPC+D7XNfJiOGsB0JxSogQc6q7JaUKrdykS0ru3ebYBzIHy88jQSqoudWiwdXT
Jg2YjEcYFMEbGpm/MOGnupdc0p2/I6Sw2ww/1D+rZV8kddmNNH8KmTYDMmIa8P86c/4dUK5n3jtN
ePKd8DpYX84NEAeQGcYFPtvYEdLsie9RIAQEGnUQ7s7seUWbRr6OoCzGpQEFt0bJTJ5GFSdQYD1M
NSZXLh+tcCjQCRjUMem8My0Ezxq+gPCwgPyDkcw4TQu0lCHGHEXiKA2uMRcnBeDE+zNpXGX7VUgq
pMk2b7RYRrhclE23hmRDwyhAemtYU8JOim0525h+Hm4DLD72j6gIe1GyYNT3el6E8lf+6zGn0PrE
LCNdkQX66U47B7FTaw2IWaP/8xn1JKNIRFANg9BdX1FABeg6ziHfHjaF+ESSmQ//yJHksU7YghhL
vFOND/bleWUnN3/UCkSXo8MhDtBP+3LR/dvVtEqYXEHPvu7oaBV+CDWHT81FR4v1AL/6ZZEWdewZ
suoi42rphwognehTi5QcZc/hCu9mQxlFcFlDuuOu1c2m5+i/dEvXcqqRZx89UJHctArX/XzyW8vh
OK7vF0+1dJlDZQYEFTqIsbXezvcm2rHRpyZMx/tr04tcTnaDJ9whqwH2TnBMi+LWmHjpQum44NKm
DeMkqfaSJIjYupuAEIIqwLosrlAgo+m05jWF4UXj3xfiOQwOhMCqQ0npvNh/QgLUPkLnlMPuG2R+
iq5NPXiyE6kWmkzcvKms/kh+39il1E2hCgsxXZkmjNTXHTCtG/LZA1aECe3jdKNrV/6ts05to9/9
Q2O4WA3qstIDec8AiF6ZXGNMf+j8uRG0u5PZ1VxICyNWoBPB8IqqPjJ6aY2T1EIOvSFEQfrPZaov
+Rqn7boHeS2mC5yroy21wf9e9XqCpBv5cFmoEbyKbA5PdO7Xk3t3MD6hrjA8Gr/X/iNAFgn8Al/3
NjrCja0hwrIL18XMP2jlvTdR0OrdLfGzR2clLPvmYqRCWMzjQWte2D8iVfXRWVgXz/6s+aEfrgyO
SCNuX6uQ7Mrz9wNB/c09omMaABK9VY5VBy0Yei3A5+mEbsGX87yDFeUyfxwbFaUaJc9lcPyzV6+/
gFfG8prEutj0FjOOvzZhuRhW449dvbasasDANs4xBZ/CTPMUCH3m1T9x0SUbEnaq94eJXJf47XSO
rfPvxtWDSfKPeKFauUg2oSXA7nQLfLaLN4WBNnX5Xm39tN8gUUjQrFboFtXWTsbTkDlT2/rHqE3G
FuI34kYsHB28pHFAMMUM1cQUG075/4O74wXMD56t6CjbTRtdZuFkteCUAEcbd0bb3p0aLNCyoaPP
2GwrkfNG1/yikJfP03QoK4YZacEaGvaxNDuFi8Hg83D7jgpyxptdj2+lPt3aU1NEPWQOOENGTOqx
gw0mRakWZh27pVLA2a5nH0xQwNfHOmEt0ZJz7Au55DnXXFNlWurlhRYJ9EXnAWmdqkk4XK3l74iz
pemj3JYLsUBZHfIHCBOA0jZfCdXhFDgpfKW49nhJbYsdV2mP15xJNaHyY1wg/4atlULMScCur+Dl
BMIZCazlQ6UjcmJ6IY8DGouKNlPce6RS1gNavJhm8ihOzf52Y/g+t4hdAFLUXxyGghwtL7m4ZxXe
S1Nw5OX2LZ7DxMXfkJYj4JuMsxXti86U9Ot3kVHgkN3ZnUFoTFBnlNL62bLlpijWjJJUT7Lv80iI
tSselLx7jNfJJ7gwyAoNt9cn30UYY9iu69odogJxqcrJ4lMj2aGE+wJEVaf2llfGOU+C3ZeqwLR3
UGbwp+NXNyiqOi1z6hqbbgfo7iLWbufQVzZdZApkE8tDJdN2YcvaRGMil6VWYUTSuQaL0WTTYSAy
4viKQBuGERgbICBtIYQyfObEwLxp+Cz6QC0oZ08GFwWTWZX6WZapTiGog1xOmudJFk1YcsiSOPwh
omLJpa7tq9CAl35odfS4B+u7R6y2tSiK7Cz0zfxyuSp5W6zhGXV9O9co5mirktEld+GrHxVofShu
m8HIJIe2I9/cnLCwNQnNJsvh0QEJenw7GhhG0Na3ydl6eoPh6RDxMVS+1kGs+JmIHKeOs/DgCXlM
hFjSzTx3cza+waRnMULpaitarzDcDYyatS/6oxBo+pApIM2kfn1Fct/vuI6BDfkPGUlG2xALVUdf
DZngFUJ4AoQFnVOx1otBmReow93D0MISGg05DwMYI2bfAxbFnBHZKMbn0ZSUedSSpr1nVI9ruYTO
CtcKi2SLTH8FcMI9bBktPmeoD0J48NJUwBZ5PcRCUdQDXmdGkVaOa9ZXVHS3b5H6degoNNsH0Ods
K7qeN0qTUDbRIBcPpslydX4bxRjVfxWNb45NNLWkokJr/QjOsl6n06PCIdSr/k7e16J5Cl8T+DDO
T9ctr2sjjkReaI4ABZrc+sBRliB7aKKrHUvuI2bUC3L4OuXggDWiRUS+u8djSSAOTuXLr8VfmeMa
FKSXtCSO9LaC0LgJYLXPV5a3gw5ii3DR0zBerqXVhisZtzFd4Nb421uV779b/stR4nFPTvd/qhYF
Uj6vppDHI2xBuuREHKr4eNKqK8xU+aZuXUEoou6+VgEH0bMGxTFedwfwxQ6dHgoGebWntxAFFrTL
U6aNxyTbJzu5fdJGWzEzjw+Z6A37jNP9CXijTN+K0j4irwD21InPofilqdK272/qBESHHRKtQhi2
cfV8lpuPNcJVNz3jV51lrQm0T1B+40kNrbnc8VOja2gQKa4PkI81UEOiq3enJUw1CwlwQ/RaBRuR
+qeUQTiP+i4u29g9NzV5UYRFedj8QBFNIK50DM4JhL6T9CoZLoG7yioaP0WN8Ey+et3EqfQn5yz4
MqfHkY7+ZbleQrYSkOLlN1a4zgYf4v0i51KN8jzBe/cZlSlBCYHDTF+ZNCJ6Ni0z6eJe6iZP+pjQ
jB5njTP1P/tOJpLe8/6SZIBWKcDKA3Tp7EGQ4rVovpqNHPUbuT/7Rf2yN4Z70BS/ks4Fe3PUhMyY
BALaH8Zl6t/ePVAo6d7vNZUgRm7/jfsY1ZRXYJxE56PZBW08S/wn6ybWr3lLLoKzv2i0wsXcXZr+
7P/S+q3FjiVQ5YJG+TznGYQIF+CDpVugQwc6cNsxAQwxeVnd1Jm+p/DWHaVTW7urbvu7MNsSj5UM
DLc9RRv/EKdgiSWshb2c9q1iy8+VndBhBywefrLAlTFc73LeCq4HgpeFrTnItLVWZZJNBcjpWQk2
5rYzDrt5IIY3BYEwCVdNQziou2hVuQNifnM9xkngXZzHis2jvxN9u8MyQnLhf1YqQN8In+XAcXmU
7NylrS3ubQH0gQQukdUEpe6sy5b9wPfkEQG4IDeMytQft455jNGdRzGICT4ssU5msNsAl32em4ox
LeY93QamtG3g3BXbM3YjL+CVMrF+nelpLQKTA/lG6wJiYko2j6q1h8EMT2Tf5J9oJEoEr/P2PgYj
QtZ+2cDHgdheDqNNZ06Vhx1KoFUXCOOxG/Cf57gldtEWPF16f8e0/QAnamif+OtY40KivNczHDv6
UVR6HA42cOAmLIeGde8Gbb5vX0WGEzbF2uRODEMAJQw6Jya6JYVgpvCl3snLJ0XTs+Kl1DrQNzKv
qNAKJO4l0xg8DggjiZgMiRyLFpjKD+FKZ4NpqFA5SyOFsujG6YKsLommKYny0mT7JZz8UnDUy6gK
s6Qt+3RlTzOSos2W4Zk30FscGg4nyJBVo32h5Ga4neG23z+LLiDCX6iNq3F5pCKaAwBNyedWgJPF
dAJUxgUsmxklIyL8J7ATOR+IVYcRsTfQSSneDoOTIlkDdfk1MCLVlicVwa7VtONmRSnugcla0Zdf
ovQl31IQukA4geK9GLwuzJU0VZtVmVTTet0liPvP73CpitCCqDAMAjnG/EljNBzYfkgNTREhPwjx
wIqlw1Qhmii69POZE9Rjmhj7GqgmXrByBV1e/IJUtE71gbOC4fBD49ypHq4Q3juSBy2pIEFgFDfN
mdKYWR8okdZ3nyhz5NBXYMiLSp6dxkpRi9wdwNXkQoXYYCo3p3m6MdJn8oSdL0ivaizvwxUz3j7f
Gg+0UMJHxaf7JQ6NWMBxGLKBVDD5hze/p2I4bW+/3Xoi4sNj+QZI31Dl+GUMZ2UIy4OLlcgfFI81
/WEiRiI9y86raozIMwGdi2uoyw1U8ciOgbXYykwJcAIjOeib1Q/Anm+hj4q43KI+oW2cWFkuXnXp
OvVYCG0SEhGIxDLYxJm465S+XpRwNY82K6WsuSRAn5eX6B5GjrfgOsRZHr1zcwvGm+Jh0IW4pawV
UdFzOEzWyo96BFy/DIU4ran0DWedwZkWsVg/2pACuhQcK0b/g1xkDYVeZcFTYD00PjH5flYrfxNq
VfUVloIjfHdX8eRP/8+mSchhfrYRVh8ime+EZqrHYB6bFQVuZ9su/Ej0H/+KhwIWVQLuT2FBPBZs
EFDYexcMxrEVgGUMu8kWuMfuMvuOFSqU808EPYBGWlLqhQbGbQ61f8Y8Dqaxn/waIuEj939fCrMv
+gLOLHr9ujNHHbgnTLdKYhlEKj+LL7o16YvDXPlkdveXN4sAoG7rfxJV3Roa4HH6HDhPqoHrb6Ej
eQACm+5Th4MhbXla8nActEZ8DTDY3osADZaT1mXjbYKBz3fMZHdmHOV5djIQIyH3mXw+dUWbLDK8
0tbGutF/p9oAZzs620PRjm7PIqmGT4+eLySuxfDlwVsGWwIlxFYELBSTWqpRd2pc7dHWhuaox3/L
PbZjZc7/abTxxIAQegK8gPCcytIlPs7qj+3bPuXWmICezflIxY71cTtAcxSHukgNeeUpSXWc4T/f
5Bilp0cIugOrjmuLZW31C3qjPQzjAMA8qQzmXtWHsCh+7dZDs8IPz5xxCDCvXCFhKm4fGAQT172e
4eKEZjfe/dRDTFqSqpco+6IBn0vp6Z24n0C2TRmBrpNfp+/G/IIWnq3FcIb0P7Gn4PyOQuvP4O7k
43WG2eTZl9OkEmzolXvkraS8rcfY7hp7t6dzsknBXa+Ikw7ErlZjdAA/zs15+iT3KAygLKB26tCf
Ch9jHogiqr6tVNyIZH47NcEuMmCBu3o8tDCOUs/urEAizNHLc9FrYELyMl4mLgSUboMeca3vYhl4
o0Ly1jpZ9gx0VBckF9V3ndok8W8jpKvZhZd7R5vobWqnG7d8C6g8ebZuiqt7LwEZeXd6P79Ix/TX
til8EfpoSxdNeRs9uWCdk/Gcc/dSDI+nUDaA8qiMd2Hfi00HFOk+77FKNyWyJDRJwHFIFa2Rjyxu
cfX+xQjY7oMf0dIGRoU73LQUp2cJCXJaRhnT0jat6/pYv4wbAQZ9OjX9z/KC/NqarR1QlpCu/RGd
iYSYpt+1XsIJs0x0Y+aVAX/z/DCeun263nIltN2Sb0LSAutbLVf+XdCKNyXzt8SzVgAmKpaSylEW
rZ3uJAUGArpu0YlNTiOJHXs0uLVvUqHgyYg4RIVWGdNOxHFWHte4t3rwt/UbIx5dKTNWMEGt8sXp
C2jTyAVJ+hEIW/XhDTje72c+9aEpRr2kBl+k+3iFnYYCtMTjCXBEyvvXYWj0Jetqj0RnNzMTwoS3
H9RKUil/hZ/Uri8TegmH1tN6LcRx7Y754J0FiAKvlwDDKP8Ul7XCKj4uxeOjHIqaqvz9xgGeId8Z
Gqzac6ASiMVlM8beZU9hTk8cikXY7KNs/gGO8om5qPh4uvJ1+6BHbeCRA9zqTajJyQaV/U6mS2wM
osiXLF8gdUbwBNcELg8eGnbOFV+WKJYjt5pvRlDDc4W0uLO9DjXaKUiyDnaM8LpxdstWL8df7cpO
AsSQBMtmBg9ztm8c6FE3dQfn+w2PY01YCJxT+9MFcQ3xdM6E7zuYSiCddzQBbUwEt9cE8xmiACOD
RTD4TpvdKYLnYTu2b/vOCeGrTEkEpKh3yGJdJxfUfezTdqN0gUDHKB8ZVB0EI8VlqmlT3bu8DgGt
uTAmZFGQ+9BugMdbUEChENvI+O2QSxjtljEr6EBPNqaO4+3C/KhFJUzR5rCFAyZbMOAwfda9IDNz
JVl1XCqnQ24lC3FizZZ9m0MI5iTchckeFoQszHnWy13XwLxua5Qvo7FVTm0MnVu84cJILNRFoTtQ
umVv5kcxxW2BZlmX/B32nTuSG3819elSmS10Im3mt8C/r/pLOA2+BJ0cOQr7KygpIW4mZto8dp9s
9vSwvDmA6RhhsQiT6s/FUuaJFgqPuYysnIGNmf0qOKJ9U4UVrtdF3qj0MLjN6jdyVe9HLlr4HIE/
psU2BeB8arqZuBsBbBgRTywksbXUyD+IBJt+1gyNLXFgVSuNip2BbGx9z0YFTEc1oij4K1gFMzvP
QilQ+fYOKPd/3TzbJshArhHHqLRKtyZZCSjB66TPmu2L5/xieg+VhivyE5tTF/tLoYc76+8FCxbd
OMUO5DfInx4lSqKrr4aVDX101MbR0Y+8bPncUagN0MS+m/ghqTt8nNsRlfyNC5VhiKE6Y7PAIVJ7
ljshUbris7MH/F8AQBtPZv/bZOdPBxA98lrzV0Kzxe4VdNu5WcQSAZ86YTA/mTEj3TxdL2YmEoJy
0Aqb1RT3xTOKHo4Dfjca7LYcNU6xy8OenGKnzlZZez6iGF7Eo3gpgfyCE/mP29MweVz5I8e7vu2o
YnkWaO6ROkbB84Tz7wRW+iGYhwpuGh51hSFOSSbZaD/7GQmUtGACptDTNZeDgVy0IJnC4T7EQPEz
6EXS1vLlmWc0fkcJn4Zs+WHX18WbKxlbBhDBOoDrcGyXCGZrBOT0dkBc4bCRAcT6WgBeZz8xOY8K
MvKGrkmqOxqlUwC2F1g3YaScyHHcaDiqQal/arJ0N4/ajOv60yTQtKg5FRvSYYoI6L20cDFPEA5W
LsHGg6HLCE86Vbn4L6vn+pWuVpWoBcokJVVpCJPKSnx8wGWRAUO8lCSrWxcfEC6doMJGhiVO4Bwi
JLoGXpGB/6xM7h9w/M/JCMTET0xdMpswfa4DiNBtzFRp24dfFA+Lf8Bk8eRo0/pc3NCoD+sVUymo
zboQHRmEH1POcW1a+7oyB2/Y8rT70gObJwGPH1slnhISPsUcud2TzQc8bjJOrldSgfPMtm2Cy6/w
gsgA48TV1R/g+u4kmFQMLJ0WFA2WibeohSxzGcUyrAVDLMFbFLsqLgSdTnnqrUFUk9pQXzAd+3UX
gdlT+gJyAWmBuGuOmcdFGl8XDDHj/jhiBmf03M5byAVpgxDgZdT1wn8uoEbdjcgdvV1Jz0mCLKKx
Y5QZz0zCR/1tiT5Via7dwgJIOEtqwUg+ZTPMme1hh9/iJn1EBHOoleY3T7WF3Ribb7EtetWver1t
BEd9nSossG7Af3hFyf5mt8rt/c8gsmzTAoEPGQir6vHGGt6gyl4AfZkdmff56cpZh5sO/cyhmo2i
TxYU4PRQvom3/rzMidWgAdcp/FhyJ6r03VujvefA7ERv9QSSvvvnfZHcyFX/05IJ8uoX4Cw6I8u3
RDBlaNw4SRRZCmGo/7n90a6VNjxR/sAqncU3UI36LxNUv67JElS95ORaI2+Gsd89YXR3AetWtB38
/4BbnNdtpZcMm36usuJxfxLfJSY6G1vXZ6rcbM/nR1HayWJBVsNRR3KNLaBG9ljC/aOtt4NwV1Vl
LmH/KKiKXfaRKx1OBnwHSLQGdhFBVGC+xA/IjV2aBmY7qnYJzHa5u2EJrQjJajJOW/DZKbboqZGs
sdF4LXhvAEL2JO3yeQcFVehUEwbMP78fYhgY6s1OWRNlzZyYblnK68GLVlWspzY0V6wg1NUmBJ4r
HSSsZxA78KWuUaD8EkmTMWufkRVhtIh1xQXTE3d3OmNt520wGtKG62OEVjakBbvAteskJ/g27WYO
XHp+5Tld5Vrkjb0ue2N2rI3KwYVofxTQaXW90UbFCSF/kectswRcrZFXyg0V2ZPuiEIE7HON6dmC
DzTVr7UQHh+aE8guGHJwvxpTYDC8BtBHRpnA0EJfl9qEaLwW+LSkdf2ZnNqg6mgVMsrZLThAal4/
KX9bN66Rxada8BkRElIkb3FHuKRyrPDURyo9juIlJzUfUSPkMq2g0kuzUQUvryn0xkfw2+DpJ7sx
3Srde3jSP2y+IySSqLM6iSmoUeuyuYO6f7nTS5HLRMQPfQai/fPGs9J/GhQh3tqludIQgcBINoC3
oBiJIqEZLzReX3YOhmJHQ+I0TE7L8wdUzB8vqz82V2COgV2r8zeg9ZQaiLf5P7gTnTv4Ub+VPpce
fEWQqk2ILZzQrZj6V5xiN77HwvlbpsI1Xz8YpH0S53Tnv3t7mwzEL5L9OCZgPIe62R+RwNujv0G2
DsdhoAn5DS873jed+yPn1WtZIdokcCS9GA16YJQZsk95NyEjDJ2fNCav4V5S33eazIDZOCqvul6z
UhIiHZeQL1JVwIlFZwbJ1p3NMps8zvaq6fFbh2c5Yq7VH+8otdzk/ZjesafY3MwaOUsRz7wgBKsT
XWu3wAYqy7EwnQ87N7GhzGTnfFQfq8Lfl1keFFwLHxpzyE2xXS1quPTP6byOsIxS8U35WkOcQQx2
rtBHmwrp0mH5Va/3gS1ClAAOuKiw/pkJJMC5YEQRdm0jlXPgWOLOh9StNbxQ7VKIHAl0Gh6wIzdp
7BUYqSDllWjhtntIdzDoxGkWvI+WAw730hPqxaybPq8W8mL6MoG2Ve4+4URa3Zm386yImrtzyW/I
h/ToW+PhoYfdy3XRuFSWRxGfuUnTxF8fB/SfCaRVLz5ImJrRoj1qOyhDVJH5NfWhikJf3Vq7uFGs
uV+HYrGvJ5WUX0YPhzBDgu1VnJPKZpvdvdMvcGyDnimNnJWrmnTe3c6ziNGKacFnxodAVEJjZ0Lr
mDOOqLDe0eYcPuoLWNZXOgwLlxqvLM+W/k2636X7F81Bzw1t+/zkV/VuT0woJUhGNq5kVOh9J3v0
38ClLAt0OJLe4jo8c8b33gVVXAKnbyqO0UUrm2qTr5pxB0hWhYwStTEMU1wKhfAtcb21aUHjd/YB
F2cZcbPrRnCR6nCIM4ac4B4h8uH+16lqQxlH9oyu9Zu50dYfoKF4E5mieTmYBYSrA9NBDwS0Fdkh
Nq/uJy1G4A9WSyYeQegb7KupJILeBkIiX7kgjV9piverN1z266oHp1QeIG7qwQnHqXNRhdJDDf1b
m1c/TG0Xl74wH6aCdh8auLnYMOAH1lU7IYjzwV4SM2lzDHCivRthSricBQ4yaWmP4xJ9BUaVMc95
kTp7aOuJz6861elJf9V9jbQMWm6uQuwKTf4hfomGvLKmqYmm4KHNvWlQZ5sAU/iQUIvdDrt23t6s
X55LgTuHafqQtTIMEPOugFkO8q/4Z7Yg/q5O7RnmOeiiyzmEnIAtBo0PkN15+nkw3O7bUBINuxwx
+NIJwNwOpMlTAgnsoz4GK2jQ9VwXvVP2DBrycKsZr7PaRenWQyUiZKHb7BpOfGl1XD5UXrYyBb3z
bjAuoc6ciXnE9i2GNXZe5K5NrG32oljPrCVPHX6kIvz5SJRa9IzXDBJKl6VfOsd/eiyPLJgYVWQd
nDVHr0iavWwfCCYJXMzXYLyajKfMYvKJA4GKIeIdzpKVq1MOS5Gy/STKhqJS9tUr/MqgkCtlbNdX
LVQsUi4HISupj5R8FFbZLqZbA9w6hJj8i07dt9aaaiEy3c08g47SJRwCp8Jt1Xa5UdZQ92WH0ovV
gI06hY4CWpWKeOSu5r6J5iry+aGLRwnYfqaPUk2HKqiCkx1yQ/4azBn9w+JrpiYp5ctvYmnfrRi3
eEUacyF0BQI86pH88zGXgGTcHuG6n4bWs6XK0IO5QnZNwE+j+bVQAwuhrpbq4m82yIpuwsDt7bua
05ruumXUjIAX5tR/owKwjwtVvfP3gcWYm2ddwBuhUY0HMeZA6nEgF+0LTfVospOA5mhLGESHCj1+
zDzpqGlKWt18nL/X9FgtWC4dUxd2h+7Yx471JXqTxoZO0ELTI7yHU34lAw6baAB3+9W0zwLHsISB
1RVQpib83ITzHYarctJFIjOb389WOAOZvxQMOuB0VKammiwZt3LwOjf8SttZebfq0Z6yCLDt9Zh0
UWNAJPgkRHdFlpjH+eQs8akbHYMzqUwdyvZZhpTovPJo8QWWCPGx2mMfs9+2WW0dgSJGCRxpiJEX
NiqUN9BRD/MYwnVtY/zCqz/r2jHfbtt2Q9OA+4XjAQ0Jctv8jstUd0fTeXmWV+9jI/tp9FJPldka
0AP+DA/DHFHYdMfu+xVxvEwfKlT/oE+BPZCoAfV4fPAwDGAkSSNR0YsYe/YQmH2/7Vm9WmtZaaDA
Rp/h3x9n5tMJMZixf4IAYQZD7KIpLaQa0Bv75+N+Yu3MLemR4JI9DWnhHeCFh72QElnIvj/0CBZy
RqGYiL7AbRotCTr9r+clSnwyWOvX8REUOkovz+M5ZK8I2Jl289sq8Ov17A/CsiGGYhuFlyC5XSI1
Z85Jk+jFfVnpRnB9gb4hfJab0ufhdI7j+1DGgkOn8LepLXE5+y0A8YuDOuZ6R9/E9wIGJ2p02sxO
7nFdli4gbYgmRAvCEaicuO4XrOPIkHrTszRCET2fcNarlcSxkVlxcJtAP9b7/ouVgnAGeEEuPQPR
/lHYsvnBS6Zdv6Bx3UNXXGMdDQxDu2CaGuV48nTS2nwoNfmF27/KC+q9sWusQuwbdDxLepWja+Np
y7ToMvBvCoQnLZ4LHSESgE3Kx/QB4vy5VuWMafsy7A8gfEDxzaqjvZjU/iNXAYjkNuPF0FvlzwWv
jt6+mDRGfwjzOtYP3uD6SYz/glRUWHOwZ+KK7apvmXdMHCT7nyM+cXk+oKCcUzDNX9zQJDvJ+bBU
+vbpi7m3HrI0GrkI08IzwEawMkGdr4Key13m/HKZo9VajwC8Sc892i581tbhTITpQlKxdf/IAaOF
RyTDddlTQlPbN/X3B3B1bvzFJWRu56RkOdZNKvVgvN6H+QWvSJgzOfsgMWXxPfE9zYqrysIRtnRs
lNXyXQ5NhLFt2cM9TdGUxXFRGg6BnZpusJuitVuLTqdB142GIDrUWJNag8anRNauEKyzrsUbGXn+
kyKOXN2jTw5aI2FpEJjUNqs1x1MDBh4QCAezshFvOJMSIrUrSgxM4KBCjK8zt6++QanPAY/ZjC4G
Vbxx6ORu5ZRFfRlDugQmYTMybkgYzuoGojWBuLFLJ+xKlqxwWg49jf1vM+00I8HL1Sb2i7ap3mUF
Jql7Fkk4PQ8RzHW9F0V70NwJMeyA6zU44CcQ9oa+aqwvMSHD1IkB9/tUnaH7PxnWfw/AYOzBBasF
pjRimzH0Ze3iMF2gyTGnxIMaKc9bUjl1qlDh2S8yTToAa2Tr9RqHA3fO4EzAvqJfKbhERUxCBqB1
pZgtgchWz7/d0nPJtYayouP3hDPm43ezKdEzev1doGOyvj6hJe88rR+ZRhkXJ5eemWgrmuAFUAqS
KsYRPkAdhd8hcezScf4kFAMRBchahH6ePMqIqPyjscNX3yNgqYrNKiNLox9Wp4JN+F9oIbKwjjJt
pRUSOGVky7qVRM734JaWcXav8EfVTi3Jzh7SR1V4eLC/0eLG7DfYe78utd5GZbfcl3hQSXn6IiAP
fTy9MuyNrn2y/pElMdNf9dIPEGalUXki7BIWyitas+oQTEJVz7kzP21LtWzFfpcgT6fEeN4JNpVy
yVMSDpqg6BbmY2AzJwPOfbiP19CRQ1OTab+u/9CBSQsSfiDUftCwDKLZIkFufPui+Oq6gy25eonS
NZZdEAOwQxulyR9dZbdAY7QsKmrrvgsRF1MCGsfWkHH3NDEvfvQoIKmu0lWK3TVRlwE3dETMyfU7
652K4Vm6lnXBXQHnL3r9PhmJKvlrnrCa/vu55j14wKjEFLnlslB4WsYizmVQKSFGT0PkKUNchTsr
GZNZjabsjdf0R45QiU2SaQirj9NJcw+vSbiRHmzpMa33ssBSyIp4o2CuydppiN+QSsfWerEDpfzP
F+IztWFwLoE17YHXG8D+JuOrdliyVehS/7OO0pDMathnd5o/juyERtfaweuKlyptD184cksnf+nJ
3nXRE9ZFJU3X8F0+Hr/siYtgwaII/t4H1ui7xpQVJs0R8Bag/vYujCVcmbXm/feRN6tWR1Yjrx4O
39Q0bvStOGGx0A4bILSyG7ZvLHriJkF0+JzxLmB0shoSuI8yoLiqWwpDuf0kJ5vSnPh15PA3hIsS
t+dZFwZzFZC2bKkX90/pbky2/K2FjlAvhYL+ODDf6tze7ghfT2HFl4NgUdi40DXKLKnkhddX8T/Q
GRUrFwnhpD/ejM8ChztcvQMFMZAcYjpFhHjr8N7znGYNcArGqRGAU8dSGSisU7ZFb1pDiRxZzdKq
QSIv4GPIhZaY7enmG00I7xPTYw/mpVwRLXYQuq5gueGGHQcEEaA+Bm79ZeobRqzL4uShu9FIjt+h
gfGRdNieRLQBEa5/pdipqe0fnWocdz0XuZeFF7kPtv9p3ZpGJR/r+OAwshWgDmkv1e58wpBZQcc9
nkYVRNQgPAi+RQCdweMzXnLjAG//F4dNV7drnDldxXtAbGDs47o1B+JnSPjjnoz94pI+wb4ICksI
iTbcaFpWgLiks6Wggtj6kS28V9PRa5YoJFyaqbh15o4W0cjt8ZRZNMzWwMx+IYcT87ShaaaMWuao
q/GgHK7exavqJ8rKVVUMCQBZiTqa5L1HgxrDDvQjacuorAyWWsEAgllWTIajUHYCwI1mwzJVSA4a
6FSmXYX7RK+vBk/dvVnzOCozVr4g4xw2sHdpIiTLK2IgLMPSADMA5uEJ73M7K9NPB69OC4iWSJgt
Izfpzz2DerEJD1zxUC0ZrOUbp+IH6aYQKdALOpdkXUEDddqAfp6XMPd+PDHMCKyHk4iKm8/RT/vh
1Xf/yzUgjw4j7pjYiIqbuKpah9Sp0S9CrjQfJ6a8H+4hshYVDEyibtpTH09S2b+6w3V+NR/0nVMH
a9sS0Yiw9EijMU7Ipbdb3xTRkvkGiDnuajtsu4nhv4/IUjgaUGEpBkZJIDnf1XBk55nVKNa4uD7r
EsvEJuRIUfFv59pBlULeTZ7bwzXJI7iYbPKvfF41AQIyqQUEYM/GY9O04EYwA7DlVShrRfcUpr63
1TIz7OuKPhUM1dyVKwhZCIzK9EO9Sx6sP2UsloUlVYN4ngRjV1nBp3OuEi2BWxp16e68oR4Tkg9i
ANn1ThZ1G1NK3Grb0Q7/vUwolB2pfgmpwP+MWx7pmm5o4nezkEd4BCK1Wus8wEyWe/QR2QgSw5q4
4QzQMiXYVVPTMJgK8gsyPH+4Etri0tMn8kyG0/PcUv1ImEXQrvxblXdMx0WuzUXo7n9fRBZ+pE6E
LvI0nKeuvJuz7+/CSNAogAl9q2CEX+2Q3no+e7yC1CVh+NORtaLTaQjTDoNxRoUnV5MmexIQc8Da
9kFPiwAVe8VvgvQAmg6BGXM8W+SWavJ8EzIK1Hokzeoh97diNpUHrrExfmoQuI2RPap4UmcGYsg1
tdXLs1BgdXwwx8NtO9e9aYGOM92laHEaEmMSBdT5gFRKhlYWRZoPFykIfSKFCAEwl9K3i+Lm/HN5
iqbtNce05rawzMAwFR/7hYeutC5mtSSFzHq5cGc4qiXrDRKbodSyi2IWkE6Q0qSrab4cwUZu6kri
Oq+dUM7443sM8EW8kJLTVah/4vH4K2cPIIpt5QxgRc0k8FZlLMjfPoJEVXM83ijf/4EHkgKwDrm9
OZgYoA1iLMI/fWuGu0NRpZMMhLQ1Z1dsToKVCzEZHrExsTg+BSXIwgAga0xMiYGBMiXhquEtijt1
WY1s7aVVB5NtW+EWcmvryUdQq4067KuXvvb5fhCHf/PpD6ChwBCnCC4E5qOWuH75fzL5PrbRWSJR
ybuRJA/DQaQisUhmipeuIRjF8q0l1DCXmSM2CZXErsaNdPUsIcoW+gnWUn6rcZ3aCgArd2K7Q34k
GMghnvLlbzDGGKHgA7+5oldeytD1JKhtRceY14NKp/L8gaVurMbph8YiFzszRPcHevjKMRB4nWut
OlyAvWqIYS/FfmcwacbJmrzxagwyEEjuyh7eh7fepM3yZesCB/tHm0ir1esi11Rrg+tQ0UbPIbUT
1hPX9ZcgA+aj40oYEp1opR55rNuFVgBSzvOGdeCle94bCPzz2uExIy9aDSYPUgIIEbag/BhPlNb2
BwtINHrW0cHipSZh438Dca+KpfFNeHM4O6b/LREezQGwPmnEiBryTKn+r0axPtueWK9NQpWFmjpG
obtXU3scEWw5TCbNybHay9GyNTWB9+HiOnIFUwcLrbpzoCjWwxJVHtd/hfuti+CUPbYIPKSRWbtp
2AZvSOlEHBD7m+RvcgDCfdLLWTCZ759XTOsL60exPgtyqsFf7qgG4PYUeAlwYNPrUYoX9hdyI8D/
X1uFdX8W+HzFXg6EfUVa9Ifw3oZqj2+leYCFFTKc679RZUNrnmhngtAoaexpq4J4lMGqzq/+7kpS
dvvJfehahLsEpe3+o48IcGZ1k+133aK/7TDGJ7J6IIY3fHNvWIpcFmXmNrDcwe8UbGkU6McQNvIc
RUdgOsKNPhA/rEZg4nYFJsmw48yJaC/dsewHb1vWt3mPEX1dab1phHHj17pPDivuqyBLlIhMsfOi
QVc2cy2N0jWiz3IybuEpmYKPO4HfQ+0oWgkMOQnBCjT+fVJDiZcIJrYLhJ3ayE+x347nM2K1qRhG
fMdf5ohpW9NKqlX93sjossZndpV5tEfi6YQTJWEvtXiydpydcCw/Kn+afZum0aQV8yymbXoJHzYB
f60mKVRR3vGXcE0hSYIq2u9BDhCxmPR6nf6nqTs2gTOdsDIzTyJJq7wCIB8CRiI6O+v2gUGR9Nic
jHiWqCrkLcbtyypK6mw19slUHpbKyNpO5l5mzgwx5Tptu5P6bu5UlMrBe6KjaYdlMTE8uPN8Fudp
rwkR0usv5DS7pKBTVgxcT7K95eoHbyOTkv1d4v3uqEoLsL1RZtZUfnt4hBv/V8WLab2hy5QX9iTb
Ti2NQvYuMTYgI1aia6kwy207yhKfSOaIxjg23rTQhAzGZ68pySAEsZ1aIhZVH9h1Yaahx106mo62
UiPgpMTA+uvRsijGVazmXPLO6a9uBtczsaohcpB0i/3lqBX7sJkz2UYYyjXRy4UXFpE5ScJCr4nL
GUiGEnsSFufzKKHC18jQ5mtuyQwfjSwcNgpj53D8hjHbAjQ2WND+O6cAUGiGl9bXxuLSIiEvd/k/
K4mPP7ZcPxA1lAGjjWF2XjON0DJzgIp6gUu9HQDuhD1c350GDqWUCkCM9rcciz+LpPKU+636ccb0
2oNO4J81etbXCQaYCUsAcTLkn+BzTwajA5YhdreTJono9cuOSn3stfH7+qtahLcGr4Xiov6bcWHS
ahkitwlw3vmgVwv+GX4GG7Ike8seKmZKjM4myJDcETnafTyE+zMJy1NOxhqsHbjG4TkmwUWGJIpr
OfTgjQjxa+ayYmtxkj6gf6sFKLG+TV+yCu94f/pdYhEbMor/VvrIKKnzcXOWLDmFlTfmalZOEv0C
3r09UWiLEyOER0pv0bktSxNT4wyeZY+x/W0iLf9CSlK/qxBT+FD/NBMeKnrD9fn4sT/HFA49MXSJ
7DF9BOpXpJpRMjOKbAEtJrVQKCwZ7XWH+ZZS2x0hSU83cApCUO2BDAFRJ5vFlqiPvPZtksXJ2rEP
YbO4+LjIknQ146aNJrizscbkvfO3jcV0TYUs4SxFueuNTPeLoPibvDqVIZYIqvue+vFzEZn74Iod
Y0VL6EWXnjIzNLUsNj2YTZyB1+H10X1rNxChhtTdEGUh6Ag+GpNLealApv9SbZJCf5QSCaeV5mdx
ThDqSQvwayTDacmxeBBM3OMkTlsX8ymvLJ6j8qh6iNH+SidRsMa7VpCDt9LmdtThE4AOSN0cM5Fm
PndPc3DPhrEZ1FE7Ip5we9gVzdZNmJmtKAGuUoppJwZ5azBg7vHxk9ROpw5tRaGySv4LazACC+HL
okj8xMWnKukc9c5tuh9BcAT+W8j18LVts6D6hwxW5LA3epK0e3W19gjEI+44pwifIpi50cTip06Y
u12dqSP926NLgJx86OtPVx4Sgt8bjkhNJCsqR/mvIbKt/AKATxIz3Ee1AB00T8DLoAVoozM0Ityt
3kH36JipLGES3Pj1YjOOL2NeI3g4forML/6FWoBKMD1uxpc5bJe2Bku5sEbYXg/JSQBGceXklZAC
3QJowqeB/99DNsHnEs1IqzVOQJH1Njb6Yc9QbsfFJAs1vA8rd2rz7aItkMlYhhpp8GjHcWzYE0/G
QOoOB3vXpeiIf2YfkLbfJHnE2UMmaLFGyIGb6mwCCFyNwloPVe+qN7noW+Aly13K5g7m5g/kqodz
mfYWWUdnULxxzz3fQRGJqBpa2rTdXc6vAqrjRCeilCFqOSDL9qcHOxqj6xWtbtpsCNuIp4mtjfBU
IMAgtHH6uT/XbfMDOD89/rtYv0vXslCVVUnpHxjxm9T0859aRVB/yDXArxEOCD+xyhQ6ywE+PFjP
o57IjQjci/VRDnVAPfugpKFWJyKjAInDtZFM3L5IbbEzAxndQ6R6c1qy9E6zvNpzFlLr4BHf4b00
a5g/j3FhSWR5SkfPfYUcB/mmjQdwoAYXK+phOm8OScbC2OmG/c1U3WFGozj6UOoQBwf3N8u2zIBM
bGyG4EbuGI9NtXdpJxNQBTgNPdJQbqF+/cP66jhYIj4r4Ff0bSSs7R7Ogu5d0GrRwKmdhmayd7L6
V1cjDDfDQT2NuXKA4srSOfUv+q+2dC5PYLFdA4bDr0pJRaVfV7+tJmzLnXR0l6G4WDuGGRj6r48h
/pMfDUV8KcEz32cuJzjgpsdwTwJTfoDfqnHSo7dvv6ebJ0yw44f6wui1P/7p6mZmpL9cZ56Fxu7L
K0BprDYbmU6UrbiNg8VSro1u17ZD2Ghom9b9Mweivd31uiB2xGU7VNbQK7Aarhslqaca1LFnnTY4
b04tbi3mNRXezstw11m7wu640nGBCWh9f0r9RZc6B+qjROU6h+SexsDuL4xq81VEr9T4HdzByoD0
UxkgTBbyPog33qsvVK5MyUZMRKu+Uh5HNMsfvh2NhrNaat8aHwAH+wnw1X4UmbS+eyRFf6sGDv3X
A5c+JAHjNIu7UK6RmXQFaRJmPckEs9xWoYeyb5uSaD3qSEvZKEUtwcA95kNd0Yicn3cAmqjX8PIx
N0ZdIJljC8WLrudL7Xxj+23kmNA45BBNM8OPf1tT17AXsjQ7pvxW1sdDEqdkjzpkzHW7sNWqE9mJ
vtaeNE9IcSOau4vph26E2KQTuVqCQ3lnnk21Rb2gNtkLVAbHknPSvGstdn1pCj/vZqUcs59JaxAr
+VrDlXFhIswVNs7fOzEWlneIZbY78WCN/G1uEGtEUlMjKgzTO7Xy9wC3xgSFVZvUe51V3quHyG5H
QIjDvb8vo5Ryzx7lIo05rREtYHQ76wqzHJZqfv9148On1GtcPga/8bn5pUceZ48GrivjwGIQK7wK
Cq8EZl6qGoLmtvW72gvwgXtGVFy3LW9UvVmMnVmPxfhaGFW1qXxAr4HxrVB109G4wRQBRTvOc32e
hNnMnKBbxmIKnZ9/2lZnVEFOnx+HWk9w+Hiua+rlYk3p2m6zAwJ8b+It4ac/1jG6V7diU4fKdBO9
N8l452edzIwnmzMKm4kQAIe47G0I/O3vv1qzoAwoK2wmpTXmfmhvSaLBjoWVX9J6qDCH3MpUITA4
tbWY+LMclWtV8CyOTk3YV/2QRSQGmV8J7xIhOjaNP173+9iZ7kPb2iKeSskwSrdrG+ZZ5UM27TZN
GfOjVlwyPn08EHKCdwLz5melLYAJJslVlkj/Z5NeAaImSwXjliG7B6wtSwN+TK7ebwHHihJy5fGI
yTtf8eVMua4rkVW89x022s4AOy9UzxCQC+GsMfvfKEYro1eQktJFnKRMCdS47h9VRXQUykbYs0dS
JJnydVRp9u9ieD3/OUWyF/iG2LmoXMJdIFJ8ymAh3KZvy+dEK90JYKr2EwEnmmrXn4JhsUWJISgN
o3sBy8d1gLBFpbrx5BWWvCmv6YPGEVcdu1w+ZFPxY6Xa1XMn3CiG4rOBGxPfkVFKK8+kNcU6NvQv
K7ELNDlm47u5nZLYTFoDwigMJjCrwyBqgwMWDSzK3LXBondoTi641ARfwV8LyFSj9RhgJh/mjP9B
7+de47gyoDDJKr6n62TwRoRe9rrgdfaad8rrLfhhzKZ25coJBHCoYn82PpyPLZaWMBQszmN5/OLq
edSMh14K2n034JS39n9A0jtJy0FnHTa6jBWs/2wcx0u5FiVOsMlNMTQOq0N4Zm6Vk+r9DMvKeUCm
IuKWVuaADwNvKPKfzk7oni0zQOkIVyutLGguhTixLYmgMC3EZRW/wj65DirMDRvTRqdKkOrntVRa
HXLPaZ6goQ98TFBFHhlego64jAgihFN0QPBGbdkSMQbRizmlNuVXePm9U6gL384Aw08/7Egm5o7M
OeyaxVFwo+zoW/EA1PxqeCMM2uz0SfgN2vOxHQMJWfT5NXmPh+9zFMgfk4TYBGVgGpt2dfMxB2KP
XqRYC/M0iEb0y477Pvknn1+jPba2cP2c+Hl1aLZtFdC01wG/XpnqxxU/c9Gl5CYfhHQ5KgzPy05H
6VA9r6BU532wGNzNGkCslJKKPzsz3MM71KRAVC82HZl60nrjkq1Yuxw7+OVQJ9ojpfa1RaMzUW02
RKV98j5SGh15HLfa6IDJgxvr4ySxMzNTOa9mYYQ812ZcXMoRU5/PG9drYs1QcGMv8Q1r+vIKd0kn
/KY6vTKY7xzB65zMMmu3p2vizo0AT02CQc1fYQPM9tR4LLqoKwdGwps0ZL4LmbjevzbGi8f4ceCQ
VmfGufk1k0LvHrmeLoXtxVvhsgiG/hDJSju6U0x42HkI9nSObpqWNALfmttCh4xanGOEfSnZvgUq
otgSXs5+QAMLMrxvfKEJ9C4LTcYNlYu14Vp1+EVu/nh93bD3GLUfx4vFlUi8qh+VBgp/bIC1LFvA
7z+YU8a2wSOn5UgLo78Rkbem7DjXRwWMWcdcdKa3uHetIQbvm/+1L3zluNSpjwH++cs4M1E3Yy2G
DAOgKjtQ7BpPWv9rLWEMLRyJsd8Wr2bMEe4vk2GT8VWIJ0fYZG7xXeVQXNz85GOsOMBkbhzEWwWG
fP+DDCsw2xZFxM2BPjjSDR0LDl8Y1wI9nU4mzqaG4EHl8c9hL6G0LRi/hCO0PeTKAdqph/gQsjBJ
3SLKAuX7b7IS0uif4CIQVP1ujW+JYeBjPKlpw5jPbd78OdR2A9bgIcdeljKixMIvjyhdoJxsX+QH
TZGZh2YJFMNebX7VUOAzDVKm5qbbMpxI0FlInArUnRwXLjPgbkJoWCTCpFw9alIbhtKbT05UG9WH
4UbgI6vDaP6Lnu+06zeu5Uocn6fhG8tgE0lr/+OFEb3r/ABIgyrDMZdeNGHeCziPYgYFGcojr/ze
SlvtmPNR9dRGsRb0RmX/m5k/QrEyfuNpBTad+iFF1oTc9lDfLfoTn4F84E33V2kHdU1ELKDlpi1L
adKcGrkLf5q5HM5VmRoCis+YJlmN9s+GbpKs/irCT0BJKKYD7RV/rjEKFZwVMuhCz7GZ3V1vlAlr
r/icUAHCo7P3DMGThTBwQJtJ+mM/nx3duvo+RDV5aUD2WLnKGPAzN5BQTgy5L8Uchh8vL0s41f1b
tOSMf3yH7c0KGAxDck71yOOTBJcXDgTCMOTW9fj022wQwfQJ8RVUL1rlXdLWLIAlYbgWGR2TEqmn
kewmt1mkti6pLJjFEJXDA46lOYjkw9ZYnTC+7qS/BO9vsVcXRSbhARBvFtumK79wyL0Get3EqOag
xwvvMdRWf0eNzhyjxoXMhKs8vli+Cs0kZr9NNI0ztj3qshM7p5bHWRxB0UvUBSG+brtu63PPT9Js
9LWEsSX6s48XgfL84KF5CEVM2BEVRnlelA/Ljefjsb4+upDgj7pkuKl7IulE1z1t+WYiCXK+qgfj
beAVv8m76Guk+FX5aPEN6xeU9vnp+G3f/29GBUxuP9/W1PpuNfzSa4MvOENR4xpgyD4LqfdtPhto
iKKoAlqxRIJL6MrTtv1OiMgw+p6BLbNeqhmP6o6Dv8jd8osWbmxZ77bonEF485dPEeLxVpUwpwcx
w1Xi96mJSdV7QHj/v5C7BFmSNqfSSbwoIHUkYgzqjofXUVNh5NzLCYUC0qWV7d653oOlRDD+kda+
60bo1CZ2uwIim0gIL+aBcIjDEP6zFRyUTq+brIUf/jGrZz+SckDsqRmpie9YK5s3Ol60yu54CkDj
+hcHo8zqhV/pCkzfURgoV3+k01YjbbaZjNvsoJNEewcaNDSbIk9b/9+LhODP40NpxEk8CRlmTEG3
2dE2hw/ksAYZw+0xYpQf4rIZrzXCk13gOBMNuEyLCSBCUqYdft5PfeX7k+f9KjmmNGXGCDcH5gd8
f04xoktzFcLgzRYRrKtaqByn/Gc6boRWe7qn5qi1TjDhNe5lIIbl6Gj91zs4LSIVoIKHOz3lm6fC
1cofiB2ZntXnOigFLhpbbAZ4YT5FQwF09pfhry/ZCsftgqrrhsYVadoQIN8r9BUhz6nATskL7wXo
SQbsrhRK1Cx7qQZhEvaLIbawzAquq3u9ODu9CM9/nVhmWc7dW7We5Ay+khsULM+6q3ezbA3LUvog
nf8E8uemfVeMGiUKqMDUQI/yjB1REqy3JkbYGqWNRmFx0sFMBq1E6opiYoF/fLRRYQU41ZJMNK1q
KYKVHA1AY154MorkS1EqlhUtXYnjaCzWNmRgOicrFaDnVulp6FV7W+r5q1x9ZoK4XTmxJIOMXKBL
a/LRFf3daVFP8xHKFisPcnUZWAkUQqVd/r48o+4+PrLz9+3ROYSKUylDgVq1ZmOvBajOgwghYJNs
XqIr5/jXU5WTrc+kbGvIO4xXRq1Cydpus5ABl0UHpoDWK1q77AzFFfTxHQ9bLKGkkkmmmS3eTQ5u
n7k+D4WbtBhCGRq/RZVhAFUcamPEOUd3iPjz+Up3lAarf1hkEk43amXaUni3UuTC3PrXNKMJrASK
b359B7yG+2b/xF7FW27rrpRhyrkWHgKvTejMNSA0/L7Y+xy2SfOdgDgPR0/3VHwLGLGuu5aw0twk
/IqObElfkVIvgMzwhoFjMwgatpkJkFdX2mYLILaYXMqBer5LhIy4tN7xoUMVh8e+ATjC+6f33q6n
3pxIZM2+0prh2mDeRgYhhCMib4jpRRa1g0SFaVX2N49cN5VrqaMdwFGy8p3C7glYbRpq7d8MDcCK
LbXOgTlHA69AX0TQDgByhzDVkWdAcds+OhyL+zLi6AXzJREULdYeoKSgBPYgiHAuHaTY7mYeKl+P
jfp4Y/L+xspa3xtl7hYoFP2vrrc8XYnsBDcBlOeOfwrqiOFoOXjo9NNtcXj0Vy3d/fyoCT8/V8pL
8R+et67WydCsjxkNX5k8hXZlQAAOFp5XBZoqWIbUkB4CspsaZNQRzylzRxuyCtE+68qVOV8d2wyc
Mg/qkGj/j0jK8xBCs7YXF2BWDlh9u2iP1f1P59LA1wOK/kWAdPphWvVXCC2Shc4gfIZr/VE04IbI
SeacSzdNqN4KlqzKBaU8NPqYevJbKVUI30PUjCbva6J6HV5QdleTaPljNB3YFrp+YIh6LBS8u7QQ
K1CyepkHvUPcF6eUnwqRbGOrtsR1ue4NTcozFmND4YEUouzIlb+wDol3AN335sVyZA1lYWz2so6u
fEhkRFMuIYkFzVyBUwjAFZ1cTtkQWedWNpuf3TqLY9KN6qlg+0dQxv9wCsdGp5HZ8bSvUIgiCbng
QPpaTkfA/FM0bMd+S0MSG47628I0Y5eeblPWY/6teqc1h/tl3avKayc3wSdZF7ljpir7mmKGH/9n
85vFUKxbwftJXKI0aWhArCnOONe3XtK88g4AB3/Nh/o4I1g1Y0iuc61TeamsXcw7AI/SivQNSPUl
fJAdkFOef97q7ulhzAkZ/O8v76fjTYqdFxNCqAwxuySrNyia5xOpWWXth/UMVzGly4mf1OqSkUf6
tpJTkqec8yCfBfv0del0Zz/oCXeTagTVDE+f1po8/hVi+SPyJbFYEloC5VwcdsQ7bXi5uTwKt1Xl
c5xKhkxLivlAL11A/51VgkRDUuByi3DhF8UAXUGBzLYwFWZ9HOiM96QN2D9iUzCz0v45Jokivmer
oLqwv0nlHfxXBCQ1GhGUBvrZZ/63ilNQdgov2WcvxD7vMETasFpomr6E1fMRL3KooRUvQg+/adGS
30BnAKZg3nRR7xRa7euQL4ikQd/9umwwxx6c82BzuEWd4Q7ZYZviOJ6M1AI4ACHvCgyhtNk/0/JM
hxcxA87hgPZxCOOzBRVEY87lL/ruzlGs4vu/oPAQyWxPVSZRrhn/gUnd6M1R9TiHVIb5lgv5fPLn
U1gMJ7gCoyzIAL27zmyKncSUcvplCRNimKpWyxv4uutsEamEZ1psLIX1ORPlYx/TnVN9XmaAS3qE
e0/eEkFHd4KtvK2vUYaTQshtyhC2YtmmqmXsQSnU4ySQRVhXA9CKCx/YSpH4rT4QMChC5BnsMvkC
VWeRR1ou7f35Ct//tXiGXzyxZLK7qgQjKoXotKqWNLL1jZR81BzHpnf7YAmtDQ516tYtzKPzxeGu
5MX/vGkVpdKGPtvB/9K+G0c5wg/zaNtJEBXf7g37BDfwL1/S7VGmunibtjj02gwpZ7epvkmSIf36
VUbpdltQ5XWXWhziwpsYM5RifBEZuyVSZ4Hwcta6HupapPIgpTQLmT73t0tX6t38wmz3cdMArhH1
+K+tuBnpngf/M7iYSjXBGVMPVHc61lCaQa/G7AJSziaBgRc7kN6llskWxyE4D0V/HPMOWv525iBf
8Ij/uaOckptArb+D7C6b+o2KIl7A5heTRfHUSgWmzZCVc/72j4v/5QyekPat22dU2eHPGcg8QzR+
5cCTRSnNoBNGbxVswICSrgtp2uPf9v/cBV7eerf31bOAdXM+KK43NPrkO0kTnkAR3pUERLCNJJhG
eyo6bI1bJqn+K15VKz1GUv++CR4LxKhV6pKIHv97y6J1H6qvR7KoPE0akgYxFqmiH2CzzTPwZHRr
zQeHrEmtKQG63u7PAsjBy+o2/pvyvQFOOe8SXMhCflDAl1SWgpn7IykMzWudYDphhX3SZnVCEJur
Sg3ZZY/UTeuChpGxzim4MirFg4n7BPfnrZ6FFyOQBko9yQf03ZnualR40sIztw/yAb/yWk6XRPQI
5L//46ICFOOMsv+LoSXKE4/+LXh+ltp1hehxRXuE/hK3DrAj8cVBCuizjfskiO8yc93yNbFvTqkm
pQkdOTcKrVPw3tm7BQDXR0d3gTMScZPBk0ulc0nujJ6DCuZ3aPqHm51cA/XMTOfA8uLA39wU841A
t4hh75AUgOO77kVDmBdf5Z8CWLRcL2uYQsx8Srr8sY8+EBUkSeNSJxdGnUR1P/vrqQrpiRYvkUp0
d/Otc7E4LZjCFdCNLFkvbusCZHJTo4SzoJLX5dkQvprM2n8RZf6A12lWNIHIOLTQe7GWpjicR5qy
IkrlZBf1EBo0JqxkubQntrie2NNs1n8ISJiDf7RhEFrRefN05TIAJJhnOs/JGXUc1scQUvANTaSt
/JCwmeiYgablIbSeaPj+JQZ15Ijzs9vJZUXF7J1D6/Ck0qT6SBILTRWpr6Nw8BEPHdyIwnPflU6k
OG1WQ1nIZ6hX3CQmBTloV9mHgew7JmLjA9N+d2aAUoWjHQe1JvyDClkZlNrUHNLOs7cMegdO/xFz
a8mORT+nRNVscehK+FQbdQuaNAuJOmls7flye0tnX7plHb6UbA4OWJhoZnZsauFn7zFpcQt2YY6E
pp9DZYShftL79FrSx4QuBwMgNaabh7rNzsZBttdRDTffnDfmPsZ1Gb7eiikaxXBthRdKtRG5NuE4
CZUJuYaNQ8CGx14abPa8GFL7DySsbn5T2id1z7GlNO9DfvODXmkYLnwlm/fdRlZyqI6qTBWJ93dm
lPLzuH0g7ARxjEYZ6LuD46jq0XIZyVze1u1N6p/Woe8JYI91HVSeLGperXzJ0SfQXRBN9gdR9xBp
52A0HBXpeq/mVtfz9HXdvD9GL8/SC8/9acEKEtS0jf3TylTV5Ze9wAHgF3pH4gP4L75pIDhQPviR
W4M4uh2x9B8ApIHBF9YM61kb3VxTltZygv12AMcRn0xfE933MwcxgNYm1X4ft+dNaiMmaydjYAeV
jVLQyDag5f9mvKTWE07A2VslNtVpg2XuF0sdF63SvPWt5t6SOjV1fzHaYCardgtdyF9BPB4E2uC3
7ncxkxec+RgPF+jLeEhu0xENKAWs8KGYDOxxd+IypoKv/0UKPXnw03um3LWPFa/9vlIGS4pfFs5v
VP3gwDtwHWxH8YTpkWerBwERqJD3Q2U2REUWeLl9OZ8le1Fw1f0BNPgwyQ9sqejfQM1g232HT/f9
X4qjK+ox0OdLIsyBI7J0exr1Yiux7meSeyxvXv/isbIS8qGlANq0NbCgKsVDsNLQSe8c5ylCtiMG
T955EurKJDDZbm2TtOiK4EfYFxe5k/Z0swakp9qtJpqVgw+RAQIYk3GkuWClXqZ7/jRMVQrny57l
SfAEeobZbjvsniaDLuXdx0d8pFubnFm6Lu42GYP2N9WOhvA3ioAPrXYMh01svzJwTp85OaHSrLEj
efQYR/kRJ6QVDRfhKOSE7e9t0M6aJ6wR92MrEKLXJ08eGmpVoi9w5n09YCkZdvmgCcKm+DoiVOhM
l2MB9x9L3/2pSi2d5vnpkB2UKLyPOqkpHvBjsRL57ZGebRLivbsSRqT7cGXgfhSLTRfjuwYAXHOG
PTC1CwIt1LpgBqKSaqqG4IGihfCENK0/8AiuHJcB0ybv0JHis9K8yzemejq3eokfgou0lKDydZxQ
YFBuI4D61OnDrZVWfMLyUbJQaIOrOXR50cfyQOI6iniqBST5vk8reaQ9yYLhMFFzJSlHSBG+c6IU
Ys/n2sQ5ct2mXLV2ZoS2dxgbeIqQeIIhz8vfY0g/KwPzwsoDy95jx3ZW3ROKDKzBzsA2nWNjebet
3QJiXouPZUo2EJhYteRwSC0EwZeKWUa67Htmvs+AvqfmjYIEd7xcdf3WtCB/Y33UOrS+XzPHqp/O
OFJW3DclNme2GC1kXQVdeDz0pn4Frerx/kR09FyQqJ2h8LH/gmNHOx/nG6X5qEDVjuziVzzWiiYn
uDvuw/6CSAzHeJYgQpcVVbT25Cls0/Q9Z51XjH6y/Uf1XIccbe4d/ysKHZj0F8gpRDwG/VFEDQHY
wR40LQ98WM/uz00Vfbz/L0oNvQsQUmH6hJ4y4/kmojofOg0iArmj4ToeNikaBbQM5s6lf5L+0X9j
ZzwayKZZZgbsBJ9Q9wVt0tctuLTG9rF66Qezx760EyVjzq+6vaUQ3VGhu3I5B4oqsCw3g7DAnpz8
dgXiAXER+uuajbVSN7i2ZnSssBdOXNsm5Izf9mghuWdxEZMB7VtEUKNKGBCjNi4hEXKvlwYShWcd
y3FntlOs5rOoda+gfv289IraByoZ2oeqSkj384o9MpJK9ZT7cNdlIRVW6CUiTdccc1yERj3AtRtU
ZAzr+7bUBDZYNwpZMGnXsmjyvjgOx3TyYbfdzE3ZKG/rr2mPNnuLXev9lbKGWNzAEdqXsIM200WI
pNv3bPlfpGQ+2oHLUgMsHCsMf8X4qGxyd9grW3GQkKHPU37LltbPc5RSV7W6RWCL3WkqVeZvOTb3
E19SRv2kLRvtdJARcvpW74Vat6czIn5gXXToq1Yvdum7LpyBRCD5Dx0yp7N2eCjKqAnJbzLh9GZZ
1Se5/sGnx+NkiKDViBqwwe65WPVTkJGRkEfLS4YIWGfiOLkd1EU0zrCrgagBdrsJep95rJF0WQek
AhJkKGsdL3XD3WMwP2RJQ0eHUCrPZ3bYUZNqgoa6lp1bn5FYoNyeIAp8aa0KZ2bgmMt/E+oh8l0J
uMKtK5IpQh4ASRXc4zxEyiFVSDGzPOgugKlDmI5rVJYT7+10qzc8u3cncV1/UxaeJ+Sh3DDpEtHD
vqGNNGRzEafVNhqlpyD3520sOd5y+vQT2Lc729pBr2WBC8HHh97KfqWRR+nV9h1ZC9PHrTCNQjpN
8eDSJsqWf4GznJl334+w+lgfwduVKxHoQ/NpZbwX7AJKTkzI+dsK1sSqHqSU+XkYewwva862uVAG
6J7694QnX0QiO8bK5zUCuKNaP42NsSGmKaw3vlhb01WsKsiHj2WFnY68VKj9e9KWSSAHwer9Y5pZ
NgytvOwXdVVAg0lw0z+sAeBMkWfqN+FtoZ9ooAyCzaxOEEDBWelOteTsaEgFUfGeQ35w07pL4uAZ
5pxWbb+cz7Ev9dK3BFBVVRqQtjhpcd6u7xRQz+Mx1mVlzEyngcrcMLUMacLy8NaHegljvmZPCPA3
TbEJLBsZ06bDY5ArFI4GWzTGbjPYQNLt4vvRprsy7WFkLCY4oCWZlpL9L5HTlumnIXRNmlcOQmP8
SVm5NNwFiXxJxnKPPK+R30kPlMxx2SUfoJ3+d0xfv64yjLUoyzLiC5Pwf71ELGyXHTVyTI75hHXE
tmYvo241CoWUJFutwPf+0IP4kIXSbHL05pZpWB6bqufhej8ki+tLmZfcRlik6GYDSx7dhqzjGcLN
s3EMFzuqN0LDvJPmhI6L2SMz32FIkUj9/lyLWav0yigA98KF1XgeGmr0CH4vuiWhvPybaN78680C
5JLxKtdEZlm7i8mzVEy7cptXK0bhozqdj8G74QL/irHb8120sjFli6+J6RgXTIId7eEvHtOB0WuI
cVxj+f3IzxouAJSTQ2ARGdYmXrcJp+ymEFiPGXqqiJjoea8gHAiptDblVnmCrf/YOuhPH2VCu5q6
lQEXoAsFl9tnShwV9vOu5s9m/h5F9hQAJ7QvPIlGW351Wmb28PHXAOlKJZWdtgdBnOG1q4xE9ckq
0T4XAFzWUEb6UKCyT2xynT0/wTwCN7bZUh2vlRnXWFWuhfXarxSwv8+MDW2BItUZeg3H6YSAXjng
ri8zL592ZLTSArPNgGtOrvPYHg5HyXAssY967Hblp87cFa60QKVGB81wNDOsa31y18Q8vjoKmJt7
mZ+mC2TGFiZxcTbIhqDSM4GsxgWlNHDGutT3BlZy9p49caVhBqqquyMZzp14sW1knZARS6lj2XmB
APyaYmmRLpqlJyoXCopMZ1b+PgMS1nBalweB+iYXVewj5fqks1DWqqzaV0i2YmuZ5Lh9SFu+eYJ0
Iubf+CSX1RqLlJTxZ3IYsfxFd4ABr+jpDiJNYtwSUXXQwXYyxWpKoZYCbGZWmIgLdkhnzflgTEO0
WzQODH5/A1XjUDeiIsogebwvM9lSofNWNKnA5etUlndWxIQ6RdyYvmKDCSLl18ARknCncTCwst+O
M1qkvoUUqWkfUGy5ywYSb8Xkt4x7bAsA4yluVMnXXHlFoUfyPv2j5W5u8m8giOv0iXJDSvmwjsbW
BXkAdpJo09ffppZ/AIa9l/OgmXyLJN6x602X+c6XobSma/hSvGgDT6gXir7IOsSGf80LJ00IuMhK
Lqm++BhHLaNpdQGWie3rM3UDo2lWCte2ZmIsHATsCgMUf4Jn60ruKp2I6VGJMpRezZgFrR1sV4pH
Zj4WL23rg1AF1Xs3/fqN9yRBna7a+MfQeqm0kS9eXskzZs3BXe6Eb0ZtQFexqNrm8UGbHP7VdVAZ
hwMuLtPg+hRkXEkhUcq67sBIISFekekgJR3xY6Z+3gufFn4Fhk9P6XyrDkT3dLeiA1MGa345uIey
F0lFX6N9H3ePGhUmgyljkJPC34a13dxZOb2cbWqt+R2scQR6Ym34OLDb8WKvZRk1NQigQtBjzckV
NeFNksuF9u7KK4bxeXYij4pQu4fgpfCt0lxjqYAqKopemSPMGtjc5KYJKH0XMxe2lgHZ1tPAFFXZ
1FmbUQgBE40GK6eRg+I+I1lV7cJOXwNaxcAyFq0z64jCLgfxsLqrbJN989Tv2lqauxs3dm18cfmR
vggL9aNl42V6ZxBPZDh4t2+aZi7iOnxHsgoSJUDPVOQt5GEvfYEvIY/xUBiYiczfqDJQN7Xcmm4x
KRh0q3OgXxkytjRvuXfyObLYPdJFBIiim/2UqGoKiN/nTl55B2lsOVdPojZZGoGB4VTdtmDap4iM
oBXp4vq8VEbNjMAluMGbFJypH0G1Oc0eXW6Leqk+CI3YyHDsyaxyRdW+DyZ5oVLLjeAT2INePKxL
R9iveswF2foB3qVREioZ+35+OVYC/W31nIByCcktrBvd/fpkBA/UE7TOBHgFpPl1nFYIcawfOyXj
+jZeKb2b1nRzW/9D2b0OeEUyO3jCDO2e9S/sr15e3jhNF7yqu2LVQ1YMiKMeOFFy1LizsBJxYcQL
U7JGojnMwIodZSKAc5pXlzVoPUm95fAFRg/21948k+dnPlgM7XMoNUeZHfYljtIJFScdTKVMVIr3
Oy8sAZAbngmt/eXDN7X6+o+iKc94TsQ/cFvjl6uFojFRrxvfUtNtS4OvRTs2y31fsZxGzifOuBLz
CCaJWlzfmz6OyFF6LfsnWrixFfxF1QOF0QjktlrRIiZgUB58giZs2hRxn55Av3slnO90DU0SplKh
yKwrbq5TqpappY2QYeFl4RXmFu90dBXHBznqpV/clXuCc8ukSaSGvP70klB5sumVi+3YQZ4fgXwd
oWox/RGbhPeDq7Irk5nWNYiwANSHWx9nzqt9Aj7U3pF6ikLHYTtog6AsGnqpSWU7jHeyrmK6b/5+
RNIhjXtLdSJz5Gf5ORQMqezfr4Y3ItcYwx86yGpo42k5Vn8LfAdGWW7nPIstHgf9O3jiowEKSDld
PdHVfN9G1L55QMWAnubRk8O5GcgGUc4I9lc89yZggOnqx7vfagUP1uY4hq6q+mY0dgPyTGLMtdae
nb1gQI5vS5rUpMxsN9m2W7D8PvIV4nESK3rSg9puM7nYSk73DzqbR8TDvn5udaS2y/cLzuDP5sHu
kh4T8Gl2wfU/f2Dlh+JaTv+JjmrbdMT5SlNXNlJQjR7+wNySWDNI3vGmPOEtm8fwBTxvfek7ZC32
ezEXjYK2B4aavwJTgG87E41xD4KejGoGBGOSQ7DilH4QWvTRCjzp3PNMcfEAUD2z7bc+sV1xAvwA
LKVGqh5Ef0DmQnYgouYx+sZl6cwqNTlN4rus0wdgzJhDo/zlwLGq7Az8rLay0/71kn4E1fHIEfqK
3jkI0km18HKcoDgbXgiV3eLZJCsaYHQS+85EbALMqCodbz9EMXO3oBT1gtRcEi5Qq6jCTDm3j6jX
42qadiZqpMtOy8HwYRcr4JLP8m7dGcmE3hB52iUbc8ahdYW8BRYMwrzLj1cJgmlW04VgCD6oINBH
ZsPWQPrw5BN8jR+0xjnMc1edsnj1NN/2weAuqkG+t8Sblf/W4XigEMcrjR1jjoSfWYMCxrd7/az9
zyIF5FII6MSLbcj8M5vxHSp+jO3uGx/zmxDMuSOGeU1IOBc4ydW/3Xyop77IwYpzsTeD47duCz2E
poh6qjWdTPtgXUcpqObMdA+9Lp469OY1gcGqGpnfaDE3tuvjN1FJ2R6lrqGqwDBBB+dG0mFP6uFa
P6fsCnGTGi92z1J/w8M/J99xwLeFycoHYMKEjYEjM20mvQu0aPiDhHE9M3B1pAQdS7YrovV9HKca
Hgbya54/AiLJcP3xy3rpQVj8u6K75B7nfwsh5L7HTMFogGBhu4MEbhb6QzwbybXji53kxhwM5ppU
4XC7Vk9nHuUqaC57oUlyMWCGlBpRmWxQK6yBQA4582buObKaubSezQWWgAStUouZdZcUrYFcPR56
tKMocdpZUjcHJghaIgKRkPJ64uNNsksV83jlS8rLglwKIovjY4uixr/Ej5bkyEuiRAuTR0UYoD40
mkTvV36WGJEAI1i6YZsjYueR33PIuW2Npn6luwX7bPkfZlpHUII17rFliQdyHRXGurH5GhgUTFwC
0FF56CvotxWuuIm1u4G+7/2+8uTFjoaR+X/8enFQz2Gb2yxwXhUaAUxMjUa+hFkT2uCUGuRYOje3
WoQ+5ED0rq2sbCyATNTJloGJwCh12YTkXDA/3d4bYtP7m8f5851hx71wQYNHEtrmm3IDZHyIanw7
S5M/PkqjLrzZEqgKh+RHg3N662Bc2GRmi0qowIn06KfZF6Nchryf9HrTvFUHUT7Op5Rm3scCnHF0
w6z2+5vv2RbTbVjATkyU+UXBvplpbyBtifSgpAMuolWmZf79PwpPR96b0DapUjZtcRairx4Ncqmb
K6h5vXi1zIMOPjifoPWgPvxTwVZhrV431jm9EGCKEcnWSa9ZDqoUDEAzcawFeiqBpD9upyTt7ZFn
p5/L95LkQZf+nyM41V0fdcnH0MmmtKHZiR8oDSUj7dBNvKT7rTjo1+a+JzcWA5mpJwKGB2E0FPuZ
GbQ8dC0vvIiKbWjLw23cbC6Yb8mGBdf3BEqI2J33lDWv6SH0zxkzDY7571I9HQ9/kaDIfNn6HKYJ
lmQOy8ivYGiAl23grr4QJXXAwjqvolBb6GO35A25rSxtOWnYjjuile19bDw+dat4ca57UoxNzlQA
jnSrwf/lA0i35+XkuqnbbPi8ZVn+xOqzz6LpxZpijKxZYyY+rzbbeZ9ZRCImIgwvWxxtc2/1Ujjs
An6kzILreaZ7T97nrWKhuGedhTYgdDhKguJgy0q++6NG1hyTh7Tok0rq8WiBixIqwVUb5ZqbHgTF
LqNdkWnaZ2HAxcHtb/aVwjvpO4A6+iyAr6S+YE3ClpkJSC+lFyudreaMbHtVibyUHVBVE2NbkTLH
kKgnGy10yBL9gXfP3sH7sXLutRj3kkubBVWCA1zCao0VQiJ69QoQq3ceTS3eIsYk1NfMXbBNDLAC
BPnaiZz2x2J9Mxop9V7nkt87V1HirPk8xLfuMbEYPVBIQ4Wjn+v2OCXrls3F9PWRe6ti3aEg9SVq
SB/pZh0a0emcBsMxJ903V9K47Ll5Fd2UjOiLqPw2k5rDwDWLsoLVB2rsvbU9cqITac+O1khzWqxu
FnbymEjOAOgFETKl7knDOV/W4GGR4NMG0+/skNZnBfxLE/XaLQIJJcgjsNApG9m6+3DQJEKF9Eoe
OTnvVmS5/SH6d8olQAkV5j2n6UXqdvrLs9vL4zt2kReHul4/be7uqLv1MhsZSXsFra7cxhwV1x8l
uOi/xUv2WUphCiqu2AfpYAsPKShowAVSTDktitGCdndVtLXbJ/MKUdAvetxDNWlUA/VMDNPuUIWO
0v8P04g2rfLA0fnOSuT9S0d9ASDt+eI2HyoKXUXIqoAcqK3u/jUxakP6Y9DojHho449XYYctFDk2
3TI2p0uuK8zLuN00jbSafiAF6VY8Kh/+NbB5hjtvgMtFxrNwTErWG41H25MEbFk7kUMamecYcvmB
nF5drsaFLKni1ZXFF6VToSJL4llDOSrD1fq9lfO0bwnjofXmtt8YfJggCn9lzDuBSOkomHPQUfIc
WDS9se3Fy6Mexa38Vq8V+gIw6j0R9J0Jf3TEIZ1ZaAdb+F1zMDpcnoUU4GfoAnIYhaavzNZayO98
m20Sz3XBGVrcppR96++pLpac/DgBoMDg3rLOP395k3ujb6OLyUh7WPiTcULMheqizPHPnoisvrJg
08aJLGeM+AYPtF8USJg/zgN39BErdrXPJiIhAChRmkQn5X/6geXnQzdv8YogKXH8tZmjjyzvR3Lp
KphDvSSoZoX/G7DcebGYuzs6K3jDHuTkUye51n4EJ5ofVX3xoUZdc+NRvb+dyyDkpcimSzGe/RnX
/t3VDQuPZxxAr6/MhDyA3+hxPtsLsdtMXJHh0xdyc1hLvkWeuM0bWMqp61mxQ6nyxm89+cL7iV7z
SBisTjZ84jtUpRMu/+UpVAPD1ABEzTxEFE/zYmdKu3gIv/vY2Xgk8M4lKr9rL7P5EJwTcyZiMt1l
EEMQbVgWfDCyd0gWaIFrPg7wYeTmN+/TOp7JuoV0Gg50Kd69ntNMx2RWwLBLTRFrF6vwLXCm8gcJ
Yp4dUGRIEsEzJw/4aw5PRv091Vyv9oPH06059CKpSkHVcAa/E9b1por9SECyYtXGknVLoodKOXm8
RlgK8Bynb9FHo7ICYv5q8TfppE+jGbN3rRpihYAl+UYykDn+fL8ZMB8JWpuVCO3P5ZxjTGdWUZaX
okDeSccw3F/73CfMk/6vyd8zas2I9nX+/ihdtKM/rE5UNrD35q2GS1rPkSV4+KfCFqkIZIxMwjZh
G+UpenUdFe6we4itV8lcfCLvOIi4+0j7FZw5frFsM+ZgT9zMv9LHcAiz1RaAwwgJXiVzAHuR1eCv
qUr7jr0wTUvkabpKelHG7nwKWu3OtxkNZg0AVvdexxcFbSwR+65icUjjfxWEDQWl4CdB70iVKFHf
g4SVnCFA/zN4kI6WesjOkKcwxNv442YaPi8BDosU1YoMmXBMF75XjK1yoJxell4/ZD94VSNdFRoj
p201CxMojOhOUNhig1u176xXUnHALgllgmR2R/Ra8+6AHtwY9PLTuK0yKEFpPCZeAixdPB3XhryE
MbWeagNvsCW3WknOqiRx74e9HEBFeCAvRKfHRSt+iQ7VrMLw04oq4yDm4A+w6x3xLmurCoLGaKrn
ePCVH8WC0E3fA0ZkJ/WPWURJvnoyyBoffGcikC6zBIHKvu9hZL1SXcsX0sILqGHuCk7h7MSS+DeI
FHinVkE7rFwXBMh12ofuiqr6jJDpHYulBp1qSKgDYRdqaPnLCOujRnTXpCGxBwR9+EgcyxNV0yRR
pcQwqg4knOfx3vUbwKCQ2HTsybLtKI1DzrNFBvK10z400ol/EqMLXCp7XuCBLQbuOZjIJIPXDCkx
fSWj3NlOafh8eeFVlCO+Y59LDgJzI7uKHBzdela07oP+wOyzueHnIW8LUF3LH07sn66aRTfUmUY4
lXnmitTzw7GJQi8yS1eX+dt7IDT77S6QHEEW/lI5AAKTFWvnYUoqBHM0qZRMQ29KhCVJkxvMTtnG
A1qgDQCNg2mOJ2j5ppyWsCziVgGSDD2XZC4tc/A2ttmONEHKC8Py7HtO1w6ZE7YabM1t1E/12X6N
Qgmemv0wL0R+IduIwk8p5gpGdD0F40vbsHmOFp1FhvH2gzIazuGIjU/X8GAEZ3nXfuib3KBPW7Nv
QbqsitAx+6nCTnBhOVWkX9aaiN2bc1/HnGBAE64m41dRwXUfenrARNxEMMeT6G+1Z23Q5BlKzKYd
vrvwgmBp8ERkDrzeZH8fu2qxlclOQJGLeClb9plqOogsPwCbOTsndtDOzOlPx1lEF6ouMQSyF5ss
UtS2H0yFsDCXdM9aTT6UdqHye7Hel2XqDZlrka4CXm1r1HnmKZZLeaqEJ7Wg3PT1kiz2YyaeKWOP
f84VmfnCM3cjaBF+DIYyvsi3pU2MyH5mjgOLV2uu0B6Fy+5lK7JxCMkn3pdMfYa/prJUTsuhlbB8
6Fg4Kd8XrdBp4DO1LCl+U5Z4ZqwKdKMl8VnvExbgJq1Rf6+5T+X6rFhxNbizpWa7sKGr+REz1ZPs
b448J7hSruYTBOk8FLMMsDVyfOhEMwAV+qfX2AD7rCeU8zLtQ7LKrDImutDB3ty9tUiyZZIhRQJr
yHhMAUNOu2nrzpq0PW7jGdLavFtOP2k2BtsT236TGWrEHOTudMnYRQpXXC8jSX/vNKqybjRMw8Q6
mhJmkS5hbWUH+s6Eu0DHmZl3ck7AeJjwqiII+Z9PF3e5eh+d6y8A/YuD/wxnlqBqPu08HlDxBUu0
29hzQboKyEEg4zBlQbdQd33KQ99yK/8VVqBWIc3lq0tKjSoZ3SHAZOB3O2KKfmsReTnjINB6vgfw
0cW9sr3tQOzvd0uqw1qW5AGCo5jkPnXrvR5MaTa45ggJ5BcE6y+9fqNpgsqOSNmf63DfBCiAEUEp
6wN3RhtYPmU4BUvUJ9+3wHSfnwOu109u3dijwA7cCGsAVQ1qpQx5fzjO1dm5NzqzOLqSc24oAx2l
H/yrYckZh0e06OIiH7Hxm/hEP8Je/D7Ia7JlYkzWs17+JpoPAGQsCPTC44E21iAyGmdrRp4r68PV
QVIO8xomWZj4fHCzNhkUdqs3W7VSpZazFV4GOTt5hPgT4d7lrV6F40etyJkoZ9elNKBe1S+lucOh
zjI1uAnGMz+HxfHtX4ezSGnHLdcG2vAHWTgixlClQUEjZqfA+dfh1JI2h/kq0Z4sM2bkGGcdO7Li
1Vpm72zudGTmFeET8G8SknpRQER3xIt+LxAEEXVGUAf878WhtV/teP0rrRRRLaVshgcHVXeXym3A
8mG7Q5f5iFfDUyjMzFr4r/35TdxthxBrbjQT0cOvHAnwKl7M9lUC/a/UdaaIo17RYzO/uv3C30Ec
PuS6u+2x7ngcAbEzQPoRtHWzVQEoRA8phdH0ClmOoC+yd5zEfAEUsuDh6wpRo2pqS7Qenm4EqZwN
SIrGqtPM4R2C6RMBZ1AulQqCySSlKQ7H7CNmhv93kOmkPr3czuKq3Nrop7KhsWRCP22nlfNZGKGk
+rgXiWu3AP36LpHltzGH/4R8OV0QG6NcOH5c9UPWyjbfzo3LjOPQ9JSlfEdUO1TzvDxqOyniUUXg
oLZqEyYSLJWYZ1WC/VU9dGhxX0eLGJKNPOBscVDgHDJo0sif1TWNOplnFIyPht0MiucDWhk+/Oil
0bQ2Gm9LFKdW0U4Z/p9ZgahKVBNzSK5iBgMRsPDaeQu/6jU5kfTklCRfWnyNoBOAmYodz9QyUw0l
5smmYnxmH4JNoawvZbqqXcxsod79coFIEd8AtPubNHa10ejaNAsobRnD3kNtpi9bcWoNjP4muB2k
oEy0IMHxDVfDn4lt8euAMjM8zojIWzZpymIoT9AZyTMbM//fLtGmcFlMoViTI+g7wj0HQqhyIcN6
GJzDxVRDwkZP/I8SqKyJICAAwLak8uV+bZRaPisQzHZ8NGstVjdjRFOWnX9D3KhS/0CBF31+hqiD
O659KgoBXqWnaS9JclW70aNgTN2uQeLx6p7tcQyJzcc39vPh7xgPRDEF+Yku1/48cvR8EgZHfKHi
LnnqEZSphT+jmdP+0J0naxuQuPgmTZJZjsYyFskOCyPcbjFCJyKC7wJeiiq5f3CzCcOSX5FMgGPi
D4Tb6Il0okkgJawsQW4iRUDphZbNEKAm+D9QlcfU7n3N81gYGp19HKCKmZqNMNlV2VJ+D9OMabGw
6YcYQBYRGv9BPb+l8HhzpKOy6jRAbkBYacztanRG8rmnbtRQxM6p5kC7gsDgpK6cE3l1q+3w5CoR
yhhe/G9YVJ2UgPJM2aJ/5l1kkuAUtJYZBqlGNbbwaeq3Hn5RNK2mu+hq07lG7BqAbUvoVOub+ARB
hYCv3sX11hLFU83/b/BlFe7xQ9QY6oA6K3x5YTVnvFwxUt+sjpE8bZpu4ZvR0Oq+S8g3XuF9SHHd
Wveqv0KBp/8I7zPBMtFBUWthovvzR6oBedSa26zS1WzafqCteW31qnD/Hk/fQhoXXCi78jCAS5u5
RGfwQ6QZKbuzNZHlKvtvuo6b4zIUz3IPMFgEXOpNkdqj64Y6FuHuACtXx5eBAeTpRTa1Ivw1UwQv
22SKDlZ2SkPk7QZhvnm4f4SLvo9Ia3NEv6smvZlEDpnDHUH6tU5yPwQu+s/47xYDsskZQZSLhn4z
L2Wee2E6BKRbrShZ+Fw4v/kuU8C+hMCPigkGiogj3jURyRsfBNKVoFF+hiJ0UQo4c0dhzorWJlXX
Fc6nZO4v0tPY+2/QbfEcs7kmjsotJBgp+ptBI6NTv/Gl22j6NMnFzTO2nyY2gvSizSyPGOzPw0jZ
Xzxyt0r0dLa5kjADe21m3j5GViMK0vv3HxG076YDgVZjXLBHr0qCx4qIr6ucpc1m3B7WQJxccANV
NKWSVFf16ww/5NSgFz0L5BHvarFUw+AvBM4a9J8hY1re45umfVaKtVbsng0ELIJEU/1OC/eymYhR
5kUY2TPQ5yzumsNlyC53+t9ixhQbPv7XuJpTBkV/cxUpEQShltirPQleUkHvscAW8SysLyyzbc2I
w0XmqI6EZdZFzzwCC9zHIKSV4VlKfe7vmiL7mdhPyhn++MZHmDRpzxUM2zK4HPSBDKC+ouLxSFBG
C7ti4tpoOG2OYi8pdf4oVh736QZOGqzAqJGeN772/ZFDxPVgB5cB+l2922yaGjVUu9b+JQLzt9mC
hlny7KaAHWpFTh4XlnSnJzwobaUJhD8yBpe8TljGZo585hnnm8GwFE4ciRW/U9mvvTM6lvW28h5y
gppWFfF4aNJ0Zae4bOCbYr3yjD4+pC8AIEGUYXmGSA03YedEdV3l2aNf8jVb09U9eD1yFLo7vDx9
VgQNBPmpKtRDFb5iM/mT4OfYUeDf8u8aLKmZ38tm2a/xYjXJDhCKbH8noO00ULffj9tZLTTTWApX
ghT5LeKRQmmbxX/4Hxv5cyG3yi021OPRfHWRJ3Dk4ZKRHSh59wc/4KvBTUPhcKJymJlSmdFg3OCl
Dzwb9B6KHvc6mTdb+KfxFzmlclbhXCT+8Uu2RoOODI4bqDfRsuTZCVECfmFcWSJnfLCqbc+LRS+t
DWS0bTCnTYW6eJJvHDyqCeJmytKzCopmAkN08KD1pQvhdNPyVFGh3wHAepFloZtmxAqt9/EXauJh
hYbAIe62vdx9v1dKLfmMOB68jst793FS1sJ60qctmfu+aW7wnrY5IQqmWhgnI21tKIW4wuElF+ve
n82Gb4vcmpUM3DC29zIQnc69M+stR18qZwPO5DPAPtO86J4ChmvV0Jv/Phe3XrTSz7Dt5c7Mi2Bb
JrIniL3hdEha+8gnhRYb7dhWXgbthGI5mwCN2Q4GE269r7XIKmU7P7qtcooXODCCUdtANAwWIbC9
vKLvpArIEUcKhrYyNFNlDzEHKXbVPhpUdOZgP8Yrrl2U3d/n8BCGjTSH46Arc+3oYIVaS8NIR0B2
scXC1NvOjC4AUB0Esh06ZSTXqOcrmcHpsDmvs6dqxU1/KV8cB7eOlKX2izHUqFcIG5CH8mPI1hlN
e3Icr+l4pwaXTJhg0VZ+sXfqJ5/ujnxEmEHX4wmLFtu0nxHte9PmUzyp3+6/50B49Ddati/R2zcm
y2Qqk0Szi9Xc25ieY5Rqgq3TtUMuJeI1gYcKmHb/DXwDfciaEhQ1EeDZXN6kLWY1HdBXpFVCp2WJ
IcfNLB7B2BoNZWEP53FEYMtlWJX1gxuo0ndh2k04QYymihm5bslwBrjatPCbQQyaF5XDyaN+hKs/
AQHC6DApghupYQbFq4P8hfJ25FFlSbWhZQQUoTidGWQc77gssi7pXl5kfjOz51AbpGspjwpZqNt5
w1TxIPQ5pa1r5dte1uisUXGXIMjc6BAvUg2Wg6uKW3iR41YxAkvbR8GsUs4pDyOUtlnjXO9qLCU3
I6EpvkzjbVoe0n8dbos15dC5dwjuou9QbNOnggc4ayUqXhtaKYTwnFaqGGjGwodW556HMleHMCkH
GLRh47rFDTI95+RKdozWhqcnrI2ZQNmYXBUwas/f/+qT3tWvcYfTbWpA2V1cDdW33fYwj9dHht6M
NklyWOgT7+mZbTqthb15XJhcvDa/LulRoJQ6TNyWCazSas9O8L3sjLZPm1UMklmtgZSg+3GXHqhS
pzwo/1mhQhoRQ4tyizoN7qaHARiq1UYEujdoi4nkiYVnP1vMEdurWCi9GmisgI9flEcKr2WlMCS8
kcmP6lJIHDRX0pL1ThtFIKNNr+k4S5Lc46mnkgCIGEdOCxk0x+CADgFOiuSugNOqm2TSkyhkh9oH
LGum0bKQtiNkL4cJCkEDzxPddSr180TrwGDubnrpKQQwsjVEv5gcK52Egz0hQ9lkjt+CQy6WwJON
iL9WKWYogkOsahbODMePioRzrVM/9JRcITfbul3+lNI+T3MnCIjBUdUVLxDvVJm0OZ+CVv5AQYdO
k5bjbbiuHibpvYNZoLnbRc9y/GraClxTNJteyRl1uhIlPT1ao/sssT8nOPTf6/7bjj+q+B+7T4px
bQGqJurSPcsmBLnbGp4kv9preS7EGK2HhnUR6+aqzff7vLuWYBl9Jdz1mXFMpQubcnqFr8mTnL9k
Ad/xACH/XceH89Ul37R0f6G2t+4ORnVdJh/HlXWWqU5AmcMDzwdjTfOjKCi/uyKwwr7Oy4bxN0bH
lqnKwyH+vFnO/4yzj/EgQfhISkbMseQul8OnSMNdJ7Puc/2rtdn9BCb0N0k0AxcNEfmsSZ5uGmNm
ZwvS+hOYW1fqEE1YAZr4+FmFl/KQeJ4gStGVIyBzL4VGoCY+dxY8FwMxRhDR17//5SDkm2/IRYiG
y9lggD5EZ6Nmrus8F5heNFcJ7cI+/g3ZxRVSikkrq3DDIrU0TWZhlpW8+kYnyd/V+bScH4DJUFx8
9gx8UsK+5SaI5a7nQoK0sDBa839MSFsxHr7Dume6uG4pLDCd8SHOOVlm9O+0IoAbdWICXKryY59N
6HMb5SYoDlNlL/QWr6QGfrGfAQ3KWDVmxzjmVARwUs1lDZcaXrHGPXeQJZ/HjdZNifbm+23rsDhm
OfKxeXzA33pkk1/GqqKFt4Ad2K45UqXl6iuagGLzXKGV9Lb1ZSU6Qi4iwfdgZX6nLnCNWRMmF/Pq
ySK4I8bZpUV4nK3KMrGL9FDChzm5xNrMA2jTfg9g69/qHy194oAYr1M1/yHYRH4Mxgdmu61VrXMi
17jupcRhmb7u5i9JXARJm6/nkbeZZrk/4wmNl3OBqCdfvp2jvUUg1m+qApTmfx/dhOcV8E0hogom
xTxXi/Qeb+LVgN/rL9enHk+F5PpFFInyfBiMf5R3zgWDbtu2ecTrNi+VDuq/0k73pyzjEkQDd0qT
GJMYwB5IIAh2StYEHhYca5FheIPPEXKNyfMF1SYAqt8/dqVWdA84ll4p6vGhtl2cj/gcaM62EvJx
ozJbAkgQHkg2Q58fHqfF2Tc2MltSmyLdddYkjGKx83rWYrFGlFvIh8RdOEOIEP4FtcScX1/si9dJ
3lPyF9OfZkXxZG57mcsI/GgEw38j+kFqC+8Bn+ZkwpYE14A3Z0TESUMZt5gwFiS6vKLmaH0Bq/vr
SnIUc8JrAGgmYx2wQh+Pq/DZIunpwrMQeITOnZ3wkL84EfDL4lpq1FsgflwEYJ+5W8B5aukymUpN
cG6FSvJn4bmMTn5ApvwXR/lqaz83h6lJvOj8p5PTyUsH4MjTEOxxtVocOXJF/V9hkKrSYinRrLgW
i6u4G0SF39ZTt6GVtkn2IBte9eqy4p6scJG9Sc9DvlE9bPnaaeFNLQJWgotG3jR7p+Dz0XtONs9R
VMMQhMGGwRvnvtsLQxVU8tMDazPsATBTA9lrY73L/DAWrCYuzOPmO+wVjeMDPN4lExNEpeVit2+o
0h7rqB9NSzU46LgaCWCM1srN5x33z3TzWHl/nAYk36SniOev312u1PSpqTHX6tzSYm/MAl0Z5xe2
lOK6lMTtvUDfE2AqaeYPNQSydgxHicy7yzuwb94ymvRL/X5xWbqiVo+o+LUnqOQcXP3X5nJHmoKA
PdAOhQhYSgslh0v6IF8qbBQLUQinBZ9mpULqIbd8tkzuZHYJ2Aces5TXMapbz94PD2Ih1STLuX4S
CHYJrqYdhk4hFeE37Ns07hl2IymLx3lcSpPtfBh4thF/G68bm2bqG82nGqIJZLuQBPaB4qi5c4W4
C3iSr3925erVyV00tO4TI0jRtsZpiXITMTc6eycg5wKeB6wHu0+pKMWYBtthN3QKsQ8DBdKcuKmg
dUItJH+CoHthCVw35oikFcckynE4q9MgxtPxNO+r/t7ZOubMaHvRdoBgH1ho3m70A1WkdU9S7Fof
m8ZgM7s7gGZW7o4HJs8dE3pahl3wnuowUzjUola3p5+QRi/P1FMqIQIjGnMLWwoHzxnp8/y3SVZK
bv4lq/3pe6oFOFpP1OVJq+nMT2Gpl74Gp4cVgzhxQ+iGhLrsQ+tngmq6rhfLOijpohbiOupiq9YH
KKeIrl9xYgFwocU6Lzrdut8h/9No+M+fv9wsW7Yn4JUWzvUaqwngGGn+JiGTqvKVpqenwtfFpico
fonhJoi715KfhhQMwfuKNu/x77f50eUNUQNdH07qsj7tZuc0owq4Y+XafeeiFxpXDBTpzM7j6+Lw
05d4kFdBZ7RobQi3RGWzUGjWuEyOdp/VNDOB3K7vQEjVHhUO9FRwfYQC24Cfqtnw2LaR0V/KkBvG
HNOGW7dBNtQn/wn6ASx28c44sCa1kA/7A2OHZ0AHaqTeomtAVJFM/D1+yE6y8sRFAwwc5qdmWMf7
erJY9C8Tj7D5KHazRvPJ9eBY+QesD1bTNnie0QdY6DrMQmeiR0y4G+2mAN2YarKA3tUATM+4Jx1y
lj0NQ0F5YNzxc2XxE432NlgzcHPCphv2vGlrwz6sUGcrYxLJ8yVw08sDPVooiRmrWfX9mNp6s5Ic
6FGxkNRgBy/t84OJLkoI37A2O4VxnUioqGlSFvRPoQcF/7EtwKDQCOthyUjMkTWq+Ki+qfc0MRAJ
XApcZL/aHT/RBmM80d/6+m16KOhgDm+WqV/zL/ZMNX7L/DzSR3+ypyNgGE67aVGoyz7h1YfTBuCd
SAVKGPX3gHHokdm9LFQqUNSzx+zFor52TaBaGpJkBTJvmXMV3BpdzXR4lPxgcPJfFf+YD5DzYvIl
pdbmFHlPCQgeGe5VUvNqB0+UZOxslYUGzsk6CCzRbbK9d5DZ6j4Jyt/adFGokf9QQKR8kqHkYZso
384FLNVRwY80Vl6IbYPifubJUCgjVOClmiW7WPPxe5cvvUXChgPi4KPXzRsa/8vH/LOyJ6E7gUBS
BBWzKxR//KBjPF6XN0bd9YkcZwkUhY2jy8Rg2reouLm5lZ2jw3BqfYBA2dAhY3UlN5wq6NwkDCqO
BQ1pS9uRTLI0yfjU8bmIylC1FyYQUxR00AHmmBhyi3x4L1Fnjl7Zt0qgnZ7+d9iT2wcVWUjwvLVe
xXqVW6qzWZ/u5yAXWYuTZPAzmk8Q+NXTDhsRuUMR1nLuOpKQMmFpOclK56vj0YZF47UhV1ZktWh7
a4RHzq27lSUxPDri/Ar5tmiZRSbHgEkod8brswWWbq4dJcO0GG8FBxkQUu8Un0XpxXq/y5FGDXTo
zEnOLsKX1iD8/h86AoP7jwtNPJQcfhrkeSuoTLuZUOeGiUFhK10uFBT71zDQh+/exDPE865/GwH7
a4Y+IcS9w7A3BUMAjwPfoSTIDADk8D0KvQtji+o2PU7RWsx6MvkF3fnJK3OACAkj4ISfpqqJrJNR
LxYGIqI3xPxDlLlZOQ8c20yI8hhrYTXMWYCDsfZzwJ+ynv84YhPtBhA30zahs7XvU4gsE/tFS6ui
xmdkoTXT9CgeuGowYEfxRX5Xz9Tw48n/DAFhpsVjG+m3jus9mdLGCp1Tewy2EnkZfVkCX39kDKUz
zMAo8xhkBmiJWtaa3pdVLn6vYUZTdP65qARXAAkLsFiynUthta322Ao2oyJuhHxPMLZbw54GqQGg
bi+a8PkRw1pbFDUPHESbAB0cyrpeanv+yPyzSAMwqd/UghumQ+8ss0jFC85LgEhtkoEunDyfktRC
BBntOQbeDYDSYKNC3sw4z1mtSqqNbMtRN4RcQMjbICHYrv2lv9IaMlg8ZRUj4UEvAWqFTUX3LYbe
cZFi/XLofwaTVHoiaAe7pOlj3pSqXrPGG7XPGYDfj3sUMvFwKmlROQsKr6daqHtCvzuzmsbfApAU
wGfYjrgWYJL8s2grGLkAHEdp6hcDPK4/ynW6LJKzBngAy2ol/TkMhvOnOBLzMedmHFO/9u/SGNFS
HH/NGTrRyI0T0F/PQ8ZVw3cckgYDOnHwLkfhg+wAKYoicgSlcUSRMLuRHiecdsS/1YJZfEl41VcF
Z65fl3TNTAfNwSLQcrdEqKvcdjBYax02pyZUs/2P3JWvafv/oeKjJQMfWvIOzqZRljKeQA3pPsQi
qEQWrMj3pva05+/3BxsHMFHVz3TYiS7tNeWTZEeugRIKrn2QLNzcp+hl7yQd3E5phyF8Flhl00vI
bc+xp2U7TlPaQ9yBe+h6GPL9KBACscWkrXzB/mJioWQokA+SrJkThl9KY6tuvhDiaMFRTc3LQJPN
9dMMvnIBC90enxSKDmH3DBsHEI3jacgrGFdop9D5RoHuuDMTijtbrsQQi1mJxTijK+4lNd5F3hA2
aTx1myi26zNiV30iDZBiCHJMV+lNFysf25SSZebAave7beuh3+C0MEFH7P0Yi5XsPRWfF0tC8q1O
4mDPlRtlBjCJQQHqBjUrtV6CnBR/85bZzLI5wbVWq2es4bvjTHCF6eoDVtO9gZfT9JXJtzZhVYVt
B3QY1wCU/Q0Elrailhzfh6E8T/23lr+2EkvoGpBaMuvhXvRxJA5M1i7UROdgKMXcFvvq+MzzED96
fyS/SIC+QMwDw+9glrEGVr/4FxIhICtYR+Zqe16ug0kw1vDi/Z87ePIdoPLPXcFXX1UBQ9cdnay/
C0aUpF5QJHGSCt7i4cLBNjQeLY/1Z6x6WvJBDN6lIZgaWNuSdTl/gK9bytTGoUNrgBJ1jKhkpWnM
wWirPyG2qNIenDc+Llj+vgU2O3vtP5oU8jkGgu00MoQpj+UCvkfxK2wa1CbuqiPT9ta/XrG50EGw
hKtgceCYlUJv4LkibzMboIkavbcVtkMNHbiObLW08H/gDLw0GQBZTPkAwKfKA027RIuBW++ktJU4
kvqUeeQ7bTrEDXmNnIKhGXIKqiYSoq//yV9aUJXs9zeV67938Fmkw806cL8MNa9W9CVdiNBjMhdw
KpCm2m/U7j6RXGAF5+CctGXSk3Xb6lwI5vg9hYA9XqkwSnDyBUz85wcaSwOKNYLW638vRHgA6Mtx
tm+jQ1xSxnu/uHEufkZlZJbXX8dRVFFwHjU/HNGVctfvSqx9XXdE6D4YKapXkEvqszpxSrgIcsWL
iu+oB6GEK7YC49wodldyJB5JBAdBvNa/378yqNEfv13apcBinmMM2Xn/m/nKNYp2xRTsiCIq44Ud
WOcWSZqBG6Wzry19wpuLYn1DPMvR+9ZL2OhiViiWQllaZDb7pHOZhftjBokF+DGXReh3T5S63bXH
qcmmKHl0tXr9GZrXgw4eApoWrHscI16xASPAS4X/wCOOMwQeD9qZHJTPHXVP25jzQw+IysnsunsQ
70HMvAkaMWhlXBmDAvQww6eYFarJsy3g6xY6PMBDJg2bzCgcIqhwJCpxiGC/uOCzcW8n1Z/4MXGH
sZhvtHeE4CxzefX1taGnO7C4aXMOYHK5pe8i2tE5tNj/+BTCUImgq90hjvQQ38jiUJBinJKj0WF7
i4sdvj8ckgZCfmJEQNVd0WKTYQ8t/S1DAG1ilyXKbFiX234KnGklKjuSFcZ5Zdn+1Jg6vVlag4n/
cBjgHbSyBNf/rBSJLg75FqKJHiVK7BlAGIsuBYT3Maskz8xyH8ira1X/6xdr/AHRRaPP3quGvAEJ
Gt9+Gp+dXMUBfQewxsLMpu5zDXFnAxfUekRNFsQIl47MCz0OqZiCgThF4ljiBhlKy5zZWFEehZmC
MKe+kJAcxA7P9YC7CUbuv1bC32xuzM4YIJfLZGXjy2V1yb2jFP/egmURDd0bJykeW0AYyvIhPFnz
mw2ASPUYBYnFBcnDkGKLoC2OOCi0U5GNEm2j7rUq4mZ6EX6IcgIr3xbQnBF8uFpB1lrfeUaNghL2
9PODffsig9EGHTK9MSI+Ee7D6KwXw/dVv/OB6lqv0R6QqHhfvzf8fndfkXeymDg4cvN86p56QETI
he9afjN0AvRGwvG7S0gT/sSPWGnEjRofEtDC6YyJmQnFXwfD8wXI83v8+s/DmdNf2KKEkPrTR/mS
YR06x3RK7qoySe8OEdOWxEztAJjO+Swc6kgMi14aOJq+KeHn/zQVy/SaXkgG1rR4/rGwDHMNBsEf
F0X0kBRjB5Ucj0i+nk2gJKfM0uqklPEocfkG8XxT3gL3z3D1lmbQZS27viwh29aVvW5PVWVb9H7u
IbXAR8OiZT3BNswMCo62DS8jxLyQGQo7k4nvy0XPRuEM+OALJgG0nBZjvbfV3Tj4kJAsNCUDgbhA
FL5153IYfqhQDpYAZVE0zdUrvwh96HRBNjjXqybrbir7E1xXTQ93iwk9dhdaXZIvu8FKsSydRczU
RCXuRt+QQUmgR1I3b8OTMMGI2Nc0Dg5/y7jZB67zXjNN7pWv55ouKk8EEHE1sxLfjjMOCc4h9eKg
jMz/oPHMnLFGuJcOsQndVBiNENb4mFksyOI4e2ZdzNvGm7ZzVrevYk2R1FjN3ZMN/fcKwp1Gxwj4
oJbQOZ1xGbkM3MRo3ZamWE3ukG1FyuGPZDLTdd5Qe3xBWWIVV0nPC8rNuLAMRAYsFW8NItMpuxrI
LulQ4l1JaTpx5eOVBw34UN+JAXqT7hs/qop6UX8bHmkFIM3hAhhv1/Py0ZOhwsO9mZWHt1bmZlEH
Nd4qvtQIG4Qb79o6qbbV/JfvLWirfMZxLpTGXVJkGlvlkRIYSDFU+A5q1fsTeF/Wu5oieho2qBdD
vBjTDaH6yTiaGf9LH5e3dHTw9ZwmPmKJcjKG87IyPx4eWKAfMUEsclR7l9iybMy+INF2F1YYytyh
OageGVK/INSCVqBJ2CMqot1NyErMGMUc6zxurT1RrIPoorcmTvYThnrZsX5GgjiyLNDg2/fNc1zm
zEqFLf4mk8UWpg6Hl5O6ht5aeF4bA8omYSBbz0xjW3Vjh2x0H/IrTqko7i8KCh0KI9mvNMG+NfF0
+crWuTJTjEEcZQSZZid88lLF/jCgGKUsKIJqBQVs27XkZqYaUC5lVROIvH2pp2QkkGJWF2uPAZF7
R0l3I6bMkxMUOkjxNvVEIrb+m9UaIMPLkAr35+9454UeLiURexmi5MfloSO9h5Hk/850wOg+TyCd
tHmKw1kHmgqqYsyCq+XpTEF0AajkB0Jqk7oqkDzlrEeFU2UT8RI5XSLWB6RGjlmrkxt1zdDeW0Ud
GSkRNsMyE12uzuK3qhJ3UpMTcXNqPHJ7ogUtsZjCDGaaoz6AeMwaT2nWRa2OXLerbH1SjdC5f8Yj
gcfoe+bIdEyhA0m6QbwdJ/ZEI4VThq8yw8/39kLVGle4JJWhiy+a9SVlMoCZ0eKCS3F/7YPthei8
7cLHMgCkEZsfH6RvPsg+mdt98flxSzuDqzTyJ2ViZw0p5xKcgFxU0kjMM3W6Hj05xRCCq0p+Szkl
B7ILk136loce1TuzIpDEp297KCTs+ZXM44dbmDffAe9OVdrFOrwIpg3TlaZc2jEFD9fvXTKKoz1P
IeOsveAT+7sXcMKzn2kN7wQXkq9o4QUeI1Cr5qvKoUqgQ7Yte6bwLPMTGGuetieRot97Q9+YpsA0
0nVvKJbvWMWsrVrhRbT55hco0cujWKR2IN9SbotyrWIY+3/qm1bOLhkh0EhmA6+Cx8Zjm9iIwngC
pToMwPj/zNPXrB6zvMH3GKNT6YxgaOVEFopwK/+1gyNtNIOME5ksCcntCd2UpgGz2TrEZNdl9Ins
M318JUxSxs8eCk3bNP8CW5Xjys4TLlhG0yQRRGziKY+EqkkivCnvQyl/Zt1g8cNIStqwTKU5VHbt
mQ/GEQuNt687Tx4+SD1TISjMtzoV8OHMgev/vmyK5M7qUwGEil2Wdw28l2p1iuKjynXNfUxhSGxs
mgm2eRtJiMwbz28EzQ3prDjymEiyjRDhLB9tM/Uz9zhV3ykPxCy/84drKwR6fQZfbCE4zB4b5kZB
jpXirJAIiqpsixSYwNyHSFi5wMTc+OiBVceT8EXbzDT6+AWsT4QoEu6iYZi7I8ysi6goFZowqpX5
gpf225+wnFkHQcvCT6bLvKn0mDDDW844xXVwNgp5syzfzmaup1j+4hUpdXtduerWwvpqRVaA0Ijj
mmcwVX1bAq+SeVTYbpqEjZx1zV/0seYGZ2zHrHXe38wIPpdyngrgzgmHrqM3zXWbBaDp90HyQZ9q
C99N8phmAe8oCqkpwx+PFq89kz135JK8PogsInSBoacPQY+VocW09L6xjPB/PTftB1L+GmM5fJjb
kYQADWJpemaYkNdninj2oClNZsT1SFBXAuYNhM/03xacj4+9PQfh5Qef1JH00d0+qj8FJ5pzz+IH
wq0uLPVXExn5Ki6YxHfMmg/XALuVQvG9QNLFRitTBGMTJvfk9UeBmkzn12sXAh1YghE2akfpUvXS
NDjhoasAQNuP/cxLTknhxbA8ja/YjnMgxZxDBBUFysscSuP+JFVL9z1hrErB+JHp+4TBiIoJMpWn
5FMP3vjZdjGjeJRG1yVphsRnqQCQFiL/wxocnB5D8zHsE9bxxaxrkIVIJlw1Vnp/W5I/hA+N0TDX
csvQrqXDK5jw79nPLXE5rgfW2gk8Iy9qEhvrQBXdRrNU5h5xlVHTbAYJ3BmX25ciYLpupG0rmb8v
v/9eq28VdJB7+vJ+ypaozxAojrpjrDVDSeMDq2MekFBoIzlpbjqK9D4L7AdPIce5YKycX3RFEdVf
vhwgx1O/xaP60XaArAnkVJoFii/0+eur9wpm2THVGIXZFFV1EcbHZLnxRCmBIG65Fh2r7oXcw8Lb
XV9vV8+VQViffa0AZwXnwfM8bjRH2Br69gabVozo9g497n0Dkp02xaT2SjBQnVWSJNqS/cYMUscG
E4p2jNNc5n7vwVDrhw3f0iS1hJUq1ztSY45IPBlS3/a70u/RaCm2SyL5YntQLSEeZUxMM/BhaZOI
imfk0C+wmLtbwAwwGGuzalAXckpL3yMfguvuho7Z23Svx708d/PWsawmis5jnlnxuF6Gjd6GbBi8
cSCDPY7+Esc9SxT3qXkkXW40cLqBYKSlmDQoN5IhluSH43ew8HNl0W5dLM7HjOzbuulnPC1G5mHv
pWuJc+CW7kdymC8QjwQPf5mNcO15xELVFZq2zgda1y0qfIZgJgmJDi0sYGPC66u9C+xi2T+YUHfi
xzoiN749pp/e7lwR+iBAuntSKHKpxUDSof0VfN+NCp05qo2Q0iK+MdMUmqrhjtLmdtr1z0F+gv8X
2O6RuLK247akfvkUkEaCbAGgkhs8pPfRiyZpAXM5jq+dgPBE98DKm6uIPmd1J5uS+QoEDzPaOJ1V
2ICNu7gpB8arbWQySkya/lZkb3nOhbr+ayYRj0N69BKvf+NrGEION8OcyFzOVjibfBH3Cpod52NA
h+VxFgX7EYSXPwnuUP1Hez6pWMBpapcRYbxplKX3hBCqhjzrP0KcIj2jF6Oa6TxN8EOP9UpxuUjz
PU5MlFs1xdKeU3JXhNw4sTQilwXBk4p4ePA6WYCDbL8n5J+oZeYr2nNdsmMetN+uRyRIetIQF/+g
4O5nCjUK+edVDXE8GLNhEqvNQN5LbG1o8px0n0YHSKbH1ht6mrxjnM856Jt1dHRrMFwCY06suuXt
ClvUbtDE+TDx//2+juHelORLzLPPXjoHrkEQF35Ta+h9RwL9xIISzdhKTEs3el0TSk6bfJacmpFx
/xrAAS81Z9jt5u9mTrBiz30NrF7Rf+iXSu/JphWdmYk/9pVuCfxAX/g0Ou+5ItlOWKoMMVVNOAS1
qI36Qtz5GZvAIXNqfUTSYgCK7bKZ4YBwggSEJCrQ541haD5QHFK0yAfA1XQ5cg2d+LTOyeUJIkSB
27ZSbiue8Pqkb+ILmDVstmiLcmO+cV4hsh3YWV7l9ryAGYPeb082qxhyGla9FDJ4i6AoLJ1PPrNZ
khkCk0lEeeV6Pjzxaz/HijtXfoUytJ4I2DvB0wCccE2dEGZBqgxVXO/eOkByxG7nIlX+v1xGR/5W
Mdv+ionsr2niJYUOhttbxs+nwB90TQQTaJq/xTJnUA+9biDJSdotx6YE8yJccnrSVIDkcQDaQFvm
j6E93d8w6sgVMLMN/SQGUU2hIyRCKTqXIPHDhiCzYqJVpfNO99beqGNPnX5alhy0jo2EHQoWXXx9
kv6tPx7Zl67zKhnOGzFxzPpi5caTNyySnHq8BijxyNOzXhw0mlsy6ixFb4V+AMxTpE9tMTfukCao
OV5Q9CYOjEVHCknWINHm4I96rk5UpIjWddgyhB6bfMXbTIy0AP3x7uw4/6YGFIYol46e4HwnTOba
z8v+Gk4PtthyknoeRP4LPwdgGoTfiKzu/NVkAap8XXYeH5QQp9oC0HP4bvw2Nj/AVrkKdffI1un/
m0mO6gHrZFSq6WnevHOR983spSHME0k4hd+zUK/DrIWJB4c62LYIB9EcqkYKBcLEmA2wYZ9ahHFe
eD3AlvVVq7l6XVTx7Be3OKFEh3oZ+qwkrJMBeTi5HOO7w1UgszbbuTX+3Eu173c8T8Ggl5YQQnM3
fbce5JPfWqy3HY+TeO+Z0YDhpIQrF18VrZxAUfi1KSaqEPfrYMeQb+mISiucvQkZmp3btDOnRmx3
FKDdxqLab1kGoKHJt1JdZGjLg/skXv/fwBt0jTs7y5oD4cTMiMq3oU9Gzwc01cFtR9AM/k3iupr8
/kHetDgrYrgDnKlhxCSESY2C+KaJW+ztgpnHle2SIOyuXYy4UxNsvzge0YLJBleWwzT9pVvAWzNx
iIfahP1PmtIiZEz+3BuBR7lyWd+00lTsTA9whuihoEy1o/dvRCv3WONjlXpEe0kblsz89rvTDcGQ
RF5vsyCeHbN32KFIFOIx1Yj2TfdLyMkV5qmzbSN1hc4IulxxpF/JnXTzuoJSe90cR3irEWHCULsT
63aU1Ao4Qq7IJ6zDeKFH3SK8eFX/KXCCUjGKdUpXTUEr8NVhE+H0BGYuWg261KJF0oF9wXd0uVnb
BQ9qnVOdfR+glB43Dh1IAied7tCNQiQ58BQfHSPfPvSQQWLA82u2DRk+Q9Z2rhx5IPRzamXsYfUo
hufLThHb+6+DN+syANWNyDxJg0RJrIxvpmjuQKT/vipe6aOtPvSnb2VwYSriAVgjLpaRa4Dl9+1B
UKR5oms4SLYmdzCvrLSaZ9FIbKy8dqpv33RSLQjjJ5ecpcu/tohsPosI3XvuVYLrtjK/rLhMBbN4
7LgLX193mCcgt6Q9GNLxI7nLdMPphr5YDcuEwFH5ghhKM97l6UjmLyID2e69Jm2hPoPe6C05I/VJ
pvwhx68Rcp1VeabGf5G6O5R1HxocNEICKaH1/zw80qpKv0FtJtLrePG9gY0d3nPKZlIcZ5hp3gWn
HQuLMvT2qzWBWgq25J1w5QwA/chwlwKDz9gVBcPRXXh2cqtzE2ZODqeGsryQv3y6ga8+KCnFfVRY
H9w0EdiRCi7y5T48nh6EU+Lia2pb5OdRFSHTCu8a6Fqk4ko200oUnpjPRPqz+zvZCh3Ksyyz0RyN
YT6qOiS55vI5ROXnqK67O2wKz5tL5PkfYmvHUHx1opUzJ+dNywiPFqKCu25s4NLe7NjpZrPqyfWC
8TjxWwgcYq65Q0xFjfZlph2rh9ANH3EsEaXSWaoEd6jpginIY8bqFtPve4BO1h42LmPm7qT+Nn0h
DfwNxS3jxb9t7J7mIjyqTXZBTXRSQNg5iNLJeGmwPBDmH3QjghnufF34j/UeDwvsN9mCfxN7M/zN
0He6VFF21jGR3LsAIetN/LRQIEF6NQGfQ02Im3n/IFI6uUpG8XumksJ+evORSbtizsw+DrQTPT2q
2Ydelt6DFYw+ZB+jX51U2O9KVZLTH6ySCreuCVsopIbRL3fKT2a1eoEuyHae0IdCjofxEdt8nE/a
+hl3+npi3TLEYViAuToi+VfpBK9FZXXRkvd8/9tFrB8eHvzX1JdUoOkMgWd3wwrozdM/3GFRmjGQ
fozH+NtcEcggSMMA/ycGZtKeIo4zW1vJewg7aI4isZ5Xp6MfuvLUG+l6jQTzhd7EzQCe3Zh7doEK
eIO7+xiUPcFsPYFWgqcPVpvMrecO8gUjKnObOLGAw6kH2RM0JIeAGJnCrjh1ohWq6NQs94/FxkhQ
Opnke2MoGf1c2V1pB8b+Pp+WIG6B22DtCnGNHKU7Nx5NMNrVDoTJP7aroKgSf52tauZlEoQpca0J
M7PPND1wzYw2sFDR+pazyBLKWGNZAnJA4P2bNOPxXOQbgwPfmxzXBfnzLBtK9f+upwyuTIWX58jI
xbrA6vkXjEDn8UuyWmKUybLfEmB39fkEJBTJ7nbmfBA/vkDlOhZENuH8kLqbW5aTxo8OLn0X86zD
H/e6hJ1G/V1HGyx1X68Yb+Z1B3sWjcWmWkBYGqDqGQOjevt1m4ek2/zPnZIfBRiAYfjWaQZF/UqP
K4wOZ/9DAOYqBwwNsH95IldzIjTNylXuRD+kyrHaM8uH2IxI9eAnqYs8xf+nckPmwjPo2yWekkE/
34aDffE4lripxNXm1h1ipz/QuDs1rmEGk3u/XsL78YibAPJM62mM/URvzRYmJBRCXg+Lpw2rZATz
wV30MaWo7M0uCYQ9td5R/Yfb+uiN6tYh+jTN4eq6erTlWX/+nptp141+oPRr4u9xnACfe4g7vNF7
cyyFNEwPhEEg7UjqfprKiz16lYogbGNZWJxGh54bCw6luU59k0mLdIb+jRPKKANQwnrhVnUyQYaZ
VAY5yZa7qFcfQXzhtXN6NGZPuUwvOj+zKDaGGW1EhImAfUAZqhXVB9y+3m47fQe4MsGxbKstT3e6
4N4AbuGdENIfMwevonf2tHnu9dvgBQhCG9ni3GwbxPfnrt7AQ6+FJB5SCpN90ePnRMftEU7fGvUk
DPyvtVWG/SIhWo2h+6iL07aFaA/CeVb4VO4Hamdoq/48P1VyKTE9by1ZyvdrulV3RrBCf5va6Tf5
NOXfdPuT9WwlY5IuZhTSzAPuAgwBGo2RVqa5JK4jWUcPEJ2M47CY2/JEvJ3n4yhtXaHGpJ1WcUCY
0fkEz5mKDj67HHXBwjRvGSKiM3VbmpiHZEKVK6l89SsFiJ4A4c4wCy7eT/WGQEixclJb+8xrlrV3
qiFg26uidtt3j6VTglj+b/JTdENrufhEBeYzDpJTlX8evFptoibNCZwWYYsWD4GPMRzb9BP893OY
gJrDEXmrRQb11SdpqN2gd82+oK//0WIlVqU1UC6h9QLRMlzx52jIjCEmJbsSTrrH23J5EK/+qtG8
pTgBHITxcTSJPQ57/dxfnMrxwUj11RoDmhsvjySiXcL/BTcT1Gs617+G5mChYklFx23a+mkFt/ck
MezDS26+vljzk2ZRVbyGEHwImblICOfGsdS3xGrqvJM5+KU4G+LIdPjFUs8+2wlz9xFWB2xUKXQG
ZSVjCUtCXDkYG74Bv4gbh2kXVfo8MQzu3eCiho9jIV1NQNYt8KQZ8Kk+nMLOH6PSc5iBnOHrQ7Pg
RN6JhRM38hF4LIWqLBe6HSldgaaiX2V5TIYcJeQZTKiTDjfV8RZsQdAsmS8gp9pGfiW7ULEWSU5C
Yhezk/nAIV3Fo5FipB/GgrROFHqRuE2xEkB5Tbtr04VYJeFmbH8VoN4lBdAf9jmBThUDWtXUeZME
X5mEKato6EM0ERcDnP+Kdzpy3rwrhfy23ndWJPNBpnDRVGGBDukc+PaJgO7n5BqHEQmiI1HW+BrL
/MzImLHDsp33YL1KdzFooJTZEERGcghdCv10IHhtwQopOJKaJ8IrCjcWvmgOeRzvGfH2zvCAr/sb
eaxPT4d/HwxexW8EuBj/DSPl/Sus/iRBEkwIAegQIM0NNfIb1DnZhKiDA2uaFcs1b97zDSjjhb8Q
1fQJvMkaErBnDdxRQ+XsZGJq4RVMUYDwwMzvXLnRK/J2WWBW4WhHuJ6VQN2ANDW3Aoo8OdQEVi45
LxrEhxytkwzSnPXHoQudSpWAbBAL2jRw8gP1hinqqNJ3gfyGDgOMm5GlrFefxnlLpymgIMyUhbrV
Vm1z1Z+bp9nGXGFP8UeeQWsI0XZHNgd/3LG8akBKL0xBaw3covwX6nKIv10OlG50m/ODaGo=
`protect end_protected
