-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
X/mpAuTIbpFRksCZcO7ZkPMq+yOwKaZtwo8LI7SKolTg4iPXAm3h+/XFSC/rxmOX
zDHsUArqQaCuiQnsiZ0sDOPA2YEkk1NxqAa/YEiR0DJY2ZZSNYy2P5MOXd0CGoT8
O2fowXBWYMD4ze3o2d4BC7ffH9OkGtlxcS7j4mzzKzo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 11534)

`protect DATA_BLOCK
GmtV++TLkjWSCIveeVeg9IqPAzyOlghX4VBY0SY5g5kExrgIyyiehXXTaZiLmWMB
RE9q7hFhO1V41Iocd3FqqDQ2bFw/iMtmkTooVCpazSxz6JdZk+C5LN5/1kJXKEfP
fcJj+UKiONJQ8vv3AnZ5WvupXTDBIQNONv+Kcw6WjVO9+oLphcZGLnm/WHrW71vN
saEA9QP2OaCb1JMIZalBFUoJRisBdUJ8LqTpDTT6eHpGJY5wR350nPtwsaLmd7Wv
ZvFCxavGlAxkHYWC2JV6X29zDQVmveG4k1hxQzxWHuhFPYHrRRLGesqg5PaHX7eJ
RJjokP3SC6gqnK8heq5K9nv3PuCN2Lq/nEmIg/sxbVhedth4mM2OVtSV6OvwGpj7
YMWMvypBGT+UH/d2G78cuNlPeAC0FsTou1YznY5lMJj3ejfib86I4yj09j9UoY2x
r9T+KT73q1YASOUOs5FAwyhEwHQNKYP5mChU5xJ+RpLbJ5zPH7fj57t1v1AQBQpr
ldqd46+mggdBAe2ry3YrGswYkgoaBl48KD5BvozzWRd5Y31OVVLN30sW0YzKb7Zz
lj67T2S/I9n6XrF9dQHO1uYYrtS/RGzWlHcGp9qcXeqkF+puSNDmqKl/CeyYteZd
12jt5drxCsk1n5E0Tvs5PpOn4QiIADG7zSZja2vpYruUaYZCx0M1czaRo3jCAt61
vTXu+BeN4MZByZMhhtm2AYdE9f1idNsHSXKOHmKV+Gl5TbOerkzQN2ljmCqWKuPi
dTDEklCmQDBMpQGcP8q/jgSt/prpqJll7K270HOuosqWsMnZfhjbY5UQ2gO8zkCi
l3xDKfIxPFk9EbSKy5Mu4UttWYjPqO66nya9H6NW/Co/OyKg8vfmAAnXK+5c1z9K
xvVJ8iAWFPIC31M9rGqJwCnnb+/41HsdOJU87z12vGj6ApOv06v1lr7MjYlejp8K
pw7K3vUU5Y33NC4QN+IPZ9ZKZBLlBlLjfjPIX4sT0yWkUq09tmApkwf13sxmhXqL
sDRCKc4pfh92lzuRvD2FLXMuHhjdviI102LK2LncDmxSI1nJ3hJZM0l3NvtMk2xW
e4MP662m0Go0BXsM6nEjM28pka5RRrao+npmNjoT41/Q/GpB9zlxoFRJYBMXOJJI
M+iTZ3soUxAUzJFWRmG61v3/+B6w0Yck/tc5TkXe5jFFynzdJA8ceeGexE9FNOaJ
ggC57mFZ7A2ETePzTcPunvORvRFB6YEDCGqvykPEizJ2NTJb7diEa9SljdMqabdp
ug7odIkaQUP13AIWDcH6o0IEdfkBb6ys8IVUB83ZOOdgsLyIDLuYSj/QeB0Nk6kH
Px0MV4tjI7Y/tzDcqllSgRM58oeZfb+iY+4GOhdGt6q6y/bEHj8xXVVpdVmNhQf7
Wy3eY1hCSu6h7RSsJAKhXuETfnAjC9pkZ6XnCedzQ/cCu1QhjthiDITxgj3rPk0H
kRQ4LJSZ+GoRpWVOeFSmSa7pQSGjZ5OdUih91IDl8hNshoqqcx6LeiORCHWA3bk9
BPkYGDB6Jb5V16wxXbsJfkD49Jp9NtmOqa0iAyhZh8kGy07f7CYuCbG/WlXThRRz
hpy/TdQmQjGbb0nYcOIaX8VpBDsrjj8LN5rCRIQAOpf5yJvTFgkMU3TnyHbXvNDs
tgWcP8fPqjAS0ogXKNZ9NA+R3Wutrf2D1OX6553tziF+w8isWu3kM/4fxCVxf1B7
CQ5bbSZXSwb8jdrSnPr2vAagOWPiVxPRpF/byMTkbz22VdYftK2xbIafqhoDVrum
iehAtQQCRvUBSteDP/Pi63YNEwb6JM9zHd7dE1wwWzU3xzoOKUxsKba80cmhfJjM
Xcm/EFmZyDbYhcoXlKUzp4wL1rRQckH40VZQzUJGjuoIdNzyGmbQ2BmjGIGPmVCc
dldTBKDPgFl0o91tGiEFn12n0KEZS6o3jngfVh6YjbjhhupH00Yqtwb4SOD/FmI8
+LajTtW3p3cCSYPvK8mKXlASlzhvO/liOn680csDNeR60jo6w+80kLnQjJHvgUHd
KBFAcGNo0RIxNQfIHl9Vvo4V8Ym2i8452Mix72KV4lIdRoQxhm59LXdO9RPzWqn3
kfy3EE5RxEATfVDrx525LXW8bk0shKgNq3h7noF7+s76R2fRPcSp++x+TsyHEtFC
YWmgSbv1+wkfAqSWKbz0EHa031tzB1zlUXziPsOKrVDX714dk/gbzqzjb4lYNdIe
ZGbJIYXQH5dnNxKxQwDC9QjPjc35rroXN7Uq2usvVH1v1em/n8xEvOz7gg7qzMHd
mC2nongRyUl6zZ4asJxfS2E3DHIJvyHdo9qS6fKX6kXqlaLSRiuTUPSzBQf3TkCV
fcca3pbs+GUxctOXunk/Ql+KC3qoQAbLW1ZcRl9jrs/eaO1UZrLO9xD6O4S6oxDK
To7ppHf0F6g0cW2q9e3OH4oTjOfrUgkIiNRC+zAG4adIA8/j6vqhSd75ui/XHPkY
b2d7EajV/ClwpJ4GiVTRaNbVUFuHfmuBLjIz27OBZNOl7AmqKPn4MbAE+MNBh/gd
QsrMBL3EQD+NRk+BjVZz0KXw4JwtyYry/hg1WEsKMralp1rDM7NBPRYEoT0cqmAi
WEK/X9esBvJIdyHjzjeFMuBY9e0HItDCW4BtEb9CtIAUI/uojYZBjRqfBMk8fS0n
odzEEcKBXUXlw4pS3CWyrTOJBnBXUdcazNReJEDHTJRxinOfP+lIKnH/HNy2mBbi
kXDmdETtDlVqWSYcRZCaexxtf9mrmLIpG8CURAVtCCEvfK+iZlq++DS6ZYrrt2lF
KymZoDtak2/kqufE8DfPUWER6xWVcFr+90XGd1fByJOTu6xUUsIMZg51/PEJgTC8
eM2vn9swW81lvKKcX68ZS71g/WAt9S0OEQV79fjB0Nrf3KU/RQD9Ykdl2A/P2YBJ
SjDXicmbgATPA7sJ+OdQZrMWd5tEyfHbRjexCqXDuzoK5Kks59pC90b/oI+5fYgA
MsGqXSb/QxI80dAk2m6qIZoNwWjRbxI/IlOk8tnJBUnfhuatwNlwR4VLU/5Ev4mO
CPEUazT8lhNJJIAoZ3uxjfX16XS1vCSFc1OzVGc0Bo+V//iZKAAY6tYmm/RzuWeX
Mc8FQlHaBlxa5XOzkceU6eFRFi8LJrEeW4wGRTELCtLty0Y+96M3kJ+29SGwL+u+
JSekIE3aOqrzAOl/7mYoP4hQFgYEcap54vMU/7BF+0a88VrK8/nCtJXKxQOXW7EO
tx13GSMSDqvERF2D6ArjsWiB9lvD0be2SHzdRhlgjJbhQ7qTvuOLnJcjWgY7QAwB
cbij+YnpcB58WH8ncZq49pk/U+IXJD1TURDJZLlZfC9l+0kzUvMR7a/HlxdnLA/q
uSRAaJo9xO/R/gx6xox2hAzN5tHb92kpFtT291dZ3LVHzk3CRWDvJT7Zxp1eCq3w
iZ4Bs7Qx2v7XmnxyP3LddvLe9bBw0RTt040JS3yodVm0iMat2+EnFosHfwKlU82K
K4IdlwJzwqHVn2IZwFXg+5O3TfsuicYu9lq/UdqNLLctXNlyhZc8PQ2j06MjwtYt
fGndDAbT9EMbLdxY14+vbtcgZrBAmWn8cmr7lQBdH0LyrSjbaxyLMt9/16ght269
8/aB1d623q62tIrEzqYsan01fi3qSDlPhW4scRsllSE8e73+D6Gk3mcM8vFeLCuB
/ub3K0virHIDmLCNq+1EDlsDhT8iPFy9FWg0vvoCmVQ20ua6b8Z/V1261QEYO4/H
JvWBRTGc2cIJT5esfWvvZqmy/aPYnRtZ5FScit4GhKUtXcp/kS4iKtKXnJzPk3pY
tc/ePRrZwjzqW4B/wmh7geOumTlVMi2YUlPmcdY9ImIvpyaKGRz0kp5pLqzgdA9b
NCmIKWnJCI//oipvISy1pTRn0KaLTpUpcj27CAAeJuxZQ8aiZ+jjU+7X+PwoOS2N
XhCerIBQp+2caHkS1YigLBIUWo2IH5CNTlJ9CDHQQR7lXo5MZrn9Yb2S0w4bsi6a
Zb9cuKWQsDqoWd/RJQepR2oogWiBPyvlP9WvOaahfwwT5f1RAmSOcwjLXW5KhDKg
KKiWqLNMkTnzqRD1fmeruE4lzihm4Wf7urdPpwCXF2m4Ejo9qnmX1uwBQqNaMaRp
mCTCpRbv7QOS7ZaTb7cQv+52rKaYYl74o26i643C+D6V9TZTrHGlLle58Ac18qM8
B6C29F/6852t41UuNf2NhWHBC7UdlhFMKLkBiYrSERUaOimenIfNGquGaDbwsGyC
oe5BzHmI5iahqoYXwYNUHscAdXxVndyNq2tlBhNnemrIROhDh/GvEQNUmaZNMWM0
LBHJwXz51IgCkfproHoazbBj8LmwLgv2oVJ6nIAN5lOe3NBNvKDai/oyWjwjzYPI
p1DSk41hLES8ScrIRJyfxpK6HorxdcD7cXizLr6t3B+uYmfCY+qIGljMDH7lZwrL
suWqTczflq9rYVweGLtUQrGS3hTWU5WmXQ6s9h00RgkP3AIDiOIr5kJ83mOZJF/N
cOy/KLRzJHOjjKg6wtzlCLOwuGppKUC8Un0YJ0Rcjba2OMb4YBm1alBkaSllb1I0
V6ePZbICwlAUITHiZU6QwTvSrLTv4JCOgB87eSlTrK3jT0TZq8c9k7d6vmRqGfII
B1vneevmtp4IZ/DXWaTHpUSC85CjnyXCkZYElrBrzWIXkVngKMoojacuWirq5Aex
VxY3ottzaw2Y9A+t6HfXyLazaeUinxYy2uIGbsZhyu1nUILAopxveKERM9mGeR88
GA58ralDkv4+kdQw4GSx+WQ9bxf6hXTtNFtVAkHz9dsW83lZW3QfMcggtf68WmlD
99UkWzDN57lAlSuI3T39g6MgYIbc4tUYALSszYNtjyjxtk+oF8ubNzdV4LKN2aBW
7jdXe6kNs6du9ar3ySZN/z18UAXKTcLvsfuozvf7g1VOO4YjENo5YX5pZtU+Wd+K
TcPCeo08tEh4C/71jw9u945ARNsryKrjNf0BbQ5pdRWTJq0svtty2yqADxdelzwg
CbrLivIz/5/eUpElfod0qDmnm5lmiMztT2ax+mSp7j3RlOZsaBLcxI7lprLEgPN9
EhJtCDzwnKwGgZ0MA1Igm/jDnCGT5qNyaZ2ND9W+TnH0nBx1LO5d8v2Vsa9nvDTw
fl8vjDaOzRWj+Wbw6hQzUTYk8rmz0FBTWs2JzW5273xtq8rtqBuw/phiddCY82lK
rsm7sMhtAvS3tp8feyUFEjKnq8I8JhpPrccz1j1jUrTzm6V5qTQqndF0dePXNA0b
og4lglLhGFA9KgLPAb3JhK2oWnQn6H0DsdZn59whqs5Qm420XGd5Bxc6/qVsxobr
WZk3e3/nRIpFEG1ZoJTJqSpynjuuRNV82kamLZ0RLKBedWM2oNEnZ5PrHOkhv6DR
jPQb9tBaxmGrXn7XRb4+3OGU8pN80uLckjEODpUCL0/USZDwry1mq28YOiRaOMNg
638++TK4G8TZ5SH5fhkpw9+HugeucVL7wmGOWp1MaU3SuhtgloETn5m8yQMNGOJb
iofpctTmTb2N8vRYx3aaT+Yym/tJ9pxWqhWl1eG5dvsHlww/5pFr2FkViGUEeJca
UnnjrU2om3pw8RuwkxC28fuhF7kbjR7eqbpyg5WtlBShn+7xCiJzfIckmE7HTy6N
4ohYcB6U/xxAoaCzjJd959/idIY8X82mpw54OD37OvKNF4hYXp/wd7CHCoA+QFCC
QxUk/vdBJd/ck8CSxDIhm2AppcJphvQ0YtWjxbj7q5C9Qw8VD9Qh8E+LMjFLWZM6
P1spu/guAqJeH2ixzRWWj/ebvewiN4OQUsSmIA1XWVA/ULJQx2Fe8VXeCnsY7CP4
5gAoUajqS7W3rQDS4BCb2eyQbb3IB9SQCo+pdbgAJbLKhfhO8ju8opmNM3Azz2iB
PHCZE+U+tTEGRxCoFY61ubibtT7tNTi9jCGGlgoANSrDxJWysTQGQ9zD6Vh6epOI
u8ZipyFjFhh6DBAgh1Xm9vsjzPgMVHc38Mu8pAge9pbxjCwmmxUMlKfUWu++cwCe
MYZdCqAehWQ4tkIMoggYa4XAS31XZZQMmY6LafcT8hit+qVIjhWTeQ84Th7n/i2Z
Z+RS1htoOi7t3vm/4AEXuWf73CH2d49aXCUF8kh/pnireO2ku6SMckXsXCA4/Js1
Ucp2dNA3tC1CT4Qf7FTWEM+BHX6+7T3JJfUvOQ7fCwmw3/y4zq+kF+vqRrg+TDiP
Nmi2PiZY7Wx0gsXB1n3GCYTRyAAvbPCJu3DMovoFKYCNoBmBimbL1WGAxwQOvtMZ
+593ES3VSZCuW4z+3TtA3ejpynuhdUXDyiV5bGf/bJr4NgIyA36uN0QJeIkof/YK
S+6NfindlXIy2qBmaGD2EGqmUl2mnWjIubfoWBS0RYDQuh1bKxFTvUVU0Q2Kvt/f
eUR+17s+NowQwZTD4SucjYcfgYNZdeKFrMXienN9Y0b3wbQy4RIdeYrTpEz6kxYM
AJukqM0h5b5o97fard+whceRAOFV/TEUgB8dVV1pw6kI4RZ99QvXV91EUgLrtYt8
ZOO9TaueQ91O1ChInNMVwPPuNq7XPXy07oNKh80+T4f9ESMvmJXrPn1S5p4E7I3b
EwBD4+Nyki3auqiW421fntxHccHz7m1NzPn6zIALdLSmhyCpPSEIq/aGBtIaXiqr
lciJDvnNzmxqLgY1c1oXAbIIyw+1upesopKyFJ7zJ20leLRrwbdubNW5Kaq+Gx7A
INHcSkcSmsiK+sAkb9XPn/yuNwsIlWJzICHvywix1L55A5CXS72lC5h2R7Jc7wOj
fHjLx70xl+3Hji/CrcrP9MJuPJFpD5HWkFUiAJ4/SpWGYR7KpUQjZu5mMRx+hT5q
DVf//PJYoNnOR8OmDein6bP4leVGtmZyhgAPGsWTcIiZDdSH6DEMLwGmzAAjceEj
vIawpWzuyvfF2aLFjRyS9u32W9BX9Djx+VBI1rvzxIXfu+US0drJVfLpMvRLrwD7
rYMB6wbo24tdBAELyzvLNOUkUzQ9qKnTK7kAlYiaEm1yMaTMFgOKTctFfcJyci4A
2JwAdODOe8vnv4sQe5hc91hd+5EVYKJajMzeQcwGU2OFzp1Li7plCXiE1UtTogMG
e877x8hwIRbPk1kqPgieBZa4nCV2MnB8VnGFixUAbQpbDjWflc9jiTqvYu9slgxK
egWsOhIc9VWYxFp1urmAjA4nDMJFvnSOEkjDWcVrq0f9K4+F0JH2/k4Vjz0cj169
kkBLKkBELyb6CKXTLxBhj2qixBFm3Xj3NuM4EZTHl0B5QvFttkUdGXdikXyCcZTA
riDkTfsBSq1TBPiuEMeiFz3/jmAw/7sBMT/5//Aqg8ko3AZXGOXa0EcREsJG9fXy
6wLROACdpOdgOQAdwWmrrVGGh/ChUHWZQAxr7PekaIGdYgi8iI6uA9zvqYF1OVNS
vH+ot2cX5Yp7ECybJ/11nU6NmDOdlEtOLW5/0kOOy8mOTu9V8OR+kNr1RIp2E0Ao
gKYAQq2oYG5FB9/suPX1JrMbeUi9nxvjvMCfFdjYoqOKk88OgKYQzX4GQ6QCQxuB
M/lQnLLsQsWEzXrobEfqv5s6qm0TmOBxZV1MgNsVJ/D+LsLp5QmgjSSfZ6gzTLh2
Ms3oLWyTQCCropuUWI32yTrhui1uxEdtgpjio/6gINlZc0m6kfxl15kWGUbQy9Jh
s1gC07vsuyA6GsdTLRKMTFVX1TT1MghPq+nRD4+EOrNYUvvEyNQgzDTjXXAkUZDM
+YdV4ocPliJ09mZBgtJ2RsChNxXkUQmOPdAfLRk+ecteTkIUEuiBOzmbhFj14cgb
V5h+EEoxHBArfXydZfm2cv1THVAoZK5KPZqdwQOOX7bpzT3/kqop2UfOi641Y6U8
yKyT8MFUCc9YhP465SfvKSHXWYUzD7PG6tl55LPWOC2NY5B+wystqOfv/QKRkB2y
oGMz51gyVGK2KquwE8Xcbu9s8qSVDLUl1MKeOq3Zdlq/UJC2sP84mHU8Q3+UXFL9
/y0ObCdhuZk0LfArCZlyTNbaTuLxUHiS/8kKgbv051h3sluaTckjN5xNJozTJQyd
DAgnJwSkI2M/o/97/nIgt9F2VZ6A/bMwK1pmau1QOb89Qt0jPetcfJclbiKbc1A1
rLzNi0uEr0/b43Jo3IXkwLPA7OI8aYut7PvcTmEuxSU+4zF99InPjH2k+25Bv1P+
LYa/z4J8dekxSzksMgNFpRdX2MEQLaD0tHlViJsEcHlji89oGAYAaTwOE/qq5eSo
6f4UtDh02O2eLBi9R/wEIpvJbD5XONyaN5KpFHDJtPoX5hcu9l17SDfYUuOfIUeL
YRNZEfXYQVdgAaoNEkSdlGZK0olL3AP0xTzK9GfoQxXA/IYSFkq/z4eOyegeFIBZ
CxiHz2USSrfCSP7NYV7Sur5GX/8FI/nZ3GaRwA/md0BtUw1doWPh2HF1i1S4828n
/A9DVHRVT30dmoa59CPZs2UL1GYxOD8W4tnK7UB8nti7AQjUU0zB3itPLoPqM4dN
7drCFg+FBsxeX0moNig1dae4HbIyg0dO2aruD+FgvKQMjz6ua9ZlYs4OLDkeZW21
qat4hDx37/BUmcFnewpNquq7CAkITngsyrzpambIB3+0Rl5dlYHjeIYlX+8lRadC
Gjfz3S64s6ZXoCtLTfsOj/M1lHvVI+rxg8zHnECJeTCHC8Sc+5WiE7nYK/uyrx6r
uB39ZzgPmzDVmmUEYu0Yh9ME9OzNEYafH1ZR3wHbWiz2SLCi9jFzVWafdBKH90Nw
iy1zxizw842S91qaTJ6wqliuMO8FI8ZFt3oc/3lUkvdtZYwy5gqD2V7pcNeolTOl
A7sd6kRXqC49fMdgDwQp1EQVvLnlivWZRJJPWpzhx8BHDAXpP/BME4eqlmydox9X
Odp00mPfp6q5I+r96cBIkh76qNOfg1R5HQ9GcvsCZTy1XG92+I1e2t00yWlZyRjg
DbP5jz/CbuxOqILEjYZXbsFEBwF64WB9Ow0ksJeo1tPVjE5D7yQ0O3caqUSC4YZH
Ilc7lTwULr83vgYeLKG/Zl0aq3kJHJVW2jihsrCN3GlP9vnHN9OpyiqU1fj7rHyQ
j0nS/7fktCBtlZX9NrHP7XyugxNRHlXab8gQpTyJs42wii6JpLs0mx5qQtU22zzf
VBqCy1UrA8XzrB+hChwYjDnRku0oq2EN58N8M4DOtwyyBrYAyFL0Ie5+06SN2dCl
/rn/TJJ5FcE2gSy4AW600VeICrsUFxpkmrYllncDtvbiYMUUWynkKZzzAE2kRxNj
FfKpREEQmHSgVpuPI/TWJov5DX9Tkg5xwNBoR9z9aF5NxbOtJvkJAEw2RQZNXJ3+
4vjH2se81xFG+AAQXNZJ1sWUT2iVbdmBZsxzAa09Hb8YKLhamyi1YEOEfpcGrFo5
mMUPZRgu5SB7qk/oGHdNlv9mZu+ly4Qf8XCCkcVgD/1DiJVgI2GUoSpSgAi93y9i
jJLmeMfCWYsTkOMnziQPTdqsYUa3qcP2GEg4WTO5wnLkszBPZm2zsWUPpycC94kJ
Q7I0Nu1IFyzWBZN8tcPa+W0Psd+h/AVhUO1BEjlM0tomN9Fg2E3dNNiQh1TQMoy/
sNe3Lp1I1A+ic8a2jM31vOsXbLwSkKhfMZwygZkHJnpTlfJCppFbQeVVEvVZhPWy
eCAqExpu07Cl4qm4NJsxlKfW+flo8Lfpc+k8rqdgXxp0ZOvkjHN8C3dYxl9f+AyG
j9ovEhvrlIqb7zFIpasQ3muJXr8/02+PQ/+NfRtGRDom3p9ns1wsrataquFs8zcY
lFCV3GLa48JDNrmOGesR+3T+ULc8SDAiRzchD2tcGvCaunn7G5MYLsY6KpaRRt2m
WyMlxS2ZiKp9ArblXEA9qkV2uF7gGjCsIceBZivvTVh1/AzTStcJiTS5cNbnywo8
LP094FkW9X5shKJ2nx8s1tHnsesZ9ro3v4c0etw3IFKg3UmEidoy9aNkuIUnqz2x
HU9fiqCU5SyBH6QYr8zkfjtQ2jNZWLuHP6pfY2Da2sc4Dkgtf2TbAxM+3EKdv34v
iwAbIStHSbFJNsRSJoT8/joDagWB4MMhEfupUI6EHsGboE+F59n3Z/q7v/vjdD5o
JkziHVOCsZFU+PT2h7N7YPwGzpgJydCZFL788n29CXD5NmRqjGE0P5kQ+1LpPskR
uD6vdxsRKZnTqZaL1gjA7RieXhVvYDFxRUNf33ZnO+hn9I3ahU+3bd51hauFlFTi
HrgwpvXLRaXFXneY9fGtZXR+O85ZVOWN3+2UgEbYIgzFo0Peui0MVv+lALVJIsAf
WsdhHhreDywhU4kj2x/83lo8bX85s6Vf1kHWDisHQYdq9X8jePwKfdAH8ZBdtUuY
5FVtJ5DFnEK8zM9yOxTaTFLiryliVPrRomyXqfrFR8+YRJcBCwZQx5n7JKz0KH2D
3y3+BhbyD//0PaPnVay2fodxMfnyip6hVybQ3jCRYjesKQR1+O/4keSCTKPu3lDg
efc5DATKQfNEJIuHPdbpmkJOOCaj/bH5Wn8ZxjjRhB3biScI5aF3YfrvRTtt0/y3
CcUIdGKSuu/ylF4kQ8de4CGAde8vFcDlWOs5NJF1PVwcHk1fbH0cbV2y4+XEYw2N
csk7/89yKEoSbDcCN32zB7NZxp4b1YfosdfEGPLp2uF5coQ48NQhINS2eirjIick
Unzq7UIMFsLw92mXN2SajnZ7o6XleVSQNQyeeFwXzB9aJloMIz6ChgsMoBd2EEF7
9+r3iXySSmvi9UeHlNtnZVwwF+sHBTRaLCuuQU4mGwMdR7z7WQK40dy3nyAKrHlf
5EiDGedhsbDhj69shkbcbo6ndZT/ctqAPB4X1LhbGd2RNY5UXA2OWhb7uftxspg0
ukWx2xQLEHF355NPwPqhYbqsJlzn1m0oq7Kk7h4tmRZ1KPh1noWzseU4VZhMZv4I
Mb6sOi8AiLeOKwj503KVQHl9d2yDJ8Ys/Y9x+B4g5NgvB5GZ3KYwlA+0vV+W2WSu
32MaeiUNA7wBG2vl/EgT4YuV2J4fJk7h7SVgUgNthBZJInaVpCz/ytZzYkfL1MnD
PGSbiKcvE6NW1022BqfMHd+4Yi+PvvPcOlWbZu2uRWBNuW58SWGiqHZ6ioAh22wx
Lrv3RCInBOnn4dRCyVMf23fS+tRzyIqaMqcD52oHq+t6OCTSPIkau2edvEWQ4HzI
1Um8OhOXnRJlvdN3rCKQOtIkQooSsvkyvg5zDkmb8BL/waa/nb1EEu8YohiWWM2o
reoF35Q38W+qfoRV6c8IJk8jJLuAN/9z9VJNwRkR+xpvYHCucgFbwW7LBgDpuUTh
9hZC5qTc92BvxGPPoBjBFjoeniCYLyqusa3ER4mPuaV7o5xs7gJy2SCp1HQxLcLk
GM2Wk7Opbojgf5cZHMgiAPrmg+EHUgOaopT4IffCeDu7LLYwzU7xZiIVTuwXo/3m
g+hMeb1B/i3E2OunA5RwnGNGJqUsRmCF3X6cgZEqvH3HEWyyIAHwHMcC40/fL7Ba
ewm4OMrKgtsnibxYRp++s6kZbpDmHbcZBZNgws4zhA5MObHle50ECAzPTB/SZYNO
P4yUU0OB2tyTvbrg3Ey1lWQQqe9EtsL6D4pnylz3ODHbF7ggeXuRqPUbJtf4Vq6Z
WZsDBIWLYL/qMjDK6UjIpl8gJNEg6YiBEF4QOQoZ3tVRKIapjo5LpCD7Od74iDJ7
WxkV80WHXUdkEZdQxnv4jr9PdAjUdUKQ+8Mv3yi2Uq7reJiF6CFQxO8v4nYJdbHs
oowoWdqU83RNLv7wPf8ddVV0mb7yZUwyc2k9LOP8/a66R/ynBlLbH6GUCV3wGhao
eh6aVaisYzljZr/hVX5Ou8MF4zT4aEIhJd0blHiagxzBpMU39RtE2AwGAzgfxoNq
KtIPVbZ6p0e6oZlTPthpYPWkqYyXwgvtxvK9lL4V+hFvdrKDtChqeu4nY6pOLXlf
hYLZIsvY1296yHBwg0lReNR2Yv0hobaxGQOfgWRz6giWLJHczg+IKlWq+wD0wBQB
7yFWYGi922OIcbWRglSHOWyj7UW02DlsGW6pcW3PWJ4uF9XFa4uq8LKoDB5A7dOp
jId0qX/dTOCBayIZbrm2XGBo4LsVha3NvXF83Ooh/sauaNswDKbGXwseRMEUklds
Usuz4XwXiiuCwPhfDdn7xChsdwyzWqAkLHWdeBGR6H9Ux0pYR2zGrqCmoJR/lIGy
KThq/ROuEBgl28ovHSdjE1hlhEVsjXSGP3X+SOi+6Ia7rWJWhmEN72Z+Q7vS55fq
3HHzU0baGHIvrhGCzQLwYFibCFwWS6kF8gsraP0tXoHsPqBZe84IMU29p1zJwEjy
vyLTDadmjQGzUQWkdYV8OuEUCTxvFPNcN/HtWfP9LEtW8ebHJ+/aA2xIpnyprgt6
P+B0+m6Wu88OS82K5IizJs6NtF9YBoM2KnBctF0UCyDqp3oGS1hmTJ50UlJM4CYH
e7ungmg/wQ/TCZqdFR22t/3y0CufMuxukZ3fngpBZcb9M3sLZXmPVdxsTkhdCKrJ
GwCaRCJYZTJiQyEMINJt/DokPHfL5vfrzwZ4LWUDXWO9+ghylFYTuxwXMLRAp+xq
tTLBA9jFIvr38IeccrProfL5ZlS0pHuhDQzMOgEuXfJ+/P3lnFb/8y+in23CoXSZ
lpZsxnEhdONIzg8o+NOnB5UetVr8x69egy342Ig29LAxDuOaSN1tKA9asDxNRemw
OYenMtL6lwtjj5zjEVK1ldHs9QkA5WjhrNFSzU6QRgAKRftB4HylF0jjwjBDAQzn
d8ETdgPa0mhNyFxh+L3lnkq4hxBJXmROSpGIC9VFoKx+pFmo06OGmRcaHq3dr59A
atfpntKTuLkT/GLa4D0HK96MKeZyLU6L9Bjev7sHP5NyhfjXn4vJi+YvPhLUWmb9
cYi3VWudKYCkxjFcUI+oxF/m6ZimeOIjAzblxauTWkFuQAYV+8Wm9XxCFfJXpFM7
nQVKkQQHIWKTWAegVz3jctcR8/5Y31gs2FDqltG0X/6915TBb0O1vNq68a1XaP2w
VBG5VsJl0vLeskpF/PMwBsdrsHgcxADdsD9ybribxwX7jOtFLBSam5lRLkRgaYG4
X7D7Abw1mQIHrJjHd9nYDqc3P3RdNiM1OHpPjmxcNJDj0r9j2llx21oTT/3CrIlo
xr1birEB5qLhwxMeIb+j7msp90S90+uYr/4BKgzRgjS/efuNCQlh4qWcAIszReuR
WeFP2Cc04lM2Bwr4ZRMVT69xjqYHdy22IivNy2F6yRRT24WJ6TVJmwK/ts1i6ihT
fybx6nCv81y2vpUYzNGkHMvXA5EY+n4Zft90SZKhuTppjp6PYQ7rRKHYtxR+W+MZ
UdgtqySsazbZ59cN43IBjmqGsCfzHYt2bfKd6+VkF4DYrynylzSJvo5s+5t5QmZw
Lk3M6SOtxmKtrSxgkC0JZlnJ3LSWstJ783kFTyQEklx9J+tRGPCEpLeJeWlJ5EK7
l2PVDDLZeCKbNZV90YlBV0IrRzFgCVFU4WD5bQGuSTihxy8QfAuEQDlPfd7NWhru
Gy1C5dBg69SQdG88EvsD95KJ4sJpob9Fj0GK+XnesaidkHlf7BSMzrMQ5jsWISMo
R/S0m/L+8CPhViyZ/+9HV82Wvj+RbZEUMJsg+xJ6FCIU1OZcsD9QVdMPXJbEVkyq
kv83BuqND+9JiR3kyixzYXHiRCR/ixbiZychjf2Oavo5ABwz9OKsqQfM5ZHnWOtY
xZ5z40ZAhBiHNbcZSacVGhQPk7p0kwcjHHf2E26ni0ZwuZiZrmpEWqx3wejPzkCi
7QK5KXpEUVDc2GbrvUsem2KNYfhatSc/lIclB9o0SKDAPTFPBrp9IK6oihMB3mtf
qhLm2EGsr1YI7cc0Ex6wxny57TMRg7PEe2cDJbxxLvCBJcYYhxwtxC7RiryaNyYM
kD/pfPptfHZK33eTEySm2g+08MK8BQ8D9gBfZijBu6dQWiInw8RycaPPJExQUNyU
piyc0+WzemEyAmF2H5O2xO0nkvC6Mc0IX7gaB87sAgK0fFDFtHdvbFxek6o4KNkU
AOI1jQmoFJaKUjP3AiaDcrckxP2jQqVinGIbwLTztw2REddbjsYfAJfgc2qFdi3W
894joiNvm6OXJyqAcWy/64QozA8UzjX+n36Mz7iZpVq9GAUJiKC9GesWDlSV4jTn
Y7Qu910G1ruMj8aaDVkeZod7D2lkLa6aagfR3MRVCJULZ+iZZgjNTU7PZMNupjhO
fGCcxMn6D91/t/gF1dDu7zXYdLee4amPx1NUlDtasOgRqf3U21IXoaDSRPs2NOZa
qIWu9O+KnPGTsm8Klh163DeZljUwflu7zUligtJDeCYmUg6c6OrFPzJtXqZGaFbb
EAjOsBGzY0ZvG1mm4V9O7l3TH5CAusyh0jq/NW/9HK5r//b/iCfmYXPN9tAhtBuf
HSnENLOxj6LS7roqWO3/ic9Sf0dzV89FI8qalJAGrj+zWjyJOmHYR6IyfR0G/tmt
Z2qfutE9k/y/pK00O1zbS2Cad0YzM5scLJ2RFxlshMTFlpLuLXTxFn28jgNOpjH7
9iHdhcVukD7nUJPANMYeVBc5q8Mo5feljQVBarAihfGwXxjDhjMCc5sUYDT2rSfU
Yh4WRE8im5WsobZavT6M4T2aEkEZdMAFtjN1gyHkEgLMduMOp1CI+Kq01KgAjolu
CBSzqXM6vyU0NBf6m+9DU7Q+3APXrUh15vjPc0PCsHaLycQfVNvHSRjwGNdNQWUz
m7RVkJwlwXvP/xiFhHG9bps/Cms6/24hHFEW/hF6YuPlygEbQcJEzHS2ylm3RpAN
OPeqw8HO3LnnqPdf21xEtHD9jxlGojiBnMY0oBNO5/A+R8fOpOXdI/m6hJ7WwGA1
5y+0vSFsGbk3acqafWgYNGjP7aCNkeZcyMJe8t8hw6SLG+Auo7BVYL57jiQXwGLq
wMzgsU4Yb0xj0BEBEATmogwZ66KZ1YfZ58bsgCInwMOKsBwYUOOdoznAiY8rbZYS
ZkAweaOnWV7uLNaad71aFQExTVVC1peOj15Fe1W2rQ3KJ+gsOGwrgD+gmZ7xf8fr
CrGJQsGKLiVTNwZ/l3oV8JaNKR8UA5/uhltfTy9gPG69m6pUZLiYSkqjAdwAHKNb
u4xDSLuF6ssW+JDdkMWTVeDJKbIUqXfCZjA6Fi7R8W54BBFQmdFGiWDG93BDzjuL
8tbRWYnYWHBSYhlVxrK2PpeVsbir6IOLtHHKdlQbmBolocCUwF7in3HKw2Cv638m
qtToW1wq+cuPWbp7Pg7liWYDFoIc2SYcR2Rz7cVBHJo=
`protect END_PROTECTED