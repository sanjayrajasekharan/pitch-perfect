-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
YuavL6fQaoiURRxhU0QKzlhWLa66PRprdfN7fLUsbcQKdQtjiFGkjDnp3Zi7rXJ9
YeqFt1EMEyseFzSVEExWBC9RMGWK9QL1oXogewToSEiCHOw283h67j7Xj45ayOeq
Ng+cND7taZtkeDy/cWPNepowHB0r+rWSA7Ihth4ypVU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5584)
`protect data_block
WEZvOema1BIUcta3DVNURiItn7Wg+jRYPM1hZsyBaU6Wuc2EiMj3WYUEzX2Nxcsj
hu+cS9xw5YmmCMFYYgr6Vl+/JdtosK005yzpHBcTYti/VamNNXyKkmYJzLqwH0b3
xgNKKZpmD0iUbdjK+LM/plXtSsq36ov/0mjsQkFpj37PIV6ZSIbKjdSy/Q3TPgeb
wR9Cm3FE7FQcd9mM1djvLQeVlTvR/0DajekZonkm+rO9G8ZW6wZ7IGEyZgKRcWqX
S1pvVUdcg9SrR0kD/uOznIZMRDiLUrsCwXooRRL6DOtUGLhyr1JSmDJv+tr/DUu7
A/anc0L/EKmPI4mFnZasBacXOi7KiG+q3aTb+3l1GXwKl8Hd363KN6ELfi0TIYQ9
1BHJ23tGCMzX2Q2UDTXeISBgqlBusRtVTKC4GW4wN6imO5ik+UTzJpfNAgeTxZDF
UWNqvrpDsejv4Moz4fYHrQOG7/lbAdgN0c07pwB6a2JRzKfVHo2Qa4VPZhmXqr6F
v57dz2RMs6ryx25wNR02FliUC//K23Hn83rDy+HEGgL0Y5fdh68F8dDcl/gJFMnv
oUjNXRts5XDBFFPoi7vdurK1WdIfQSPFBeRgKS0ga70QFfh56WVsHcjeffU96QAk
RV1KNI5Ygu0Lq9Y4lsvyxFCNf28vMnFBTtgS6iEYJPJvgI/SZdfXE6UP65aDqWpa
omQ1kRi3eUsho+8gf7wnAC+VJ5omR80GZJGBnhsMpml9XDsCgF+w9zVNEbJ+mIf6
Fw+V9QGVgRosRebU3PaOvz2y9CRJJDl8i/JmLYO0IE7Xl3OO0N/XtPOFQNDG8F//
WvmphISyFdfgsVm6RT8ShuY5quLmqPRQ7xQWjpH1/bx+xbYLq8cN/+a+nCGK7oR0
ZtM2jwY0pQJ9kE2W8o8lzD7eOhET4FZH5VW17A/Ta3kk2aelq9EfSvGe5vjaJj/T
gns9bFwAvKHpRKogNhU4vl2Tdyl/u7h1KLSuspdDjScx3pRIDVJOMQEi5aQaG6ww
jYTDsZaCxmGiP69mwXjx7w4TfqphFUpWuj+B3DwaUkEqic8GTwMBmq/+Fz1vX9Nb
XuyqlxfVGBbF0RYCJnHXzSdgiGZeHSJAE1gUfH9NIHYLpswQQokNVgmSFr2X79w7
Nb3omtXHYvqavk/+7lLtpaGP9Gre4gpAaXppS7HJnNmJM2En/q20Ugn8G10wb4Jd
Vrh0YvDNBIr3ekkRawhZwwS1HaxYMzw6apfQVwO9x5YDvvXTo9FGiHD2DEZaslRe
ksA+My8Zer9x+HrZX3qn0r67LeWMdqZ9kjoWYuw+22QvzPftm5/UFR8R7mUOCLcq
Ja/KQzSbAESplRDi8bydupfUSZ/covlfgJt4m3aSqcUpuAS8BXVBvyyelQaTiBi1
w7/s60O4Kv9AhiAZHB5AO5ZqsKI8nEjPhJTimt4VXR10LqmzK8imITl+YRQNyu7b
TU/gOVLJwf/T3FkmUps3J7NfD5IQeE0060+wW3gqM3xSNJVlfIMAKxSjTUwpT+Zg
g8DlOVqZ0pdci5hABygC9xpKb4kYxQY1M+BlxvvPwzGCGUnwvYOY4wziH7PWreW2
ZuTbzPpDmD+ki5v5SdSHceDA1Im68Pd4FVP/Wn+IxZPx+0ufoeDUSU8GhLBc6aDS
M5EEeVJlW+eRmNwhfHk0ofzjvjbOssACM/Qiejo7NayJgXdq7agJo+C0W8BgAkWW
n4T2Tw8LCy30CtRBiiu095Cg462hBNxtdUpKDynVxapAfj/YXFCiUpP8Dqww24ki
CPjzOsS80ifsnRRPL6+ZzmwL70kSOx2xsxvn9d7ln9hNBXLrrtiYyB5MdpGm4CLH
4p1r3fD7qiIrAEwXOT1gMq+5BZwQeRaz1iPO6DiAQ2mi3IkVa0oBt/85n2sX6dpe
ZIMHvVLK+FoLyHaNwXvZdZugJ5q7YKIEwzBscT9qpc/yiH/b2mBMau2cJpffWyPy
0qGzh1Eb3/VF4lNd9pPP/TLo871G9xXQuAH7gHjh2BFdL7T8IYdxBL1N5YbpHJWk
Ii8OHUIwtdjyWybnpztOcdOGODhFQCRkRl0viqcHq4bPWxcaETmLhfkLUTEjHVo/
9SwngD4O/XoaGiKC1hezvPxmWOtfFYrjpYWJvS69idJN7ztON2kkt6H3ylc91xwU
2dTvGC58jRcQxSZ8O7CJHwXBBvW20li/qH6EHC2dr12ai1pdaC9mvGlLBa576OWY
gmZGvULx3EiAlbxRB7EyFa3XEO+JEsRQhorwDA2MrUl3WcIfrCNbLKgpnug7qwvZ
RIk4y0KRrVduJ7Dv8lVuxTaqiXzT+m/ym0XnRz7yzaiVlHLE5ccyjRhu2Yq8RZJy
uXLTCuRxwbeO8Ucfeuqm5UAA0LONCdN2PzkLdA/f/F5Nqx6o5It5oD2IIvP5HeOj
AocBivn5Fey58HlbV17q1co8lRehGFMAAxUVXjiHm2iNW9I72ARrwzMU1T0qTrSd
hDOhHkDxEyf0z4VMvetB+rLw5y12QtxBtPwFbznJo4UD73c7iQX7vCJvWuwJM/tN
hbnu8a+uapR0pVBwZUeQQrd8JMmkuwJZx7jYste6x9RLr8liK81mE3eZU2Q1LxIo
YgzYd7RqqteiLTUGMPWCpXolIjKNsC/QblI5IufqBWCMurjNgTjNH+4AHwwWU7w1
QpeXOZ0PO4R0n8MyBcvInc90fPTgWhxsKDL04VRVPuDSJyOIvrut51WUSyX0ys7Z
m2qTmbPVwqrlyJoUNTwhfAhsIbR90/ZUFN83dg8h7TtEvOIzm4ivOTjV+1ZDnUb9
Xp5/vFwMmDYdpfYI37nf0BgiyiNhWsDFuTvCieEy7tzUDHZX4ZfJeOp7yY7m4x+f
5+GNx5BqdvSmMgHKyr7cLkwBFdDaaaKwDsosX061k0OMtlpJtr0mmKWp9XcLXmo4
s+0YrA0SLY+bwrEJmrAClL64BUF+b7a/twkxvDhGAOrLdDzuCbYX7RSMlbaHP4Gb
skD6f2soKBHrRKwmF48v4fJO77EAWU+xGN4jVH7zOg3B/JJ2QXqFxzw9Gpd1DcRH
NBxgIMBpvik9NN16Sm/PS9oZEK8T8iMtMBDvnlJp+I2KI3XVIhNMeHi8hEW6pF8q
asGU4gCdbXumc9zBOflO7COKYw0B9V/R+xjgOF1dJoFxfEKYUuV5K+Ql8GTL+4tO
7RmlN6W4IWwO+SyEpvy8N9kbi26aJjPfPGEhrjqGRDrgWUruPPPwnJLpu0PN33v9
EcHHyzfYxtCTZEBOkraN/1VFoPEBnE3KGxZvyiBPC4nHT0SEXzVhp2D3hpbMiBaX
8Vl8i43IWe+SQr3KmdNbSzZW/p5eeh52L3RuifsFW+O5EKOZx8bLiGSWDgoqWLcS
nlxqkvHIN8PbPaJal8eTItupwXvSwFdtnI0BNEnEJJCLtyUngEx0Fri8M5oOShN7
mxaOANA6+nVlZtBSGpgcR0xSwpJmQ6rWGKcrEmh+OK/WzKk4pwpOrFhf8cbZ/v7A
8grur4GeQq9w5SQvCZWHhb+QuCD1ItW2ks8fpSlaOHdJF5aKv2q7g6NVKPcL9Wst
CGKB8hWAfsclMJCklEn/BW/8q6XmvmDFuR56kvZjmUMUUm5B9YSB3xmQexQQ7KAF
EQIP1LDIuZEgPN39wjnvq/4G9dljeZcT8lwTjpeesaOrbwpkNLeKqUX/NaNuamEX
OX4nhvLMH67tEMbuylZXeufpHZQt0T3hfguaCZOpEpCZjLg3jZdEqyiwqeUd2HZb
d6WOlVXQZC9HDIaz9TGxYDXSmu6twgKBTxFpxZZ8D+5+7y4mGtmhjI2nxGLktXyE
RxOdLy26Cq/3xaJrwFDCWUBNG6qrptq4cl/lHhdFZ7LqPB5JorXmG1vsRR0iO+B+
Bv3nuJMV8NN3NTeMVAzhWidHu0hlhE3kFlKifDA9Rvcl+6rT1MHjTURsZAtx5ODD
4PxzCmUTc/euevyJEi94OzVUwi5CEmxKSqVzJhZlkWP8Sni5QGUO26sEsAl1FxaT
2I35nIaIUGvqunPkHozvl0O4o+dzcP4cbmZJMlGlWDMJ9zOMEL1GSZKSlhF8rYDi
t9h6slNaHBbt+EGjv7ZG/WXU7sGGJbg08HTdXPxfL6tVQjuS8PUwJZBjM99p/7BG
bAmEbCbyr+3HCy/NfYFlP1qtJauDjfl1eXgRhfLT0bPr3UoZR7730OpO+Y9cX1Or
lHE3uDKWvo2EfURGcCVH1Oro0K/gELHhNdt7QUL/J3mZydQJ3hDvv7F0uVwECfE9
TMMzOJXRla6knZNTYb8m+qFQtOMGLtZYRJc8GIObTMVOdejynaszNiDcc2Wt1+Cg
/kdWD6hUsDwB3XuD/xuk2jhmu9L/RljvAc6Eg8RvHD8mygBBECATKdAVHmCBsn8P
Y9DxLFStgZigVpZoM58DzBOW0ftljS96A/eKlJ91hD5JOtZbLP7L7x/tumpbpEh7
2lKfDYldqgIGSZJSRpiooHZ7FGIheL4/LZgdUiAfhNaRv7/Q6Y3cKpbmHyNhAUga
ktnp8ggvbdOrVChbWTrQi+J44MoMp5RKIPl+x5QL4MNDNo542LU6fV66aLcDH2fk
xmUlOwcYqCRb9RC1tLm2P+vA3HxQGQnl+BpUc3mLEkHQTOiyRqxe/IxeVOBteJwO
JLOuSqQR7JAFgS5VkEMXLdvrO8NagGGFotbyZTCu6NiijKDRy2pwqB2UWpI0ab0e
ccdlR4ebTAruOT8UkC2Gg3n3hjFqhzaGtjILoM4NfFWT8KGJut/mG5mTYAR3p7E2
6d7rY2mML4uGNrwEt9clZVeEmsQBkye6Vum5RvB4DoAN3PqBT91jEURnhL+cQoSc
1e0HTUQwsIu1OvvR7oc6aGTtgCu6gdCf5cY+12RVu43OQTquPKg2tUC75nX9TYLN
07BSvpXrZsEZysqkPn+RPjIPb1MI2geZ9RrZyIf9uZi9AeCycnwa1569m1d6zVhX
1SYgg6Y2RofjjeHSg/Gp41U8Eq+nMWPpgqYToUgvTrwrCNPbFQ7SfLXkwEfRBy6K
aSCGrheePP/3q8y1Uyba8DhiHV5der0+j6KV59TB9AXqaIn3Kil3FjnC1BferWz/
JTZVNbIRPs4zai3Vx7qQzrsptKtJ7/IT0bF18bAl31t5faJzlqw3cvJhNluU1OMH
WDmTtKv9drF4U5qIDwzqGhxO64tbYZCd+tHiDHNVH3kOLUm+znYY7Hulma8fEPox
rLoDcvAD1YdH+SA3gTpKS4uPp7uZlWL5+g8DCCc8aj3MNYEyx3tz7ZoYezOh781w
bl6NmU/YeX0rYrvr3O2ely2FJNF1rBr+oP5Cfe+TSLj76VSjPSorQlxjiMJtsMP2
aGysP4a2PxVfdk1hTduXTjpXyxkBeKC+GkrSTHW6FIx3i1UvNElytgUGQ7YueFzY
srF6KZMVIm83BDIAh0CYCbqT3UV8aJ6N/q3buoQ99u8sO6q3nsA+m1oW0YrdXxHv
2CpbkaLOCPnDTC147rrtZAeN5qWhMTDQQrixgkELCrJROgDgjZ5Et1D/MFcm1GgT
iTIoYbtvXA4+mLtsisZ+ifrfk64ivshH0tZvX3mI5LfBH2HMx9S1C5YUJABV5fsR
zIiDK0/MoMJASC5i4N707NjBGK1kYNMKZbIxLDJ2RzxXsx1AJimXbbwwJOWm2IDz
ujgtRyHNln8xoqnGmhpFHg16KjB8J9RkOl1UZddbbBVGyjkNPrN+Dfb4DY6cccvI
HmxNevkZ7OKP7hCxQzT3o0Z1u6FD62AJIRwOPqTFcs0A7b16a8QCBGt6IY+75RKk
7UvYWZ8VWowl0Bjk+eERKcjAAJImxYe8iqHSNYQQPva8+954rM2oWB9zH+pbs+9v
XsGsZUlPp5dB/VCC8Y093Tg3k2bRI0cYTrkOhZ8j60NWPcRSoD+A8gny8s/tjTtS
DtxIF59cMqCgNJQy6JGRZjPt17Qslpfn3zmDfzFf2ViWYMRlrhLSmFOTPMpFvITK
xHiTQUyvcF+Enzc5hpicipx3MGBezr22nxtpxrt/VfFh4665ZmluDZ9FRMj5lsNz
Fs39GJ9IRZ8z8CndpgKFkI6rjPib5lMurI8NUQ49Fyss/SoLZ/KkbQITDVgmOwvR
MKn6eR6bRiDtR55KPzGemH7ArMdCTK4Biq9CEgPJs+gpxrwTYWBiQxOVPk0MDIdt
mM05jhuvUBTZJaASiiVacbo1OUbuwIRfZyL8SW2NFitmnWwyM2B6/OagjuR8RryV
vLz0ebUmiKTytQ8X0JQlw7RMNPSjeIlu1Spx1mrtReYREXvagQ19KkUKvG6B+Bfq
mTJXqO03/24Iivw5OJt3pnvtaMcW2aIqDqHQGy3LwxLMkxTzk/wtop6GYfajdHPR
snK1rg7mR++4dsXBdikzzRPoyxhd3VFzxD/YhLV8idoNFD5tz2KXdgRmUKICjXSW
Byu22N5polY6uwYuIY+w0tIRjOY9Sya3AlXmhq6SlKcXXJIdnX8okrZp1S8FfNLW
cM+FH1ixCNV1Cwu/83+CyIff+CMwpVLuDS/8dIUaKkUy1oJbtbJipcDz93ot9vbC
Ciibf1K9H5niAuutStTX064H4pSyoTx0EaQ6x2y2YaAlxbTRc2QsT3MthqPuUjG/
wbnJr+H4VKjs8eu9t/tlUOf1xaN0zilAb0rfPwl88G1ZrTVB23iPhzLztIdQCAes
GVlyDdwBqXQYyrz0EK0k/cJ9AJycnZVzSdGPIY94tuyHn6UObYqC5oxBkRpm9FPn
Y354HpnPmgQhym3VMAr35X+x3aRAGtaxsKaGP1rJB+maWVL7BXFtXZmOQFQEbuWz
CULx1o1Xs5RMFTsBUxhe40NNXs2bT0dluOaPkntYJlE1F6PMXfuo1Mt5Ds343R34
jMj7BQNILSYCL9rTbmDiBVPwLYPZq7mtdAGLbDGqH0NsRQs8NJK7kMFFPSQ8CqZ9
+cNx2oOAPvsj7xKyTib/syb4KxRpMEMXXkck/TXjJjlHOm81fJrUnLcoDwJPwnmk
9Com4hleBULc23S0UlSGru+uNx4Q4TSZ/VwBfzWZenTPAcaErItVYdRl1w6/o+Ck
gD0S13g3HAXai14VpmimeDTW/WD2ZEuDzWdHFwfcaKRroz/2/yswr/5nInMJV5YG
4i+eAk5kYdC1B6c1y5DUBu+bnKM5ZLqYd8vysqRmefH7K7yfXov2WZXXnKSmw5yG
L9rwzyxcsaUFwtoMehtDfeA9HUj5gpEYoXNQJ1wNo5O60g0bDPF3xQIm2ML4M11Z
Lq5C6OW5+A1LDFMjuhzCCL3hG3G2veuZfHGKnmvW1dg1o9nPTLViDtxgyxFL0bc2
qKp8c4dfzV9QVi2pKzLX4RD9wmIE5SXTbyKTHRUZFKrY364Pd5rIM6vy0fy4VVCP
eCfkAKLEw72ENqU2UEET2g==
`protect end_protected
