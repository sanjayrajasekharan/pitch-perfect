��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x�O�=w�����v��Dwt��$�c��U9���f[W�`^�A��2���z놕�Y.]�c�3 �%��A�o�+&�Y�v�y4_�����:�Kw���U������B���ï���^��WX��MG���"2�!��`����IEx$30�f�(�@E]�3�ީ�~1H��0�=չpGn�`�h(�u˚�(��Sb�����T��~�ӯm�������H��^1R���7�8#ĳ���Fj��K� Z�%���z7kD�ME������вn7.�����ʆ��r +b��-{Q���*&m�6��R/W��n��	d��O��E��&�}�tf���O@Ff�������-lFX������gk{����=��]0u؟��+������+�D��ݯB�p���� ��1�UR����50��J?#Ӥ�P)Z��(�0o4�bP{�b�~�Ҏ
�(R��H�|��u�7�b�8����QOlK��ZS�Ң��f=��������3���ѯ���������ӂ��4�����)=��w��dN�3@ɴ�#����6�ٷk�Ogl@#��=b.��f����xD��+� �a7������̲a�S?�nH�j��_Q���Ӵ<俾��&��ǘ�0	Ǳ��7�b��<o�Y���ձ�8:b���D
k/KY�E��̝�Y����>:'�w�/6b>
�]% ��œ�"�^8�*��*�J%�[Js���j���UD��Sf��f��RN��`�:�f��hDd	�T��g�p�������e�����P����H�sT�[��T�n
��&vs-��#�=�ڛz�74݋���1'+-�_��h�����cz%)��Z��8�(v��U���S�x��;]��?����O��)1�&6�|��C6�y�~�i$��h�qïK��[���6�P�~�����A#z|L=# f��E���4��@�@�����A��)���-g����ܻ)�~'	�O�f�v��,��ED�������Xƞ�񗀈!��n�Q�g�Mt��՘9��/N|�r���8Я0j&�A��l&�1�bz�+��NPzf�=�7���Z$3�L�V9�X��/�ڡ�,{E�"2�9Q�[5mٮI�oB�@菥6Hˢ��UF2�jߧ��i�|!c::!0/�*���T7l���*l�V�HhV�0�l�/q��Cz3\mR%�fɅF2��F�6�ې��oiW��%t�Y�E���.�E�a^t�L0?o�x��:řC2�;x��Ø�w�x�+s޼�~�u�W+��yq�G�WX4Y`Ƙ���AZ=�x�!OA�x�U���l�ш�/r�n��}k;��=C!�?��!��}�Lwh�R��7zu�1e�ﳊ��W��%�+��0�������9Y�R�ly-�ϖu ��m>q��M� F��nN��o#�bu�.� ��j���G�)������Q���4$a2x�&;�)
Τ�I��C�Q������e�7��R�T@�?��
����f/�ݎ�C_EK�L�-a�S�bu��V���T�f(*BkM|*����;�=b�"�S��NZ����E��m�h��I-%�ck�T�(jV>���#����Kw��k�xf*�
� #�# 98�����؜�؁C%��/@{nn��Yk��K��5aM&SY�3z؛��9�E�|Iw�O��������O�0�bᑘ!R�B/PfŝR��;N)�ס���� Qi���:�jp�af�͑l���v!�����%��RS'f������A�S"�����,��z\l�2�ʺ��i�����)'[��B��(� ���o��n��c�7�T�ORi�Em|,�4��<�B�;����M�2j��.��۟�����P�'��0Y��5��<"j�a�'<���T��[H#��1��g@N��VTø���"�����F����L{���)�r�7��S�w��4�;+ar�^���\�a���).;*J����o�ݨz^	%WC�7Q�|���}k�e���WW�)�81Lf�A��>��n��Șl���x��E�;;ъ��tK�t��a�m�#q0�xc]u���d�36[����y�G����;I/��'�cdDZ0�\�U��;t�$���%�c� �u��gx^�z��~�:�wQtu�J4w�k��G���d����t���k*_c`^�Y��Ϫ���>�9h,v�)G��g�.�@o�t����?ĺc>�+� ��͐p4���*Z� �9��be���lT�����̫�6�6��m���E5_���a�*>-�j`Y�py�5Ѱ �m~��.>H�3n=���5\P���ۼ���N@�(_;>�N3h'���w��&$��HE��hh�/=jr�I&b��K�_h��<Ė|]g�6�_J�H�ou��bO���nE|��Һ��z�b귺M��ǁ�ģ��Y�*ρ�L{r�\>V'ׁ��yʩ���`�̕��D̏;���E��7���˲�ni�
��N	�sA�\��ǹ4�#M9�3����aٔ�I=RBhp U�����=MrW3�9�%��y�Q��L�{h��8|Lj6�(X�T{~vJ�C�<�c����f@���Iv��@9��!���nFy�����Y�Eco��ռs����{���än��