-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BHlzAvH8I5dUnLfmyW0kO3+vN6qu+nn3mPimCqN4mCBuJD1ww5eEUcR87EnmnekCidkOB3L2dhUF
AHVlnuuz3avfjGHnIIAd6+snGT1mpLMRO2uPL762iGF31btv46wQpXfmK1itjjgLuiDqfVazlaqp
Zgj0MHBVGsubIzxC95H1jKu6BmKzF6LX7HWWG9aZEEFhr2mlzweK0GYW2FKcqk+RpGFizS6lMquI
3pfGXQ2KaTp8bFwgi2lBFnXp/MVXX/nvyT/qCDYbUefLV1fmIpnauf8fwAnyIFq8FHfTGh+qMb0P
EDq3i/96eIUnNlCPg6eBIHkWnGIQyzNwmaQ8EQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3520)
`protect data_block
1wLmlH1bj/+3ZNqQKxSgQ2KYggSDWCWGokjXgHCzujyirTdpZ6K1gA8e1o2TOdkUh2IxSRk3PmO6
6ZFNvDwrA/9R8YCcMuskHHTIOsH+wCstr2RfUboNbJoEjftIRYpxGKbe5KTGZjWMfTlkl8EGRKxO
i5tC8dt+2W86qxjppmU9XpZ0LIRb+N4+Q/NhNr1My43jyBnbaeW36fgKFHkLnDv/+Afvh3mvNVeH
BYN7e5rZWNnYm++OZtnSNzU3f9xRQ2hNzC7Px1MkN3+nd5Kf04pAfZhPneVi7jMC1K/c1jOpWMd3
/ecdwBFrtpTb6rXCUH7XbxC5KSAYzAinz803GfNvVmOSLMZceJ+8JjLH1AFbAHA+RpE1LG4ZW/WZ
MTW4eJYcKJullroYxE9ca0NpBiykCo11HBUuWBwCsVgQdYD41Bc7eVRZubIrWrHxy/mJ5r8Y5Pm1
/Doss/8i7RseDZOG040xZN1/f7IQ8QMix5kfnRo/Hpg80HUf5YDALYQVQMu/Hvpw/DfxFNCVWnhk
csFtcpA/FT8204B/0H12SqKV9vJb0JFikwhyah4uqJKcTdH2vBI2u6HUVxdex6Gm3Wyk1gCbNuiD
8W0pb6Ka1zo9msvq8UibKDYU+BXzJxf7mcwT35aB07+Dgpv2od7MpshioLderpCj66ky1s1rCmVH
CBszeaf8ltbvq3BJ+Yo6KaLJ/5WT5pVhvqthQ9C2RBG455tvMogXpqJZEjJVsfO4CNPFGqFWc+X3
rPkMtAeC/qEJPiSf1xiPZ8sBGop7ODMzdiiatcks7K7N538kgaW+iDPWzGNVWaT6czXcs+J0YD15
o/8oKPjYKrmeLJuPL6SqDyDrtUfpvLgFSrRF/aWb85WWMlnq6mp4+jHvUJpTN4rHZre/LTDM2qb6
0ZDohP12BTeLrofVrRO7mILKqNV8hRdSe/l1DUl/bAAV/S8XnUlvfx6jwj2Y/HFYuJfEp8ccuIEe
pyY7OyEO6MLym61QaG35Vw3oP8ctfoAoQr3s+JTb56865g3FO+uqT75j4uJ1h/wLHDp3DcOOmCFl
krJ07E47PFuJIyUdFf++wBWNjMku9X/XVCDnaRwz/DKijIlq4M4EvV1ulgH3Zok+axl/2AonOmTN
gjidXxeVVcuXRkHvly5jf6x4dwf1UznVlObDn+/xaUG2NJLlBaD/BZRFSBVFrLUfpV1LAwigE//n
BYgwd/LHkvmHhXf5Ovyvj8mfi3kuId8Zc5YcvAIaTG/EJ6gK+xEPz8jxQ7eEUxAqPjmKI3kfvkY9
71SM9ML4zM50mZyp942qrs1FGid2yUdVxyRaCbyEbrxDiGkxxz3ZZg32YMMqSPJAxOi76U2XyjxS
OMCgj1jTkHDvPjgkRobEt9HifpelVkhBQYU7gBd2H3kAsbHYY4PylFlPYnw9luWD1OVRl2DEGIuJ
FDSGnfqJix/0SpUG/FvC/sesYnkjmjUW5yVe3nOoITYjJyCAHnFbsoUVQaAvWXv2yGPmpO953MJY
iVxUAr+3TzqTjIxXuHULyzR7jnW7IvemFjuixYcG3KEVuuzkrTAM3zbO6uwzIgRBEml4ukLt9etP
2soXTRM9vJ69t4f9563QmQGmNgAmGWbvUyeI9QGH4DKLcbISUZLrnaI4PKOdE49Gnn/x09uwPPkU
FXGDCV+GXFSLK5/PXSq35vGEHTFIlwA864RfX6STLISfEsje9DQGKFCP6bMefhNFLzWp+bAwthXz
5Nv9nNAnr1bcZF7SpiTW+ics1w0f3vKklCcfjY0uBIH7PWIs0CXpbdvf3aZzV/Jph/qQoccD+F3H
HHVeuCNun8pdMByloSbcyZc1Arb7g3DNmNpXqtan3G+T9pEtCrkCa+uxQJDIJuKPIQlZNIf9U9so
CfDmtcsR/XP+d+MOy3oxvOStMaFPYciRjDRZCugXhvVyK1/MMiNfN5Ce27Xoz2NzrdzXyXyzewW6
nqz1cLKEfpXVuSPaAaMb89vJAbXL8znvcR3uXhLyyMBK+ynA9zQn2MCROnJ1RIciMNC/OpHPKtFy
hSjq62/TfU0iw+M6OMVMoK//+EY2M8fS7s2GTEYk7GAObAONg8ZBB1dAwffJQkm0kldKDnVueB0g
YxZPHBMj3tyC0r0DmuFmr7XORKApcDS+Oq2WofHOjs8dm8JRGAbi4l7/JbrO46so/+eGEtonFv4G
YuTCALruyG3FpYucKWXunhvI/fDf8nyCZc/DQ2xqQY0GmNkmhQEBgJDsXrkzmQamMyJFLlk0FbCw
rN5rmc9iha/rpFer7h/brnUYwCDRvOFEQ9AZRlKjXlNCkdP4+MvTJo3S8xKj5ghEL7IPKT+jwMJT
67Ben3GPqGcjhFNSAbIgPTOjpxZ67gyJH79ruIc5XZsYIy6UwVvN47ICdhOcxF0MsQ0bvOlBOyt+
qp26IqbmZF7PaN/RvjRFEytVr5XNUrYsv42K9o4Ezht78emLbBuKjiGC0UuSKZYFUFF3g2qA5ID7
rT5soVljA8cThpWIWYJTtODt8f+Xee585Zj9Ri/mZweaN6He/Zr9CRTq+eQmgIqLaWMmSF5czTfD
V5hJ15Fgd8qgMFndemby2OvOJ46aD2tmvhVQSCA0hyywxT1YsQbxXU3dhFOV47+c0qe/fe2JJlSv
yilb6hCNQuCofhJ4mGHJ7uGHWWkp80ttG5B1Nfp06oxky3AXQVKPiBaSHS6h/b0PQ6Zxwuwt/uDu
HugghIHzSv26N/ijI64j0hRZAjuiXnS0sGzuHWriMY2WARXGfROdPITm3wbsyYKUyA/QrGS4r8tV
ylTv8RuQyZmKlopYEpRvzaTblIsug+orKSYOJdesxnAnidr2TwaW6SrYqAKa8+tNgteDkuSECa8f
UIR20/kaFbM3OlPULOxQvWpE2Hm9Dj+PjCpGYBCiCxo/THW/5Z6rOGhXHSiILID2QMoZ0p/OVDlw
mHSxSxWgG/+NtxuPZzkOJZ6BQbOI5z9wtkrLA0bpcrQDRnDNa2A9FDxjRBDZ7qWhxpZYW8Qgzb0G
ArLqybZZtfLZFh6DwfSKi/LB2luSdiEgHpSBzZZ6yN15dhHu6zc8Ni0q/uDSX2t40jzVSRVU/HLq
p2U1Apqi+DrI9zOlqsu3G+/SLUhuzLS/U4wIGkBmWfzNksDuLg8KtBngZN1HOiahJ1mbN/DaR9E9
5Go+iEahA1E02azKLpvOHOnM6c+TYUmQgpJWXCRL8MvdGSFutvpNjlKcAeW1+kpW/Km84tMoJAmt
Il3hLamYN5AXOEetp0YHjpz4pQD8RErNaQKM9n4G69ZsyRF2sT9LVrF2DurqTywH9gN6FRF6kwMl
bzUZd6opuUfpAUDaavz1pTAKkZPJBb9SowwQvlQDvcus+k82qodKpEsuFjTctXUPxAq/kWNfEDkU
ReHoeGfCp1eFCEI4/7MN6y4SLWZEqL7VsO1+qHh1DYfChRjmyyPxT6X4g9rlYD+W9/YsMDgKwZNh
OrS3DExVxtvYts6BdbkEwPV+VaYs4xqDSy6ZHzxZSPxu4S7KL1SpsrsBDfLyPDLyZXTOokWhfcDT
uf1cF9TwMBZtm8bJTxe9mss/D5QkxPNJqtQn81A+naR/nv4NclCEYxyuMLgxmTotFwmUdt8TFT6y
6l/Rrm5H57rmIwduw/Ggly8Lj4psXxooK9+jChjh0PROqJE8Ul5H/7sjFZwe4f5BnYnjAOf9zXlU
FV2/OCvfj8bhOb+BrV9On0xzbjDfqNwBfjn4nb1hG1MHjLGSShLhG7G+awitfoJB43goLMtE5hKY
Mn2tIpLD/aE6QRMeneWory724U+Q/88FD2RDS9eC09QMLbJWdixh2am0ofveDiWbZi7m4GMKMCeq
IPttVcZgE+5pXobAXdEVr/9lMHoofCqpgCzmG5XvHzSQ58hqn+lkqwuZev/pW1MOeR6VAPRjJVQ1
8wFpgU3RvDKQ5STJN/LEfWb8OmHd6J1Wn8oRI+r3YmX1Y/Fjy8PhUO6sLH7c9aTWq/xkwkyB02M8
zN8EH8VWnuV6g55Pzb2fBiRCQFQIQsF6i5T6uNDJcQJGNEVxYRgMnj1CkiRVm9rDwJlP6w39K7QI
Fz6AeOpIuUjb0VTs2bF/GqI2Ge7TaNKOtlRWgrkMFywX9H+RPWUWUw+vDaAsFhhgMUhPAUFz07Us
YUVuji5CgIMpJtJgba5L8v3f+smtTUG7naZ548/y/HWNqVrm1qHz0Ux/kXw1Az6TT70gd7iwDifU
9JUi6lOZHCt3BailmF049BairwngAUH4mTek+3p1oPJe5ygor1Sf/g/QtAMXm7YERPUeDPXxS3X4
RFHX0jqAZmxN+hclwDKcQSDi7lXQ6yn4T+Yl5VmE6i7O/vdXLc3WyTp4yoJjp7dBGm29qp3Hg42W
5encyHXP6xj+alQuTe87wSZHAcqiJKV44/yE5kwwrh3a55TZeE70AxjZo5r8OvinOlu2pAe+G3+O
YK6XWYRVXNjzR8qfJjIKzR25LlbybGzZgILBYYjd2ENcmVdLUA4QwholEoDhxuj2kF6yNONUTw4v
HYiRJrxHklNI4tB5rWSg1fjjzbX/68zIwxFoTkXpm56dxUg6XvJ7l55szQGzZ31FI+CtUnJ15f7j
kbdOn7aohlHgnTCmYmgcWD6ozjHeTIbTpdbGIiPZ+cfE8kK0FYRW/nOueQ==
`protect end_protected
