��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki=/�U����ef�\�����0�d��h��f�>�__�Y��0R������J�)�4˙d�p��.KGiʝ���y���S�k�?�-w$s��M��?*t� �b�h��]��Ms�&���I�(l�f*r����:U-�� �s/X��a�`}�a7%�2D�I� �|�B�	� ��'��2��_lX��7����� C��y�;a�e�ojq�ˁ�18�)�J���cmǝ��f�P��tǓ5��+�Yy��V�q��ֶD"��3��+1��.Ĭ(�	��E���±��ߩ���VM��]`�<m��5�ꈻ��G�nĮ�k7�\��X�|I �oF5�;�܎��؆/�N �=�L�ό]�9�1��"�%�Wo
�R�7����`����1�g�$�n��%��8E@O�"l�C����J���zw�s��3�#�C���+���
 kF�G2���ATWP|~l�6���W$�n��N���h�Y��7b����x�F�'���;~$¿� ���d�[3��G=�)x�]�Jd�Cx�X�1OMf��($�XͷjRs���"����Qݶ�'��RA���ç��������̀���RcE"�.1k�>#Hwg7�����?��� c�5����&�$�$Ͳ|]���A�.-��5a�����Ĉ�?�3�A�x��5�	���nm������؂:
��2�ؕ�ϕ���c��D&0�i���Zk��q����ﳃ�X�Ύ(	Ӵ���o��|X���Ƅ��GN�dJS�z��QRdY'ܲ�.:�9P�<rA~Q�)���cԛBoP鬋9~�d��8%�c�랂v�!g�=ͫ/ɣ�7����m\�,w�E��G�����{�ԯv����R�S�cMO�5�n��pD�
V�_M����>�-}����@�`�rf��_�5/6���p���az��b��%�L ��?�p�m},�O6,�d�z����8�`�s~�[ d����J��Bi��3�V$�PfR\����j�r<�{�z�0��$"Z���:*�zz��"g{����V��?�ܔH#Fh���_�ù�ya�T�vm��G�)�A�&_���ݐ�W�	e9�^�7TY�z�L����1n��@/��=MK]�a���}�6Ѝ�t+7%7��k��2ە��rTޤ"՗��B����΀w߶�O̕h�B��F��w����~�iqa���}��f|��KIt$��l� H���ВH��]0`:@@M��kL4i1c �)!��{��,��\H*���E��DM�y-���@�-��T�n�p7��������A]tv_j)3#u=��c�i�p���8��	[-��chGVde�#���^B��&�Cb��-%:	@�8��}I�=�_�H��Î4������u=s�g\�@��|v���`�+�}ݬ�͂ݳ#��u!�0���*j�0�l,tTd���{/���7�WV2d� ��KMJ��py�Ƀ�[�7T>���B�;����h��\Rl�䇰0a,�k�&KJ��h��\a��rO���;|Zi*��~+0���ێ@S����r\�����V�pz���Qfu5��q��趗q%$ﭘI�^��n����;����8�:���6�vC�����6Ob׮$z8�e?��Ԕt!JX;���m�JdB�t��>��G����-�|�Z��Z��%���Z�:�n�
���lUó�\�q�2��z=**5|	��&^����0�8�12Q�h��d�a�g2J�v�n2l1��mP���O�CQ��P����$uah��9(�3��o���$��}�my?5?��Q�4��ޙ�r:D�fҍ�>~J�k�������*�A<R@�;���p�D6Q��tBô�xG�1+$�6$La�U�a�(�X�@G�tUL�l�� �x����{M���Lҧ˄�l|��	��7�}�W�[��?`�72��	�ۇ�u)���TE[�e���(�a��.G�����Zn��vJ�VM�:-=�4Dǃ������V����v�cE�B���5�yE�T,��7
$�T�ͪ�ɢ�RNE��2{�%SO�q" B�J�RB<ZyW�`q����DĿ��4�FpR%�%�G��Ĝv���2�ZA-PmN�Ds��/���F�b�4W7���~A��nk8�N�B�ơ��/_G�ќz�X8��'���<�7���U2��$����0'�Բ��^�{��a�]�}cy� @!������5X��~�!��_F�d��ۙ������}te>S�����6��� ��X�����*k �ꋪ*�n�%��Xhi�tg_���vp�����Y;9�! �Ul�p��(Z��� �~a[�`���V� �ڜ�@dl�ߒ�?��l��k�/c�O��Z���p�4���/��K�0���bD�\��]T�-׌��W�N��{�pRR1V{��ؿ��2ޖ�Q�]���X�0��,Q���I����*�F��i�l����j��@U�Y��~��~�\�ż/�n�<�%�Q$+WMg���(^�鞈�}�w��\x�C�3@Xψ��/ &Y�_�J��� �7��XHj���iU�'��A��V��p�U�4�5iW�h���@*����6E��m������7%��c�n��n�UZɍ�ƫ��E��n�0�tT�Ҵob�R��붾ʲ'�j<4�yF0ų��2�z^5���
u2��*	4sU�������!ɁH��� �H�(vԡ}ʧ�[
2	##�ej�Mjai𤂋q_Wp�2a;y�RmU��Ns-�%��;W�Q���4�«E�zM��q0VO���&5�`�7Z���ᆦӕc9���nRyp�Ke��eUY�M�5K�t6�=60�%���m�D�Q,2�ȱ�s(���#zN����[*�~s��S"�K�O_?O��dc5���s�������2�Z��'6۴�U�\���K��"H۶�/¸�]=@����Bd1�Xn�eZ�v�K�u��H�o��M�
W�U���ŀ����:��0�UI~��I��H�B�%�xDC��m�� ��4��J/?�V{�H�W5��]���$jU�)�0��������9dG�N������Vq{�h
�^�kuy%������^�Ec�Lח/��O�+�Ê��:
��9
ZPs��Y~�ηl!Fs��N\odD`M��
���"�&N	кc��ht#Pr}Q����E0�+���;�#162�ĥ�g���)���FV1�t2�������M�\!Q��񲮿�_}���)�����5ʠ4�/�5(�қ*�Z9=���&}�u�I��\|̨���L�&�$�OƐ����҈�BB!�"�Г�&l�"��� $ב0���B���b�|�h��l]<���~esɯ]�����"k7'�T�G>1��
���ۆ5T�+�o��}���Q�@���gԢK�lq*	�ÇU�"��U#��\!�?��*S֣�f�
J�z|F��A�֎Q�!�Q_��d����f���4荎z^_/~�`������pK�!�O�F��bW
WX�^�6Sp/݋�����>T�M K p��R�[��{�5R�b��ym�m�\�«�zv�fIrO��	��1�\ g�-�����zu�J'(� �ł@���r�%I$\���	;w��"�Z�����G�z���%��^x��4�mXi��~�fi6��lz~+/�-(�w��9F���=;�OE�&���Ak��vo�]n8�Bd�7�p���r5�0�<%iq�mɌ/�c��
-�ak�aU�W�g]W@��"f%�&�8�H���|�8n���ך�Cg���-
�HKy]�GB�Qγ�����Ɖ+�Zp�+Ӑ&�J���#���h�d��7nWD-��-���K�G��tP�!���u9(,t~�o��m��A��}��O	8/iL�>T|{h�S��Ur\��(ˢ��Mw��s�UO�g��D��w�s��m%�c7VHjD|0��3?��칭�Ɓ+J�������?_�G�*��Lh�r�Dy1���/G����T΍�����@�����m�/�M�<�T����L<u1�Al"7�#��ov�sK�+�<�s����v5̕�΍���]q��:O��l�)=S��U5@o4����C����̓����N,�T`��k,�(��^� C��qg/�`�)]jD
�%�[هt�����0��l�.�H�2�0�QV2V��`������-_X�ߝ'cg�>^���"9�g�}Be3�R�g�.�?�3��`���_�
[�|���-3���d��j�L��A�}"�?�C�m"W-Nw�}=�bP�xO+�L��/sӢ�z���p$��6�E���J��}��$�N^��5qs��t'��UP� -��-��&�-EyL99\"(���]�H��m��ϢUWI��=�ft�p�"���{� ������M�*��4��&@�%�S&��ڝ(��5���w��q�44|4k��2���dm�͹jG�}Ϋx�S�.J�s"�����w�(!���&v�n�|�g�H�ok��r.o�N�a-�̽0��(��U�)�i8v�������VT�+11h凙�}�M�
�j��㽍tI�b�$�#��	"�H�$
]e3-��4h��6r�:����J��5��&��"�����n�T�/٧n�#<4������$>�6)�l���ͥ���Ȫܓn�N�}�R��=B�]n���J��_�8��ǂϣa���u�=�اOw�����¢'��%���
��ؖ�ƴ�mH��#wQ_�fi��:�'��e}�I5տT�J�hQ�����;$g���Nf֯�7�`�6�B��Jz�T�9��JU��C�r������M}��Y��L��q~��f*G��5���+ G��h�
��<�y6�$�al�CW�e<D7%ё���N���θ_ÏQ�M���M�,?����6.�J{�b?g#��g��f��%AzM1d^�o����bC��+�m2��VB�S�����f�����#�!����C�ulYBƜ��,Nu9;E��݋�
]��3.7�*��\���h�l6C�:�;��;;]N5u�+�l���`>�HA�NQ1�J$V��g"{���:�IS/H�3���j�<�I��S�OY��?&���1�v
�e�j��6Q�{��W�Ϧ?��k^ȷ��5i�����wEM����}PC)�n@�6!iL��Q��4��ĵ����F0b�Z���Ih�_��s;