-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
UwJ2dTgLGw5d+sv8LGg4T+rsIyksYVLNyAgpbWb6mnpAjf01dUX2aYnKgQGGPdVi
psPLRk7TZkFnlAbnO+DN9BQzcHnMi+fMSFRwY9Ml0aRXbJbpKCA9UNLbYhx6DeV6
5PlfNmmI5XvtTHBepk/DnvkdUDbp4eSfYsugE/QGuGI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1650)

`protect DATA_BLOCK
5U3sUS0p7H+lmc0ga+Z+m8umPiMg2nBkXqDzaFBob5LRdIgvmvNkkpv9+W8IbJvb
aSputgdjF2k6vQnlTmMju1KkbcDF//tibhVVqWuBZCK9LdyJ3+5C0DeyNS44q2tv
ocsATnZhzME3nQPloTU4hIEs7pe3m2tIufdiyG00xTw0bwQZPRYeV0UklS+CAUli
ufvbIYmkmMnvNiOi6uNLEAxgupfTG1Q2WGO/ChVX6qY/iT+AD9sY4zu4y7V7Mpwt
2L0ydridR5dq7Rk7qFr6Y1c9QzFIEbV1SpMIvYN2XmXjCSpiau7P9RL+ZcBxnsSs
fMIIWIJxP2N+mkEnHCZgDd+Rv9JcD/mWMLaWqmNlBbL/ms/UJlxCGpnrQbbZfIXN
ZtiHofxk0Qeupx/YnRROPtrKDAmLtq3aRCmPje/IihRyMFRccmizMJx6rYWSDD4o
+1bG1EDYO/bFzxY8vkN+P4s0F2ql5HopxlhEYBGGw+KbB2gcDPLonlulhLN4ATUC
SgEXQME0vm4phNBsXVn/+G4kbCpGqCyf8IweCPAwJpU3olxdy4lcNVcRWzC93MsO
B/oj7F68VAKX3VJ/Fsb78tOdobMpmh0r8fah+P3jTeCTDlp/9vpeiAC7+2bVJ08Z
3rh+w5251pMaqaWMFjg1oohpJKfKfaevSq7nNeSag743lv9Yv2YLRu8zZqKHxWV+
sy43Cf/5jDwrx1o3cIi2Yli1zUivbK5er5dH1WwKMjT+kc2TOjA4L3jZhpgpqYni
/JU/5GBxm7qYWD1aDwm0fY/83IxaH7ccUi7ajDqnVSIlbOHEyGqJnv5oPx6T/Wkc
me4/x29OBAEKTIasZOhbUa7lu6ymCiyEWD1/V43HOstxV7mRJ676LGD4DQgG8gkl
A0VJ9bxk2qK2179UA/qtnq3Tlm3qvKvrXRVXcLu/FHgwf3v8P8COvTxRZUQgOrVZ
3dSFuzIaxw84Dqt49V012bVpj9oOg59kcwEUEjMYPqrXJEoTAF1RibgwCQcQ13gW
EeO2ZTqLbov409xtXKQAG/xk49lwPwCSUn2pc3sdoUh9Sg4t5fUO8DBpWoOfk/I1
KeJ2jDhsMowhPkkwejXNe9Dj78Qv2aEACYzHX1jUEQd42XgDlUa3V3lTyHsneHgn
0iPeyMV5W9jVPdGWaUqy52SwFKVspRhnBw7hOiqaXGj2ry/D2v+YzTTnX8JWFtp5
VDJ0FN+d1kgOr3266L5mszJu3e7y+8431YOvYO8mmXR1h79FIPhjlEaJYZsiu8ZH
mRrhjsOhkHJb9tZgQlH7gDncp+DWI0hNjXXyCawjTsJ1nkWC7r1lw0mDznRfPa1+
l4XWKept8rrnsYwgVmEFT+pjPKo0qq2VszAWYgkDteRxgKZSFpAqA5wGJkNK/B1I
tvwHJ6+P9tVnvbKMVh/PYvk9qJm1HYJZrALUWaq8i67btENtZ0bcKm1dGQ/q6yK3
meWqT2mB5Y7cuA2qTCyxb5/8w7opb97a6/VPjNsVKtZ9E/F4//HG1cFmWh8lH+7P
TlqWWLK4HoEDTtdsSYncuyER3tkgfo7GwDY+HMIafp9yLhGj4EKO54HKYPS6Y4Ag
AFEz6k3oidKtY9C94IISAKAv+kcKweHmYshmWbBrFgU4ODCOmzSYkkXmDcy62m7r
jKEpJAZabV7Kf/TycULaTS8H64b5E78YN58KkmhQBoq8HCw2Ttpn3X8pyyi91TR5
4y0puuvBsfvSmDF6g4SGoY1PR6tx3zSSdPUIWn5Z/zt7+zdPHArbw/AjWuzLY1gE
xUmna4j41p5thHzcNUYC99jdBCEnH7SZ8QrIUvOBsW59jTrpheFD2R55DdkEPoX+
eVDYDG29a2DoQ9ludcG0454wuMnE+CZD7EfCldhkxxF/WIxB0oOd2pDjR2epHJfg
UQO7OBN51+5KjFVMPby6KBSCvi5AuJXhEISEMWf3nOZTTyuyp43rzPV8iy8USsZM
zaQltnFaeEr7awnzD0apL1wDClhyr0aFQGss4W9KPGKosI6CLnFv3esvu1YSsxeT
gMJTHyVN2vJptq/iYdjiJrwWpu7mg4A1qslZVjmXh272kz62M46G4JgumhnnVE/2
sja+H1v7p3EY3JsIxtu+sjC2NWeSAtNdUByCz0EwfxL5nHO7mhNbXg/ebdwh/au2
uybOBEogWKY6C7SwRHYQBKRnPeC2rMt24cQuinBAVyZ4Lnw5KDaGLMwcz7EgKK90
`protect END_PROTECTED