-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
iNOF5nLHL7feIZDpQDO8ve7FMLczLleG7+6Dau9GyLt2KG/8xM5hEbhXe2V6caAm
1nVDgqZZ4AXqqSdQsAGTlj3+xWRm6cIZJsWk1txtI89UpugOw4PA2Xl8M8Xy/y8i
MjYLncqbV41nmoCbctWMZlxpEADi6Cp/B9YCvbpsRoE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 23392)
`protect data_block
hAKTdr8dIEhphXVAO6qO9PkLeBeJcadxMUJy37uM9NIp6W2erTCH55n+TY6DHhOC
l0wHF+N0uO/GXFf+YesrNValTMwL/RUkNiM1KVV+HBp/QC0A2IGPUo5JTdPP8Kl5
Jp/u+mW2fC1YFvqL7qSFetnQYlo8MEc6CMHA4CMGx3h0xhLXOEapiVWUYjSrycIz
MmHMpUioljJ3YWn2gmB1AF9CznwOaBqMG+lkc+xuIlLL9jWUH6jXMmoDJ4ZSZGvD
WYNMi/LWFpTD7CP7bujJ+mtzX/BncngPgoWtP6GOSy3oPYL1My90XMS7RUUTtXQE
RE76KyNQ/t5bCpaSFZHLQbLHJo052TdIpu7ESRlOJoYSAgxYHwzxyeIWyPmLhTxD
kog7Vh/nfPn4S75Urm8FCnTsYCNf+pISXZuSeRHX5/9SNvPhwirp/aJy75vNTUAe
vsm/GFduq/jx8fiw4v4YJm17aJPtFDVjne2e8N1cSWGyewtnrRNODh1Iny8ZxmLf
xOnMRUQKxV9qL3yyKnIUdQjrrkma+OnlmGipZ34ueBe+63yH4UdZNyEmBqim/Acu
7KTLG4HfMUFMt581sGQgjaIZLPa1r5uPSQBMd3uUTGl7/Sw5Nu8gLtRx52PtvltI
OhTwgnJhLP0oRmMsDaMwHcwJw3xvTN3J6UvrAWNVdyqic5x+cEGgiOfAUdUkYjrV
85gqDXa6kvybMadaN0fjnnWcZh15yTAdkX5f9YXST/PJsFOafaGNwJo3mUjeAkAl
FVQXNK7BD8iMmdEwH4sOq+BwRsZCEti2zP32F1xqci+awUBE2pVrHo2V7LUNawCV
l74yTWDbBCZWpH37U5tJNJB3gQiECiKrlMormL/mByBevysWG5wrtdzMMxv0pCt5
+vlnq+nsp+LcIBMxnmD7isxpJCcqIhO7Zvr9p5mqwNx+SYhVL79BEn7K80sI25CL
74Gldx1TtedMlXYyZ9WjXVtg6ppVTFC08jEZhI1SaZy4bVY+OIO9EBC4IlR9Jj16
j8Lg5iQldhLaW43bJEGyNLh8Zp5n7DxQChmvYrIxnPR5QFJ7mCZgVB/UWMjp0/wm
3PZpd5TLoQ4MV6BOCXCzlBB1x8edaGdMm3H2Sh8mwsWHa43yiTT6PkYnqsp0EzI3
NIChddBdABrLUMJrtdJt91UsfAb74rJsXXBGfhoQPkLJbOqyaTHzntZjo/HL9dKO
/ZM6i2R5r17cI7km2/m+9LN6OU3K/X75KM4lCyhqyILnSgS9Mr5Gm/azSMW5uXdO
HZbCLIsOnx0xZkRiQSC5SrAPCmqhfbnBGdXNXWRERkszvVVps0+XuV0b/njiZd+Y
BB6DWYZ2POI5eNLGUwtSzPUzGzgdI8o5WLdjuKoW8/oA17Kcf2ClsYjZzFNFUNDw
vuj1+Y0WWtEasNeONHiCUgzoVgfrFyE3r/JLb5zLHxGa9ZxJs0zMSYSzieL8PXmo
SfuTZzlrSHTtxZdYaUgmr94a4d8CmvasCh2sZkXhO8tOLAcq3ZUtzduhJksN/yMq
01mqYN4qXMCHlorbDsGxpSZNZaMnIFQvv6G03Zqy2N6vzVPuO0PepukOhPO+OHFI
6A0xVsXEcaj9MNue3XGqZpJyRhW3dl58WzW/xStWdoUVxCSbslijAgT6u4WPmT7f
xoKZidTr4szJTrduy0cGSBCg9npbdDIYn3xu/YEk5gpPtJjatVKBsD6NqN4oSSxC
smQoqCVMVY2oXW6kCzBxKQhB9eC9qgjjWqC527S3b2r5tyFCDqTwjs9HmBjWKVVZ
xMjk4BqhRJeMBgYk2Ks0rZaKhKbXY1JaWNhnU/IATi9PvZoWk1Au67SBGsHb2kwu
zQ11xqi+uHmGNtDOLJJaGI/F2s+FZU+KG6Rj7s+vzCf7vEOj0e43TIVLDsztaHb7
c//jvONWy/3p8HCJyOXfmnzd8bWoyGVMzDzi3dFb8/ddiiiOIr2OeSm6BgnldKFu
ljj3pTZoxxoBpqZsyl2uL+pOsTOJnKEokYX3i0D5oxXTW8BLfp/mlNV/gtJ4+pF2
7/aOT1/KOmYs5J+Lu3TvnuGHbulTgP+2E5ifRFQS0l943JKIWFeAa5D05kp+lAIW
ARgqVrYu/VXQYiy7LsG6UNWSy6sewZmEtr1nb0b3pVM5XsU7Y6kgC9Ygqe4WgqEO
0KxQtblvlgU1ELmbnx8WFvDSKRu/rie4RI21yz5MQoctueiyE5Xh2tCDUcd5zeoX
M5EwdylxDx6Rk4g6r5n5ANMx3ng/mL0HFZXs+mqAcnktEB0EbOiWCkzwFmwbjUn5
Tg33LaaxSFfB7ZATPKQgbDJoOoKMo2BbZmL4KFVjE/Z9E7nw1qLkw5yTGQZdJKmm
l3/pi2WM926TWgl4yaaGpzguV7EttP0z8CaBhd06HBtI2y8uxZ2glmHEU/xRFrQG
45VXRZG931y6huEwD/2p6muyO0AhIEQzuc13hc06ZQNe8J8RDhidF3BcEytFOSlU
1omy7HcqgmUqMyQ68PlkLDgTHGkP28kLbzxsDUeUXx/S6Ff6HCnkzin3rNwWOsXl
xhjELmRxMQkqqnKfVkv3awrn05Q4yfHLdiJthK7txXZAN4QFb+qIID9hJhcTQOzu
Jo/RV9ZZkEOaei7/OfsreSGHr8SAWusWCz9mouHLu02UbpwbNx/MWLt1iIBgDLRm
8UuD0Nxo8MEMTX73YzqSqG5MeiVtbNbldwdK4tiYYPaKWLz6q9dKXlOs3BoE0Yuj
p4PgY6rft5OVe5n//vkMQ5Lur6Nt0tMt55MZ99uCAy+L1WdsJWd8yVLcFSpWCjmE
/tW+GUH2MSL33TsBTTkxuxutJCfWJDIl9oVzjJvvCHOJyeTj2N0IUpcWyLTnpzsN
0gO0u3MhPjEQ/cEWNDXBG414Brhmgo6p2O5j9+AAVQpzMhvXNs3Ov8uHT9t1dUq2
BwTsf9icTC6L1TpPc+jALYtWRFHnQTpLOG3zzr4ztl3p+Hs3Xq//rPyoOJLRurp9
U6a39x3pK8ZcJic2uFzJi/gNRYv4C6Iu7gZdBOwIGHBI97DHrRTZ27SkV7W0EBMR
79VBw72v4IXUNAQFGyJmAcNSSkqDghQ0XgvQleHogS/XvBdaKCFVlXA43Om4QhhN
qVRMTvjIrNM/rBhHigZ83Bm1PnPvZe1rRtlUwIKfjYWV4QQqqjAYSNAKskz4CKts
M/JoQmqVKemorXnYqqrEkeCaPtAAWH7Dxucmnh7RAx9DtB95BrmCxllChz5toOaa
o3WWk1KH9WiPXqvwbhHgFVs48lbWYH0S6euKk6qveYGwGcWO9w0K2c7r5C9d+hn8
qFIEXyiAP/Kvo2ky1u9e5owNxHTsLS4D3SmfDlZpklu6i/lKHmYeDy4g5GRamaIM
uNpB77YCNZovA+mXLvrtGkZSo0WfRvN4pgZfL67dxzNYR9AKIGjDxIZKV4bAeRME
o1kVXqOut4ud9mfVf3tugnPIwcJwLpTdj6iCAfwH7uzRbGI0ahpwM7she0nQch21
d5IattAGk2PzEGnTo9RNNehtK2GMpskM8INjLlWA7CAKNABn3ZDmKeBfDz48amcO
zPcLNcrVDEVvWKHsKu972DORibiX6HpR/PEfGH31kqahzCE/W7p3jNWy+tFPBH/f
49ylPaamqVucyOapK1K7m3As8Q8XMNUpHIRYn8fz2b6AqFhgLcrR9UkhzxPMBES2
0uHAlRVbWftlPMO5/cCDdzUuqnwn32UzlpfAAaOavTqyiYq/G5aObVnO9lBWezW0
fJORpsFHsGurSHnMY6gd6MMu/28/4JwRImlOAlf7kLJXEBYyycJOah+WzK8LFAGH
fSEE06q4vQeFW1uYVOr5cx28FFxVSej1qebBDx3Aqfhii7ySaJM7gTUHwcaSTpJv
sj512Tswv4dxs9xSx2QG1O/tUe4B6xkLomKBISq/XuOeazrntF4ZSJO2OfnqRSGY
ZWKN58eYTkALAt5+VnSBLuT11kOe6IO3KGAwCUmR5K2yXrUDCGNj0OEgxdPeXUIk
O6MtqLolh6XsQkt/1lEdGlTNXOyMmKXk9Pbgc6TUrZvEjo7or1p1F7/5w9JYdjhS
rAoKcRy2w0ec0FObGgQiHDioN7e9gHoowdhYBvXi6+ljpyuxswel6xZI8hVp1lm8
S75lxhRK09cQMsq+4bd11k08JRXgsz7D+f3LGsVzOFl0bBiEfjnCUacIgmvelYqH
xwj7gajBD5QlCXn3qoP2HPLZpJk6ECHpGB2B5/9FM8Ah4P4GcnvnGix9mEZGVbae
DxnK7vcw2gCfJwyFElShIXJ4/y37uiwa8O4s9AoMkhjihIyrF0C3Q6Yu90tydjpe
8fFr3dLIpCdlQyl6UFwhHXm57s4vXJFYVtkfddu0gLmxtIHj8cRsmKapUbMJU6wk
fzjbxn2KjfVRP6cqVlDt30lmtYxRGt5IakRG/Ul85rvfQx09A5ygxenz7EKOnyvt
mWU2tYfilRB10NGsDjbiYT5Pt6DVZZwLUF+02c2g/9vscGKsvlpk9KeTKDpAqoxc
HxrDhFTWpYQbE1JHRUhXWlESNO7Bx35Ge26Q+9V8k2oTxeod4mQsuex1KOF7f3ic
pydO9rYI+JT6cBHI7vX2Chqdt4vajm5NrkHLCXqZviho++8mjrUVDOfnbvIjVqzt
twU/JYICcuda+AzTGoXPZlSgWDrou4I5WEhAOe2Xhuv+8+2IhO2HTJEthsnz3uJO
RJ7FGH2U3L0sekcodoliQ8uytTiQi9erz0DNy9MlJtHFmFz3UQerZNR2QAqoI81B
GeipU/zST6NiQaKVYLmtB3txt/pAvcnyXh1rlMPZ6ZjoK/7t4/95bwq1tYca54dT
4U06tbpSExON3bvQlNkH8d5dK47t9h02PI06T2GhbDfK4p97o9LV5Z3KMtrMTC9j
sB6x0cC1E3khIYWlEOxTqH95Mbs0MnN/UDTcVpZW+QK+LY/8nzX93CoBhl+7AbCW
C0mY8T5McPNq5MRIAIt/OpW/XNnq3vatAVAftQ/1SNBeeuByvnm81MXzlJz3ZMHu
7PAHcAURxjEbOsgmUsurJdlPHUXegrNt/iJ8UZMiHbOsqueGTn7pr6Fi1wwjECkJ
Aax+PZSl9G9hsJAxHBJmTjZijMsdCVLr9LrTVx2VD3Nf/I0E4XKoh1c0M6fhD4Hs
vZhoUkCfXzHUXRW/U9EARh/7UV2cqTorzpS33FpMpQu6yiqkk4aHxDxcgojvsjOs
GM6DMq4tZDZLjBQAj6RGJFYw4oj/XXhq//o58pdPcnGqq2OcrZoTsgA3a4WUPnaF
rSsSChVLsjm5Vnu7Pz8oRnBueYanvjmQTf+W4KqO9hK15nuabC+lN2Zx3+eM3xTH
kYP+yDy7Ksx87dDRJNR1811tKjpDDUCkY8VSm8qbaRcmNhjNDy493JmvRzzgQoHu
Vs77Q7w0jMYQf7OiBDczdzTTUklNGL8Q52r/+kjJ6BIuo4gn6SZA6T8C1TIHa7jo
yxnWp78E3XRa9nz2+KIYiCT2sXwn9YoLhVy6l3mxFpXSnOBofYDD7dcl/Wp3GJCR
4ujPJrLNHwVQOvs3klRhbuwHG0nmsR+FqxHrcZXVfFplwjzONl/544naXu3qNm2J
TH/SxEAeRTy9cAppTOdzm/l2gPqHFXDDSiY7mv2yqWTgK6sEeVb0h9EPULXxbXuK
YsvUvrL0Kc28cj6y1D5yeiQJckPMx0TBq6QEiAQdVzasOXtuG7uKDzLJTV27tSDe
sCNBmoCKQ/ufHlNTvYWEkyKQHyFcWPhdWJUu5M+7ibuYBgr4goJTk0tB3dkqkixZ
n9DEePnZVn2dGmP5TPf7IxGfjzp7zX6nceS29oA7+9RvHp+kqeN8sPtpYvXStc0N
pw7RxH4lAmGTuzgZc5q4DNZoW7Tu6NWU0zkx8ScVFFu0Ooz/uVlIBYA7tauZBspW
zi4XXCyupW2Q43D5wV+KD/LnK8LjUo2KheQl898kvTMdqDfo/5EWIGi7VGLNILr9
16rFUwqJ0P+4IeG4V+GulqfPv4+7IWgdlro9u0+A7t87/FIfe5q8Dot1HuoEYk81
5o3GYqwWnLPsCV8ogmL4L+gA81HE8y3j4165vjKTKEExQWTbBpH+X0lhrvuNpxth
qvHLEH5HHOz41QcgqiimEXMKgYHr+RxI//VPzRJ67DvxZtdKnEG5rteIsE7gjhUP
yBNBDJy21It+mdjUcICSJhnGobcQhlhZomXHNGfFDS0zjsqp5/F9Zz7SsRvJKhB6
XOCueWEiFtuKYzLbwTi76fHOyGMfLotHa8QunqEPgBCoED3l3UaYlExLMNbhY3Nn
hIW+g/Q0ZOvmXHYo2oEQsxt9WBCBFFnSKYprVo2qUtprq5PTu1J/2Cy9KKuHOEnL
jwAwdPvKviiV3pZ2g4nlouI2vDpGkva7xdYlv1D/962rKp5+3lBxWdkZPDM8cgSC
+VkrkENxsj+ypMX5rs4jIaN0ZBJdjrnc4dzyoDfZ5S7QrLYnM9SQjzeV1JizlfxC
ZuEUHS+8W2OlmkUeXy2faQNME01Q2RQfb3mfOrkdTfS/SJoacCBlTowVfTMT1z+7
9R2fpelHeAJml62hx8e06eKHHgbetfsApR7L4VGyDxCZ2SUcGC3Vk8Le1ySRDhBV
YhgDXcpyb83+gGJNuHtqQkW8Cn8qYX+gGG31KuiW9BoHG6/lUXA5j6hmkJHv9AIm
WWuCwUSwd9nAKwBnJdSaaImugoN4w0N1ZxOzb3x8TRJiP/h2ZZbqudaV8pjYfNNX
RKkXIh3HJSe1v99uWfjQ0lRDHnbUtQhnmEsgskvfGcv4DzQqQbniBEpX7V3qech4
/KjGg88wOmQvJ9lo0X/X/dPdpUOdUdAWCZNExNOGfbJAC+Cd00pWK4xS4T+RfIi9
CJDBlP7aINhPbOL9Fe3c9z/ctDtwU5IVFyhxbBF2B/itZSRo5tlmqRkjtvYVUjnV
8tvPV7Ngv/YkTAVYf43sxKvcSjpR7nHsHnoEqD6M2MtrS6vyURySEyJCwktPSPQG
9xmzriZ8IgUatRcRRCTBt2t2GUTh+oJNfjyMvQKnjaJLsBMQXKEKvXbUNcBxSjxz
uryqO61PKcj2IHHJ6QQ5n0ob86f8Dbx9KL/mXsfF3qDz+EZoLPEaYIXNIeFi8QP6
fLzC0198CNwyRhbz/sNc1gJT+1bVE5Cfp3JlO54KwSAw/u/WVq1nRDSPYHscFATM
cNv4MuHgYM4jaI6D5ysrBJxvSLBi/9QMprc+NTDGZNoA/9VnudWjS70koEtkrr/e
BH8ubhZd1IT1OcnLVZwDCcLPRVLPeMpeN22pb5i+qfUw1Kxuz6XJF3+8626vTh4O
PrpA0S/hTv9KNYsKKybfjeo9FQsJCGH86wJODsAvE12kTql2qsxVFc0EiKhhte5d
msFE6ZE+W4uA8DsT4gFWdR0fQgXsGmaeTpdYdFmFpvMkwG5clInQz5PXVqaxBsgB
VgfXyuSxgfHtTyxEkpMCyTUyGz59xv/vyP/uc1a7yZ00AMFEt3eM2n43CJA4tRNi
unqttNaBUmtFHmvyHgxx2aommVesyIZA/EgV4T4Je7I94+QQbdPofJcA+bU4L8Zv
cLHhPsT64VhAK9mZ+r6tRuBZLuqSJ5qkcdpQ5PM/T7I9G9pWDUZT/n5y8kZw0A9Z
/F/2ack/Se9cvM+N7x7VKiCY9/pcMI4fQg1tBqRI4leYZ8GTr7Oui+ajZ5mNQrRa
o8jqVH7kiB/wG1qFQZZlfw7srz64bnxfts7Gk9EOWKyjnjpnI55yIG33pJKBXDtB
LuEpijmWpS5epaC2DFEgXhsT70VBafv/4n0Xv9/lhdboLDuaOBjF/ai1L39DgcMY
TPC8CGjoszbcPi5Cme1nzrmQPUtEgIoLK8YYMuVLeQoT1KM+T1jUgOlht934UFo2
SLEmAbEVIs6zJG6TWA264lySs+/E86U0/H/dJo7om6gxZ2hFQ+5aZQrz6jogmA3n
1v7UPXkeu44064cBwWr+fH1m/6pc8xAP4E2Zc90mxm9igX/fecLOpjM9y6aTUwWV
Z9vvKnybUnx3iosUFwEf6v48A/j6Ds9woO5nwTtMlMG5nycD+uWIVszLktxSyHSU
ZcBMk4k4Is6CXiWLr71CbOSBfRosn6k5Dd/PD6XTOaJh77OjS+9fn13pGu4d1URC
4mveNyQS+QIKFdTLjNVLL8eXMe7BkVDSAfHgTSYUNMTXRQfXcMg18ONMKUr85RED
tYQYNgey19xgMTHSszRLwYygZPlQJV/YRoS/RZjU2B3UWvmZCuRnCEEOEGLcjTYL
vtRBZilnqF/DHum++8UaUOlDwyZGTInGz+a6akwG1KEwDX5NzlbbG7lO3FUYR1sF
JBX4eIe7732ve+ZhZha00iEczZbMTvFFbJ05MP5gI5lwwVVJ9jW5EpTfwO+neb9q
R6Jc5YIoZqBLHlDC2RWCpyLSItESHDt/N58vGwy7W/d3R1hf01u393o9izJFi6sA
LmzeaBefLq5wlFP6SUipZLGeNmJryf8DJFi2sNQp9mmDvcem2O9q2ojwyEr6m5Qc
5C+3extG0qYWrOvM7dUWBH02ciIzdMMtSNqoXMzo/tsVeucOVfnJCVP+uSu/1QrM
zQUHHAvZMr4aBzWYmnmlDfx98jnuYYJWwIaJl0ps8pwnbydzNDfSnZJYnYbM3aEB
F6NE9rT5guMMzSwbKi2mhfoQb3+gL3cuLd9CpWlmtgK1NowaRwvKfDvGBo2N0KRT
zAHfNbWqhIwi/9OwrjSr2r3a2+Lm9cBBqbpdA/r4z6uNZ3etiUIDTGfLg5mz9HQQ
FXBDCBb3hZds0EDUni6+ejd0SuhQ/ckmJ8TJNdRoM/w/3zMYhr4nTvE+Ecyq/WZv
Rka6ZRWH1p30hTAyViQuJiQ8904H4nUwktUtkBiYBKfOpJc+jSb+kBC0cPCrIEJF
bPpXkyLWPK1l3X7OiWjBjEddq1E56+1FpuBWN4RfLlUbyM8hKT9z2OVcD1dHoRXR
zE3sq0U1lbeIBOTti4xVR0fQpDCdmWJDxvA95OTAfOeAx577ivWC0a1Km4FAHwul
dv38CCUUG5qQmhp7AVWPeP3Ko7agGopkWDU0a3A50osE6rFVkWQCpEwy6vNgXZVg
B5+DJtFgcR/GQIjQVXFPWqN3Dv5J5LQdAFh+ps6FoN88UtuffWv99WMf9+9kebOL
Od+DPYsjRqbQmnbC0nvzjDOGnnxlXtwWmb7tT3NyIuXPJMv4pUgLfwQgwBijW+a2
CsktJIw42Zpzy0CmdcOzEA74Ks94zqvb11FoBLOJZii0cizCwtFGv1gy2g5gFofi
R5+W91Xne4NDLWkqXYs5EAcIZGGSCfkJKj6cMg8C577IIm8sC+7AdI90Lcny7CN0
FCbIQRkL7CHMNoJ5dfKWbgT2i3Zx6godJJoTsSpxLkUaC0h+HbbbptcZBskhsB2T
gi3v8+nYK1OQbnZ/j/UCSOwjXCBBXtgh32Tf98BFi0uzPTO/6DGpJP0juEq4jrFo
JPr3gEbCIf8VDE/+1p1nD7nyFpsNXTysjZCTDEm/xITnQVAciRF9te4cIpV3jqqF
/kBkXK61KrEEDpUQ4Ze7TdMAMISGX6PIGu/I2vfo89ITEXpA1D0dDHg/YNzoTECs
hxclC9THrx4SC4ikCI25WgKduVUF34mTTFU7ZLpV6z8jJ4ScaOmsW5TAMLVdotWo
a1y6WsC606JAM1Y/thxqBIvtbcqRcoUUWw6jZ9NllPBJu/7HcQK3/wR/+0UxP4IE
oECXUeThRj7Ix7vXQll81zzetxCKls0PbzN4CY20J1d0QGT0F8/uTEXnPahFT5+P
hq9x1mb2xPk19hPv9146Y4IgSGjbhSq1q9bCtVEOSVKkFQmkOSf+Qv18r2h3V56I
pFdhUqmgqGoEpAqBhCG6zLUqyrXoPA3IxyTKOFaOXRVysf2bilqBzoZ4BmXZ5kQ1
ttqbjmvtS4eHHPQvn3DtCG4NdvvcR3fGdauQhwSsXPATTXVAX04J4AyC02sV30qr
cZp2a/8W1MIWnJUKqx1vvIAofcTfI1rVKda/LbjcJy3gRG7qdPEhblBYSHEQ90/G
A2HKOxKOXQYqAuhFwXjf8mEqdgxUcqCqNU4dJqqXN3uCgfNZ566VMmouFxBwqcLZ
7hjBLVPML7MNLns/u1UMdBoXADVGQ7ryMPZ8nmefPzGLDgoRU9uqAWmFzsihQcmS
XcNkXrwTfGeVXGZ/KL8ygt0WJaTo4bny7yYms+ETdbkFVgYT51h77eBW1R+1oDlR
GPzTRW9cgBNhGrIPjc2F3uCE0RQqUn7re6uRpsbZ6zdNTDHvcori87MGvVeNo4xX
ppMcBqiXrqhgPDZx/rZcVsPMSXgyeC6GefmzMlB8yS0SOEvHGgVuhxzUYoc8+5Fk
we/KTucBGydko23CPEpVD/Y35qbEZh/002ZUeQnsQPaj1MEg84MZ2ezbEXDXf7OE
7NXyx5BwFZ6YwWv8JmEbjIk78l9LEJaRsdQ+JAPLZlZAzNYMhHL2yENXASVYA2g1
hd1kvh3+e5NTmWdi/sfd1h+CxNk4UtkqhWhl8PxIN9/n6GjHOsVwKuyM1Vxk+aTY
hpWIorcJyUjdpThL5hLeqCGMHgCU6yj2hnEfHLNagr8/ifBIwXavDBucedpKtZe8
5uFSxMJZ3G0f8ISmY8qevQFtPKtMbKnrsB5cUvYsb4tP+FxieQ9FvPW9gQvGGoXE
wDaVbvjLCmR5Ce5dnOrwvZknRAyaPiVp9ha8gUtSYI36r8DZTv7W+0AZPzuAvvKy
WcZPikkyfRr9lnwwHXNvjnykos5NssC/1vdtV/E8Wm2C5qjzJyzqorkYg7zjDEtY
7oOCYNQgtqTyFWUayzr6ffuM71VLVF2MP3GoKczrFMb/Q0laHTGnXBIT5Ue7UyzL
nkocAmD3mxX/L8z3uV3cQ6F1iLOEru5Ophui5SHI0XsxuP8FM9Qw0ZSQvD2d81Cd
xvKyZQCfJiacfAZNAC4CJjVcSEphgQquGTTpBDmQSIpx+eeAi5UKJYy7m1VfhqWg
APkcEJrnReXjb2AxaHWKsckZxXJ8C/H54NUh5sNgWPJKJYRZaPQT5su8BIM5hevf
WIDSJMo8rKEHtaZ5fE790qwmULLZcmqL1lUln+fYALITfDaWHB8ya+LIJl1trpDI
mCz8vnnOxPvyTFLqmQgOHXozDvKvi6V5oXB12OhByQlBbDtcuQBhxy6w+t8OPIe5
AXpWeVOd64alLhSpw77b/9i7b8SUmW9oBTlw2ticKBQj505agzUCp/cB6gNf06v+
U7ysm9SKJP04TtBCs062jhz/bAS0hobl8GAozvZgUVhk68ranSXmfdabu+0vFRF6
48Ucfk9dhHGYahPA1muv5GUv9xbpgiDtnKuDWpfaW6+Nxd6nP99Z4XdPGTJXtI3Q
rRRhoUVcOeyXxCTDKXm/r3B1Lilv71kaw4ZgHAnu+y6XPRcwpxFeHReuSsGyoI+Y
PQ/XRjNQhlRSf8ag/QqPEB1IgjQ84tG3UCnyc2qzArTqzbThTbxw9joyxN03/qzE
LOKi1cuq/kHFXKWGs5Mx9uPOg6C32fkeJ2ie08MTi7O5ipgBpCYUcBD2mWc2qcV/
wHc5Imdw5Dc/v1u8xNxpDVAjG+TvgYJLL44Zg40QOkRT9q6cZb5B4kQhiQwaLhXW
67iodjKvM2Xye4K2/Wx8/orBZPx8kN+Vst16RHfOSQlQFAfycl3rafVBFIK1PpPY
1j0PhKYIeLyodWLrvD95KvC6AS6pXBTlW9pqFXJwt65piJTWA0x/FYT2fIbi0irB
0DC3xS1gkpcuidIGi2KgvZsQZwXAAjZhwb21nKVBHtPCvFcMqMZCUI3qrx+3RcDf
GQwheUjNCl5NZvZbg4cycK9JqHmUZGjD3r4L/buC/oOcmusrdHVzxiwTHiXz7IXi
Sp5S8pqoJ8O/4LMYDUh2U+0FbyV7VeZa9dsAXh0m6Y3Cw1jwbR5PSzdbCo9TFxh7
QBk9m3eWqp579QTGW7CnHoKdJtGpOxEfw30POQc82GMBjMox4fM03clAvv1tcpRq
rtK6cOziJi52xaHq6fevsJKgg/BqJYytdvbddHqiAmIeYOqKrNWLQKWMWOSgb0aU
+4TzAueEcMj0fhbJ3WxefOxiRCYbr7vh37QJTBt4lxxvg5TFuwEVpHOPFjuuAAHh
T/uv4cFlGEdbHJ/ASo7h5gcnwwligtRMvIVT9XXhiSh84IYejQwcseJms+2Q+GRE
2ZrxehPrP1nd+084Fnx3j+8fcv9IzKD0wpnMWke1xzbJLbkwsQS1x5eyfQ4PBQ5p
evRN9wjPpVessegZcq8bWaev/qrpOKKrjX+zQ/t69Jwbd6kfA8lxf6ons6F8Mnt7
CQWTTJjPm+b5l8ZYoR7M/JmmgLITjgXrNo6BpeGpaxMVRHhCiEO4LVHNsa5ewxE9
k8upGHNW3FB44PUHSI9YHSpAPqoIF27a6UtM1+j7XyHgI/D9WM8e6hI+BCtGPphB
3oTdj0qE/FoiFwLPyFi6Baas/qsEaG4Ts7Yy3F3zypZdfaTCKcMCEOEBNbONKNl9
BSBGsdt1wB5afBy+aucuW++Yl5nI3lbdQMrqbqSLHzzcrgTpnZcjKtOA2Vs3FLlR
BbrjwRlqb83mHMjAl0D7g+bnBVSHDYXTsc814ct90WvAVxdAVWYDTrG5E7BKN9t/
HaDz5bJWgCk0bizMZGyDfSS8Hiux4AqJJdNAo8H1/VSvPt+pbR1ft1UW4PlFrdpl
G1ffBNGm0XRZZtH+uZ6fOaPG31QwwFfsfOsmITU5tlL1zCrio9RFFVptTT5hgdJe
SVBXqJNtXkpBWhHdQNYyL2ZrWn4lg4xtNvDMBaX9uMY081G9wWUKDby1TESIkloR
3lYrGUCq6Nd9IRnrT4VLnID+mhIJGZaxYXVAq0eCL+lSKIy3p4SzWpmbBSJs93x1
Fcv0E/mmL14F7yMEZ6+V+k2+AMAuxOZZ1Vvcm5BE3F3aGg/dskQkCwN0RYNvm0CJ
wqZBR6HMF90V9s9w6CjvJfDhqiEl/1VqYf53H9j+4FI1v+CAbaYrq9kpHYUSPBoA
J1KeppOXPOL75RyeO/fkSJuTexdkAU6ipY3Qi03fg2wwCXoDh40LwsIaAXj9bF1j
ymKpveAgzRfUogT4ZmHoR/iUOd9WiunwZUAi+zQ4tuWJQeoXM7lbrZLEWl1HeBdL
UMR6daDTM/tYHsiTgRFtTHiMX95B5go4630hzG92EYqxKXutpLFkQDx5CraElooP
+JwLuBF+aLOWC5dFIRtnHe7XAt6HlmWtasjZr09JYGMZfcTx0hO+DMvShrph41Kn
HFjldT8NcU5wKPCwkdrnxEq8cR6hL6arGjHXOrzDU9QSY9oaUY+9hOZ73DXd1Itm
0VGA5KkFKNkQfH0gu9r78lBsAHtVELWrgcLrf51Sce4IAD9k+Uxc9rbDmyZYTCEX
Pogi+idUCYp7MLtFOt1HXIFSqoAY2snwtPYh8cfvxpd++h4F9zcAUDXAaZHSdCXQ
Vo6uIhkS/X3uWK/pNlNlItKZlGlb/q5txJBGs5KOwe5DxbCqltW7pOBRVc04VMdG
zKEwWEEV+qIXSRVTJq8RFnwQUWiGH2xBaYizwPs8bGhIAAHIzUxoUhXaZKnTspRU
YqYmJ77+N7mcYhzeSUbo3/IIlfDW1HueNHX8GQSh3WFwYJFB0hhtcltQ8XZWuHh4
GYbk9uK9ooeUGFuzOYe6EJ5qLMq2YsqKTiOMvxoP9ZAhfVfRFFu1uyvYL+J+vLny
QdXkdLIKogQzOoMgb2a725Jo5IzEAWDdOZDXDb2ynZAhFc0dJsy1VYu5qLRcbqRR
t0Pnmq027Ii/5ZNowXOKfgrBD3Zb0fJxAx303HjYf1aj5V76BKIvXgylsrZmHGl/
cPwquRBTrksqwsU9lhaYi4DABCKHkVKrZIOhhJgHOFQIyOy3Xc+qw+A6AYbG1RXq
V79Uu9rAdh6lGY04rd08lIxk+ZwT8AZ2/YOe3jUoo4ZSLNfe20N03G7COnojEhTV
stBoaRvAokLXG/JhKlPBD0iA6Ddtw+O2v+s/zPadaZmJwD7KvyJ6tKgQPFBKXblu
MTrKDISOhXTc94qUNm9AhkcliXH4N03T/YuSe8oRLoz7vQsfb8bPn4Gyh5M1oI/v
lkRXyHEs4ngvrcSanMwPie5UeFBGHWIggzZMW+AxzkViCahKMwIIFCkcOFGxQGGG
EEDeQicIkbSWx9qHJIYZfaGtE3wos89NB42XwnsaYJd3ZPm4zqD504muGczo9Izc
3JSIBO0lapgrddwp1D/qsW7UJXfAHdI9Nbam3/5R2tB/mlTFZtISDyABDqerkjs7
LifE+RFulgDIvullnDvxD6m9IJ+bv99EEKODadC/zYlt8cKhM2mKG0mr/vULW/8B
Uq8198MpsNm/XIlgUSsZwq7D2ebxFMcQTm3Kesz204FVnWDzQO1RWZ4gypsThCC3
8jKOYOnC1p4jZtYhck5OSOrcGnQEgx8SOJxVJ4gC54+Wacnj19BEHpdNS+FgITXc
rreWXBBqIQZp019pWGPi4TFn4WAsCVePPOwssdqBe7Xd5d/Bh9PT34eMMOxQ7oYd
6cQm3ZFDwx96EIkBqpVcLo5NcMwiT/KuyPdW0Tv4qEEpJCwT6539UdcJwII1eA/p
kcdVfkaFWiTm45GM7imK5dJGelt/A4L3e6on6Eu3/F2PdLCB/7msE7HYiuyBV2kU
U5pdWJBAlq7f6DYAnm3TqwK5A8QGK0G2VGCMHPUdX/VNIk24ZwcRUlz8EAdKUx5r
emN0G0brvQ7oPcYJNeNjVg+D/cY7/Aq1aShDkNzf6vv1B5CqbAx6Wzls0AqYx8R4
aZ3TAoMDI5O6w0p6Od2wlu2I0OIFghdThx4TnSefbSb0/U0d4/RBWfSxT0o0h/Lt
VcXJPFe91yVPJ9dLSM8xE+LYNhcUJLNjENDttSj6LBHTVPpRweao5DuRTi1+2Tii
qCS6rsBmeQiXUbiaK72s23v7o8ZFZqepof2u2bggflpv4eMX6kLIQ0VwEyGCSmuT
pUJeH1VEcd/xcvaOuLORUVDDfiiGSHLJ8WtGmbfSJcKL9x9MDZnZ4K/OECOOqg6g
PDq6+r9O58jTjDUQctK27031wj0uReKbNK5rVx/Vghbn9wkF/DfrnupCLM6eFE1U
OS4vUOke65ht1YCaGrlCd5rqyVU0lB6lkykbiqJhfaOLMGCmM1UKligeV6ha94KY
hYNUxl5qJKtyD0LjGyDde6izfQ8mODifyKCNOGRuc6vYNEkwuUrMxWfUgakTtj2R
kCA2z/dzDXY2TTYaZAZ9HXJrnSQWEKy0yeTVIKR4dzAxKR7micFdrP4xqTNCxcsU
r7rKnFDhthrUABQ82LN+t1KgzMUYS3sB9dFCy2f5VvMzLpajgVORuYaZnkkbTcUR
5IJptOGp+If37lc3pTe0fqMalwmOIwe6XF4+SrzyrsQq9GnxUkluerAuJAsNqrZf
NJl+XwQHjhpzhnZq+k2Z71FiU0JdJ9M07LmmOmZdHZaxo4nDK5RzkhL8mJYpjNmN
XGWYiuzvhQQWX8TLkiTT3/Va2LR5Y8mS14qXVABqBb91cvPDPThbvPOwe6dmvavr
3GWWm1FWCxSKbycBoQNkfNiT6nLuYLQOR5s56DPi7boPNx4sNtWQmz5aiqhOuYLw
7l++kUMDjsQ0moXzQxBY7b2QtcGCjB6QTvsNv8gMf5fYCTV/jBiPEmvh+DlFkhVr
CHLnaiQyTN1P9W0ItrC4uVM84UZJ+Wptci9EbSXZHecv3hd0MvzepjOSo3T4aG2y
0oMcx5lkdzY+fjP66L0YfsTfLuTmZ7rjf/4zVTOQCyO0pFZp3uW3yJe/BTRX2XE7
QxkMjO5/9v6J5W9HWpYllqONjh+EWf+q9Ma0tIQW05yTYmFQSq0xMP+fmSEp+yeY
1lFCCM7YBgqmAe88wkpkJFHY9IHn00EYYqOEhQcbyP0bGZBBv+ldbDnPbnIEXBbI
ABVU+J80eoWo+Q5PDdHCzAsKWZmq2+0uS/awhSO+dcVSExF4G7/jTPzeoCxGCIdc
AwfwHwPQvkIkCpJqw2So1TCCeU0DKFux9masH6w9Yy2OAlcfgI3bCKEKfoNd8LCS
SFM9BlpiUXcBV0/2sMUODvH5cMrN1pd10hW0UuxQA/bgS1BsD42ImUxlvBOGhT9j
PVbTFq4MZo1yXDPkrCbTOFu7eCa69wt2eSIJCOP1umBnHlqAwpyTYBEw3B+1xHe0
r2b+hHdPepTwoeOaLvukQY0EdhAg40+etuWAYuhXI/YQviVYG+EjrHPaIx7vdiMz
/xvdwSKH9FccjamSYUwqNRF7Zz5rz/gAVPoGtO2EJgynufTr82P7crLu+YqdxYn6
6zPiwF/rkPnQJ+jYPmWVXMqp6kzciMMy9Ko6++rhywKDOv2L1AZv1TAeHwwUZyRG
b7qmagpj+9SYR5HVLNvXhw9Ssi1eM5D/M8mvwlCYto+G7vlwuRZhbCdfwKjQCExg
pItabufGj7mkMqt5HbqTfecF6tIgQaz/hduh5ipZI22eJIV2M2A10YS2ANPBD+fo
kOujkpFEEIh0nf2ly8TpDWC+LJ8xMppjt5FzVyln/hHj+WxyLT/CYfTlWtpT4gI1
wL5MIkUUg26d0mDRE+rtpGvLX0GiHjSoGMhaIC+TWORsHqpakAi6yK5SbshD/edc
beXu5CgE+pWm/vOuTqe5BSzQSfhDML866RjIILF8B9Zw2HK1ihOiI8DY+5y+nbAR
k95qqe1PPiPRqGl2PCpADxc8/cu9pZC6Vob78pXM1lKsZat7YH43/TCAdJ7v5ugH
9TCcbEEyxGrwlY7ERt8H+Ybllu1en8G2t3Cytp+4bKA2EW1DoXwScnONQ588E9zV
1yvSyFsH9lBVlxfd6+oQEXz0KXdxrxNrprJ7xdEGVpLxrEBVzE6bUpafzw3Bgw1B
/L3/LHOK+ywnBabJzT3Zliej13V2uUfvZXZeF0y5+0yGdmikh4uI/rwdAwvlDjny
S5FOVhIiiWKuKsy6nqCvxL0jukU+R4z1Mo+JN6Q7PnuqdT109Y3CsM412HNMfn8G
+AU/xnwEJ41bAHdhwAfTQSJow//NiigoQqtmMz91Fla8UaHwldlVb6rv2Mjtzamm
W4Xs4c0SVOjid6k9GwPrPRueXRGqfFNyWCiP0kXHhr4e9k80eDC+dLxRZ2SAeo+s
3Y0kPsKseaJ3iOQtGMazEOv7eLaHCqfRiDTEvN4L1PrtKq8wK7Yr0YyESg/s+kQ+
ADiDFRwh5aWKOw3h0RjF6DDvs18ZLEHtmYcYYw7s6GDaizvK7G7jtL2fLmjZHzRx
4iKB9Ysf/Hg43NgS7+21mmIRnlOsO4Kcr6ii5Iane5CjPfKnm5EL6iLb7475RMH2
sUpUo2cB/d7lc34GiuIvujqolM5VQLdCDIGNPDyeYmnBwpoQVOP4HaEDm8+oXEr5
WGrUXDNbCLTkmkm7OrBAI8Z1Apv0326q0ndkHc6A+Y+C/x84misufkcz2l1GJWmO
ag68x5d8Lalx6PPFb7T+g3NUdllfqrGXROKAzkppkmAeUvuOLP7BQ1hFkV2Mn5+e
Ys3Ut/OOsWKK4FFQ5e4PTWoj6LoIUE5EYRQMqkfoeLQdrZM9ZzJDtIDso5fpjsA2
kg/+1egYXOQQbKWrGn2qnmAy2lJmxmYsJxMwf8iUetMGngUkCZACjc9QMyol2ysX
1fnJJtYeRtazOzLBjtXWJUTEvXsUH69DbGN8USoNg+KbIpydltsm6rMok8NfmZZ1
YEXp9YrTyHmcR497uVT+LEdaXptdb4tkJQ8n6DQXX1lAO3pYAuW7x7XpdDOp4t85
i/B0jDHwhERwJ7C9gvFbD9UMOIlStRXnw+2kcD7vlwq0ZCrIos5shEw+d6atLPxO
GsBnloXZ5s8Q3kNeD9UUly6gnx239LMZ/bEQOfo7yR7i2t7ppAz9bgWt5rsD6iDv
amKh3u/AdGQu5ikqQCuGpfNp2p9L7EaMKTQ6wymNfGwYzhhqOdyUWdI6gjI8xmqR
EsxpKbOqCI+2+YNWxLdgP4vVuGktqNeW8RM4TklyigBRfu8Ajo4JCkSclB4ucpmM
wkhTKBh2Ev82Zii5EiueZ1q8zu6/1wQI4kfFoRn+gOu5xqh9QKruFcVMr2Ms0Zb1
ZIr+ncZv40ef9hUz9zgcCpyObWiKV1vOa7zBM7Z2Pu8xNEty71fzugoMIB//pi+m
Luua5bq77S0guXZ+kYIgFjiStRW3dF6UYBJaOA3DbwmtPi4ib6TB8YXzJhMOJYC4
S4/DIPfgXnNaihZoXjLeXlL7yJk3Tj5HBE6jHUY8XeuGE0BcgcbzkbJuk2e/ywnr
WX9xl+FIMV1MC4aOuLvNtJxlLerWxlqHPpmi7i3UGetsrL7dxbCxPOJZD8dctXxT
tZqRi4ZdUj3RwS/TPLaS5jqe+nrKPDbujgz2jzR6L5RKC6wQhDnO9j/x5I6ZRzq/
EuhqX3vj1oJcKYsaqXh4cMGNqsSX82ZFYGbJDwz9QuwAUYG+IfYN36HhvsBq7Z37
RjNSKmzENidWqAB2Dn28Eb3Hs/9cVhAgkYtWVEXIk7CdPVgAOVJxPqt9v+g7UHgF
7INrV3NaZtx0Jx8YjfBKOlijhRx61Bg+FRkmCi21p4FNfC+XDt+Fb+MY1YBP4kBF
HVU5Zj4M3ySxxuaRYWRdwFNmmzRFAEaex9dlT078d9TrA5PPPnWlzdcCM0aEJiM3
WAB1hNcX7wsb/l+eF6wNFF1RIXQV8YlmnxbnbPWCu2Jp9sMSzFsb7ZY7VbfOcBa3
wpszKOCstAZeGbb6/PMk/RxfRkBv15+Eu8eq9qUyAa4YApC5uqoSwPgHZpwXaEa7
jYPQHtrpc9emQHPWPKJvWjmkNg/adAG86H2rvUPpj5zanObFlaks7WMgfq/XzNpZ
Mq2Tr4csGv9TVQunj5yiy7h4DZ6Pb1i1Rh4/V3PiQJkyWX3ea27Mt4MPB7WGKl65
h1BuqtuksAwekBV/aoAre4wJ96NpItq84kdew/CX3h7Fe5TTF56l1kE+GDLE5lm6
vktmLjB9oV0p8af023D/O0xAWWpvE9iQtKzIFYmIyMsKVjrRDaLjdA8l4kvgaEBg
qMvJVTmPlfjj9NRh+iIEOWdHtIAPaUduaqnxkxiYahxvbJwpvHm8I7/O3AtC+Iuz
CPWv+vZ0cv8dspnSlQje3mwRUOrO0QN0Qfyj+FZNMz5yYxYJkhIYUUFCqPS0IWdy
A0UpOCkFKhayLuROg+nKWC1HjlwbpM/WsY3LUWcmF7u1BWadp+5WvTDQQUdxF12c
4IY3MwRkLdaBJbq0CMgRFPq3LeJ7L0P3HbYen4FCUAt8lY49M11WaHwmsbTwAzqB
zYxz1IV0ufUcl1uYgpD2xifXLncIs0vJbOY6gf3EJ3Ad07zihW1G43JYIwdgOu5R
16/irR7Uz+rmmNj51mjSnPnWpVj5gq1lfGEZADjxGW4KJTNOlv2IyLwSua1usexN
GOv2dbGq3XGBMEhDmfleGa7wa7O/i4bvnIwwXGXW/ZglgubnYbIcTC1BWwFCo75/
iZFRsYPCwENS2hzO4T4iT7cj/frRaEN1pJy2/6+vpkQxaA5mbAI4NH3Y46GzE/6V
BDyAUbA/fh88VRbC2oe/WSvhpnLkzkiERn5K02LWymGJG2NKjhiVkPNzPm1rLYOa
dOZnW50W12l4uQYGCAYHH9A0JXvZuKeywYw5JpzVMLxYNLLPRaK1NE8Y3aQnm4Z4
xH7Zm2jamLAKebFLY5bNSjyjM9JhBQjd+26W/O0dSBgfKeshKyZumOZN0kOL1StX
C3HWfyoQgn+/KiQ6o0VS9+1qBzstAvVs7sFcoksGyjIiE6pMlzYsgfXISjW69YU0
gayFqX8yWHt889WdhYoe/V7xRPczBjQM9Z2tmSYrkLrcR7/FkPVWpPcOG/xH2MbT
0eHrAINHa99HPBrBnxQL1O496CG5+oOlZSaSXjsTJ60ze2316j7NQL+TsRt6ga4G
DoQnxjrGYF4HsVW1Y/0kstqXRW+72CHpugcM9TY9sKKjR/W8dJCtTjPMpA3yO7ZD
Z+ny+j20yaiSXs8kuhmee4GnDWbWvsg7tfOMKwUW2t6X4VaPwu/gpyD/gcFABQsF
CPe6O24Zc9h/U6hZPi6XMd1W9xQhONIIGYIpxEgs9tZaUfKDDf0QlLNOKvwimqql
Q6YjbYkY3ZKbmqg7Ayezqe4cryMWHawnF7hTUUIYD/TQY3W0wV1auR5N9C1k3rhb
oJTWpRvvlXvLjQPP4vxBTuOqudCtYBV/AlW2cb59i68tVBCXD6qhKe7W5scIn2TK
QI55q/Kw5AgjsbOa5Ig0KR8suEXlbVrtvt6dKyld0xyl0njpvNRERv2EZmnPfifV
shGW/E/c4I59/hsC75DHMfxkNuXuy8JNye4y73C+l8lRq1Xc0Ll3cBO4CxCdSUcU
Gybm8RGDkB0RPLpH0/1Q5QS+sZWcth4OX2w/He9RYhKyDRz86Jisss5eQwIajhBq
OrDK5Dhb+vuFVlOaUAMOYPQIGds5RFB2nXoWDL06Q6WlN9cEWJfpG+KP91aVI/ci
Yiwnoc5+XBCObG2A5W3kMEhCzZ78MB1x6cDrz7pSWIQs3MR1yeNXve/IpssV05wt
ayceCoQbYLMijtm5XCIlPbVDQmQEX6++CyTIC1rHPG1+YCMvC+DjEQYDpBKTVCZX
2R/c67c/Lho1zCKEOFNic9wmJZEjk7IVuwRJ4QssXeuh0AZ2IYcqNPZaNIjvcD6D
JCf9nCeCJSK2OEwx1IQVc8O97unUa38fZQugpBV+AQu97VMy14ykVoUhfJZh3q0D
i1SHXsXWel577o4GyWCy6W/5sAAIUb9phBTd3Pe6NyjzdxZZm+QGXcrwZR/Sw08a
be8rqS+OqChUz8lZnPKpPGY38//QisJam0t+abjnwitQV+nEg2dKqe6ObXzu4hAe
w5rk+CY+6HjEHYLefwTXCqWahw8O9hg3asIFOjU8+b3AGPj/JHe/yc3jwK72IbsI
8H1ygMXCHMXP+bIUfP6+M0yww2DU7+V0d7gRLEORIqqmF3tzPSb3OKDeBoGgb5av
dPRrASMUb+gxNOjGOq6zOpxoqnYwpl1OD6DW6kU0GGMbd7TWIAfZzcOWzC5hz6gV
yuaYS7NmeO4n+vj7kF6c39U7FlcUd8oHYe3VJ/ZmFYUK2BJuW/C+nSNmjNG6Pm1O
Uf4rkoFsYLpx3AJZdAFQUZomWhTrGycvgm1qGXuvjHVx/XVQPykck1EaOJjQKJuz
PetLxA+joCvdJ1DJae2ARYuXxu6HF86c8L+x9xgdls0easoaOigUwTr7Cn2uViwW
ZrzGbg7OYJUeKLQ+YpVaOyXYxumQwGr385HRf7xDBQ2CZoT+DZarqVQt36LhM5lF
X3WPPogSJbJNVPD8tAPt3upDJpc2OMobwmq9BBH4ND3QtaJ5vQ7MH7cGPP6w7yDq
hx5oicvwOqEchBwdYPiCA3j/nqAnuSKS0a+CNGO1WJ1LK1UtJ6Cw0Tw3HtOmfjDD
lGPhH5Fk4l3PoFT3M98xwdECgKkHnUPO58xhZMuetWXglWwvuymfD3lS9Uuf8LB2
DSzUvWqF+7UckbjvhD9j0xuGBSt1MIqpTTA+zIOwzkmtT/Xb3//+zqZFAL7R0lVy
XJ+7vPTYVApXmH2g5q9nb+4oJnWXHkMbPNJHT4NOhM0oVQVIZfqqsfORRMcE35XA
NaaXeGjYCTeZQv51yHuogkhYM+7qU8Be3AR60+b4EPOfHkY54sLZ9B7q/rZRuLaZ
DibFlbQyqLWieeihDvpiRp3WWSSf+30jyHXka824TwI8zIANu72rb64zGs53q8PR
Cn5sfLmYqKecj6u1SAgmFzx6utTKnAV7DpXONkhtmhIXmDpNT4Zrg7Zqka2Q+f0I
bhBiiUoD/1vSeu8TYttKvnJrKlR5t6y3TdB1hkTDngII+U3osIxOtSnkakUblGzg
iSN3ip+kqzB+FeLFXf5lXexD7d0Ahv/uWlsnw/fJfHNKUEo7BnQJ98kC+ViBM0Ju
WArp/cBJsUlIadwxckENFyOAEXHo6pjZrXA7CZuvBB75BxoHU5pkE9WOVskmw3Q5
nUV5+7sphweHTpBltUgSE0EnYo8TPF5vGc8/cGfST2w4UIRdxe1BLcLqgwmBRw06
QWf0kdubJjOszeW2t8nWExdJ1j/lWVt/jFAD0t3X9tvis83YY8VT0181EaaaxACS
x2r7ik8fZw1HeaZP9DRc1BubIDFqEMA++j88EuSi7wihurVIqY8N+a6aEO424ebS
a/9bTnczTEHGDQuFtDFJk29tZQXAgon9nPqCD2ACWJPk+olvjCzesYwrPuBJsts/
5uWmpq+0vitbY0oYyD+bVb6YkDJsP2OAvKsQ2L5KQQ4m97X5dpYeAR9gpoZNTzH7
/EM1C0GOL9opbbOeJ1cU2t7h34f36u2iMxncBZVMnkyEKzmC5xObViqRslwb8oO0
h8uVTB/ykaUau+A65XnKgoo7eYdMxgAcaQ3sGiVVjniVT3sIAyhoap9upZMqLnzS
JpxF24mNxGdwE/E0/L61DAlwxjsim1ejTI2Na86Ub8Jp2nmnq8iSu5l5EymXBf1o
aL3rk/nioHm+NlUoM6e8szuszAonxr3oI1z7Q+bwy8Xq5cW34bMJB6y2t/bdaPfF
Dg0VufCKJk212YtGlZgkpJ8xJUZDqCz7RS+BwIwl4ZNWoCThCl+jyTRjg14ahg0R
lOxSbpzGtNHnOFCeKLuK2W+0/xxg/FUMNILX5tJLHxrUrmc5M6PLTw0r5/PrYydu
J4mdrEltok0V/iS2o2iytJe9tV6rECs6U1+hrSpYYldaZPdF0QjheroLYN/lzkjf
NtQmM0z3zAk0UMI3TgaD5+rBGy3PYpODBCWXRGfjyI18b6QCGe20TXbC2NESb5pR
NHIWMZbd5egM9sTddHfxplE+eDV65F55VSxylO3aTvVSAJHEraqs8JT3TKp/81ii
i8TUIhjxJL0wiKZZQj03T7pCcNpew7y1NyC6ygqxkLkgyLIO3hWSXT3pOrXtJhN3
Kb4TwSbDTBj6NRp3dsDc3XbuT6HcaG8OCFIyekYA9u/2sK6sH4z7iXMehi9oDtap
+lgH9XNuNub6hBeRlcQjNlbd9hLJYDHnm81ZY0MvCz066zGdpAZc9yj07RT1zvy5
ni5d2ZiRqQSvk/Z1eLLRut5oI3I5dTV0ard78pzZ3fPQLHmqIajT+ZQnxYmfVbzd
lmdCBliHZR3sqssKjlnZkaZUjzF05AOf9wPlHDmLh6Hnn74XSoPhlwf9O2zQQc9l
w7kw2fz4si3cQ9i6Tl+bqHf30yOTbNB1nuevFxSkRLOySAz28DUu2c75JX9MbmNA
ow6GbdO+q1QZ0rB9KHnCsz3YvtChodck+j6mA0F9mXwY/GG+e8ZHm0YyFfTp/YYl
ca/PP3yneJBtTWPmaGc7i2SpRWC6mbKYlbDlX49dD5v+Uz24Wc3kBotkUm3EPNNw
dmw6+XJ2+jbprkZfCZmvV1Tg+0e5IXOylJSoAaBx+6mkOWGeKlG6cEkgQZzEB4EL
mwgiVQeEl13K01kvCUjGnhUK1bcSJghDe7qdqkIkbFOJhAthePWakg5fMbFcbvXW
OKXJbRDueO0UOtRJtu2QU7rV+3v7BRi1ueuqZYEeplGSLz6pJ+9kWKWdbQ5hYbtz
Xdk/gST6km5ZxBeXTwLCcXRPA02S4+8uJrHAlXs+eYbFIEmX4J31Asjozx/Vyp3n
yODz4amiyoDS1EZBkloDSFC8enm4yUdf2HxHV12yAhytWxEUJIigsb1nTfJRzHkK
pORY27bKwDg6QQS+qFB4J8u0/HwC9N349mcNY8sMsRGPrLxSJcfL7w8mdjgetpCW
AtWRxHncCtRMpSjguI66DyEPHx/HlX8ZylSToAf2UsUmiPdfiYW8ug09ZVSHPZQy
C3PdGJMh2MIzHxK5Jnf93+7sZPIv2DLPBiSnvUA+ujIZl+kYfsLaFSDgKAVzuZ08
ozf9gvu2fDSBMGERQvpKXqiGC06nEAK/Dnxfc7eMqi6PN13Wc6/laA5jNai8pQn2
IuMAc3HpHD9SaEvW2CIQAtpQJCk5pHH0M2rkg/+3INa7RC1iG5ujxKBB30d31XXb
kHw7OcO8rUUHQ+44uy+OAoN48bwzOPA4o1iX3DCpufJa6BEJjnMsiCYe2eMjXltQ
TWKRc8POSpvbM97Z7RpsE67ivpoXlkPJidsC+dMyFj3GfEyjaoriAJsiD8YMVIWq
MTw+Mb0Jbwp1hZKn7sB8kwiWmTq/RY8TdfwiEoJpqiYa45vE3VwJQL0Y9j2iplMr
uBZx0ZJky5qRdWqmcZ42rAz6ekjNvQ6NkP4LamAGZP3SlYoD5qYaUWhS3C9aDZ3Y
HQkRnSgOOBMfXHGRZLOy/UK5RByUy613/TPkFBA02o7WVvXU33yiyO+qq2rekf1M
fEwP9waKO3EufAQRNQS854L9qwbyO4t4pinHbNp3C/H1tVjHApL5JtBQbefrRqc0
WtxO++Cf/4x3xYwmub6S+mclwQXrud884Us/yj1M0QKbyw+yHo31Q3vkzk7hE+4k
Aho99/GISfsaT3ylv4EwMEgEr38UtwAZI2T+yor2s7BCDFif080LDaaMw/9SGoHJ
2qbiZv8yCsgbHpXM0GLdvKm8ug5pkbkGjmQzkHf30tjzFUqsuX4612A8KMheS30M
3IzWj4aSVQpGjxf2dBgj5hAJDoCXoYn8zkGJ+SAyA8SFgpm1rkNMjuq0D37gD7yr
Nap+piBI2nCB/Q0FDBViW+UdotLnfJHk16FtilSqUGOf3kYb0ioNwWnz+F+V0d1B
eCiViGRekrRJz8Ge7T66gpQJnBVCbXMGGCoRgynvHY8obs5yl++czuDYQl0gnSfF
Se9U8wVQ95X9wI48oymm7U0Z7Gk/NkYaD44elRnZcOTUpEM0oBfz5ThpnYPnPbDr
JoH+cjLZj4CbefsRwnGVj1UXRB2y458hVVocKEFMUheAbYQphr/nf6NFum6Ik+fI
tmJB5qgmWgNAQdGpXgRFDNl3CaFuYT1Ihuz9rG/OBpB00ZG4noxA336pcIfmqPXk
AKLTYTI9694VBeY3dZZUpSPcb2551V4j4xogLJNVsA5iw8IxP1FDflf3aZ57LQl9
vpxXcJDrVG/tEn5wy0o7CzIptzDMXI11Zie926z42D/MgmRPhBIs55rE7Qk4F7xe
NyNGCxk9xE9SmkgnKDygI6NISqRcetA0Xdu5HIM3EiVWe3y0FZEZKEVyGSAG/y4O
oyxh/0ngzV6ibqryhbyqZljd6b7RBiHRloNHF6ZzZZPNnOw9MXsxxbgLG5v0PeQy
GM07YjNrMTrFiKXNmWKbhzu6aqZQViO2y0lc8+z4+UzwdPC3Pf3CdKbqV0MPXhxN
kKsJx5rMHJahlPQjs+cP7YRVk9NrXwPpx2Ik2wPu24RJVJ0AyIEla2Qih6tGr6i/
bboXUBE7cprxaEumhtFVruqVh42Pl3foG8uh3hT4xpnxSgKpXHO9Dsd7ejdCfOa1
u+MW0fCHa29LaeyeeVKYJmtbYVG7zY2LNYq+r6E03/kN0Ps1DvVJD3JKvUlOU4oD
rKT7F9wx+5o/THgaxTl67yT4/D905oZLyXCGkRxlpV9g2gTfSLmPINvrweyxtmg/
2XKk/oxdRUW/WxPPx9IDIA+yX1wEWVW9bkGD2R9X+DSWSE+up4ptROWuM8JAUlXX
/jMvu7TgVMfkf4J/zAB7giahKV1tCm7lBoVg7HvfKxC5/uriIyP6TChX1TK8QDH0
2/T/DZ4r3PbXtODUHdX4g0+zeIJnNMjt3ZbZubbm2s6Y6wn7+TMtW7JKTyMhGSum
O7iZDgX0EHn5WvyXAGz64wGPV3zBLPT2khCVUzD5Q3whdmx4i40fmPhKTLuECEdO
eEomVW4LpydFGEYp+XVJADEL+X3uPQRicUvB4ZgThQ35JuDaQv6s6SKCsvjitM2Q
dCH078mi00eXdSqv/lWkFK7NJZ67U/cRXNDjcnawMMSEMIOTr66D+0I2/31Z6OXU
ZEUHmu2EpES+H8ao9DSn9Kpk5PIF0LGqGQOMEybv2s0Gc22Njk7aoIq0D0Vkr9NJ
Gk8PBqXlrZ05h1YoLKWEUEco7Xizsimf5Z7kTEWQl1h/PupquqHvKJe6J4cSrdHY
HwqdgBsr+mHQZt62q38X1K5hkfJjVeP1i3bcFBFckO1zJfB5Eko0tHPSxwZDY4f7
LNzCTF0qSkQIUD7sl1O+zQ78dFjYNk0RECsD+9q8kKz54uxDnbIt9rI4NVcgym9n
Kw2F4XfhVTgOXy1q86n+n89Cfg5sSUXveU6J2AZCCsYYpL5H6ZS+FhRU0oAcKzFd
1OX2eHiQD9cE535UbrQlnjK8vYor5avdDVyarNWyabG/ICp7VXbe61dMAPvlYgF3
MR8Vwww34p+Snqms8fpulaY5hCRZotvHnR6Yl9/FiNX37PDYxvS32QMpnGwormeT
WEbLC9lWiPrwBiXkR+Tw6sU5mLqXv25wuNhb9oqgsR65xHeuu5uYw+YXpQPJVRw9
7ZXIs7e9LqiHhlSOc1B6RZxrgy0+E1Cu/01RthEPW+p7XGtcAIaZ1XZxuAU7DknK
DLndVq7CUlnZZV5Ba3q4xTvXe62JMfa/YBdrjTwGBTFkVpG0bkSSh3TuqKMr6feT
8xsSPfP2qdwjqjiJBuh34jow6QEqOkT29xsnorxYeHWC7UjeC2ABRocjSgC5Byu6
sMO6dLmt8skBk04x5xApj28sSTzEBhQzVtiUS/m3qM7CSCiqQRye0NhV0RqpDBYk
9aPxcTV69lHMKgfqC5TFkRw/avFCVdtDgxDfPvUXBzQ3GCw6CegspQYJNZgRyNgh
/jKGTkUgu+sKwLInWsrwZJAW4JuGHGrIdfhbSnB8b9QOZpNzqODWTaLhcjcskghW
9jbebgoM3fzRCYCG1aLs0TsVOm2C8cKAeLWd9NKg3lP+szbQh44bAp4NIMxLCeBR
I4WEhMfGXGMWaPzt7KS4xOAwu28bAx3t8EO1oOrmogkDw9s4fErYIbgkIlUevqtA
ofqA4QVccOudiILBjWMXFM+/+AVCeRNyFa/iyrqrtJE7UaOwUN1McWySP7ySOexm
D1LMauxl9qPa0vGRhIpBAcKhiCpJykbOWkpaSKfhbJGoVUhjMmL6v/t5jEVTX1wp
Ks0rX0PF25qU45GtaUhL2fYnXb2Hmine4UOV0vpsDOagX2PISCSMKPh3MuUJEJwK
Hgy0iUwDldTGCanR8v84Bt1Wa+Mo7FLBnnYQM5x00PVGuOznkTUMFHxM+Qzthg7r
QYzfI1z2C3erKDvrtPok87Mv8huJA+q9lYWKbJhVRJqxn0WYnsHri7Oya4wVldb6
dubhPVN1S+LNF+OFAGefLCWtCQCR4Sd7lgsGHOFreUZMmLgZOQB9I4uBYYLWW93J
IeWpxIW4hPYeQjNnxLZdN7ITPHl2tDCiRtvYY93jWA0rXgnYDepM8K8+n7CoH2Dj
OqxSBLukexCCVP//7YNUSNH1oAFO1NXMUAv9sHS5gn3aMjZMH8nOg2OxVdqpwc7i
if+g0jLyOTsDBfyL6dEQitkEtdfwY2me2sp5ce6DHfRZ4pVo/UzSjgIjpcIwOi39
5oOE5XM1AxE1JEk0OD4NnGW+Nms/+TcB3zXHpyDTf9W0KcVFZZB7QjqJJVaRSvFu
64EALBRDGeqKrdFdMHqLGHSOx4rq1UlloZbE6x3KAzW+COY2LWOLwCXORfAsCJMg
x3X8VSmHdlTH6hN3H3o+2nT3c73Too6njpbh8R/+/fMDyBQZcivoT+JZiiByfVkR
6uWFErv3sz5bb8nIkjOX1kcWjlYeSlzvuSJXn7RZfIRFddAAJvv5STprwfD3HOV4
PeGgPkajiq77ikhtAfodbW57QB96YK+0Gbd0rLYl96aM8ehIsLULkaNA3yWSQ9bV
D+nZWri71/qy8H4AVi/JZ+77tvHsi4z5EkR6WoJN6oTQwuAh23trxvwQ92axry1x
ocOuU4kcROw4PuAn98o6bU+6WT+9GWqhKwU5z7oNiz+IZQGn0cmwEC8ysLqED97s
Vfppg3G20gltAKcc6aOaRaLygrIId3c1Xj2vgnbtkJY9I31DgkCXAbjuQRF3kXr3
ZA4biAWaytMjL/k6t4uGlgylZ21NJcEmfuiVKDYMNz5VLIh67bzpZ2hz6w6BfWqS
thMoK+cGU+HxHyPNk2fCBMDuX6VsAiQtndNDsLQzSgwhqjC4Cu4AyWf2LojdlkBS
NpDkYYh7WtUTJempcg7psg7mi/Xcp81014eA15p3MYDvZKM0qz3Go4982L9mXhb1
IuDLiIAn5ywlgobCBtQMvYsS7T3hu+jw/wcK9HsT2GwllIF0k6ivUvCRXK7wLXvG
tAqceFwnrCDo9MxHc8tj1lRvrcafkvGcABqEQM3Drd9LfD5wPNWYFcAP0hj2l/VM
0rr6PviG9oID9qTiw0bxwDikl5axQSfUmXKue0PSrhCfWwGqAiYHac0bj4ZUPauT
HD+6J4yMcICcGiHyvB4bjPj/+hHB4MxUQ70X0Mv3dO/Nr5b+bHRk+jvW+m9+319y
utXgvqpD8HlnFeGAwGCmwMLC0SI8neuJscP+37sALY5zxuKHOoYI5U5npoxPaTWj
otz44fYKKMJp+FoCvSBfwZAn75ozAHen8PxO4z3If6Iz5ip5Adg7If8O+VOEe5wf
kmAQcjN7UMfwPWyDiNkDS4iuRp62BzdU9mRIvMS0kXSRiBTy0cbGfneoxBNomVt7
HzsdaxVCiIS4LPUeY+qG6cZWgaWng0VIHmqN1WgswPwBCjWFHRBqMZQl0eouoDFt
iqOBWovLZ1vqxFkicizUCcys39Hg+NgK1t7PdYWbLxTO5AYHJCBnAuBCWBJOOT6/
A599D/dpE6FPOjlS4clIEEDW7otmKKA6tkeRylTjDRUApBILRmas/Wni3xxIwwjZ
vrbDULfy4fheSNicZBAc99NOv6H+liTONLC73ERGlgA6m95B9M7seLOHMDPXK5Go
1984/rNOgwWY3HlQD/coydLhApxqPHFrrdnD77fQ9nnD71trBgp1KPLo/h39eatq
yqO11xUJB6jsVFidygegGh/47XjOnuZa/bwjedYMObMtsIJ37rxGQPGWybnLFtvf
4gDZzaH6pwBrE8kQ+p58rxGTbie9W/o2kDz1dHpBHRHCG+wvALV1LZEmjSJxnksY
3jS/54nzS6NbqjuXHyNkPbIopp6EFmzkFPR0EEYiUM3F5S6xnXW/xZtBrH5y8KUd
9hHQuRa3osCfZ6Yh+CsGW1r3ILG4VQqi0ebVsMPECxO5K6PHZoyFzcHYvwbCO/kJ
MoOOQDdytoY34bH4IYbsYeEWAv74m95dTUQfK7g4koynwSNdU0LpGz2LYHEWmcaS
LaIDHuiuF85t0Q5CSpAIBHBChxPxzBA3WaA3g8MuNxXx4x7/spHHvkz+HUmX89TO
vp0i46AxnvS3NG5swCR6/25QoTSW1mPLYS4eD0E1QcgIVtWwbcin2i1dpKFEsXMI
K/MLKCG5VQYAANQIj56VJUhOC654F0j4099mBQjlYLy689mM+EVphujsJGhaT9J4
fUI2o698Lb8m7+hw/sISAnoZkcKMvQHNYg9DMa2D1Hh6W6ijn00EPSYqmKFyuNYr
nFMinaLs4e49b5UlLK7ILtKQDfdPggVXWYHx6MGTz0xqiSpn2aIMvSYcA6kPkItl
EMMneC00OWbw3NNOVvrLoVnvuGaHrZ1R9KlFd6BcJOHVVBNvMjbqAvsoR2Ib78TJ
qpAaIET2Cib0l+0+zuz2GF4UHSV9WF2KB9NkEfabKLkMKvTU+mtuF6fN4cVt2QsH
AGmTzyZGYtPQd2KgN8ALYYMNFlPki+FwrbfAL1iMaVp/Chr82Y0lUWJ77za8acos
TqV0kNQax30U9F/pNX8bFSTrZR4CewKfCm+l1yi8swOpZ7MPczaKt4ag89j/B7oJ
A+Z0N1fzWpBWkhbkkYn3axVIqKWdt5NW4k5dJfk1oxnc+yDq1iL2KA6DXUG+j700
P8T1ewv0HdZLDS3IEoFXprF/Zt50gNzofcclZfsUyHe+Pa/2/7N8+Xk8513cg8Rc
TwFjgjfcR/ejNsUm2YUg88AZPdG4F/t6Fh+beSJRu4+bslOAeckiCH56ofZrFEB0
0R0QCYaEsYO2CbC3N35sxvqjN4/WHfU0lmEx1l2sRa1TZD0bAwOAn0AdYYmJVTIY
TZriaQbLr+2JiZ5MAkOJh1TA9zjMYTOppJwvNJFKEL7zjVeJJuXHUhj6ChA3efpH
SltBG7plO5vJ+m9M9dF9UGtIPB30WEOpRzhy1xS0PozPGWsfb5qSh//7qOyB13gm
8Zbu1JU1gyXdIzQxuPI8nSgemMSfua+Y5iya1GGqqn1BPFr2n5F2deLCaTNgHb1i
/itbBoLte7UljYlaBBL5Ld6Lj6dUFqUilltie9PGcj8UvoMecefk71CTvUpMEr5R
OTVpNtcVNzQRL3PYejzBWDOTO5KmS9i8Cb3W12Znb5n/x0ODaJQRZZ6JlGyFQ7eJ
tPFUq3SD/QziIn4YkxHnqosWXNqb4PXw38YXFzkJ39hQvK093cmpCZepT4mdDDc4
YYDN3Gl9lqU29X0dbdSTb7Pc4LNkJ0+Um7/D0okzX/7tK5a945+hf/eF/Nqpe37M
vBdLUc7hgbLb5I/JMlABWQxDfs75oVEgLI4JWYmp/APtvkmwUdNxjhcUOZ3Nqed/
fe455yTd2THP2PlFjf3FVXju3U6IJ5cuAbVyT4hymt6XVvVN7b10KhfCi26tMl4E
2f1zjRN12SGR/qw/VouQQCLn8FxBdO3W+8w/gnqhRp7tBRn8xYtpQUC98QfnCU7l
GPPz1ZVa20GLwo0xED7KI0jqDiGOXDiiHwRbZ3cIqolBPpV+fJjJexRQKiWan6J4
+wnjsXYmR2x4EdoPC02gkogZG+M8zB8Zs9A789nRIWnqYOUqehCA5tJ1aAL3osOw
58ILKXcWzcBmMMF3BPmN0g==
`protect end_protected
