-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
K4nsPobTTL94nAKx4uACL77Yi91LU3k6XyFchpK0xBXP0Tk+D8SqjzP5Ia2xM9/B
b0nuHnHXDJkjZGqiwOqjb0vow48s+/chz8cAwZFibgjaUXAAwXu+pPAMWxZZlPrq
AxEdgyJbHuOygABaUMSRtWm9aGx3IqH7dM3n5cpoTfWOgYdgFHGKQA==
--pragma protect end_key_block
--pragma protect digest_block
Nz2gqX26wyBQeF54Nb4s3CV9sII=
--pragma protect end_digest_block
--pragma protect data_block
3hfJNA2d5S/UPE4TwRBXrjCpJIbRZ515sNfZxi6MslXqG0jOh4ZQ3XbiDLOPLxvb
4/2j+iCZbJMgZ+3YXgOV31rUn8VT/8FrpFVH2qEr61icgjm6nErIqtvzheQQel/K
T8uG1qkC0qV9pdEdU599f2wZ8EaMuDCvmvHU0LviiYrnQEpl5ef40V6pxAuZAzb4
0wkI/Aqf7BG5Zyz25xH6nrvhdLAq+F0YcSlnyxCuIa9aw28INdZu67sBGJZRZqg1
1cidTvMYdOUT9LQZr4VrKBSyLAZn8gC8Iza5LffeszV3l7ym+qObZ7Da7Y4b1Qnr
d/0F0nTwYbzaZVoYwvTbMtElpy9M+tKBd6KWQeJBy8t3fZWpwIyYkDtpRCQfjAsP
O+ZGuqESolpR4rUmsz30lqs/iZEuSdajsUKtTO8XPzPOrkiifjsnO0r85/vnH7N3
fAsY67XprO7Mni6kSXo2O1vpMmjctEZsAqBwUtNfJbqMirVjx73RnhIq4NPgoDEp
eANpvIN7Ey42MGPpsLJd5Q3o7wfs/oBKcQUSvRhhUNARxA8Xy1LswBh1QViHLcJc
0uwsQcMo89gndYEvoGy5nxaasE2iFzFKezTUMxIpgZRsMeM1X9hsOWBg8o74PSsn
MvQjbdQ7quqVcQIev/4AzAtQdJ6lbgNb+5b5GV2RQ9tvxVdCE2Lbecnx5XUj9spa
MhVbVmwAdfGm87YLemOT6gg3W7HEPd2JjxoLB74CyBwYfvQSq2nD2div1JUMU6Dl
a5nKK7bY9vxfoFOosh5mUr1ACHFCCkyJcubyiD3kFGZtILQaFAlPzz2Xz5Qps5Yv
6WbtFqOzkhLr/0WGbI7wzToMS1okYlOosy/yv11uu7fe6FDLEGo0yfWR4d3pwTW8
V83ywhRkbsUpbVrim9EkGywg8A2t9vOHrKS50bKI0vY60dGnBcle9OytQPvowZrq
OCdNWzKxLoRiJ91AsqxNbq2YtMPo69vssdhsZAV0BACafbs4QOoOXxzHGztT7n9i
n8M99k4d715K+FjmSrjpgC2KtnsOTCwfnX5xvx1dt4l/tXAM33sMz12u9WUkqP+v
CLqKtxBS03pbiiJ6eECoKZo8J8ujm0+s2syPukaYuFZRoJuOrbJjxdMDp82I9JsT
obNCPynvLibEMmMhEPA3sR3PT/tUCsGQC76+HAv+TDrk1Ws1xAaJMOIiXww3xUxJ
k7/IUNkGXHGM+GKqgd9ovoj9yKXIiTjrycSuWRVvou+6kuv/H3UroDC2semqzhmq
r7mh28MHCsHtLTwmE8G1CxT4ypKxwJtQxsWrumiNJGlu+EeYKt4rtjdh7afgWXhE
aev3bHSrHbSxWVlRj2BMizIXKG4BqR1p6kn8XOrLlTwymlT+HQz0n8nsxXpJN4QU
Dq97LyeslCd/K3pfc1vqzaa7ZsUFptVQR9bQT1qSxumnEtuTZbOeBNdGDku6EUw3
Dm9CGiTPQUDPuYAIS+PaolMDwDUgG+BTF34toHtHllfnlP8QMsFYdCNCKNpsAhBP
c3ttDsA32picVhXejtqvlpFozFX99OMTPIJ6WdttgQ76Ef7lVOjWaRQeAEBdEJq1
nWWqn176z3ZQoyzEeO9BAS+Oyg4AjL6bVvoSDcQWdC4nsXOcyPzI/vSrFYT2/7Es
y2oU5tR/tblAcoHoUbo/aPOabmM5tbXVnrPLiSuFpbfVGAWrDAx9ur5/Z7L69P0F
BkpIaBEqQa8NpO4yOB/1phxY1/+Sp5zDXJ4mzAhOBU7S/gpKri6/NelyWZlsMSug
akjb9zPKF1TJpogBsl7e4k6QJllFK9dymGzjMfd/ms9hUnf4A0crjoiwnDaBLHXf
r7R44RagB8gzBSnhOKcZnL4IZJ94I7ikpjxrtOaLvt7fbq9YjzJ3394CUihUwmBd
EUZ4z2Cz7w4zb9NH50knQq+HrK0wIh2+tkqwHT4sofRjtg5/efm9stU8JaB/668z
2BoPpxLJSfgEkX02sUm6dsSGzaQ3a7XCeDoSTRsL2xsjvsoVGOP4heDcZWijif7p
w4jorg1snk0htIj5nRQcur15t8aXpLOh6GJitxMEbe/QmXoojWQbYfU7aHr6s8bS
e4Dv/HukDIgPk/cnRVPGHnkHKVnbtfJXxS1h9kuL56SWVbb7W8iVgg0pGhpKaBv1
+/DSgabbdcnN8oKA8RqkiHfqFApF8EFkyuxP4bP9j48+fHu6axg6d0q0vx5LJpUD
26iSXloIEZRxTUdh9YaIvzkZI49yOH0Fjr9TP5DNERqdsr6QsPHnyxWq8Kg5bPae
gKjNvkzS84LqL+NlkhU3/jAQcvQztCw28dKWdKlOKztBOY/qES5d12YXww6rzc7p
pQVe0iUPsZJgifQ4Rn1qph9Zga79mFuCbhEhqqjelUPZZxasgyZ7+4BDshA1HgoJ
bXa5yr+lBRe1Y95gpqwvhUaKFQ0rvqJqpvnKVcsWlMzGv2l0HbUTLOOpc4a5wu+2
sYqF8dszAb9GhS7i4qNfendvvS/dXC7pE49j7/LwNi3B85u4JgdCpF9mWptdpVCe
NhRRJEdDcnOiYZTuBbm+rUPnXw7X5DwwC9NfxBwVoRujJRdK5phPd3NuQ04r6GXu
jiW0TARhz/CIAIlN5XFozPJ3J7IA0EKDNifFKVgJENvzniJTzOI7/Ie6caFNWoqg
NGHlyafJclaRVM7YnbZKMI7hed5Da8ACAiSGrlAeHw3RJwl1VOgSp92B4CyJhdbI
o3m5iWO4fqHyYi45bHOM3IGz522nOghXiBygtAbxYAo6a8SwUum73bzRx84Dbdq5
QuJklmt9Qx/b7dtPsgVkJADI6kgyFEPLOoPwpNC8PTVM7p0P1VJ+wcld1l8Nyf3b
glwu1bYH01o/On67SutRrsw9PFmz+3qqTi2fm+o7U1qfToZm0k8J2299wYaxmY67
n0cHc4PlShUZF2Z5rrhjqPkP5Zc+bR/GvCf06myWOqzzlB87/w/0RhkhLynp0JNZ
2CgmaHBh6CcIeooNmPDGaozjN4SFQxdD69NrHpQ40pq33imHoMsskVdSQlmhoQpV
Nto9IZwYVO4mi8oA92lX2yXlLpvo0WdW9tyGwvqshX43fo36vBNMu6s39zjegRIE
rAg6l2QJypzwIklJIaxHdM0Jqn7ug1JpOVGX2IflvbmTzO/ywE+shTPs8Idpjj3w
Swypo2ZRdB7m3oHKDNNSIz88BrVmcnl+c0oOou24JTgfnjJCIWcyL1vmXOlVBbPF
WtkMPTT9dMKGl6eol2ndGMv3E0hzekJk4UKANdEbgpJm1jrENgZZwj9LR51DgDWW
eSM7q0rrsm0NWsZvN66jP9uJVt+83xBgceB/dKC1OAB6GO7W67CTBOyYJeEUScuC
tIC6vdd1AIFmMm3CmdpL2s/Z79gU+V0ha1ChOkLyJ9o5piEHgfGSfXb4HHYbdRvO
FHly4jF+LvuXxyZQJxI7KgkqEln8/mZoF6qSmxHQMoZMtv8VWMsvNFoGczoZ9esF
Rg0d4QR+89+LGCAwVUn7DgiwPz09taS1nM/1AFAKkloYR8xmqzW+ES8+cNOqi4hy
HtYNfdAdL50Ik3m8AIOdn5Cl3+5UVF+Rv3b3/i50EUrX5GV2fZzeGGGU4bGcDIq2
idAR7njjUct2p124B3Y0NoWYk35fW2MhKBoPc9nwWTcmLqjKX7Sm1jLdG6pM7OmR
Z3wuks9W+eDW1MNmlHP/k5RBM/1i21h4FjKsAKne+ztCZFuvFgCFqfC5u8q7HExX
ffQhcc42pYjsCJWN3Nv63ROvDqj0qrkZX9eqFzxDVWzTTTdsIEegeS9MaL1XO+fZ
1jxiNuaqujKxrtVsQbqXgsPe3bQLb1xjE54DSukQkPzZN7+8LXNEYj118OEZOmly
ZJ6cj5yUGAkOPQv7S44qUnrksFvjuDJWn9NUBwXZGghFUkGhzGn9cvcv/e/j1cbG
i1Ql4iN7pB/KS3PsKT5pNviqABv6O8wse8lQ4MckSBexDsn37jNfXujw/HB//frv
b7AHBr6hjRbOBRNLDFkV1gY/HwzMEoKl/idilRG32FpRjmT341UvqsQd17daSaAJ
fSmEgeesdRBDj7i4cinwu6J1ZUtfdFer9uSps/YcA/qd00vo1gm7L+Tgjd/PYltR
f2jQQjg0MCL4ITeaEeLuF5N1oiMwLt6FIQPpDVnvKdJPgQajK5iemjwHZzV7WCiG
FlqFXFnaHxzNz96pMDU3m9+Oh2zYJxt07GMGHOW+EOrHnciSef4fMdQm4znvUCvb
us4Te96E2rksSKUnhFeNDlw4vUNX4IK2jxdnC3lJ2gvTJedCwXz3T3spiwvewhV5
B+PaTjULnYNMz/pXUeyTH15YBibVtamsnJ6H5DIS8X6O1Z6L2xTuQAKUfjc5uF2L
FoWEKTgUZUNQT1oCvTEPvxgwU53XWc/2acA6frZ02XK2ZJMn1lyJcrrbTV7qqJFP
ARZDbO9QTX5p++6KllrA+qEHY7C2EFXOVbhbLT7e37/iJ3sRy/1oTTwEeV3IwpMh
t8dWZSSjBOL8e82O/RVOtKEXhUYbmAluq21mhbL/9hNnHh+KbbkW4Dtbk0lFVKuZ
3GL6Z1PddkHZSwdy7KaW8Y+c5dz2LK89/wGOdBuRXFdi88jk7h67PKHqHcIrNTu8
6K9dsLAD5OnR6l/CxozQsj33NVMzSZj+YeK9w750qlHCuqaBOVdmWkizNXFIa8Po
niswPGGmURwtA2nark8bm0U9/vTvMnZPCzAsbjDAf5oSi1jBpOy8RGFgcBlUsRq+
brRxkTaa4OwX5datX9+SwUsxTN8qlriU45YaJ7Q7AGes36EcV+lH/0zKH6LcQMss
OFlwgT9JJWSt1cypXn4o3qNtd+v4K+Rn257f7Gw6yujGaO6fuJzl4LELwL/5qjs5
4bVgt/mPHqMErWm0btY+QwywKPi1+PYf0+d6jhLUuPJIqR3yOCWYczTffZCZSasb
Sv0D7l0lG2yubh4e6iMKbv9hfRUm/J9oOXtbm/KQK6B7AW9caRVpFyH/0xE0120n
kHLuoQ8zO9ExxrWT7svHrg6Q28Zbu7W/ogn1NTAQvXc7NUAgY6mR7NlA0JRTRAEU
/+95hxnxPD9uC9wXRMSxeS07OnCDY9GgIG5XlbSt0sU5h6P4qWWrgsOPd4YHf9Pa
qksqs4lyx81ri44OWBsYrpN3/AFvCToJmfYVK+4cfQvY3/0/CBC+0h9z5sR+/4aO
HJss42F7QcPBQX9I+lrtqTsxocx/V+iOptmIXSmXGOVCXq4vXadpO+VsyBhiy3An
Lnq/UN/7FLjaP/jLNWQqj1Gv2BwqJZjHSliaYoFMEvBliNxcWbsfllcwPMnEJpID
gYr/K1fRyrReONNLLAHWu71LX253Wytpx0xEMUKKK+ZBXpQoYTfBHyvuGd3wbgZB
0hEKk2tEnZwRezo1KGcFT2R1lvbRaoQrTY1vNNxUM0QDKif0xgk2X+EH0JKFE8as
c1in4p4gfqoWRrz0X3/TQA97SOvwR0pG2wlFjUt4vSaoootsxa9tGEQM4jXTWaty
916f4B37HOjVXPU/BpTISeff2vjDnZZBZKBqkR63If6JBDeVi6mHf4VRdLwX2NW7
dWq7y/zt8z6GLVZuoaqoYx2fNp784NcLK3g4PHJcAPr89J/hzhJPgi4b3SL/gmGm
enq6rweWqPdtjihd7WuF5Y3WIpU3L8p8Z5nsnmXbodYL6HGZLH+3fEMnZF0QQI51
/WYHxN9FbMOZsVe5RlduJvhsH7/JXlbfU5aDMQ5uU9aiXQGf+4oMbQlheCATGdVT
r/3XftnBW4eQ9G2fryq3+XnkFTE3avhcPxuto6C6uNZ+dSMBlMzW92zn7gFKBkhO
nA8KaozdgVQHuqqndASBekDWFlsSC52c4ph28fa544LARLdUadQnwDw7Vxrht4Y+
8raIsbGDMuqV6H6KvpvtlW+lck8JIzZyVW531Zs5Tfui7XT4DqxUhV3t1WxHsXq6
8R7G2orYbVhI1O7jSaVEnOka9wk0w9OE1hd4JazzklLs2C+pvWeZODIIZmSbXAg2
5VTzH9deqemWkLhDJFSYetG9DfHrSbCobx5Ue5U3w6s3TACJe5DaqWX1o/0fB2ST
JTz0I07caT/LYcgqksJ1UJG0zOy+19WbO82m+uh62//zTl6HVIKXTjtX8cctgHvR
jDxSg7qIfrWU0/uYGwDho8MoYwis6WFkGDl83spzGadVnfm0Pz87T6HEnOgLUBxe
ZCEv2XaatkoxjOuGIzDBTOjSTXW2NFXs4vPRi8sXLbCrfSySHqXi/JMIOVB87Eb/
4N+t9qziXUM4+MpgQTDjfP+Llv+aYLf9RJUFUsg7Zh6XOdG13Pi1tfxo71QgPv7Y
oXh6MK+atLHRg6JJuN8LnESZSLrGIJfrHP/970JhsRf/y6LL3A9R/ZQU1RXmyrfm
CWYVEf+daRWNIyvQbiIII9hmV8JVMyL/plU/id/a3t5k9V47w3hR6CApAUEOOCSm
HrqGXjGiC1bAWMBMgHNwWk8c012wTChwQ8bbikpxHCwHVxuUPLIC32SprYHPiclF
Kpwn72QGZ5kCtWvf6EXWjK8efZMYLQKh9p5EBc95SbQwrPcpyBPLl+kX9vepOF74
iLK1pNB+97Ua+kUq6SWfgMVC8YDfaHHgTpBxo365Z3OK+99nU9apbcfDdVTe31EL
4Bt3Q0GJ72C4/+mzuDbDX83d8i6jLmwpVsKf0S7dKz+a1DG50FGmOeRDCR8yCYCo
/FYOJ3snLtkrBPfLZQJVUYQQT8CMef+SVyttg6OR3m9khM9bi7CwWx+yiSNDHq+5
L1fdx7Mr1s89/rUya7nuH9Hr1kLAIRgVbs/SdLaYFfavdP9n66BLAsDCFT3Ozq1z
CEJ/RmSS6IuJ3XPbtSR3Tzxd3Yhdf+J3e1g85+2WUsGduXDxJCKYsP59ZNS43X6A
F9pSxa8l1nhRuOWHnAO/7t1BmLrvLe/nxphpJLI12vaVtVGzgxRcpw/5woLTKL1s
TQmQdYPWWQ0enmvSScAcj0vKGz/Er+8L24WMV27iwcEicOw2016XLN59AQoSbbWN
RwEyUgW1x0nhNesazXZHso5wainfZmIIgcCxHGbYGMvAz1AMv3NhwEI/JY3DSHQo
aHe+043L8bTgWXReGUM2A/5JPpiED0IsKJfG6T8XSDvK+NX0PrAYrnEDEtsMPlgT
vCg7fSwTXf93epL1y20GMXEtXPyeExqEal9BA5it2RWNPQnNVzFdFwT0oLOIL6aB
xmbk0C4R9nG19TEM+wzAGcV44EoKFU77JSoc4cHs6aD8gYamD4glDllV6QT+88Wl
x506itQ/gbnAuLZvzrRt2vT2aEr9ahAZPNSu0lNPIXFz49PooT+bizceSVAWd7i8
YNsfLKNlNCqfAk7SBp+5coQYdEO4OZC70oibgpXm5E2XewKBz2RSW53df4/EI8qA
orNb1yF4WirFQdinJC2ig4HIAGACsOsvjsTlnNP+K0Z0k7pVXHAWMmSw7gGwk9Lx
7wj+c6iaYAhyfDENquktHYdImHk7X/8XvYuOU7Zul7bHo0urBWRbNBhuvDuoWWkb
KfiE2AWsth/h2pcHmyO9elj/EsxU/mhuaNGcZlctoNHuSl4gwTx9av6oJWeyZwxh
GTXaDqKl3YnKm4Vku/LG/shp8jNyZki9ljUj46QZo1vUE1mxbEzBbl0CK8Uw9bB7
JmjsdIl1nnXBj3D3i4MtPh9PxJDwl6tboi/CNzGzdlPVjMxHTSznRa/kexANy4Mk
q5lkrBX7E5XsBW4DPMyuYBOY5exc1g6RsFlKSyfhEF3k5km0Uej2KhT8uCmEIrUY
tEWOUaxczLJBHPfNEwbrEvB/2cX/OW+xN+T6Sm50PwzTOcbou0t2XICsggCEoLiy
5HWvx+f8/tpgZE2z4+TmG+82WHNyTxITLIOb4RBeYc81Ita7oS/GfoR1n8JPv2vz
L++JnTiQi7YHmoljkBBNlfUKbvfs+g+7NHBn7sIKzr8f580WaSOzbUWhYcdwpTZy
1+uZz7Km0QrScM8muHvwLbkrLytievPLKtCXoqkzB/IqMIRj1HRLdrW5WfsqB7AN
1BeR8dsaCozabZYNj9BMnhGBHEid3QXb0XQLV2Wd1YlyqvFOviBDYcI2c/vpb24j
QNaGQ08z+J13+gmBNBmn6ZirWNoAXC+jmvpUXlAArK0RdsTUdkWpjzsxVSF++GNA
iJbQxzKG6WCJOPD/Acw2duJ52ZESveNpScpZCyZr02X5KApLLnL+o+FRUmhCW79M
XqyYm4HBjsCB3Ju7cCnnUZOpvtqNb/eFrzq3kgp4RQJIyHnIxlfB3Q/dPAxUKAxb
1l6dmrnfzi3LdOaNURTTLXjyGg6bdioSnWCmc16xCHnwroJCy27/e9a+HhZ8t9Tm
HjSf3T+R3prgZ6cIfrv8UgDI4QGGi7DWAPve9syiBUmRBFDB5MpYWRHwA0s3Pdrz
Dt0fF9QI23oBGQaN6e+wCH6sTu+63oMgZgMA15Xu8zS+Yro7bI+da7iO5AzeETlR
SkGyD6lx/QYqfO+h0iNhn1fq3b9FlnK0T5rOpU19ps1BOKynN03iuyaT3jBwHdMY
n98GLEU96GUCHnhcmsUwygNz0C9liR4KdQwSZZ2twYZqmq498DMlditysE5uNoA2
ncr02tu5bDgXcidoI3T7ZmJb80zh7vcDrzGcd/eAkXk+/Ky1lYVF+qzYmgLdPo67
xfdQtmDQq/jFxD7eeSbm0D1rIDu75insBv1UM1RrQt5Ghhl9pspDVzJzCRJS34AT
JmadSdqpriyppzODrmogNiUeZv4jpCmJzS6JU8x3KpnRqd3d+AuP5GnyTuaYZIQ+
MKg09fsFAAe/d6XKKebs2sbR9nusOZl6jZ3rOX9uAyy0ykkbZPao4VqoRwggsDeh
T72wWOXBUV52gNti2OAUE5ZjLg8ycRzEo+i9tD74/crCDZPw43YUhuMJY2vFkiXb
BhSnwnDuV+c3oheasPzWFD/9uQ1FBgJg/QVdFEgtsFEDrrRfa1D4fZqZkrnXyARe
2evBDEcxT4WJMYN0o85Ox+3o1+Nki/H72pqz5B5d4xdt9RBVlHHmD4ozrg4AGC3D
M/kStM3Uzhu+tUcwLM616mVFDUohvIl8y1UoKZelubPiQ0es7F6sYd4iN423JmW9
o92YZxr9dXRgkpUzjBEKA8QSDsi4WbRT5sJMtAPodpcTJ6sfEd9QnXUd4ejMXaQv
BP9aeK6/FEV6aWjMIYItoT+RrJPlVMsyV/sH8JtvfLAeF5wUVFTqdWprdpF3rvTu
szloObrMIDKREx2+ZGVU+syQt4TvSQGOMXkYWFbUUPTMf3LWS0jYgkms9061CNl9
8WXNIQz0BFw9NXgdaU7zkuYKuM/FDJMVyj66pqbE/QbS0+4P85GRlGZMpBTGq+06
/680tvPg0ScEptrSH96CwCP2hoyMfC1XooN+KRHse28j9mwy2KzFnBJEKJkFq9lU
ibYiQ6Djc2qIQc58GRV2keE5VOOadrXNDK5iEP68aI78Vt0IBrGmhgpOx2uw+bsr
l8b0GOXQyg/ZYwCAWfntIo8Vge3Tu7FitPyX98yqjuVGSB7/MsPKY+u0MSgHQDt7
THR1GmerdwBiziDq92i5w2sNyLj8woibiEbvZHJl9K0Tt5xAHOc3JZsn6ID/RWt6
yaRXfzYcCHjSh8YDyBo0cz8hndcSvne2HMu7degWDUPXQtTp/j/fVbBAJcN4lc/+
DnGAZ3Nsk8oAODCeZTm0o567H939EWTpM/WcdVtsv+8375mNtDcEzxjsgPQ9JqPW
pjLonS+oF18g/4aIudETUCuMryVJvFMzEiz5nAs4GTkn0P96MRw90JBwFeSow9v+
GilsCRfcd2JORWGne/jxsDZEOAeqPiyWad14pKuE2R53vIzzMQeT4Uesnq7Tvt9L
JDxjDBKqvKms78MYlvT1fPDRHJSW4XhaaRebbFg+j6tel6nz8DA1aPVamfAQqk8o
t6uXaXFY5yUxGPjBWMQTTTRHcWrWIZv3xHOpnkDuAIOCLmpAQcJ68BCb6zY5zLT4
3Mw8fzrg74Ip50RgBQnlNxzQWCXwfdEP5eR/Xb5Ob/p4/JXzC1SBCzPs8i+MfqlB
9A/BKqVzuN2o0FH1/tKHWU/rKy+0UxNhbyybZlTnJSMPF0YOhV0wlnQul8AHjRj9
8rUpBMBjG6Rvk3DeUuwYrIHxexc0FnSm2oxJSNATBaM+G3tHcp9qAHjIqMKZcpP1
QtdU4I64JfErtSaD9rO4JgilvJDcqpWBOi/nb2DYb8SUeopsGTh4nEuYH9RW+YLN
k2KzlQUiWkTDczECm/piV+RCTjKernTN0fR1P9MFml5YzUsIPO8l/7BThlkZplMz
OMT/49AKBhZpTTJdwSf0jFrR4WV6m/bI1oQmtBBtCb5/NA4bDU1G7g3HOpagy7vF
+651Y2trKYFCBG9bj1uaTvB2FupS5oGx3s7tUAOLrwXPorHwSLkeY8DN8TcpbeT3
EeUXP1vAJ4KUzTEtI25fpA==
--pragma protect end_data_block
--pragma protect digest_block
f6EV4pleBNl6OMhqXYYA5hklMhg=
--pragma protect end_digest_block
--pragma protect end_protected
