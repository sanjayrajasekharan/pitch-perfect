-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
KIZgcQpGyMhooe394dKiK8gkDhPRCkq5xJLfgQoV04l9s170vSDHzsKgLUVOTvom
UF4ZWLTns+ONunJmGPg4vVEut7aE2nvVHSSLiAv82K0xkUa+pRisEEO8eOXID6qa
w63x7b7UEl/KJC/l6wyRX4lwCWF4RGjNSaf3PkmQaXk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6314)

`protect DATA_BLOCK
7KwYG6J8ax4q99i7qZgMvZugDKwV/E+0qKgMXLV+5YpAgCof534kkFZmBWLpcaoc
c+gEklkC5d8twW/l3M7pcNzqZTGA44t+AktZxnXgCoBKe54hXRNagnnEwPwL/bl4
wxeM6G/ARmD4JsjkRBXVP6o2F3uuwLpSAiWOt/gcGNQYNzOcKmje5njCSl/g76nP
JdT91KBZ34YC0FRqwS+3QB5REmBFEao0ntFycwYBClQvMDLxvpg06JKaFunled8C
JHmK6bRIFE+pxb9+1V/bEOsS5u6vL3nKPJMXwiHfFzvIFGrt06Zt/NlkLF+jCspI
LuSKyqoCJQk5cl0kkRa57FJKAI6TRxvOcZhTAWd51/RAmXr4LvJkuN9F2eM110Tr
Ir5zK7uzymYdslFYuoyN1qJ+dFewnH+OGmCP4qM0mTTeT32ga8WPG+UBjpKhWrIK
KabJIqHWOWQ4zBb8yPZL7ZdnAnw0h493UyHRYrRwqm1zyKZXA1nBDIwzgnXze0Ti
FJj4KobOyaCeGrriZiVD4uV5wkVueJ+sX8pH5bQdFFcyo4uyY4VClE6S/zJem71N
2KMAb8D20CJ9XHqhyxlT2GfidphX4EmPyQTcFU1xxYqjlP36IovQg4Q3aTRDUowS
VL20tmxImW5Gt3owqTy7O7SkXfEMqxtTMVKzS57l4EA9gIB263QBwtDTFjajJ+GJ
zQgazeJrwdCxQK4aaLSbinWSl65wE4/zzqJ+wRxW5aja05peQrSKpzvUQ11NbL3Q
Kin01cEPzxab6uNQY0yKVHo9rujBuznD4w6vaDN3CCyRfE5d9iJIm8aXsVae85IG
AO4thz7MmNDMVt9a4LKkIQUntkfDqx8WQ+QA6tL5y/JGyV57lWLEhKulErvdiPWo
pW8HjO8t6B4sWCbibAZOIKxSwSxwqGHaJ695Nj09sBkCXxNv+eRG0iY5xOgEB4Et
QqL85haED2LpQl4sj1w79cse75BS5NSeTc+FYQ7kl0IZxm1tnljDJxIp0P3d66e+
6fYbBcEOvheLaT9GURGmMcn3RHrjKmgPyVPpaWTcG7WJ2smqmyFyVcKNAnpVAMU1
Se59x4pbKCh24DDM3rl91zf+aMknhCr2j7Y2I5ejHil9uLsZFsIp+Yj+GLbQENby
6+oq3G8d+ECPK+0JSAedrab680sS1t2r9L4pNNWuhhIl8xVy4SsQ2OeVOyg5fbEM
y4xb+d15eigr7quEz7CZ/pqGF7HOnY1SCx0zKZOSQWSEAjpT/qpe8oUKOV8LLHcP
MsXc6RPtgkMmxxsmajmiJ/z/27wZOTjyAfQiAfqfiHUvwhztTUIVSLpPFRM56MCR
41NdQ6AkxztlQdGsY+f4N2yTAl2uRlX9iGQsN7cxM0IpnhMqfI4GJIAZj4uIvPCQ
59kxqe1pDHz3OEGoCC2Pq7R3fc/tOj+GTuWNw2g9a2GmSphHfrpomCy1L6E8Ap2X
LfmE7Uu9dAjWeotwgJ5DQWfowa332Fp+AhN2pPgo8jyY+0G/EwWRoNhWVs8t4pD3
Rz6Zgdib9w6xStmfTtBYEGO27nKe6skL13d+oJlPM6sLdBf375Sn+dL34blAS8mL
7PFJryA0NhYeNbwkzVxAfAFkzLcnULzCkv5PPyTdx4NqPiZkK1eZZ+FZxaKqslB+
BERZR+hTwrg0yre7VWNWd35QMnDeT1tA6xjvib1cGDSPCs5jCHVhnVwzx/iFkUAa
NJFvrLu0lhP0IV7Zj8ijI37eRr55LvfT/eK6H2nCN/PGeG7jj8zSYRynyd4dtnhI
Q0o64OBNOS9QLgAlMAahZcb9jROoNW5wkWFZ7se8jN38rXpqx9mpzpiUdXZGISZ9
GkH5DdLFTu3S0dsivNhkUSGZw3NxJVAKLjAhr4d1aeysJpC8GHorqvICNyk9i2id
Qc2QpSiMgFxES//EwNOhKP6Kh452rS59hcV1/NSGM9qBe3tE60FOEJ8dEz5H8igp
BRy8Ap/1V5VSwUGk0EGbJuuP3/U7S/cWh/s/4S5uPQhXy9RDG0sr9nqx7nLFb3No
aK4GUBsmizq2Y02s6F7GaygrPobWC95mP8kGNn+j+vOIUPriw8B7CRnXb8npGTd8
RrSlHb2vbQAKoTX+6hBOPagWFuVyxD6TKUDBbBSAusU/ZlOCjPuPwN68N84NmY89
AmS7b7NpAImg7/uoAT035aGAXscqHyYXsMd2T3TfDzKpKApm6KHl7qzlxO6oCeL2
7sVl999y98NM0BZz5krNcqpvn3x1knfSukEJ9xLsTzgsCox2hGTh7h4ibYJTCT0k
VAAq3dw4lbD8Nzg8XYns//cFYD/ebJFYbjbkHyUxKQylr1dqJJ3YBvWx2RUNwl5v
VsjqwvSUtT4QAQLZoR6sHjGtb0wJWs/0HNTkbehXENLlgAqqUivAN6C0L6zvySkN
5oP/JqsMFOSvy01QgPsRrDYe6XmeJRNcTBdk1Bc8/cERYwc91cQf/ICqO1LgjVFw
9kTh1UmZQ6VQKM6D7TBuMK1LR/JTRSnzltAw+2vGItQm2hWa9lbjgZAD6tp6zBDl
noij+8EG03r2TcEPA1QLI0OMmauDMUWYRYZ8zKPaI6yHoN8u6vGLYaTR7MRTS6r7
UGYXHv0hbCnEEWa2mB3oH4ko7D1h4XudyNz9JHLpCDBr+wGhGx59VCFSH5sV+44F
rZdaEoBldOwJokS7mLp7mrWi3v/IIJ6zTaK55wZSa+630QNQNOcY7+yIXVsxpLR0
nnLTNNd0sTwQih7EkheY3zQNX7xwmj+M0NhK4gKcoUoreLVPaWGaT7PD7ewPLEPn
xkvbbnHc136UcBzuuTHrjIWyOqc8Hv+5ZJa0G9lpafzA3ozOFuBZdrCMhirm/D5G
t3o0/mmwHgEtMrfMCVobTerqpaPihnL/b+iFr/p860du3cKTBVJIyPEo+RqIvxur
whsiKy0ktSG47NaO3P4Cw3rrE1dB4nlCnS0vM7rWeypcvdmoxUAStTDt8c+TyNP1
g8gDDEuGSS85KYl3mIcdgz9WWIXbH8cDfDhGjucncKVukslVYwa2mH9urrrER06O
DkwuvW7K1Ic1aRZDiKQCoyviyO6p71460nqur9tkrip/jdM+mZjrlMhUg90896xg
0mYuCpyemWIo0P4IRBWgd+HUHXfEQWzOZwJY5luytf14RaV8V/TqEb/kvFvWe1pl
GJJ4711YNy5NopYQ7nLd/NyDAhoIrA1SWrKA8D8tLWPFo8Szr+zvQ6DSI+c5Xm5k
K4jOxzELl64hkfVGPFYLmXtr0nnHt81S4oaK8OMlht0gEo2vBF1/ct/qtAJLMtgm
q0e+oj5thhMX/GAF9aRv5sO/Mrjc/zI47Ra3V3Xl3SnkBE7Vw36och762ltjqzMB
Ru3U00ex2M7xJN+lXVGM/Fhb5LdiV8iL9iLmwmlaNknH/T244YomCXBJsJatEVHI
b1X8W6eieqjJBXQauqFG3xtiEurgbweXFStrQY16Vv1xlz2Z1DUW+BRpRdHRmSbG
C9iYhfHnWzWGtH6DjjNKJsectkjR5wNl3miIPkiRU1XaGjOXvyhGhGyJjh2ymJe1
+K6/sCFXAqFvgTUtkDa+QoD3ychatPSDX387ODD/W04M/iqXYn88yscb+434oo10
xlRpNJ2jBzlNP2ioLXFj+lVVg0kT48pkAudWih0NEVpafQX7sesjOWHOTl5QbnWw
Rb8pTYavqvEmqLXhqiFRoVB1dapLO/J/9tcK4CATQ2wSsrYFfI+q4WVI6jmvmCGI
GJ94QbUO7mCWkoIJRT9K7WgHwC2QT4cJgYgiU1K3vgVQzqxUoto5GfZCDIFAtH0C
a5mIRmGKce/4kNTZoDNS4RkxO7u8lQFiSgJk0nbwHlQFOHkvP7GgsAQlmpsJOVri
K+SuElJJR2zOS0sSHSjpl8QpDHLpyc1wCPIRof0o5E/2+iE5zePaDjcO/0ddYern
QonOkatKYy6TGVZ4cf6oJxCmMDvUTMd1dtnxnNXYeRHzLZw/lBXLrjd8Mt6gAqzW
iw8SgFlda/KVMqWaj8+maSAQtVzx9y/HMOGQLS4GYqCnxruifF0xx5KpP5CTR7jX
lnM7/bw9f76ij3fi4UFCWkiWqRzfwGKZBILJqOvEkTbKJq5jxW+G//bQ2VC5UfCT
0zrFJZ7az1R+9d7+E/NcytYkqIOnHP3e4hkKmA43csL0HAn6MhbzNOKyP8ZgzM34
V6Gmi0C3rwT/o/eCYNXs+WvO1oR96DW2Hl05ufZyIbLXuYFXBWclvOfoT5CjOTm3
9SzVgkmsvLAf4H8arLumzkT6BMVQEF7Qc4TjvisQmyLiLqSIjA5xE1Sv8e3F+Fpk
qZ+96Ww1cYlnvKnk5gx2Sq6gI430lNdF5dKyY/Fk+5ZoGlj4gFLVOcM1ogsAllVK
GaDzQ783odidm74v7dG7l4EUxhRi8MiUl4R3koq33nt7Cy7Dhj9sRZx6LII+uOds
aq5RJESDrZsQVIDswwGXXzPDzqj/9UgNwNUONkG4TDD9h/fATKwIcqLV1bXIarXS
9pSTm6rt1vzqQBBlCUDaJ9XYadmmrMoet8oF0/q66Xk2iC5hd9XwJFWvDgyQP5sE
hGzY2JDH7hdGQHgLlFeNm9YpfUhrB68o+5+8dNtcqMMcBXIE6ea7KobibWLZcFg8
boJBuW7DAEYrWxyA0BNDg8g2yJLNtd3mFgYVDb7OU+MSmIcpH6/M9WHlTmt/Ukms
EIvhGQgaBbPduofviayt8U32tJXgRfQZXkZ8cPMlcOk7uLovaqKsU5h8QHdd2rr5
c1pj8bxSpmcuryLb7Gfw6l2yM3TEHezBU5kaPjJLC6SjuFv2jQ5aboprvEGfG2Sf
mhscAVAR/NVjtn7OTXyoZdSqRgoOhgaZzuMFr4UytTv8Bg6mIWS4L2vsgYS8eqOx
DTOuqh4CWEZNHX2Dsrf5K4dhNut79RcuYa2cQKaDqVelr3WnX+UE+O3nAV9ZoQM+
/GGUSm1waGsI1KLo1tMmDRNK0j9xKKPElgVyzRowlfDqHyAKSiJxAOKw6qb/R95b
rROl8TxX++GctOdLXNkzEmpl0ZCP2LumSdUMZQHybIasVfotlMR49sfp6rAw3mK3
1aB/JnqscWPUofOKMpCbYZJJqCdskWU+WeYVAvnDGGuY5KOQMu+05DvcTcSP5nzk
h37PA2GPBW1Any+PL7n5Ilk3i5f/I/GojDdDeW6Fn4O1F6uXoVX+ntOVr4sg4K5A
r2l4stoymZZ+y5AuGJXWS7EI0ENJmEYnqN/Qkm1mlVOGVAMOa6/OX/BSR/DQoKXg
/VphI9po5RWLarbtdpDEeCJPcoOn7x7JQRluBtJ8QsDlLl4kRIt8ZdO4JAAe4h6X
ZBZd98gGFXxfiefjJYF/i7t2E3DDOqWqP2MfIzNLpvkhp5MwQebmV6y7/MgyYFFO
29UhOVHGXevifRdFqcfosNsCmTHi/5YibOiKmYQiYLWdl7r2iPuwhVMHOZZX3Y5/
V28st0VKQBJJ3weeCQs60Kq1GVKRURWk/APzQSdP6q5iEce8WfrrJF21S696SxKk
0kR8USPTuflFkOBjqPaNynV1ci8Wny23LMoBwqgG0IjpKJWxUpzG4CtS8km+2OIk
RMapnub6DBSrGU//Cx/yBsPxz9I61ELIKpauI5aEP385K/IJf3JjayZpPuOr20y6
Y0NNwgpW1eLPBWi478rO/+srwN/aheHKSygynEFT8Xf5f706vwaZ23sUrPxcDC+a
KxlsHwKsfrwd5hQt/RzAyvmV9l53weZh3BBjc+Mk1EMvAn/LKtDYmp7rq2QZj2pC
/doZDvkFDoS+EDwU0LnwX6YkNph2ii9Yor4RtOW4G7XqQlpvFGIBf3DrtqG2FIyQ
OAm3f+GykgOYqBtnnGaQLOCspcNbCmFJB22ZN6+VDyeWVk3LYaSESqnPwd0ft62C
Q7V9tZ4VHf4vC7+IN30Bg9HeU5O1SVvmItWjKmQLYzb8XW5GFDapvqJsJwXa2VIb
ouJwrRoMXXmgdgZX54GevcpRiY6WkGFK02hMZtuAabqzPC7vopMhtu9r1s0QLw6M
QZ7yYgBjPLBQx9BGTmS1goWGte53jrNDpgZdrYd6kvEr+n3Fir/Y26MQnjjNPlSj
ojpWh1c1jBP7djPBl8aevNlWGG8kl+pF2fjtad3GAofH+Bi2U/NBjaolEgf+f///
1vTQjUHIF5DeUNccb/RroVd9Iv3igwmTJT4JpuKklS6P+CJeUU6gHV53dR7dfel2
xOS6nXVyZa4FLkqYOm4+jMMZWR4ts+ceLKB5eZ6hCb0r2e8YydwpjvQkY0hwla0r
WnEbQm4T7OlkTQlgKjnYVgHwHC/kJAOtOK9haVW8Rv3I/vdPpIfbxoVDypVzEyiq
IcAH30XaXpZQ8utQx/VLpxPNKKafivhhcSfCGGGP4QTFMRwFu/S0DFbPj8oVSDIn
HIVmb2Si4e36ngS1aqftjeOGwE4/iPdLupNKJicRCr7eLZ9pprKtuKa2on13NEv7
H1yGuMTE5cfODqUN3mMe1EbzPSElTbpyribIq1GUxmgmrRcV2pN03wL8s1KsG2c/
3oqnxW9NJQq6Z0KbKw5NEsT0IPPmhbyaPaLbBHCX73F7KTkup4y9zEiWWgBQ/cD7
Q9e5X75a8qpmLd8nzsR/Sz1Bl8lb8uqg4iEjQrAfNGPRbvqC27fJutC35DIk9R3a
d/Jz25iF/dZe63M03MgHgaKwE06X2lkxa4gimRbD2igvM5ms5tT8BH7amH/HvnAw
HgzokZLAzzvw7VWnj1UbTqA9FbYquAWOXYnpEaM1tXWrC8BHEYwKc63KO842AmVl
F2htiIL0iOv70fVC48muZK/1NqUJq1EwGpeFkzVPJrulRIrsUQXksWekUp9BlVeI
6CRX9EmoXVwkEtvfVueIFsLMh8t6H2qLw2tmlQ3hCY2S/nkCREwPIKWOqEhKDYEP
HK8LZl4uXxBTusN1OD5o+7f6h1iNKXoZ3TbvNUVpKSt/BS0sxuvPLtttkeTYv5nv
K+u3ycumxDlxdx35EJ24AuvWXv5z35/auIT5f2ZzhYuD91B5i/VZvL9gA62CnVAe
b9WRgR87bQq+4FMtAZJRpES4zlxEbbnMSN+g+rNbMlZxc183zYdjSOyCG2xySJdX
ZvHyAxABqofctChaRis2ExB4Br3pF5xu1RYxnSgO6eBc1vWXdjmDd2ajgbZIBlDG
5uA9v0D2Lt2GC6OYa4iJ99kJSUa7a3JkD4jhvC7dJNipNbCnBta/q7lt3wr057Ub
eabTayJ0dLAnd6H6/41HLbDmqSHvDM+tbgZeVA2TYSBLXqeo7ERvf6QsUqtGZT/Q
picx+rJK6UCPbt/dAQs6U25pXSyn62LZ3TK/ZZgY0I6u00AxoX/3Hb6rDsmYzsK8
/FZnsPsJrK1GiZb5i7jkZ+mpgfzDKNAY/HY9xHDVt1pGjQMxzsBc9U+ickb+n+M4
95LGlgM+IA20xDbw7EO59FVmN6Te/zTqJZsBMJEdWSidfg92HyU5T0G0z23hUmW/
/p9N06Pft1dIqSE3QYcgTNlL81EPo+/9HHU2UdISryN/+h44AM+dAr6FUHuXxnel
aYVJQBJ3nJ4c2kHzmyUT9cG0/aFxF1TVDHAVNiUpIQHuUqquJMM64Ws738sQmrrA
EpTik5MOkwV0I8rxudu+PzdQsf7YOqnJyiykIPRU2DK/tLEmcC2aFb5DZX40miCh
II/KwhDRwvdDhWpNHdYBBkkuCFXeKvW/d1krLGTdC2klmtulPD2PlnQ2wmwu/2hM
pryf3rNoDHBfW9XvMnr/yj14OSsRQoerPDhWlUVTWhUw2BUoXlyz9VVgIz41hUTK
sVVemLQDP/XM2MKiS21nc6AGqa+R4K20Nmac66QhiASAKbo6fdPal1UkcPsyVWMZ
EuRozgv4X4+UZIs06PAbHhiet9U7EPAiV2TKEyQJOV/iXg2pB3Pr1SeALBmff8UB
NdTmijH4Rpi7cNeTh5SkoE3hsxukGEWwJsx+4oPeHUXAEjhtFdwa1shE8zko/HKW
fUcehaghhUCB8/FXEu93fK7GLBJcbST6cLJItoVsu8XGQrHeG9UnQVFR/GaczmFn
B1Iy2ytWT6iuctjbgxYEhpYlov5VPsmOx07Q8vkSPZcpu5IL/uyNfFTV/+j/XLvl
va+JDleLfUM9QXCHU8tQztbVJnGeTkAujyODP2bzvCK+FyhGewHUoAO8xl5C4TnK
H7hsLJEEbGD7ihiJZkYumjBP5/aziCFxaVy3dkuqO8HULxdatMi/x78XjlusqDsF
2VzUdxpfQHNuKtJPFwIKpVdGhzUkmG3qPCBgR+aoi8xTTpXZRvd8VRhZNaDsLBYs
UU5o++xxxcVSW/lZDNEBQ9L06ZmeKIrHFR3Uk0pyGJ3hnS8RBoJznY02PGUuAAqh
`protect END_PROTECTED