-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BWcZCYR5/VJX0jP+boTqkeQ++ZZnfO5dFTzrUZqfaMc7zDAMxWw3Z2VIgXvvXEPTzzXWPTjprTo5
etuIcRUa2h3bkOjIRuAp+wggdLCE9FUHZ52YCYMreMkTEJuDwNtqOXVcaX/7MlmbhKlGjWUk4J9A
RTYohespUHT9dpY5GhxC1AU05W9ZW/vTaVkMNVQ2l/f0TGlLvBt9GD9cFWO1xEIUuZDCsizlh4rE
7UfvxLp4vATtd4RaQKUeV7gJeeHHvsgA1tCo1g8TIJJbmJuUt7fdrNoxfkD82U50bwshNfJ7oXCq
ESdQmPx04HALedJkhFdPCn0QYxSyu+zmYukehg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
FnP6SipWmyF2teOAlhpJmwqJaZTXQG3FhBEt6q+frJD6QOo9m5gQrIi2QrvmSxZqhAcYkxqsrgNs
MFPljV+6i/uvqnjcYSp3tDjscm2qLzcSmQ+hSrsBEQHZpwP8PKx0NBMX1W7ZIsrq6Tx0msvuFtX7
MekrTbSBfR+7Z0sD3u3DBIo0wkV0h4zdpb4UrAFV9ArY2yYaUmexzUIBGGs42UsRBQ/WXNFdp0SL
CWrMcU4qj9z4l7S3NbCDJIvrBkhHcCtObxekbOvshyy23VHhYMP/A3XYyqD81KTa0MVbh0dBszE0
cuXl4HZQKGpHUq+IqXHvxG1WVCXT2AWrPS3akWbDtFK4fYwvQpkBIVHKzJRyEF0McGQGOwFK3ymk
JlNCU9aBl1Kz0oUjQvU6K01mcSsHU9adPRXommvkNFf+fQMhJP/mjg2aB0rb8Lv49tnHqnSZOZNI
whHwsaP6uc4FqBWz9/S8NKevrmV21a1mZ7O+4YyqdY3UtlDf31MrR8OhgjC52TouovaQgPMDzmJp
khVwSZXUyvNTznlMo+cAkUwWN6QlXczYZf7f+o+VBEat9Om7nLMSeBOo+pOb85kYjCxvfLlOQiRX
ewJhvExhTBzkGK/klGaSzwCdmH1ZyEAdTdqzwGJGkZp9nun0Xo0EYqSJCiRW+qv5mdWx8OzgOOP0
gTC2Oi16pOQ7ID5BE1tlcfRz0tmfD4tMs09tFnEccyp7QlfQDaJAi34YB4i+eFnUhu0f6xCnW96s
w/Bed7y1+cN4j1lBbVEMds6VY6YfT3ufHZhjOhdK2F+cuFUmnrE7XIXBy8luD2jP0qrE7Adt6huR
qRUCzOwK0Fx2e2wwGHIxiYwXi0tDRqS9iv8zWSe2ajLUmsC/lVpGqQtWZ//6eyLX+rT821JEJgEp
0fP9rw/gKXpKp7KFGG3WucIj5ffYMlpI/thoqydIb/PWmbpHnt47wOTWio1npMF+jsllV3AgRVKg
W3NfkmHiArzWryjPpQ2UTqZqi5MI7/pBqj8/sPHsgxpuiNAtMEhCG17w3BIyapNZeuUoQKbWLm1B
hmSYg2xmW5etjW++Tkhy5kD5UxUWDyVkF7SeHpaCZKN1TNPk65DS710Cq54yA6ggZdhQ0kK9hOF5
n61Y7rib3uEGNbvtU1hXDMHWOtIqM5OIsPU0UgVQ46lOcN6N/Bv9i7izilXR9cyi+UuYu2TbD6W8
US5ExmKPS4pzoXo42Os3SfoSHyrKVPWZYUAlMLJA4IpN4we6ymOSv8qtwZuHG0uFFnVZ6UKPGB0H
CKEANgWGE28TAeJyveHSC1vXdA5Ej9mToILmLWVJ7YdJpBkP3cWx9sIaPznc8ymERIAAODOaxUd2
9njLzcxNJmgpVX7lrYx7htxTZ0CYD7KC+VS2umUyqS9M/Pg+mcRI0G/c6H5S6jK4qH9ce/SWt2dG
kYsVmEzsqT37U8QSOSHwPBJCE93NutjNyECoHtJy8WetMy5J1J8F6W/vL9vLNJWLPnQ7iVqrVm74
lHxyDqnBNDuRONRVdyTh/KmAIIKiraNb9pwgafNFAMDoG9o1Zo2+HbaUJZWdXfUwE4h4b4Io/7k2
UhtCfSQU8lDuR5tJdPthNbEAjn6Awvd/tejTaQSpF13hJ3NqIz+Bw/+5MB0YGyh0xrinI4x22QaQ
4Ne25g2WgahGnj0gHmKtu974yAB3WC5uN3WFhemx+C3EEjrc6ZOVKmZlOapu1FG3MXSE6JOXa7EJ
lVkVnfGcdXxWrwZ4GfTe/t0KDcxsjwLyz1qeazVLxzVlTO/RR9Ow2YXVZd7KjlwpfletWIbO6tLP
AZWOcXuyxGWYFpjUOBcTnpMqx3j5Im4cZKqiyVefEHjHAU8B843A6oBjLWdfbJJf4EBskCgO0D3n
KUwEke0oIc4WgebKQv5Eqv9MiEvhcGA05j8EULSKd+pa9ypCeTiG46g4UmUB0yKRrOzHe171mE4Y
Jj8gcpWrFyWn8eBi3WidrIifG9lpFlROjNWXyqVjz6+JrE9If+QYs9lAGM44sAOIRpVVAfCnpTEM
Gswv0LIbCLZWHdvyW6KFY2wMGea29Qrk7SjeMW+FeB/xYgPgHu+3GBdYx8fn0vN4A8/5p61qYigb
vbs54A/g/nnLhdlH9YcTPCXRO6GFcSsC6dJe4GRHyV0wNnwMFT2SuBwsT8ixIP/QotboKJiPlhM/
0r21a0reUAym9DjTD6Q2lTOhXyDrEi9nxBxX086kzDToaARZYi5vVc+189biN1W7t4DJKjfGVkkS
j9gQi65u6t5MFtaTT28DHSrgNlLf2GhlQ+rm9VZlESftNgREmuW7xBovmZhfSAppE5nOiFwSWlfA
O43KLmvmTPZuh2vrt4N02RsQBeruo5s6bMCnh4x6jXMN9hZwikSEcrEMLnU7wT0946/+KIaO1frS
lMbn1VqfoSH9S9jsb78vg2QihSai4QjZzWHrCd4cskQML2LirkE3omOjjvOTdZaDQTyQVIT9LACm
1mqr0XGYa5aSlY9jqKUhS1lVakMGwrY6GP8n5kkjhTSO/7bWpTjaJ6xcoMc8i5DLKeLkWA6pP6RS
ZfogyHChm9vYdEpJAeQsFOhHB1D1w0vaE6aF7QpBcVIlBo6dyt0WR9ZFWNScjTQVceSE+cqCehMV
kLJVd6Dv0iDiHeXo/RmrqfKVAJscI7pkJQDagLofl3VbI7e+WUMR22IPANyR4vm3XKLQ1+RmD1TJ
LUzIxjNmqPlFVTUuY2QIswZAw5Hx1ij9QulsxrdgqsYFPK/dcO576ijytqHjeCffXabEbZFDer3J
hQ9I8O3XiKn5bR5J2MxdB27G47vSONN5+ifQB23GGxTHEhWNGlDRJSIz5j0uwgc8BCNbFxmCKkf/
qdDlxR9D5YocgvKjy4F65B31KHQAlA3ouECbH+RZd+31gS1oWcqOerdCxnNnHkJzR7oH8Ac229aL
QY0eC/KBUE3qIZNfetjCCfeiRqFjDi/CwyvQe/aPRZ9CY2MLx0wbJI58KkWUDcBNOZlXg2DhT0hP
nvPVggLYje4ZCJorGv/FAyv+ZSp+ohHcxbsSg7QCljumKZZhrrWHAqv4pfOmJtjYVmPs3g3jR/mI
qBcVw5S9vhSRXjh/DZp61pf9mrm3llrETI5+Cm11g90YPv/nWGyHX4O99BQjHxtTfi0h7hOmtjCi
ufh+QrKIVnxdD1jotTdECHHcgxwAfXrMR0T/T0J4ZSw4wxUEPVBYHmhh4ZlUbqAIBJUtQM/Z4/eD
NYOc72V5NeJfwF3XqVnM4RZFOjc0BG/1M2/OUGusWRQmEhUI2DGj1JC9D/dBMZkPyq1yJNjPXYbw
EQ4IUpCBaLXl7/TKUnba9MmGNyD/yNvx3DTi4jzFKJR313w9+CWCNRXks/upSrm16wRYFGFCeEen
bdSVftGERKWGzq/iyKis33B9TjaH46J30pEUDKErOFVvsvjRBwfaKnWpqekdB8ycX4d9lOMj74oR
sz0HI/Msz5TJ6+kin/hZxWBupnA2UFKzt4Ww/SLIZ0L/mDuXNsLYEHlMZGSfo/iHzDEP7HItG2Lx
iyJDmq7C2Sw8JgY+GxzBA5jgljZEs/EAYIgw7lVOVOABHlOL/CYU3HEkS/3cSBfww0gVHrVW1Hc2
fNkwiFThKZFcnaz03sqGb2IySd/VhHccXuFuNLcnzW9WakAz1FVvN9xn4a0CluopC9FGO0t27ANK
ZOJBbQnt1IvD3vteu7SiNllq12UdjqNvFimnUeTlhn85DUvTo8H8HQQaydOhxN4eOBDqZl2SHiz6
RGWAG4e7/CP3BH41ZKhfs32CFcfNiSZLXZFaC93N2zrdj0pw2ATHPeDURN5RFOIpewZBXdSHTbie
3SkJ2f8F1wpT7u4Q3pe8i1+aIhzC7ZQ9R0uq4/62OjWt3r4E/2lAmONC0ort8pLioGKNFgU49qqy
feMqX37z6TamRgsN7MLP8tqDcbkJ9ajZ+JeSZ3iR+NBo1bHgzCpSTJ8gtqFKIWqq6cYH0wQCRN34
FwsH4LCIjNfnRJzQx0oweLhOFtXABbpnYFQAUKZE3JyhxVyce9VxQ+isx+c2metxVhu00l9yjn9T
9QLnI7EUXMxabcn3Lrp4AUISDtJuEzi/Fdx2JkMnM41SRCkfe38O1xqSjrKvQOYYf2ReLnfqqTku
RT5xJ86VLr9Ltnd9d2phYpQvT11azSf5GnaNfTzvL7xhmuKL8awuksy6ruODNgsSa+BbYsUr53lc
mvzWVDnG0JpEi38ojnINJXWjmmb+KdsyRgvsjscBh3MUFrk8HR32G5/iSwyp2ByZJW//9B0BNP9C
zsfJAV8E0JHkie2EeVjPxM9cC6pgE9sywJxWLLhixZdB+HTDGBDP1TFwrgJMKwK5jvf+jprMyZV3
H5sIP8iMCjQ+EqUEMAUZmHkGAOCp4brsp/6WIX3HxZtFF9KBIMPZC5TztKCCqtIskfqQwsomEyl3
8AAUU9vE4BC0vlNGO7bFMegyIrRgrMnXEPJTZTJFY8+Vdin3Pd7ytKnByM4R0QbKnv/NCn6LRkcZ
7/YKx+JE3/IKQpDA389/+LQB0B93K2nSGJhilfnmrL5gg+gNphcsP0ystM9k04SxYX4KZ5fHiGV1
TqOM4oSagYs6aAXQ9QRJ0U4JTRyiVELoCJQc8MW0NMp1Wpvldv4mSSfMYKaeGg+1f2aOVJUD7zsr
cSVRExKFvXVLEEKNAve1aVdL8l2BePajrt4o3VU+6Ls2B+hcdgWhoUzwyLWTZD5DhUKscy5JB0m1
ovYzaLuZyJzGWzscJn3KpjDdcg/NrU95VvCvgN4MYZDDYTrRxPby8HhatxkVxZoHXTgMsLwLrd9O
+OZ9QsXO37aEIKOBMTmN2nND56wgKt/ixPdbdCQemY+SoMDooqnS/i2ZHWKtjodZXEraOV0uMwym
CgCBbWPGwUH1ppUYYpNf2d8K3bJCreGsvYQmX7dFfeUFLV6K7TI34dRVIMpDI/oFS0pTJ3XE2cUI
2Yc5TBhc7/+MinDekv0yiCFP0i/Q9ez92/Y4nO3bFG7zXmJuniFFVe685LHhd/FZn1WpxpNEdWqp
spXVWY6X0WD1V+Tt8XJ/845jno67DmhbSzMB4GgndUmMmxTn/HtcRijubfMopUfrebIIDPg/kbZD
yo27CnrGSE/y4J0Y2hqXPCgTNdKtFbi9YqIrcvjylq6WzXOYh6Lp7x7Sec3mbFfj60519IoViHfP
IB7yVOHO7Q6mLeoNFqzOZNR6wjiwlkbEqLQzLgMFGs+MNMZ90qNyPld+kvl4WykVNlMdJ1fIP6Y+
b+oev6V8EXmI2gV513AwjhIUKUvPssFixkt3uiuWXs+eyuyNYeeXWYUdaG85Q+gNxtr6roha1nM8
QzHWPdE7lQqY5spVlqVmNNrSfvJ5T9AJH8LkGNFh1I2U29+kdJAUmcksuc88VI4QnlF93v5Y6/M1
vCv7ZsgWF5PnbAJeFvJMDwxCZqw8J+8BEO+w15lVcYrinISo7wjeZTv15lKhu5YP8dGfQfCxkO2i
O2ghBBbw57Gd/NHX+FcEtW5fH/fd726RkdyqC45cCkOqEdeMeWDoxGw6pFkS7tFFd6iQfOcH58sP
YXAhIEyvmxdsv329IHofDCDkkNirVVzNplc7ynBZeqaGb4mmRWzE2hPhdw1mrIKrEDofQOPVgskN
0Z7/ShBF1egIYCzWZSgVKGCn2bpIa7VwtnSB1IsqoV9tXdO8fmj+yosW4xTVfaRYvvqSCqosRh1J
vyMoFjmv7kBD2GN/304kKIqo16vZS/WDPRMuChtBjwyUP7oft0IEJWsOS4GY6X5Qgok0cblpjoGH
LFZ+VBizaw6oJJiiavV3bKW8HsYllsNWHk8M3cBMqWdsBGTdCnpZhyf7ViOmQYZwh5kvFzt/jMrN
B9wocoO4G9IP7yeVY/VXOHeI54tyhqEphyjwYIo7u2sXZc3U2w8uimUdiva0WuMDYQY3DLX0cu3R
bmDJlCFOkW1YOxWgS6hrZPfvhrXEQeRjkGg8tq1CUwN4AHspw+2/x61kOt5cc6y8Szr6xteAU7rY
udrp6XJAh9Wr2qPsDUBatEHfS5MNhNubooV1GaCvT5Ig/08Bupn/frwKWgBobGIwhhtuUgedXm4d
yhI95Nb7SEzMhAawTYsNZxIxwJhWa6a1ydFfxFNp+nM7v+dvB4RCGHSFzdCnVnCSPHPValzgeCou
wVVqL6CgWlJG3qeBKH2TRyvJS0Y+Xu5PLaGVx7z9yS9E6Qt8nzXqaR7xpitq+ftf0bOxcu1glX+1
BT7b5BymMaLOQ4V/VT2GGZ0AynsBSlsXxCBGs7VGlM59+rhyzWE4FtEp7LQsxWdzLX6mBJ0jlHm3
v69O3nhN2qEQC90gFby9psbOypZ8QO71L+OCARd66XF9ZGiVwbBoACFi1hOAR4636CYwB9KLHyrN
qygsUoiM3GRyOyinMElxO/miLmmOL6o5lF5zSQWGEntRKSyH3B94aXgub8uNvchrHh+Hb8NHd5A4
TquUjS7zXto4H7bdc3apsenLBXYjFZ5VfkTe3Fd9X4VlbBnVXF9w4rrjukzOA6f5iqZ2R9aoWh6n
3HdFlb60+hc3osZRirBj3Zz0DY/kL+BaD6QyELkuzINWu7J/merqSbHwTULGQcOk0esRuh8s33Vu
eiS0CdsfTSXCDnq+ieZerLActoFuFs3FMtrpA//wCbkJEfg7i8R0I5SQCctBKZUkWqvcHYfDmKDe
rj92xez9RTZzvyFtU/mN2KAOmWTOxiUDPemhqRaK71O4n9HvDAL8jPAAVUfO4fsqtatVQBCwMuH3
tVDk5eQyWzfmfln1GoirUVbrQwb4rimqLtw6lj4Wk16Nz0oLcsDQRQpw/hMBFaefoJYOz3z1QUvY
3mFalsKEvMHy/gIU2oOhnNNc0idt9rjJF9RRW1bqajhQNHV/yqcEtFbWED9EbGGT3YdHhFH963SX
/H4RSvOjPKUkC1cH+5vILaOjWeZSC+Q7/S6/cJ6Y5i/EpiecznztSEE5O4aFzMWV+wuqq/LaovS4
q9IfWXTiOHdrk1zAaWkncXMEZ4Z0YpVCa/v81cQKg8lU1G5fAm8LoO9dHcJz00NJkIGUDZI8yr1W
4qGthQTiuGYdr6jIB3c6vGlqvCb9U0cu9SKWGA23FtdK4WxgJv0QUlmpT8XNTsBY95k7+WA7vdFa
pqiZt9/BIA2bY7taYh8tAHHH+eGBMJvZfEqGecokURVPdJm+Uz9pX4QmjgLVwTn17uuV9owdQ/1s
7m3MxxihxLI5lKCfDGTwjNBY/h4gI9fMFuo0OFzmEBdqgKBKseyhNFzy7tEMTo/V9Oozb5A+yQwj
sub7iLclxzNKWUauT55aOEdgpdVZeVzMAZ69hcw3AycvBW4AI3c5K+jdfT0us0bpCYui2AI8FrW2
oj/vAf9+SEFQXqq6ZqjogEdPu5sySlgoFwpl2bdpoidJw651btDaqSCpT1XWNC/jaP8TG9AmE5fF
E50cd3fA+duoT33cy4+dx4KBpSFbJl+1dRB+LAsR7KYrrzyV5GifSxh+gjlE8mVrpESL2RNCuUyT
DTSNaHsSbENrU7gTo2DorPFAnkY6JbbJmpHggMcf6lToA4DYt49VoJfaNvLcqf3TlMbDSnhQo+nv
553tmQ3VK5QYi/FIw8Zb9DwmzMf7P1sHtexijJ25Nh9WzqxKk/XMxANwoZzWGjKDWlAXIpFKNVUO
K3X3TjLkEJ/myxL+e0e9Clnr2t4M6v2b3RHoF8As8ZE6lLoNB7dpSXIvEbs7QrLiCbMnAkgTr6JE
MU9NL0n01+WQiwUHSdHP+U7+8wyt4FSMYNAWxwKX2rFam9qk3hMkAQtz8Xk4cZC/h/Dr3aebwUIV
iRprY9EBhQ4iMyfbs73xcsfSO96wWLkLLBTdiymHVa4cKHJt6kA5p414sJ6zQPC8PiiPgfj4mrWo
w6LEwhLkQz5o46x5DvQo9C2fqEa/W0KYI3FWn1yqZPEHAbH3B+ZxIsUAoSTdvIXZsBLZo2eLa+Rs
K9Kn0xZcx6Ydca1PJqMS+AsRJLhQkvHObvKKGSgXcCjNGx5suZw+x82dDGMxurFuBCtrmiut/GF2
VIowAD+r5Pc5cnT69PyVC65Ta8eN7mljdoxT5KRKPSlgj6R0rZyB6r471oBMtu2CfW7gd4CY+zOP
kSKycwnYYBcTjMn9G2iWZEfhGWm3uqVKDKZsEG2TEVYcav4bbeDmC6/+Bjg1Sy6xM5+lgE0bvfAg
u8+ecR+LCp7C9JdRCIee3QL7xEbbx1XCRrlnaRlZm3qh2W0ayQwtjGRwCk0JHjlYb62qFZc1KVH/
EJWuYREiNRr1Fk7ag5cglFQEiIXSFyuj8FTbNUcoCVfof/TSAUu+C8i99qBlgVcorfdJ8fG8wtwV
aVwVNbnL3K0xHUSTa7b8tfYMKixlo93N2xMBtrEsEJNzUYvOSuYqfW66UIGlvVZ0de4fhstUgO/5
dSrwsvfjyWJYqXpOMtmqWINyMBKSiU2+XlIR9ZapWU7bwM+sRC9QSK5Le6jcL0wdCgXu1OnJQbZ1
nIAAQJwIHdbzVZmEmleEUJSYAWLvUmp6GPBw2LWQMiS6/lGuLn3jQULEQrHzQQhTzCaA8kXTalsk
rldp5SGtqLT/e5Yx8yAXvZJzyW4ZyoFjZ/KS/7GjmsM6uZkUpj/7XYkuhC9apM8FKZm3UivPDolJ
a2f9Zgn94KM6gUkNPxn7QOOaollUbVdOE0Nus1IMwr3e1GAHWmBxEM0KVZndSAJQ7/Qb9F6i7Rxk
L2T4SQ4V5OB/ijAxXaF4UEPMLATvX+PiAMkDRCOl/7su+Lu8PQGaBkpqYztek/ahQd6V45Uf3ncO
AmNf21cYtBOoJaj9rONB3xm9u9q9mIPcQsRLrW+uBCqSiUisqC2o4ZAsWlVtvArN6iEYoC6XiWo3
DH9p3j86LSoHFPAz9wk0DbKREpv0jUma5EV9HbYWwZpzPuX8EaOInlrafW4hqHsSLrmzrlYDRu/j
33s3ZXH3m/HkZpCA2WVrCRim9ebCPwTOK8qvNpnWPMSSW7gjHX8WlDNsC/qBIStlJ4i4OpS8LWHA
y2zr9nZ2KRLV+g7Dnk+MPUw9OBTCDyP1Ip/EqN6iATgRloJjSNHCjLAJ6NPuQdgB+QJgzfNpYwaJ
pvlR7C9M4JYXlZn17FjYK9g/Xd4tSHyYjnHMvCDOHtBnx+ieDYLTCkbNN47kx+IQwwzdl67sZDWa
l1xCswCG5uaepvBy52Z3SSwyWwhIbzXklvN3BeoDKQLoVjDXqIfqS4lgO32C2eDWRM8v1hYHvjjR
5iBFwFWS2iV8CkFnWw+Sl90YPbNB71E7KDUvRQIPaEk7FClthlG9RTJtW3J5mw2JWJ9ZcycMlgyY
UMA5CJJ4Py13Xzzt+wdDrkOYN8ixp3cm6Ui+ZmkZMwJVOpyQJXESiNenMtOphm9UhoYMUZ5Ie87Z
hpF3myZnc+EnwARqMgs4e2Wtbu5g/YNQSZOtRJfmTLrzFpSA17D/uTbx51Po6q0oQUTS6tYHvaob
nO7Zed0osMvbzLwd2HKMq5MrxIh8KTGm5OZ7gtnK+CJ45NI9CG7DmCyKe0wqlRHMGsnQoEpDgUKf
O8XPwwhigB7y/Tih9RQu/kcCCc6JYeZrgdVNK0DRFFnQwLHvFvJ5wT0tlo8LouA4888rgEsnJOgG
85y0dcboErgxG13QXmKCxQTZ0JvPB3kU/WZmj8YKGKk0iEwP4XD1H68vGkAQl5W442PMPaXIPffZ
3v6ICp2vGrusrcOyHU7K8BcfsggTrCfwXi5XXt5xmJC4nvuzk+6WvAUevUU6GWPJ5iLmlzGKyfYn
DJwoDhm4PqRTaqsB+a/ryP+2kqsr4QLVIElDUidMLMj92t58zPgEzm4u0/LA33oyKYPlAs5IN3xJ
r4dVAoRkYBu07trc9X/LwWImmVKL4xpF9sTi6t5SWEGz/Qv9PLSIbwGh70VHk7K2Q+UGxgiqtqOY
6ocn6dLmcuBgG/BcSfUhcjWIzYD7Oiwlc00fLjMyS81rICX9Zf0osoDRx5pzZLc28OLr36HTnmtz
kZQwcdpJ8ta/Ujh4+8Iz6sWR2xLu9YVHmi0D+WYfB+1uFyIxgt677cHjzBgKI5pSP/4OiKuP5JxR
StnVSfU8bvhkbqNzx587akHa4980l+8UotJcUwaljQQFs+iE8sId/us1n6Ucw27YeQvvKHwj3AYd
aWKHDWTAjE57ZDDk57bQkJ/LMe1mSKTiRyeupK98sC2ACb+YUg5dD+V+oDVKpDNKmvHKPBR/lPxW
98Mo8PLQ0E8UZASMaqrk4NDPtioLB2leqmkUYkckieD6xomkfd6a0sSlKfPMaPOXwJLnMr/QH+Ol
34OTEu+BSLEEPkOGCf6d0WjzjNyBjv+jr9/EVKwLgiu18ycF03peRZhf1heJEtrnvvIQBI54a5lK
Oct4LVvtbaVOzguys+tyJwXFx6scZm6ND8YXEVb+UnUaL+o8//Rz8amZ/NOqs8gfHERwZnn8LIdt
9iNaOEibNERf+J/KBtZ3Ul8GOFa5UWrtO1bWGXqtm8/wHutLM2+L/pb5i+5IqXNZmLP3Rih17MIH
qDqkDK1VYaV1e2ia+G6cGY4C95lyczkkVDuwH5HLIwOy6OWz0pbQ2V1baCVDiD8cOZA+KzCsmQiL
j3HG0kbNIAdtDQvSvxMQHK4F4Uh6lqY9EJqHc/uRdMx7EZhl+KXf4Cf/I6Nt7D6AVuNcy9oP781n
oK4oFiflqOvo0q5QydQsKsZX0VqL0/nKFwij4sKphczjdVQY5qtWSMDlk/jqZuzlr4yLBYCOnjNJ
9Q/WUj3gza4CHnmbRFLrzjhhAtpTk4898Yx6ssM88/oeibtDXa2dChYvT2VCYbiubg87e5cT0tsY
G4bC5i3X65IkI6aEquwPg7NBeH3quF616XC/pxCmQaP/7sfkH6x4eiPVeQ7bk4QToZ2b0Fr4gsF/
PDjxZGcGJrgjk/r/YIghCNYhsGGBsJTDOK9S1woqwBI6l7JmQJrecGivgG2uyoTuIozkXlbBrPsp
cdGTIC6wSJbswWhlzf9YOSKQSv+3Pe7QexjKUkWPZnM4UodH+XINbgoiwSovAWvkfkpt1YbLsU0v
0/qfG6tXniZ02HbvJYLxYnlGhyHohlf48mXtKQ1+QYWY/Yx25gFASijuvonIP3GTbhj2SiBNtXv4
QMWTDWkWhlhh3dlK87uYXYP8WcbONJOwBkD3ZWuaX/rSPh10ev46pClcUXvngsmIQvPeykondUID
9QlwG5fwhYtZDJDLVnxeWPbUtHXSGukopi1ADVYaoUUGpsQVFM0jEYxHKgh22j4+mFAskYl0ENYw
VAaqnxzaxVvcjIRpt6qrHMZQoS+YctzmnsM3D1DzNej7DRxk5/KDfcQCVqGJI2OmqW9cwA6Hgrqx
awxfbuHuEpEfNm+OXLmQrvF05hLMFVQdr39DlCjhYtIzBGOD+Qd7tq/F7cFlDJwtzS3o1f426imv
nDl17IdFwmY4ysJtx1L01dScUq10Wq82GjB1Gfu0cQycviVVUhsUCg4PQG0X8bv591sBtRKzSeWe
RMby1W6TuctS2CA2UdF34xZgSG2vlt74rDR1VPXF/w+mHEC9SXbtO0mmsl46g3UI3hVFEzNDbtfd
XV9opmN7keepEmBKzYpOVxwbP+BxVB8HV5LUXiUApsrTOT0T3x7tg4NmY6DLLSq79HmKoUmh4dr4
j+ulfeWniqfiGWT38YpP04l449sd9dbRDxXA262MyC7Y3bpupMlSVqACDSHoJnmkp9nxO9KS9sAD
gBMzktY5EqkNVpTZ3i9S/0xGI2+NBkanFziaNxpOWhXXLJVj/ec5tCIQc6MkIEoly1wMkMkQuSOy
NpmefW7pdKgAwa6inxfNuf9KcJ+6f21isZKtwlB3xE3WmqnPLPdTH53RqSWJKPCz22731tvk1pM8
5Ux8zGx31NtfQ0fevHP69+xlCVz8nb7dtsOYvK75m7SDEKbtX+nYwMHbhCavPqqeBB6fV+Uo+fzM
UaisqAWIX+sDixK9wO817xi0cJ+uvQmLZnpVLngQdCbXocFrgDU6/rdnisCZfJ6eQqbTomCIk+IW
9D7K+jYv3AnScBRGVonHPVLbRIusjXt8zKtC93hXBtHVXlQZK5nNVEKwCjdVF39H0tcBdFI7LzX4
QXGKScQ3QCsgUuqlEy4N/f92LxTIOtxgZMqkPcyZvO2KbQ0Zo4LGj95si+zSemFGTtwy9z/+2dDT
F0KaXEOduMKClfC7EVBaFRucQHnZaVW1DAQKXirdLdMJ4+0d3COUZEw6MRf8N3sCadqqGJddFMzf
or3XTkJ5aGCLJTWzZGQ+7BRxSq5HqTdMYV7VbsXghsKiDutL3saJkOf6i+P7fkQ4HMA4sh5GC/1c
70FJo+9f2e6LbcU3OfbEhT/AQCV8yhp8y2H06njmeof76zC7HyCyolN5lu/QY30QdYHqnx+EwUhe
Gqr/2xzXc6BnaiOtxRKFMNDcuYC0HghNfP8M+tdoAdOdene4HfDKfo9c/003V8cTybbAC5K8tGhD
dwEJ2TZobY4gPkoWXXe5PjIxZm/aDsuEXWctfI4x3OYTO0rdGP4qcbnaQkB6NPbhYTf6SKDTA7qH
e+IiWYBbrZmO4k/f6DgeiuBtZT5XpW0YSSlgf+BUGzrOjfDAeQhejJFyp5AswkuhQdfH9//DjRBW
QOTEuLJIRBI/CjzmHPXSvN8JrfYUagAjH4bjh4KgmItswE1DNlMeu93X8NoZ0GKgezjvuRCFYyUb
dg2zhJ0VPf7+1UwwsoHzR/bA/XvZzUmNUAtaaXv5Y8UGUlrV7JHoxIFJ7rUaC/LRB5n1SeHmcIaQ
O7nbkLPyEMLEsxaP/G/nmHFWjkMZxJe13h8SQluOmcXmko++s+futDvq2hLdz1+cgUKMMBy+WFQA
37KuYYaCGaMIZy20+Ey7enoAC5OQ41875aTjDH1B6XRmYC1dn1+vqHfteOcNF4ElIdIIcj6FDu7m
tX6P4RiFNTxog/VUMp9qP7v1rHJBLbKhKTp9igzXR3SrU+AcvMNsfJp17d2Z7o4IgIw93C3XVAwA
K+6smf/OY9j3vRFpp4g4fv6H5K6VSMocjv6ykJp8aNxk2L0zLgAKrOFUtmCm2oN3yuAfIrlzwXUg
72J7Ld/WrqrvUIMIxV3imt59bIvA65y73ZXD3tk9CDSo3HmFgxgsOESbBy5MNpc8jelrl05qtWlS
VN/tHhLb1aCSb8ah3/H19F4+ceu3EUSehNCi3I6/FA+NCutueacsdtIwyQRKdXHmCHGp7REwxI4H
GIMUv/VosdUiuaDpk2x5PghRJuwSwkUBsFbIvjYVTVDDeb4lk6c0D6Y+04i7FM045qMMCfUSD97I
OKT77PkTq2WXpSzWdl6+GZ98niYXaDXpvLvZi4fERM6M9mAiyDzWdYQr9op0DcoMbTaXF1QmOMvZ
0WWoCW2ZYzj6zuh1ZEIgzSFY+89fEffOHLfXSHZeuknntpf9n9q+WYLWlnURUU31XFZYVlOYp5KL
fGcBgDIH947/zWCkEEZagkHfYK3hPSfbdilDaShjO79c1vqS4j5ob4N8Sbhq7rZ8CZS9p+xzM6/M
WnrY9Uwt+ZNoChMJcjsyWgwTMBRfXedbz5lIV5TxxV/ncTjeDdnr6ZxAqXwEwG1XT/fsfOG7ug/z
hMyHCjeq7CvtXqRmpPWoQOdVZX03wVkurZOomGRFw6msarUIa3A7lztu8AChbo0eon8pebkEkSrK
0iOkNCYnW3ejGHRVq6c0mt9r9xRpt4m+NInXzfc1YgyWv8SYtLzdhoNBB81WCqqkK9ekcxvfCsz0
uLBeiw88Jy619joQoCYk+L/3w7fg4ZFZYOdLjEo7Pfh/3hD6HTg2tnT9xAdm80U5mmFd7S2TzbwC
8QNMkLhah3fREijTSxpRRYi6n/Em2l3dWw617hCHx9Z3FNLjo+5pfiru/Ji5Q15l0vjgaf9CG+qm
or0qY8i798rpkJkVoeU8QfJIJfDdTAU+yi18nZDxMuNsvNM7MEgLf+cPQSoQgDuOKaPf6XkuBVNA
bT7M13EXAzUJS5/GKsVwmNwZwp0tD6+d1+yatQCznRKaMKhziv208fvBenJnsia2SmKQGTZmyUtT
0ZWRgIpHQGhDrd6liLSpDU1Ax/XiX+FAjjLDEzT7gPvRRZ0ZLpqO+LtDbrDkCZxJFcYddzjvwhxm
HMOXgBvDO/HUpEB/eFBJxdBD/Dh18cKQiCkP71FUMo6uFyEKSobq961zPCxoOzdeHRxK22tCy4MJ
nAz/9DOCKR6H1ZpoPsFdDdsB8hIwLewutwK9gRNkVHIAWnk9+JxIzuXj4r6dziS42UYnEps2xwJa
TAexFzPksSU7g+DAemN9iECih6yjPB752RhU8xtfDql7FHKYPnABKfDudq/N/F0s2Grbx6nruXui
XdFe2AhGERYPUVpn5CqCTrew7ai5qv7d3PLw9aynKQfKjPZ/1cT1g1AfEAnR7ji0t2ck/QiPZAqU
y4RjDtL1x1ylTFuxzuGNrQrrIQKxwPmHGHvVdZYR987rcHa1ZFqw3THaqfsFaICSsj70cWmZ9bqA
Ilgpxh0dBZ2uOZdrXowH3TWIEiiLp+quC5CW3yaKY1wKFSPFIW+h6fnWWqp+ZgaQ1RuiwAJXEgNH
NuMfkBsjEx4Uf6Y0vMVWRl6OM1Ao/RHftpoV4QCaSVVSE5rpfY0Z9bc1t5iY4K7/pPorCM+B/Hf/
4FwawrX1HvF7PzMXB3FihurgCeTX3MXpibuEdK69w8JL6RMTHXLHNL1LRToidhf74Nm6kwge0KX/
1MWmVpD2yZxiNMEdc1L/TrkZk6KyNI9wUnh26UuEPGjKg7tQrDAKzLF37y0ZUuz7M5G0KMVYnOcm
idCVVbIMyPBE7IZ8tMz3siGp9siUq064VV82cNIuQ2iDNh15H9ai/bGlSNRT6v4S3QEHRcBlVM9q
NNxfNd4qEyueraeY/ONneErwtF2NgHimegWQlZqSqwfMacs06lgkkNIKO17eQTcFjFX35H29xcUL
VP08WMcRTeKyNUZJquCy2EAPdXEbEHGYbqiMmw5Mf5E75Vby54TpLGlo6Lh5phLlZcyT/ebN3+e3
ugGvSfMX3X17zMIZfeXCFRuMgleOcGh+hYCmMJwhRthS0LujqsYGjOQxDH4Qs2InFexhXrTRLvx0
5JrQW3b2xe7ffmNSrc6Vk7FTDvHm6GlRgEMxW4E2bFb7k2Nop8j5F79oxXIqocvq5uaMYF3Idjd3
JaE/NXceppiM9rJ1ToTyF9nMvMN9N4B1/5DgGXoiU2pkTOFT1pNFUQqBdbN7JCD8wMV4++W8LF/7
B7VO304c13n1xzKxIdJpT8NqUhW5evcvKZ7zNzVStTS9yD5zRGfUB1DHO7gJ9fJQobaPvNgLnmOE
MLp1kFFPjO17NKkiGq5CTSvOHZUWv+XV6d/thgVwJHqkhu95br3yJ4YdWnmLgc8iHbj/Y/KxQ1j8
0T8WLJ3wox7/KChvxJPLfxW0wlnlYNQCy0BHMEcvitoagU1dbHVJyqMRvrgXb4U6O+H9HOUCG+yX
NfUzEE/wvIrnwBQ1SGQXmNNJ18yjKtW3wMIqVZKWni40GnpCJs1uzR1qnaXFqSyMxitjyRj5B3aP
nRylMw+7EKT9ndDtrvP5VMtzS5XiRZvCBqCbB3CNxCNU+gyXzWPuTNHUvZ4oqNBL6bPTjLN9jHIs
K4dOf8+2da0FiKgnHzHdaDAwN8dlSNEgBhDTS5Zv3bECcTgx6taGZVQcQu47C4thIiEpSuLx8Y8P
icyXGHiTBZiQlPJ3ZoquZZZPnQlNyQkS8tUtHY2puBmjmJhjNzEEMg8dkdnTMoT3ATzkEVN5Ye39
sLcT2oPLcr4yEILMtErSq/mXasaFxcADfmH0EKE0wmQtJa8m2sutdrEVuqiEYkSr8nlmLLJReCgD
5MScMW7AvaUeCIKtCYfMoVEWY208egj7Hw/vlj05gNyHIKERnz+zvnEqZ1ajBj1xjLR3b4sw9j5u
ZvIlFyN03a0wWT5YDAP1bz9piKAnz4V9xvdtyaSSknJcBTAPz2iSyUvB8q0BuXalmH3OpMJnI+ui
RMd7ssoudT7hyizOsvNTB/WlnlDzHrB+OLg8+JNkegLLPBSbBxgmlxK0wEjFOTgD8JEOwLGAMgch
RJtD5PNuHymbwlD3yC8eP5kJ+p7Sai74IDhypyRBttr9ViPQ0ja2xLXhdLLS6aE5ONnvYJf7/TUE
6VnkLBQlYjWZDThwgfcPrBaF6XD/beL0LtWWmyCmw6EJtjgci/eRq+ssI6h3atDZRKDxuZRfmd6u
26XCIa/0AOjGJ89xraoN6LBKrlGexw+y3/kfNjJCOCdBp5Vhi4fi6cnT89jQgD6gK60/PIQrqpqF
Q1RNde99Kq5jGtej/LCVsU3XsttEePJbvVhMjT2GRGnsLIo7g+t0COf6To7u+oGVnhwRLjuH3pwy
ObqExheM2XNJD/kmMbVnxEiStL3rKmJt0mggxGJR4H0ARAAB5UheBQzP8PT3bGSm5/BVHiV6aSgk
ywrsQoCcyiXwLc/Z6RZewlc+P+1tH5CuMVeOjRDIbpDTBdBzvK2l3iEMKrtvxCdqBW4EtOjdCYji
zuDTwDQWyxh7kSpIyCdec6ulnXcNNzFMUGpV6QGxjxd5IvcX2M6xHilZIIsKr5GcuvmaxCntofNc
1WAfN+0kJV2nwAQn/XLNiTXdd4Xpd3PV/br+IagnsceZz8WKkIjcgC1sDNKKYlCHxX9s/b5FQ07Q
W+KSorjbf86J5uQfb3HHJxm9S/O3cfWYDSuqXzN5/RpV2RbqI5QOGngDvPgOw3/uEkIBahN82BD4
/iHvh0lWFJA34o6Tb+FuASf8ACz2vwRTVDP8Egby3rJ2oz2UIso4SfNOJT2VF4MSgHCS3AdznPW7
IpJ/ltbU9bqcv9IQ4IW/8DCsW/PbWA2ypo/mt4NOqbffCPk0hlFgTkCHxI3E1VNLdxsTSbdvs617
df5HCIwt+q6o583qtg7kZD4iE97vdvRfhgkVwSu0UDtT9rD7vcyQ/BOdPSp8cJH8ugrDpBoDiPji
IjoQCQZCwMX8gdIvUbaN+E56pBbKOL06YKUzJOTLEtFerJRPXuQu5GSJE0WFxS0ILDNNeHFl/DqB
WDTw7VY2v01EJsMuRwflUOpWaQDi/rZ8vynVum5taZusKHgl6vgId1wvjTQGeYJ7oRlKhO8Ghsam
HVreKaJNbDGFjX2gcD250rCK8m6o56Y1deaTmD6es9a2mSQ77bJbZNT3+1H1FRK6OKdgUzfBUEXj
Q9RomCvLw5iDxYdsrcprAxC3P4kQrpsPigIFQ0iNjTHh07U+JSuJ/xUrqpgUZX+0cp2dc560LWWZ
FshvtnThp1OmSKZDueBN4u8AIh0LXZ/IvcS1NjTVBIOs6BYM7/mSAnPn/HxobczrbGYQWWqXL/3U
B/G6xwPgfD6KToGS1+1b/XcZWXF9+ze8LrUpsm9e+cQslqOypwgFg+XQYPNzIAyQ5We1055fjJSc
kONs/i9pPrFlI4B9U6fYEZ8KlZvyAZevo8padD+yLwKsbNiuYzukvwpAF3KlcG2YuzVs/MkuYbg3
4ldZHnjAuSlHGJt3HNMS26EMPOWXxdMFf+FLeKTjrJZopTD6INSiK8fX401+MfEuQnokZVQmwqfQ
R0azcc1Xok24n/b6NB+8jVCErCl8BX4wc+FumVyz2bzAZDwxf6K0iR1LEcKWUADmDzPN/pE+sr0c
O/0KMCapXs1KEjiGrNcdiBqZ+Qrr9/S1fF+uXkdLVUXygFSkG4ngtFc7vgLPxIlyZCkMSC03gDnd
DCWqpFw2B563ItP3itB5fh7HYlnbidNhcUEiRR1VvZ5MCHzLSGacHOmKAmOl6xXFFXb+C+3CMeIM
MI+RdAhOioTcVKuZ0oXe+26HQ48qUMUJxPb3Zpu5nhxb5q5e802zXU+ALllB9daCaR4WckT/XHzM
X5KgAfUNaKG/rjteR4pRZ5+898JbqSQGNzasmVgnB4iV/rIA8F8IQzk4QqEXd6EKK8CR7VlYsKzu
DOHzOtQ09Sivok6lTpdoFvAH9AxhPumxLnrvmPP6a9iaSxiWG/gMZWA0Cswaaf1IXfDWHz7dWO1G
tyS+AVvgvmLwC+RSpfOOQTtUsVdRKVndRU2LPHpEydF5kooFBIBaUXWXuZQt8gJYuDH6hQvf0SBM
ESDrHb7U9HdGPm/42wicDduw/3XZGqH/6BDG4/MQtyuqa3h7L6aJi+N0e8mYZPQjdqDsBL4LSJqI
tHUQsaGgOCiZNDCmQfYOaAM02KKQgC2k0zHZwacFvDMS/6QIPCCQZUy524OxPrv77ldYE5vgao03
q/JTdv2cggQWfzfI7WBzamdgoZu828SMUmSDMIN9SarZi7Az0dFQoC9dllItMUuJA5bRQEC0hhGO
VrL2+23jsUh8yGtGxA+1kKnOkAJT4N8jdiTPnK0j9dxqcFzpdPq7kPRAbzWRZbz4U+X7nKDEGsXH
Oa1vmTmIt2kNAmILI6Ej4j2RZ3rnqBbEDKGZ4flu03qh47qh3c3Hg9it948eVisXVwOM66wSbbRA
g69bD/RaDaxIWXD7lXUjfQnzvfI1cMTnqVuJtq1yQXamZXIiV8slSPNPW6tBo8ZAjXUCJa2f5ka0
0/EMYS2rPMCQEwdZPZGdZhBl8VmyPGjgtOmbxzaJwpk6wawAqYj8so8ZWcgY+JYoAjUucsyuxkdf
BFm59cu/YgUorE52fddqMLnQg5amsmRkYO1vMJKj7Ss1MCkDBpik4gw51JtPrW6Ur/aRFqIWuTDT
aAiG30jeOCL70g0kJwpgt1NocFQO6fUuVjrk/D9dEP8IoyzZEFCQ1Ktte/bNb03zsW2fjvK5VKbw
N7lb0/K80XU3mnT0aZIiDc2j33333Q0xghqLkBoL65lACA54wC8/ZVGrtPtxjqshIKLArMWsRKNR
NIn31wJ1EgVssa8kwqLl11IKHrZ2lvrTPOplWfvK0ixwHzce5LvBBiTIx6jFBfBJ4RM28+YyL9uF
guiK3JAKPhwwC0k/StyeRIh6ARHeY8q8ZOSS3GI9QE/QgJ9HieDcCG7HNYIRHN5o9TXBziz+PYKE
E+xeAJKUVmJIvQ/di+yNYFu9m9okaL58T5ioudfzfWbE68FmyK511O20eLzbOgyCTq5HRq9G4JwX
/aPUZCd+rxAF1aMzdaJuISUliboK3io+Ay5qikGREvCJqbCgPtXHASQ9rfOzlhEO2FEWTEcjTplS
Dxzfevd96UIaiNOp1nQx0c9SbB1GavQhud6lb6pjpNVdd0bwWkPi2l9H7IY02ze1jdbKoZwC0ZqC
R7aXnGu6noYe875SddnGrabNntSIIMA4t+YcrloLciax6EJn6PjuxoP4QolRhcW3BM8qYDiH6vY/
KkHi/nsue4GjN/5yNfFnmDVum/n/qae3f8pCx4yVC6S57maxdXjPSjGJKEkVWtbNhyhlqkoHZKZk
brbHTs+YtXL+nEud3G+P6B4Ghd11AjD6ZBN4WDuUx5CXSisdK7byhoTusOd7rRoxX8SceSEXYJmz
7LHxnZy5kBVxVuTD+VmU0WnmVeB8kh5PYVmHF2LH8lmt9uxRNd7hXF8tgcBmC3FAglTYMbw7owHy
HxCdJcAOgB3I0VlzHOR2IDwYfLy3qc2yeZJYu+EcBAd9B2s7j7/VRcFuog3q7S+c0d7mHrhczpHc
NBXQjCoyrmY/Shj0/D4meXQDuvpLZ44uSK2s3FvTuDrmPrOxcNlYiyJa1o8i9fcCxG3pF7uZhFsH
SpZRwnh51KlbX4OJ9q2+4aaHwZv5yVmX9b/7dzWPD4OFB+HMB5hUdnVyh7wgzmIZMhjpfvgNUzN1
86JXGLF8nnYMS/TLKkxKpkQnsHw0i4VKuo7zrrHg32GiTCiaegszbNoHDIkfU8kVBeqL06ACxhhC
Su5xT5cYK0IfGZnBmXZoGmzurBr7hDGtRTYLnvIsG+cG9ae+WHAbzNwYlVFpWagUf+vH790ZNLmv
iaHplb3f2/sMWCC6T3iWDBJQSdZubCerw4t8+m9wLHk469+jkotRbVpEzqjuEGmVRUmYOPSJm9dD
R0hoW2sgC51Dtl6l465z9luBvkunq1+b3XmhUumJtrclf1K5bRqPHGpT2n/NWa6PyFoFtWkdmxEC
whjcXqnw/2tPIeDu8vgv7azU2CXn10PXjpWD+t2qZZIbBRlVZdWS+mBc6h+4gau8iF1Cr2q/GGzR
65VyGRqVOYKznc4lSxF0EJ7m5jS7arf+WDopI2NqrEXZfOWEZTTIx5jugN3UJZIdaudLdl+UJ9AK
pbFcpdSkC2L9iAxo7D/T6D1GXL96tyq7QK5q0v2omWjCcSD3IbRhEPZhnW45kky2AaemFnO2rHfL
klwj0eEvT3Xba6PY60kcQm8NYOh/+SvnqcyupkXx4i9ekyu03dFfChrV1QGxkAsorDKEVPaRFWA8
HKKLXb1HW7f5M6uPIRzKjNEdaYb1jW7vp4i0+d2gvS+TI3gHgc/W/Ys0K1VOzLjeiLi59dzxnGgW
IqgEtBlAsjhPwZ0ZUXbAjoZoCkciwJZ4bCLn+uh5gwfMv7jLx1l1IKt2znzkIc/iFi41eTQhREWN
toNaWzh0bzQHLfONKQEWaY3AK2j8TuP3J7HKGzTLPO2hayLjQvH1fqNh5oV1276N6JB2M6KZPzpx
C5GLzzI/o7vN2+h/N9fsE9kqRNh0ZBn2vFt6IVDJofHN5sG3RKA00OsGkxnJWziZV1qisvLOLhBx
0oQyfwcBvuBB20Ly+iPWyKvsUdQ44qqVKqP5LEYdtW/Z9IcFBVV1u3+qmQzWc4FDcUpclfqUhU+c
VzKJg8mlHEee3JNb1XCQHKFEgX+MSTmOEvdOok2uV97BY+rQir+t5efDC3t/1R0B1AZPu91B24v1
cBj3Zwmuwfeqqo96UevXVIk638KBtMr5B8D2z4kq9O+Uu2a9ky06ijQuO7SO76PAAWIIoSTXl1wd
ACkX0FnqOSiDHdfb4gPu46qJIgWJUMiEqwEgXdDZkxr0lSFs3P9mYT1iNMtcWbS97RpJwIPjAp3r
kQvFBhdj/C2vKFiK8sFnbqFmUPqFtrpOOchmSkNx1D1GB81PdP+f+w0X4qWVAWU4He74NP2lRNKZ
3xlLEusqLqakG+9ux9a05I864Rd2w/64GNFJ5H2SEm8KfHqu5C5UIlUWhclxxPNQtDBEp2RrxR1E
HzQ+dvTxkEJ0vBdSdJthi3FGiWfOPI1RIG3IxRX7u5hFOeELl4m+QKiYSMH1CkgMS+rFcoPPoaKF
0cZod8y7d3Ccl2RkyygENoktwiPXilx1n71lDFy7U+inxNySgmwdADsdlAPqRYnDSF82XAkMB01N
6+cgTVhBrCYNPuE1C0X9pA8UdoGaF6QYjPaOlJUXYb7IVAmja94YGM+IoYORz07zZZ6ce99A8rIV
xaxvUJVYjPt0b3iu/RP78ND2fLupI+WIdVYMtQkgkw5wcx/3IjA6bqUs56n1anE3wbrnSZUlM75q
KRHc8bI+ZISDZcr8JlHM4InpMKD4NfZHFGfB2AvEJkqcREOD5N8Sp1a5gzATcaFepgYwKtlZRgoK
MIR7zlPitqhok20Fa/HCT26IWyNdZCy+CbV0ii51cbjrYMUyTE+27b3EBbCsY6anOa3ufUnJvlbg
R/kX8goLph2u12K6grpYqbubZmTaGMZuoapvHXsTwEwxXUiPX9lqHQ94T1SGBRhaU/0ciYfn9LhO
SKkwiROiPhbAAr3weMowSkxskjWtRO6DsJ/0sC45Bf8wLQFiT8NEpZyJ8FftB8B/G+FQdlrTpHKE
udQml8WSrVgsS4HWI1XIkZSMEQIvoQhctjU0VCxVRBA4Y6BcfgFcUsKEo3O7oxDU2MNyoOwBoI9j
z3HKK4FwkfdaII9tUkd4+FMC5KxVQ7DGUcFP1KUJBn4lY6RQZLO+JFVr3pg/0rZS4LC0690j8GJM
q87i6L2NOxk5/Geud/l932psatNUrs0Igdr1uHXbqSNwbPZ7EHDK5lv+Fyy8M7EWp6DTvYhcVN4X
r2z3lz5zRpXzWTviwhVG1Nbih9foN8hXb0rtAgp4P7CZexqdw3SIrfkA0gE6ugr3Cg8PNuLU0da8
pzxCKITInhhIYbEEmqrw5hrCD5N6zbO/MTfNiqop/hkzi36Wa40VVDdmPZJvYUwFsrFXCRG8OgPn
5s4Liok2iaj8RAqBZSQC8Y/RfnYEGodCe4Mxhc6LNdXc+6S6Wjvfxz2pfaeMdBAg8LsRM/AKOzh6
Jpa4lKncT2sPOhK/7Q1EmiM9nWShLTKr6bcFVmWVyOeyXxrRo50ZTNvA35Jj7iSAnaoXTZxvBF8/
s0YVbkjLBp4WwnXeV0dizBr1FBZjSQrpRh0lEzyc/bd5qjdk/nFM8zq/fr3yiEoUind2fIPxQF/+
uckZUKPHKeZYEAYa4/y3NAjnIUISzAUiMrE4xZDzfO5LlEf/9Krv3F9S4URF2TEOEB186t8rkxIh
6HmjyTVjBsVUIuSzEyJLHTrCgaxquHwBahX1nm9YiJFSF0pUOuP67TIr3foUCQuK6hXkwlbL6YaR
WvWL8nFfZ+GnGS9Nx5UV4dsn4FcEyR/UD8fOHk+LsEouGftD8CVM/aaPy3kylz3v0+TTjhRUuS2o
Dn/mbnyZHHU9Ld+58Thk8+Kpn7CZ5ZdNEtJMbzBi4FbDdTUooMDdpxyTpEEr3zCtnZR0eSNStkPH
tdXYkjLbpYqZfPP04C/HKdiJtBpGusd/4q8WwPhssfRDkggG2jmCg5q/rzdGvf4MvdQEFw4TeI//
f7KEq2kp2UGie9IOVjeb7WXCHdbqBDPbBmOBTv5YhdwgFam4FCSInJX8V1gzPvKCxU6E5g3foEsq
2LcAoE3iTdkZRapoXOe6Q3ezphpFFU0nqMHgXnUmlNC9KYFV38y3w0UTq4dCPlKsIDyp/yNgrG+Y
V9V8GzGQSA1BNaiCfJvfSfX37CDXjsFYSL5Q8TfuZJOj7MgWq0S5rFuz65zlvypu+X4rZMIs5a33
21C+ibjdZIIBgZmtiUJ8R1+n9wYlytLG1QKCsgn2BzIG9WQnf5dfjA4CuHAVk6bwgBrWtwXZKrv2
9zkJFUMmxGs3dkxfdi79Jl/xEhlzG2FCbziE/j3JImwu4bb6VFPs0vFlr79cNIC54wIZP3oQBUuB
5F49hWQKr9NCjS5vRJnl7W01OMrrHUAmNRBJUkySLpLqcmg3BFNWTUA3VH3AYeLOZMrDSEgT5pt1
jRPY9zmw8JOYgmj2ozqzfBfbMScZkLeTYR9pWCGVQHFvGIG6sfJL+jPN9dkML7m5VHbNIP6kHJhB
T9HVcj0gwCanCQhblksqP3ClUwuZbArq2f5PwNpnNIzMuX10BqaVX/xPUn2GPy6gUmsnlCwM0mbz
xQdxyBwU2TEs5x+tlqhZrcWBupL/0oD6hWKkrz3tL6nyEqeAihhUoUB3y1dW2UkLMFrbqFYk2Qrq
CZk8s/FDv1iPikoStGxEahqTOwid2SHZmPHNf1JE5xGDqXU8rsO82ZvkBSTsQxIgkP2z4ps4D+Jk
EVH0eyzQksgBXyGud1LKRPzMpxRC17/ztjLd0YuEZDQFDo27GpsbGjBzhfzM9dnr6hZTUCxeTVRG
TTFYlxv2wTwy/MsExfqpUH4PmgIzn4TWI4dwQYsXGA98S+WfUK2iz83BYnz/vUR0rxwkVR51TtP6
t79cCNowC19hmK2cUGCqC/sMC4Cw3PZQoptDx4R3BJJHaBoU5eGUJNzsMGvlc01JLJc5bEu641By
NGdKY8NCZgdJcA7mOBBBZjoGrzPTU2xfVuu4b3XPAtYFi5PQ20VZx4af6HyIGACCOaRz2yqofSnE
o5X9eTjVY0sbzyk56+CvP7V6wWrtuzqueD7CxfsIsDtieSUi9s94/bYSZ312qeH8yCd2f1rjcD/8
1xjH3+AqAXe9CEq5dS30cHX0vvXV69ay07JNm9+vYep93PeFR9U64NWi5oHFOp5/ajfiBrnnzbT6
4lHVHYetx7Z99Y9adUNKDbse1Mtgpm+lDd/EpIC1Or3eYtsPBMNYETXzhTLFzM3wT2eyVxxEDWnk
h3MRXafCFdHscmzyhSQKz7vo2+4nWJnJwfE30/Nr/2tCqjnt9/D+KVIgsNaOS5EUaBeUoq3Cqx71
6yLeDf1dxLj8z+QdGQ2sU+eZ3XSY6EUKqPT2G8uZX9AibHdxdiml8E4CbEduASO1//fACMiv4mk1
19Zjo7+i9daOYkKNvE0D99MlVP8ries9oxnjT25ocAE7S/U609GgRwHvpWIeKPELZMdJmZM7oQxg
co8eEKH1ESMyEFqZe9hBCWlobB+4pWf6lWF0HnkTwwyNOTcgKDxYfZ2AtQDupj4j3YPNP3XDBwxb
1dC3iwZHmx0FLIpIEi+PjjdrsXYL0Fldrfq9VFavJMTsN/3/oxoBoGw2sZ6QdZn/UkyU6oOcnKzS
ktPR6/vlI302Sz4c7B0ilMcrb+8pQAZ2n4LxdI5i9rxJxIJWWnxx+fagZqUyyCBHXDObrVf6Vjty
Wo11szvgGN9Dyp1n0YqWgJu428sWcau3MYMf/C7rZMH9LqIe6jSZhjEQCD4yGaoKfclnSa2t5lmj
nHgfi0bcuFvzC8IlNT/6am9EKEi/UZ0Tf4ZAXWsZj3NtWEE7Ne6kPqUGccVae1HV70vi0ZPUtsgI
PvY3wvSCE2wCUrjXuU90kWhnXVweNoS0fbOSMy07i1ACh+2E2UFgXJFnAeP7qXClA90iPIDGDss0
rB1dRTUSVrSFj3qbaT3Psjh3b7KvN2FPbbtR5EZVzObpwPNjog+V/8mMCeW/aRgk7w/KvNchp6lA
oVoVEBoiV3+egb3DVxa34/t9UHScZF5gHLvhlmceeQ+Zgixvi0SoHgfgAeND1eFWd+BrRKk0C8UT
Tkn50J/6mNtLOIZck7+J5yHfSI0ni5rcRaLVIecbJMlIA6o37cefL3s32Abbo4pYd8mQIdqEe/z2
SSvG63QYRd5eujjNmLQ+UrQ9wlGKL6+ERFku/QUHUwJEkxUVKEP3pv81IUZ1xPVoQfW36WewdZYj
+RN1hQ1/677xmCF0zgAEASHSGodu3G4Y+Rr7C3PnbGYNg7Q8tFTrDZniPkIg/hv7uWTtsUdoLR3D
L6T7xdxed1c8im22NeDdeECyTS1Qz2z5LrkbGJ/I0NixMXr+sAItKecCRngtAgA983b/wCXJgDZu
bH3GFBdeY8WK9goJ3jDaIuN9SOb/UfaLOwBg+vdVDXUCGP1SyxHCFta5q4+zxdCVqTqb4D6z7y7+
j9LiC8jMbe6sEK382ew78r6LR4mZKC5sqPeOLMXm97oCaIpDY5lOcvd3Vsz+HsxkBdun4Ryz8W+Q
aTMQTsWhcqj4S2zVNMZoyvMqJdSKScEyp6rNIKSTA3SrnabeUn52sc4hGda5O8qxq+QPXT4VP1lv
W1kTzyPP71W74pDbfUF6chHxhztrYSJ7csJ/4+0ynstdFY6nNUaTghbKv8BMmDDC6mEHSceUrM4V
zq04wWRtN7aIS6yZiAHC5CjZJhlbiC7m1qwoqVHu/trHvIh4ptGASv4gD3x5pX7LoGMOezwdbwnI
eI60fu3ksTHdJ5uSUDPq7yucQfKtZ5jWK4n4o8FDozgjoCzJdJaqsPiE+KXsQEX4LoG3YBmxqL6r
OzW0u/8dMPEqu+Ajk7HC7vlo/qI6c8gwkS5TqsMpL5Ukg2v2oealJCmAdKTrFy7dWF0SYlSqzeQ6
pqleEhMcgIA0SbEe+POQqT6w6CklrOcLSVIA81BNpRW3NVRCEOU/OK7qYbgypoGhwQ3gS9br4ASX
3QS8CH+Pu87BTOKerSzCasdJ0OsMSq7BOyuCTI83MUfLykM8/OsDQJ3Cgvl4RbtDz0bWAfUpwHZZ
ktFJCHspVhVVCcg6QUpGf9IcfB2cS/sA9bednVIZ9tOTLdeMCcpDsQbVE3OpZw65YxAzHR1M8YI+
UsI8UctbElYdZtgyWu5rFSemaxRI71pCYKl7JqOihTWq5Gs9frVh/8vRI/z0dujeqXa6SojUFxZ9
CqPOlY3GNlM0oZzyhgbCTYpHD0UM32MXppqSMXoXNpGvJfS7Slj9k60JTqgemqLaeE58uO3mGIUK
ott2Nv/f14FSfh0ujsFZl802apjMWlFX3I8lktV5I4f0nL8dRqq0s95dGOfncqghqts6WtJ1NiIy
xqqR3ucuNTTFulSiVP2Qh4qrhPLv7aGhYR4atqW2LIHal6ugnByy8M6mOhhw1WX5EtyqTQehdpX2
/1EJnzSL1tB59qNMM2eOU26Mc6Oa92L0w3lg9aUr7MW2+Q3BhCm/zxMasTA8CLX7dax9Rudfc3+J
54D2gtaZPe4u/d+4O+Dc3Mz6n0H1lA+64bhhM4S0NXOB94P/wv3y0hW3yA7Rnt392u8pn+REK8y8
GtdyXCV84IXOCW4M+buVABPGpFKpDV/XjBd6Lpxgk7vXeX3PnfAXlFvs/N7KLhz11B++yw9WiRl3
EbpyBiH95Jtkgzvb2gXlJtlEhSECdeQ57Sv0Jd8tcptQZ+u8SFKZcbh+ZQhFZEgj8hQFQMdViMXS
c/7lz9+e19FFetAwWbH7tb6oF4RMXSoahK15MN+MtmxaqqQ1L7dsTSUXMm08UVrVE1RzTLyW4Qxa
6mx15QRu2Hyf0D0NhRjjEKtsBVdARitTrae5GMYjx1E1QqoGJY+lziKcjj1gNLQWft/RbyY4NT1J
pFEui+mUmIM74OgoGaFuoQUWDzeWkebCDeAhZKioNRhULh7Wv9qoTAkya/RzRKs9iuTy7JZ7DMu/
IPCOSZTcZqyhI6UZdc/ZJnxyaNhtYQHZaWT3GkzPkMHylwexDAbO8BTJ8WWTwVrIBxDvIm3jPIrJ
N9RkHk41xU4zNlP4Xu4PkzoTxJvhPqvrtAw+s2MTEocHwH1kx08WDkDjooFL1Og96OwpUzvv6feX
4fbbPnm02hubjyFEGVq+iRzES3/Hi1e2eV9uj0j8l2HpFG74SVY41cerP512OjweDUpMZUMLMDbd
2AB6qt8s570CeWm6BJ1kzFlbGew5sA4KvExnAAjdyr+eWcLWwBAV1wMHl0ptM1YtCJA55E4fsBYb
b2/JH83CqtxcUBnZcjxioldt5DA6DL5WYfpXtO2+YXno0lUG38mxdBQWZ0JN5YC0TDnhPdGd8iKj
6IAL89Hg6gox8EC4wY8QQ7YEqXEXVBf7JXSuRg+2VcK7HUjqO/S3aH6G29LVpe/gRUpHiiQiavIL
iiroavAVAV37otrERsDb7IvoBBC9F/h2i+ibyTKg+trIXIlaLN5+m3IeW3s9OeGvlPMjp4rAISLX
UgChTV/OVAkDecNtgS/wOgIIcdLGUn36qRfMauCeQOW3U7Jmw/GdeohM1NPXFmdgze0IhUVmN5Dy
5CnLNxbtqh9hFpB6TQX0wxSP5/wpkUXCwgvDDrwOB1CBw4l/tgIyPLg8e1Fj39bMDygvnCKKI3Yn
2i3Jsir57RX9GDx7TRbV3h5svllNhvXoNsPwB/AOovIHQktm7u6/SZrX0fJok6lRCSRkksLXH7C8
RMN4a5//Kc0JbbAbYwBbu+uV0/x09Nng9zgUPPBL71wqO6WZpUkUnqq1iYH/vOViXX0t3DRClzKD
sfXKBgq8gXYwTXyW86A171y//Mfue6FHY+xMdFmVhHY+8pmx/iaIKOzqb2McuRA87WEiNcAmxjux
Baswue4AlcfFsn8Tdm+zmugaFwn68Q1W4WV8nKTl2UoqL7EZ9bNFvHNAAuLkf3xFvS0r8OqzRPGD
Ea/x9zlBr/a6/UsPMKEB1i67uAHop1pUPPB1b/XOLdVT839254FyKwMDfwn8hT9m44ihjPSGzX+h
5m/bgXwgWa+HXIfyzLzVSZyWBTZzW+4uL/IMhPuwrT0vLmlgmcGW0cr5V8fwr0TCW1i0aF5JsLV2
i3ivmngTzuAepmkUpRNhm29mKLmU60vySi2GaYgxAf8x3Z3UiYzxbZctPz9yfBUwq7kNriir0Lkl
8OncpoqaNqYNuS06LoejWtRhWiSbVmb5oKe4f0m7+oaBz7fkHnwP6WgosBe5UxbwQrvIpY4I4Etz
ZCxWoZbTMScd2EufxZ1oHJDnfffNclTz+bSdQOG6ywmu2hJZynmqzytgxRtWMYDc7j1X1By0WKJN
DtDXcCwzKARFlUqWQlQF3KkTXtyx/NZrquR7ZvThvQaiUKO2HsAZkf/AlB6629VVpvjZdAseUfGI
eeT1UhIf6mwcP1z47QYfSdz4EcCOwSL8S8MjlpmlRQk/HCM0dgi92XT98GPGJ0TmdMe/92FfJCj9
G5U628DpHwygmXtXfGIb7+KPO1rTSoKoMY+W3SISERO1+mseakaksV7gIXYfrFiLSYK6avgs44KA
jUX2ZGFKmr5zQJnxz15Tdxm75JeMlo25sA3KJgphYdYyuZ9AZ+XeLGhej/rQ7VpbCXsTW+v8TAlT
LmONfkif946PmpCkUfZ4NIHlwPt7N4EuEpK/fGhvlQmcuIBZ70TC1jnpEcgF9jKk0d6aPlksa9l8
PwuTVfkjErmv1GSsiTRif6V+a1/zVN9qWq/3JbIf1TJSR2DbzJOgxh9b5Pjujq8iHnlUtnUY3Fkn
WRBhetQwX4RExmO3xmrUgzf9El80IaxsthelAVKdHC6sI3Dbr6TpqG0ky7UHs7Dl246o9Y/pghIo
Ac/69A9fFPR6jAC0dDta4Yo0z1DHGLyeLX/cR7xGtmcfNtXg0al36OADVPA2Sb8XaPnS1wgnaOpi
EcPH9yVpeyIvvbT76dJO5JbKQAPJpMjfN8b5/5cqxkCOPjXtSRjlVBkj9bfnQC7icWf4RzfgSSMb
o8k+v49r0d6/PhYwWk9Wii2tAeZaC5ghXuM7QPMZJJae4P8/zAgGucIdqpXCX5VEpoXtD6U+81TR
Ke1sxrT3iaCX7tPTuwgMpIxKWc/mONgKvWLpODkaCcaJJ2hiLgnYqOSfZNw8XQmu7DYzyFQoeMeF
ZQ4Q/fmFQl3XR6i7Br979KOpjLQ+qH/Dvl9JPZzSjQ8tSRu+8Tsz8+Zqjc5BmzB8CqKbRAMmBKR1
tae+fHKTvyWy9qUrkh2OOARkkRqwPfMBZecKAfEwJd9oO75YlKc94CQZMpyJFb7XMW8EECOk2Vti
J/AuEmuZ3rFAF9t0gJ2aGK3Sr/8+plgOKf4bfpuU1YS2+I/nhCEueNjiZsvJz7wcq7VhgYb2B12R
Y47kxScb98zJ9mgoZ4Qf+RzaJcucXFbOjFz0tUba1HDCl2bm9mTY1dGmQSLnpcPRHH+bqVG+YpLJ
b06jhASF0JbI0Lf1o1Z7l0D9ARzUm3ZOtPVhqOPEXJOH/91LbhHnIpkwCrPcU7rn8sFjHFSBhmYL
h8bG3bTdRiu6QSDq1ztSLovbg1VwETxyN3pO3mM69yBWFDffZG17yDAw3r0WN5Wd+KUdHV/DGfeC
Aj+63PX7S8k7kRpqLHZ+8Fspnr+cJ3G9WNkxxJbBpUwM+Tc89gpFwpx968q/5YLSrO0rglAeo2AM
WeVHi2e/mdOdeMTKcMFuhlSbvO8i1/Uc9yPXdMWoincO3IjFQAQlHO1NcS1TVQesKp+VZunibCMU
lNbC/OshJX2FeoiwelcTMHIqxhjm0g/hS5AJgZByXAkb+FpPw2v+ODEbKoG+Ia/VV3xD0olcyCcv
MM6RhH9TBKY6vJftdrgEE0rjEQ2Cj8TbTApGfOkmRqNZy8ojzSe9Op6Cm9Qy51eBottXVvDrT/ul
lv1vAKkg/zEQoPpkFSlvVimC1O4jShZVnSWnExHKgtF7IcVcYejFFLTcHL8fucYXOSZ88VqYvNzX
1KceIbXUIntuSKtNvWyNr3x3+K5xxP9iUFQsfdCcHbJQ8G8tXBQfPbgjNbjQzv/D2rl+3b/cV5rK
s2WdPAPSz8a/bZyXz1CFRa9QG/azz4ckuYEJdJB3+M+D3Zm35JH5/CK9mzCpRr7qT68p31QLhw8P
MHFPfmETNXB5hajrSSBH6VsqoGCKvhS/2Kb7Di2G3K3YkTVx8ObvLhuzwa2p26Ev/JrsBh7cZPr7
cP3PJhGm0xVM+quWynq2qd9htv/o+lTnTpEsfNUn3Esim/99BS5a+qudUHyUdP95Y2oB4PJnBzGE
nlRlxbFTfl7uMFdqrcajx1Ox7RctHGxyYA039kf69L/M30k3b3Bnnpi8Q5rTlQpp0UDjunVhmacJ
lf3h8JAicBJsVbzQMO97UpMPZYyCpEhu+2/nlT4ZZ2ZIk3xjqMM8w71GQnyh3+jKGL3BruNbzLJu
J/Kzgmg40exZIqY6GdnOHjGLD89isK9Emb4fUfXVwu7Lv0qulLHbhRrN/TGwOgN/o2L5J9IXv/7s
sUp2Xsh5KeQY+yGIqIbvaVyGZXap3uidtSX6ximKQKJQPNirjsqVfozAjw7fd5B0yRn4MA/8Bi1h
hXnC7RWpLRPAMu47BPwI0vmdNz3J65JzdULoZnMdd78QvNAbt/CWl1VCL8dm0UnZAXZQzYWYl1mS
VBxPwxtdqb5YeoZlrOssXNfRy2DhjO7vT1+zUUHBlk5DIMfbXrYwwauW+YarEZwKp8YApvdW4hbH
c4tBeydHs5KWAzZkdGHdNrsf8TJ/Jt32SdAq82tn2nL/R3IN0quL+SsuUjXuGS3ji/eEWgz4J7ez
hJRNu1neU7ELZHnXbduzxzHN9MT03bcZXl+L8DicftSHhlXimLzO4CQSqOq4VzNrJ3/UBYVCG5JZ
8KQgC1veY/cEJgEmAANURWnweusRwWwgIezlef7yy9KXrjXB8Hzi8/eTPrc5T1C8B53ouZnrPsVr
dcHG4TT9lg90M9uxiXGAnLQ7ffjzYYIfBfmXXm0wygEAx3zHDPJai84jOT/jpucsUQg9FCyyoc1G
bFhJGYju7q1X/E6+CwOr8MUjCjeiyMTMkjnaF5V+H7m4FBlGHpZvSDZBRJUQYRsc7X9KLi4zkEzd
T2rgpqLNW1Vy6ODEMx1QkZfZGRrG/z7FYOKyNjt1EYgykDrAXpDDDygrq+xOhY2VCFhNkOq56Ush
nseU5vr55lo3AH5ZaAUH55j6QaVo+fTAEA+T+c0hOfPTOtBx48WbMhmBIZkLcQVYHJekHFQs4JHE
yHRxB0L1y5tqbczib65Q7x1hutpAh0/krG7fsJ19qgauYUWz2UPEPp5/KZDhzMjvnEq4Gv2vVZOj
XJzw2lkJx8wrBwBQwP9/Hs5+H9S/67QLWZt3IFxP52ljb72ke8gwgv52KJaSAMUSiTIbDvvkAGqZ
vA54St2RTmicEr5qPF3MChSWasNtMJ77HXa+N35TzncyMB7maWJruCHn+2OtKRDFMdUagt+w7T60
H1U5mGW1wVBOqZ4Gi8z2EAWVHj2EVAbNxmB4lMN+0PIbIj1AAJn+qIANHd1v8bDPPOIMYweLdSvv
iX4Foe1EwJWhloXnPDdvAFwzGz7JSdkk+8Xb1+0dXoVTYO3n6kzolAKwvz6/kKtDImrhneXIewBY
xGQtYOjrmMZtUEcx+yTmRqTSN8wi4c1/3RHhTjv/p8In9BZdAPCSuUX0aZRIMAsh8jprC+l+2G68
9P0blr0bi8qPwl8I6SQrlecBySXSXZxqXY5oGNgEztPqsi64uKK+ku2DxfSTqXjR2rFlyZY5kDd9
qzg7lTKhZmXj8qs79gGWx+8oqIRf4dkGaiHmmbUHi+jdxIvAi7mSBAFHDAK4JosiRNxJWhyMhlZO
CmWqZp+J7g9fdgHKvo6GFRqvHwxqlXwMwcjw1zuUI0tbUmLhRhdPRCXjqBxqsIH0E7svYGMsUoc9
5KEIOMaH13n9NaDVdr6NMHImhhpcd4B1JQZlmwqBm/VhEb6FwdasqyfPyluumEcS8qNhReu677+i
Dq/nl3uxkZYcCNPUmnjR0jzUUk1bdY0yt5TV3GSSrIeGTp2JHIvU8qETOg/gyweu0n2nWRmEzSdY
mO8G2jdZh7yehxmHYWm0e4u5KZUGoZVbY+HPjabr5DTT3THCqTlG09zYDgMVBLe9tcAuJnTisHft
Huaz2sxC9cseXSG9HWGHdtTPMCSfUdHTfoVySjQyovzNIdAulQrVtr8ZSf9N4wD1Yw5XVql6G5qJ
R1OCihP+wUHGDtXRfEygavjhxa6bOvhjiyb8fovibwsHOZ/LmEinMPLpBSpQ79ADghGct0uyKAyq
CJb1CG1wd0dg1a0YxSVbBCFpAoueencarjxU4iJkKVK4yZIXf0J1Yk3X8tTwBvx311XBihQiCAAE
3M/zad40d2O4vrQhhahgdkorrm5btngFOpm3g/d6LGVIsAzxEDzM+I++KhgDhsSNDPErFZNHxiX5
DYnC2edt2d8P8qmgWBy79lzlGp/HsMjf+1klP2MzwVd0/NDzo+LVo3EVpGuYFn/j2eKTuRvS+uz5
7BRhn11hzcW6SIZKTmUcWcApSY4sdA/Hc28dztlpR7nWQGGOdESc0UByrRaHi7I3i0Ua4gjJSLpZ
/ZS9gD9kdsy9KZiUqiyRztcB1BpHJRzF8r67hrPMuU0/L2TGjA3dWNdS4sUCTz42xLvmhuMuPo1K
lZrwtqO/Vrgxgp7xvmTUKT5oTxbnSQhSi5D0BXtmQ0+PUQio6Bv2sbrcoZRTl0UrQyqc+dmBN/+Q
ee7l0eG3nO85BZLEXlUForv5UEBa262nHYgWm0GWCR67k7g3ECyEC/DHcT8yD3X36xIP9nejc2SV
deKhKrvUVLhwZhhaEp9y/pihYkkY+Kg=
`protect end_protected
