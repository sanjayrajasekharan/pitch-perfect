-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
OUbwvHlsQvFfCJrFq6BfK3ND4bqHEdQU9ejQxhZXwD7GAuhQvUmthovAtrmjxU2s
2Fi2s3a/ooDyPYGr5NYLJcXrrjMpSjojUXL6HE+CcFoK+jg4gIz45PCTigf0PyhX
N/NqdTTnE6PHVA6YOyEIAGu6NFNrMr0mrrwHOET0Ovoy+IwyZym0Vw==
--pragma protect end_key_block
--pragma protect digest_block
U9FzHsabJm1JBA8Nf+h2NmqI2t4=
--pragma protect end_digest_block
--pragma protect data_block
nZ1hRyRUiJtljcdcVA97USga2Je3xeZ1KScM9p7FTlGR9ma7V9OfZ5E9wFOg3use
kvp0l9a28iI+4iescoxTn/1/2pOn/93xomLn8+iOi6ET31IFDJW8f/+Hn3xdezHy
54ElW1hl+J8rz5cDSzbQvburQ0vtksmEC0oUQUgUDAj1K+c0JOXtGP/pKgWq0BRh
ql/Ocjvh/mbBYmzVU6VhqtwUTdESKMNGw9VpgXEzv4c5GkHORj0Lo2s+PJ9/pLaO
OYupVsDSI3JXwozKnIdrlff22ZwbJM5ErZ2VlU2IXIVrDlXlyveYwIxHh37AzKsi
gzBt1O7QWRwxKBfAk1RvfO2Hxf4pGiRTlhbbwv3NEmVA524PBVS0zJFmJ8IPxOES
DAQwupRuNY4kqYFGmSLrXrTAqbphWudzJrj+VjG1MjClPc7/Mjgv1dmH4dI8cUKD
uxfQB7QLsNA5PS++nCzthc3qEcVJs6weexzOiO/3DlX/mlvHDK6cmPDdtOZZ86xo
+7BQxAUskYM2GWIuMe5wmTblV8+1R99DqwRKpY61AiJu6B3ccMcpluwhEzzc2Caw
ivfJkdu1vIISo5YnH/VuuafoYSpQ07bMpre5mYz0RU8CAUHz+MY7oQ9lUJ+0Y6ED
q0vC14le4WqqXfL3ldvQBm5LnlHMn6tMs07Fr5EHziCWfRhaRubSH/ckmGssuv8K
99OWOu45SfktpWOBDo6JQ86GT9erK7mcpST+4hOXh82XQIv9qA+MQYBGNZ+INZW9
1jX//6U672yUNRS1w+u6vYZLOei/p8goCaLfIB6S8pC1whN7z7dMope4Q/pIJdo2
jWSeEVPLD+O7UgtC59B3Cy2jPZGpLQJ0Vi6W8KGdGU/saMeh+CKmeM5ZTydYUFHx
e3IipP/zYkSmS6dmQkij7mc1tfFmTWXmUK0tun0KLi/dXdTzileHYK5ym9/xcRU+
vg9C12LKDWkem0nMb7eOpNrYdxjKoVh/7YlovvTdGnmdLGhUijR9ZlSPIiutlJdC
5ahLnp2y/gEpvj7XgSaIb7dg91KVVPvwEs8NtBkd7rCJKbZnmZkBCuCOUwrfKy6d
v27djXwoLptqE+G82yVn3yjf+/U6t0KWv1eoHeUfzVPCeSlDuVWfCqYBNP8AWZla
6o8kDehWaukw/kT7Y9w0cC/KEZHo2KYIxFCygne0nfkq/0ZnVSKSO7sralz0fGtw
uU5jp/ikRE4AB1kFi63e5vQK5CxZ0AQ1BvMXjbQEn1x+OAsb2ieZwXaHUQXSMWZk
fQoVjhlmC66qvlipWler3wQU26v8LSf+mLoihrrSRBbHCL2d3F1aTLDH2jff87Ch
SG4LCEK2/MHtu6roQFpnOhS6hr8Yq9bfHsQk1nHjHb94gI1afe7cuVWHxJG83hdm
SS3iVWbMnhkHJLh2KEnQ7dVQ0ILu/SN+D3u4RO3gp8Lk9tONdVj3ySthoNOCy0+T
CjEP0/bvWp1yhB9eR3AL43obCGQR9TwCO32sHxkSx2pmPc92BhtMV/IYaUpelTQt
CGVdTL6NFmZRWLVSioU9dXzg3OYmIQPatgmRl8wvm2Y+9OSaonDQMrykJuWWUg25
tGObp9UGvAfkJ0GF4jOt78cWvH2KGxIFKcPTPmwh5KdlTSR2nlekEspJvaOGTfFi
hCDFKUM2zCWDzUs2waBa3gzwltrptety42AlgxWMor+/T2pKI9ufCmldUiCkFF+U
fgTIpkdysJ3u3so4k+tfMITJYSY6yiCbmgkfzWkYF3BpmOqCwHk84fRa94RUFxPL
zrC4XprgzuLv84XhqI0neCtY+ebvJIOwnA35XVqTrzC+JvE217gBASJjzAiT5ydr
myFegkiT0Q0oE/Hf5pw0wPlDyulOxnUXnAVkw9eHsKUa1zj3SQEF9BICjsZSxOE5
yitzZLcpCzlLZs3U/gm65JYgOiH8Jsy3pumnbqAQR5fFMLUbECxbS7StD4f9HciP
Me9Sx/OHcXu56IaSD1Kb718TeKlyLEpvs6Owc02nIsT51GPoiC1o0A8l814Kwg8g
4Yehhon4LnwlRbu2XEcbzHWe58EtYIGACciK/o18Y58HTHYYy+wtvtdFIOvbdDWL
d7UNeyrK74CAUqyG164l+h5F6eZVe5NK7lAnYZJclF5ZmM/PvK0vQ5a2YpAX5t8w
qutpCA1pQ4NrasW6BihGlwrgcgbox/JiQ32uqFbRgSlgBRxNa5x5bMB93mp/RI9L
g604FcTrhkeBg1bLuVYNfNuZMyQVn6PndWzTgy0hM2rAxJTwFUeexcTXZv7q+QIB
7wV07WtwInMkOfIIYDDRhSFNWIZ46eV4L8OwgG822BRk3inePznLkRpVA4JAZRGP
i+aYokfqwEwxUCXEv+ZKrVLfWRYDh5qR9xwZJ4+C5fq634ruYGijaC7v5lPzDswd
BRNOnGl+S3RngHJtbd4M7MrPiibkiHD9FIFVUdUmECkfuENRTPr9cwUAup52umy8
czg8j0gRpzPUhXMciHF+qs6vrgjWNALpHFF9C7ibohj0hhwhmXVfYb13xp5Btu54
dOFDUzRjwveQu+3k17ds0NPg9zgam/QgZtTKZGkoEIYCS/v7vToSDiigO0agxOOR
mdhhkxe2Wic1LZlteE+1gW4htzupLibwAaNQ0hPxdeVS3cFWPhuzA85A2HwqJS1R
1EeA3WqqWbem2xFuWoxkf1YIqczibJxsDMZb7cG9JUMyY6lCqT+yVQspyV3B+CBa
o50Cy5qm19+M16witN4M7oNaejcbUESAxkfrTHkYeJUtwHhK4zpoevPkdc1SJxFr
Vi8fZE0+ooUi4i5y2qne2m1B33HDA27iSuCprCW2QdTI4pUV2Jt4zLI6YLsQ/QtZ
chT5DZrYJxiGqGsQgIZuOmdtAIEtJZqt1C5hgFYz4VXK5D73f31/EDS8PdrH44K2
bBfwpyzhKcrpM6i3hAL2TVFZ2+3dzsXROsHS3q09qxQqtDClEYjh5i7FEr5owTDX
ZcIdV1T1BbC6gj3a8NSK9gg9PtiPsvNZ1pjttFKGtmGltHH6JtdXaEchxc98zy69
jlxHaM1kdynYYECUQHhgiGISu3Dg9w+JdyOymu/duuV3hR9WgxzkAsVmQFx/Icfk
fIXeFf48RH+PuWCGriVTRMHIFxMKtem6BYiSb/89PoFgqn7IzoXAL0Z1mmMxzDzw
8gyB9pAgumrEFK8yTPdnKHSCMWRnmJYWtoHWOmcozLW+jcil12jlEt+S9zbka/Oi
Fj8TQ11fdKFC1ZN/WDLgsSnI+DgMs+8gFZqp8ODD3LlxntqL7QjyB81A2iy3/GGn
7Cp3A1JmUlPNONlmYeNXh3stSH0ki44XZGpXsdT90DmeXPCiOlD/K0toQMYJeJmr
gvIGoIPyhPLGwYU31fR10ug8axq1eY3HU68NHQGD7ja7dv5NF56tS1yHkwBBRrK1
gbfj03ij47vAJSpxNahW2ZopoXfXX5fje8jNaHHwdWDskFpwdY42N5AjSrXHDUQp
ZZZbrwExNpl/PDKprMyh6yColXi9pJsyAVoF+8JedINk71QzHFdAaBePnwfXZbVQ
oE1uTRdipzJ9SghNMM+X6rGNaUMdkubnfjmEZB6ZtYrp0qhbgR2fV1l0GbMODfci
fVRIV7TUIs39INYnsO9lOloX4kGM5/LqHxFS+HWZ0F984+eP57iWZ5cWGTxqweXM
KG/VyetGWTjc9xQZ/wAhl6rHzlIcj0xccTrmJsvXhxZGFoq2/BzfRd5flf09cdBs
TJ6G0+RbqjZVgeF1BCKgFhasXHA9PKKt6/kiaYys02TEx8OBZnmeTjZzvrievTfA
gCW2hlxn74L3Id92khlBUJr6sa30pw1mgUHqKO2yNVuiD+lzUXg53GfJSwaXyIpl
sBjt6dyDmQT3WnunlygwBf3GPOFSclf7XbtdoltZVO66tUAU/PXwmGfQC2YpOoM3
rZQ3D8F/TiSyxR2IYZCYzFfrZzKLuGJB3XP1zAU4VMhZN061RvUMkOL8cY1m+eBA
FGBundFklULHQON8YRwQrhh5bI7rzPE63DAr+VZT7Mf2Fx2tDFyNt3Gww98wFdu+
eDSWk/TxXD6zvLKtqxOJcoYJsg5ZZ+lXyhqUHFGj70BRKsV8ywrbcllw0QdRNrO3
4wa4DK3lCaSeUuBJNAa+po2rnRswAfmRnkYh0oz06vB3y9NvNs7q9xzovmpgQj2v
yymNZLyrBqhNb9G+lvINlWbfVOQWHBhiXwqpDVpY8klOXw9i9TgW6QJxT4ObDZra
rCgRTdDPXCV82V8SPcT+2EGg0nqBKkMKpz4Zzt4RJYmd2+Q7k+D4RT83z512Zm9D
o5IXK0uZPwgVdNvliXnh6GTCS+PbK5mvmfUTakCIsRqxQKIFmmxlVgctqhF4I4ZN
tI/efA9bufS1O2tD5QtHDS39qr35S7dF5mzJbhQCZG/Vojnf8GUZSKWKiGH2iqYp
ezaiPEtveNyqr1jO693AEoNzkGCIlq+lfMcZoUMT+vJ+V2weg+9G1C2o0WpedXCd
20fABowanJJ0gteMMVexah+xeWfl9xaU5D9NNMjkrhBDPirHLP02VgWmpDPLBe05
Kt9jYgHsoUvK9GWHI4HuvGwlnEU3cbZ9mTUke2nnE6UhPYqsBExpzcyVLlUxz6rH
bE0Z+Xcira/UHfjC9p0CZsI8SLLFLj0G5lsuRNTwgc0CYbg7EKyx9OqDGPPu5r6p
S7vFpTMrzw5sVUQtrWKdubTcWJW2nyJVman25dn/+8tLBw/kXr5vFW2o+0EIKk1Z
nIU+94uCPTVInrRqjNxsFkDGXpUyTZ/L0Codoa+BYSYk5sUb62ItxFa5H8YHjTh6
pab3pCvQ95uIg+I/M5tP6MLRKqjIliu1bADS2WaRcJnKIqVK7YVwlRJRdgvcIuvl
b65vM1NaXy+tYRdYksylPFPmljs5uaFlozvfBHG3MgKN6vKwTazxrmZyhUgj8FF8
00DXxoeqnfQMqinV9zkniAyzJliqeVjKXfpb/4u8lFM9cIYfsz1Rf6EmpCIL5uqY
tlNJ3tnypfGkJBtqlLM8IFI0Y1yd24Mhs3JpuSXmib7glNRUp9lX/NJh664eWtSM
q0KSbWwCzPr6KzRKuoRnfD3FT50+y61h7gQMoXFkLF/4csvM9VuxCV/xlQG3sAAT
MyOzV8dhqp9s/Z/uL4emnhieb0KeqtFevuTkT62ET/K1hKIeF7IlCYPCJDxT/96v
yP249Ct2KAMeWJUknABFp9uDikVv89PR1VYZa34cVCsz1k+RI9XJ9WRRjTJ4Kqik
U73LJLnQqRzYGGVVOeSWZPWUpONdO51JHc3jMMD4bN4DWlVUiV1dIYNd+Af0XIis
3K/J9GeWLuQb1Jq3XKMqGLPJYnBCL3aSoMc32OKPQH9xaevJsY7MI6+nOsh32CFv
S3NgbE5B7gmdI4ETViMP14eUeYSXAHs1U4EoGqFpcTi1V2b7nkZMvRnWWLmdRphO
gUJstI1XExpaxQkevu35TSvpeDXz1u7Vt7Ago5l36Ah0ROJHQ4G1KQOQEjguMXIZ
FkUQspWWLckqTQGLtYmPfvRyeanYvjAdhHKgqJPidJSWXlL5916G98+V8OeiuVBZ
8kCYUT/bf24WE0kjM7+e5RRy9yc3uQ+QbSIpB1vidZxuBp4CVEwVLL9Xc16x37yA
GNdYuvpI7dDgnLaBPr/U+LnpAC0aTIcCfbogJJ4ozQNZYc3RedZ6M7WE+rmF1XEP
7npEtewjkzWg848HS6GL6wmwwv04n7ciJAk6nQajyjtHXFGk+fThd8zwMnUp9axJ
q6jfQuVAKCEPFgEjDCADBvV1Si9m+LeXvxin3Pl1/pret6k1kkeRpPYyEOjzg9Sq
IpKu+6pE7ICNG9C5OYmvsZk6lPOKG/xLP2V91G1xQhwKSJlf32EQ3Ug5u/tdDpxN
Rr+RjIU9IxhIusl6GppSNAjPYgqGWn4DfI+/D4x4+RKs7pg93Dny/9pIE4OOniYt
/jbkFx5CaGFemPiBf/Du1yGNVLS5izv+BJTVhplE5HzRej8xnGlSiKvaygy+YkMi
JyMb78OA378fhFTpEH+zb052YquI4GzqwZ9Ur3k10nJLT5WyK944xdEC1qWvBlw0
fiMsiwUORS4WyJmglf1d0LCmlEPCHb8+4AO0b9ulYPQ3zh/CH8KyARkGeoGhLqoj
TE++yCF+bczl3vXQUnKqHrg4nqPX05zXw363RY1QDTtOsUr9UM4M9YFA77QIlotv
//WDZMpQrOidrfORbjUHdnO+bqTNr8R3fD/GvtQsUrGM+O75MRJUkgofOlvVZzCQ
ZXjAg+7j9ni5ixUqpr1CKhe0MdM263/qG7lcAb+YTs40VCJAcLHCMNubJFNUjlOr
qNYEPjOMqtUJrJI+c2pYQHRsJqFftnFfRBOfvlg7oTW/gHg3T0ct6qa86bixfM1S
wmbXdB+miQGsm+5dnJfy3n/BoUF/M1RyOxFol5FWFivabAuQMtLHDkc1A/nF2ajG
tUHzx6cXcCn9Bv8/dhB25RRrjs8swQL7zdElmBsia/VRBSgYmcKuZ6Ikz9NvVMMH
qxH1OdSu4GIfB5Ws6vIC4X0h05q9/iVGNcXqJ9Bx11uFWExsFVsmjwxl2bGHcrYI
KKOQLLS1Qn759+RlAxcrH5JoE5M3CDmFBeqnWOmcM6fBkVqM7O9h22/ew2C18/FP
Cr8DSjV/OOtpTwvhvveKJ+QwF2h4bRL3jooK+yEXMGMtH2Zlg5cS68e39JJMw2Td
5iPaFPIfpVxz5HPvc0QewnIqoSEwXug4BIl5CqD7As9vbtin7dyGtWOOTN5PMsaX
3AAAj8pXjF1HJp03PnqBII9LL2n0G5rvqkGtObSVOf1pkSGDhiPFY9jBUWO7+yJP
PwsPkvFZV/9DJxkmgPl+qzazib7r9Q6UF+JmCpgOMxFpXJcsUl189uRCmGcIf4NA
+yMoJ31D4zBEAZgYtNJkRiBCWaZReFokbLVib+QTDI+oGVuQEt7oPOiPo7w3fKb0
bD5Eay+TD4KXO89ZPP0mb11Tq1mdLtbXj0e11c7nWICdrfUK49iX32+2dCcOd6LV
vSmCSWHh8e6525q5kAt0JtOygCyCEo27lS9e2Ixcui45ceSKmCiFgZllXhplSCDq
ew9mxlJ3fQzdI0nMO0t4PS69soFuMFNH9gaOQ4kRr8A3rM/7w0G9PEkeMTlNKx+l
b9jOjD55eVVQXtSIx8iOojGmA1OQQB4PF/SS8IWWfnlHGbcmO6dUxjI+3/bmF+HZ
Vs0O50BI7lTtXMpzVk1wvtT89xt/AfqxOk9xVf7E+TmDy30+r3TXX3qDyi/YhzIc
boo4a36j6Esw+YZHt+Mswp9m/u0ywf7ZUJBSdnTMWKp1NvKEv2TSBviX4gEMm7W+
8QK7ozWUzBZh7+RU7vTeELZJAQffD0omP+S8zXJWdVOnhH38q8MnPwsZg4Mk6pXh
4SgxC2RE7VEikvc23Bw96Wv3ntCVzlh+iYtJsslnp/ZWYxehrwkRS1Baa6niTbvT
QKESSYWJgLyxhr4xxadI+X/qVPFWxCyvS4XD7vmdUIUmrNFKQw+oQjtnV9Yp/1ft
0rtyf3fM6NK29gDSUdADnRDTv+OvJ0JWrNUnNFHTMVbm0+ODOc2zQaW3RK4aWAEl
k8oAz9fGFmS95QNNcAIlWS9lw6BjNLFWjeiHpfvZy3aINH/wrHnITUhMuSvuOHcw
K0QBNjszn1j4iBS/Lr3Mn1dllr0uknoqJARmYt5yPT2OIiFUYhAJZ5yQ1JUeC6dZ
gq8mHrlhZBMKAJ2tJlV9tl8cqY3RxAlb9tnxZZYJRSxK8rC1o8Nk/4j9mlrqj5DV
GqRb0doP3GsNkWOC+fQn+X5EkJCdIOwrvQphuTjol8Q7S8KpU4jGpRaN2X+rjEgN
YHnry1JUoiPDEVuP9mlJNDtDMT7iy7wKpJIzzQIWOI0RlSh5DUbsJ5SID+oG/KRt
ZxLFauB4ElZDaQ6mKj1ZtXrbfYqeMGnlENJL5iTymqKn0hN0Gd/YutTC7XCufE1m
yKcyq/CwzXYQRvpV/ZoR6LRD/HMlDe7ZuLwCCHzPls32mzmHY01yUYGqxVTdaZ/4
A92Z35qRnEqWCjwbCQWiEf9GCXlGa1qIjTFN2qeBuoVEb5hBB3URZ+D/ffHWvlSE
uYsPD6E/7AdpFgnAK+tM7MxaMBQNAWvHPm5EScaICPjedcZbJDMrJ96t/jIFEYIk
nCRL4I+9c3PLt9axnLjno0SOQ57QurRiNuwurCH7Bp/ai8mS1J/eAky/jHvQex21
cQaNXgma4BGg1PmoOFy0AtqHZDFB7KkfjFmgr27Ihrc5D63jXlAmN4OoUUjfCUwE
u+QcFvWh0EWbK9g+iV8DOmEO0rsiT2Pswrt2xpc/FIsatKFoFd81S5Oz3iGL+ejH
ZlqD2ETFzI7OKhZSTDIMBFKVZXPUuAI9zT/ir7B5PucCHzIFng9PBOFovzoupKW0
z3oxh7u747I/AMkDnD6sHE6p116mTdCDokP/rCkcjMe2VlYBIOzkuxhRzSVW8MGk
sxKdRn2rE5J357kINLlTIwVixE1hxMvETfnzsh+ZztWKuKsWsNxS2+ZaRAz1dXT5
xgYvE60GmMxBGKWEgU/plgc/rFMCSCeht1ajIgs5GQmVv9A/ZW8fAGMMh86fPuEF
X/PVs2NxeAkfZYoUusbSAFIu543DriPeqjeLlO98P5CyvWgnaDsu5+S6Q97OihDG

--pragma protect end_data_block
--pragma protect digest_block
YH0oeuWIwwQvRXLs2Nk/JbLMINc=
--pragma protect end_digest_block
--pragma protect end_protected
