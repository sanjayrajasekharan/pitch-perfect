��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����S�M�hkF��1~� Ά�``0Hɿ��b��i�<�1�SzFĐ�48��ch�iIQ���H����:4(c��_V����&��}�w9B
��T#�_qx35t���D��<��R*�E����nK�N���������19N3a7K�0~��!�@ըfG#�=V�[��&@0Xy8�U�N�
�y��I�S���j�kU�,���87��u�:]q�Ƒgh��8�i;�f��ܐWq�Re�R^Y�˒�
�1h��{�%z��1(Q�,1:k��S�pv�p�$�듮Z�����C;�y�A֚��Au��*��1�-�_��e�(� $��d8T4���z"�������0����W���j�Eզ�$f\��W�t�(;�g���u��A�j(���g.��=�kz�7݅cִ10m�OɅ��1YW��F�O�`�,�w#{�iR�{���X%>�w�?U4�re�C�E��C&�i��r0��vf�8�ԫ�ft�cY!h�����Ϸ����q�ׇ��/j�"(@��c������mI�kru��)��2��*��0�r4�������i:3a����-�������g=���\6A9l�6ιB������:p��Y�Y�[*i�29��w_�\�&�h+!�)�v<�}�!&��V� !/��y17�&�ţ�*�Ҕ} �2]�H�,�nV���˻u%x��[�n^j^���XԞ:��
v�9Q�����3.O?����Խ��@��5�RlCN=ۛR�J�%���oP���'�̐Ӓ�J�嫃C�EIg,�	кOY�y�f�����{I��xBE��e�[��a����-���;_4 �R�y�D7f3�ݛ���N�v��{,��ı�2°K�ui��:K���5rp�FJ�Z �ca�v����Ӟ�onHa_D�ޜ>��SD̈́E�8��>n�X��Y8|���"�UҚ�sq��x/?l��$z~և��NU
�[�I�I, ��^��Z19eA���j�)������s�|m������ǃ��_Q񑣰���c����j5�"-� �6P��z���f�p����$(☻Xns���
SI��(k��ʮs��e\�Ps��@E�=4Sﺉ%E��XD��Z�N�Tą<GE�%>>��߈2Y�Ē��S��<�un22�ef�s���|"�t����P��ݸ5��)"!�0��=����f�͢x��k%g�dq�`S�%b bN�fxU�4<O�d,�Ea� �X(��i�r'�1�杉0T�̊��L#��`� {����)���K�����>�� ���"�EFe(��rV)��\�}\@UXeU+'��B�쭌L�RB���!\�/�.��<S�����z�.	-�u�q�7-ư�=���p/ �<����<.2����e�
��J�8b�uc_�.f��X��.��o�s[#���N�ƿr���n�e��ϟ��\� �}���1�ؼL�;#lAG^@�By��T(*����/l�zT��f͂2�兎�"�S�������J�'x�bk=^F�h�H۬'Ѹ���!�+���+���.�Y�W]��O'�̴Hl�+-x�qF���vnx���IR�ř�x=
�8�s	�ֳ���v��(V�s �s��C|>����"�{�)�V{ #Td=����{��1=��S�1�������%��/	NZ������N!%�gn�o+����9p�r>Q�Uy�|�Iݩ]1�[�S��Vd�</��V9pS��3Y��Eb�o�R��p9>k2�8�F
f�9V3נ��^���z&����p�{��a��O�c��A�\�-�{�L~�%�!A[;�褄a�l�4wR9㹅�׻W�s'����}�<p���ԩ�����l=��Ģ~�!ˀ���^��9�v��E˶��k��sςD�����n���7ɤPK[�ɂ'�Т�'�AM��g�Y��3;4�}��?�]���ɉ笄�jY�Yl����T�3���y�}��0�]j?�����ʖK���"[��p�턓ى܈��aƬ����ٔ�[xߘ�r�Y�JL���r�qO�8eV!$ۮ��n�{�a��SG�Z ,�����~�TG����Mx�S��w�^M�5���M?���ߑj�φi�p��v�l��3���`PI` ��{�d�3��7\��W�|o�_]�4�в��[���*^yA��$���I ���ӏϠȞ�kR¬ލgFM(��)�� _���/�U�sϖ@!��~������/:���_�%T�`rg����F�_������b��Ȍd���J`��؈4	;���0ܶeyN�?_��� @L��iӶ�K������+��m��ĳ�q�-	ҷ�9�!�ُW�ѩV��V ]�i���%�Z-�D�F�N�$�)"٫3��ƼU�d	�31h�Sx0aO��IF6���	�p�����ƣ�~���gT�A�p#�\P�sl����8�8�*��Ǣ�2�th�i����ɧ��E!}$����K��(8�(p���)l���X���y��c����G�=�O"B�	�≰��9��b7R��br��~���,"L>� ��#����B
�Z�@�H���vKٟ']�D=>-�Ц	���,G�=�|)��X�Z&Cܥƫ�P%;Ԇr�>�
W�!3��)�c��R]�,xD�C�D1�Ş�\��,�3?gL
K���݋� ���G� {�<8�������9*
��'�qk�#+fGm !�q��P�#��M�#���=��/���rڄ�kx
��ge�?�kN�+�/fK��S>�=�� ��F弬ʳdTP1��{ӺEA�q?@0������f�3�����oz��VK��k�*B\���k��4��x����L��X��6>q|�lm��������ܡq���g��j������<�v��z�n���t�����u�oHs�q�@��o�wO���Խ�btl�42���ŵ<̨��]�Q���\�Iݒ���ۤ�e_T)0X����{`P.gM͞K����
ry�L�c������^J=���ԃNI��0�&+�����7��r!7T��p�7S��7���������T�����6��C�vL�5�._�1��j�_�Tp+�+:���%a�eĞ�����I��Fz����}Զ'N8Fט5q2�粘�RO�p�]�z�ir���pr
p�H���o@_�
b�ޯ��K�� (�Ȱ �dS��g�o�0�ɦ��L�ة�PЄ5�e�tj׺�[m����Uz�+8^?+{����7^��[�t�|f�Y_�{���[�k���̲��\tR�8A�ZJf����%�����K�f/��y�V��2�t��.�툼{8��і��Ax����m��V�����7*���F�4=�n�2���V�}��\��v��aJ�Zr3+S}�,?:�H+w��R����	:���Y_%�t�c<vܧ�r�w�`D�o }(��NC�=�=�b��jbV�r�>��%c�{������Am��m�50�f��f���y���wMcϡà�M��'�HI��Ag�j�����O�[z6`wl"�1hr�#)9 �	�������"���ϲj�î���ՀIb���'	ĭ{*���y�� ��:�_��Y2Ʉ|�śev��?��������c�_^�U�d���IRxY�q��Ro�s��
)�r�He;nn]��\nj:����~��L�
Z�seeSq�L3�E�eߪ}HXKB27J=c!Ƣ2�y��*���7P�˝q9\j#�� �n,�ծة���-�idH�x�D��:iR[�>�������*SPP)(���;�� �p?��&P�f���r2�.x���+�t*�+��È��M���	<ݳ��8�fy�#Ҁ�F���%�g��?[-�{fи��F�f~��G�� l��}��&`꟩��X��ss�Z�M����8W�?"��$��|ɓ����dTeW�=%ÙETB_%��Ͼ.c�`�a��sE�%T>dY��AKbЩ'{��y=��]�� ������l��u��g4z�5-��Z̬L�/@qi��#[R�4�,_����|Y[pׂ��k.1j���6=�O(�+~��ر|�)ڗ�gk��°��5��.�H��j\%�����`����`�ؽrGM��P��_�h�o03p�����ީ�x��7��Wg��)�g\�����9=Cq�G*�����l��oi�9���EKLk^�B��\�7��$�����Ԫ��Е�B6g!��T_v�@�������fCǣt!9�`�:��q\9����&Pnz�t��1'E�oPor������gM�T�0;�����"=�����/c��w1��e��EfCIĈb����{l^���J�=�nRW* ��%�/�@0f�yh��Lq��?|���3���
30���8s�[�vZ�ߓ";��X�bh�R��=�[[{�8� i��3�D"pt�t��;�w���������hEs%-d��ކ�X�7z�>�H^(�+�xqjuJ��pDֱpx��$f�v����@�l}:G�BM)=y�a�*�X�K+�L�nt�to2 �.M��F����l����(�m� σ%&���� �>߀],�TYr��g��H��Sp��+��C3t��\G����aaT��)��I�Eg��c��g��l���9�y#�I6���q�|b�S�4�d���