-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
CrwHsiYkwb7Zi0BI1HfW12+PwjdOwk4y3x91k1KgLG4yWl3GLzYpECMZqvErs4Hb
YRyYALNzv4n+53EdG5z08LIDToMEiMESfbIjwtossd1j7mluB+QVdNzHpjHY6bOU
68l3z0qsXLXEFNXVsepE2nw/n/gni04DfbEgPO6NQFw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 43971)

`protect DATA_BLOCK
vIpJznFwnr0wL620QnatGbhoBGUaM7769AoFVdBf/S4qQebq0jptk2HkpQFdQsIj
7KIblsUaYevFPAtX575dDXFCocYTAKFlgaSFVpekGztVVJnEyFLew4eWY7GjVygB
yagADAkw8kBe2FT7lFgeeV5m3EqmmpSQSU1DNz2xEKLfByAAnbCWt3ccQX5/0ttY
BcstTEtHNJsnIJNhXBd6UdN3WsJl6f2nVln4w88Eg74gq3cnIkjPyMR5yMim5jKS
IlrlM5kEAxTdBAgglDMfWiF2wO673pDRv8zAWkdoV0Lp+HBFKXIUN4dUSIutwbfR
8anVTiDOuDf4htTgEx7ghbM9WWiJZsp27lm2Ok0J+QCJgAZZvgYeGYirHr/8eQ/Q
7YCF/hlul8nSY5E/GIHWcBgOZGfAK8rJOXRHutjcCZkpof1Y+YaS+DCM9vEXKB0I
dcLTd0t4a208LSfbPuIaijXm9rHNqLFjgRCENTEetNYLr5AyDqTcn1VU5u7qIm8P
qRsG1PR+sF1rcR2F51hsZRdBvn/bVFcDh7p7bVqSNluWj5xU3sRvErTeaAM4jfo0
7NJmpAWoCnjpJwHJpOkbz03cJtItJfwQ83iOw7rFxh4yb2SW+ZJ1OBUsD1BneBi/
5O9WOA069eJnTVum8XQDF/Ti+TY4bUb6xXl6qmR4KiYi5wjBHW6/deR3Varx3gyD
nw7ashJQxnpSpXE7J0D5nvo//+pwjSzyeihMeFmw/iQl1QXMpgkMAkOT7XqQzIXw
epb8c6izGQganNkliEX8qu6+9/a4aG7BkHkJU8QhRDhoXH6R3nLduOdO50naoKH+
ypm7QrEIaZstmSsv3MOepHAIudKTzjNM6Lc9iLrZo3zmRMyUKjMBDTCqwnRYJz73
r97miZmL5D3OTuH1iF6RJ4k8k29HlVDiDPDXn8Q0OvelprL3g/F9BoKCsGqkzShs
wiI/XLAoHs2jUUaUdmdTlZur0Ue9LQywV/UFx3poxVOEMdS4mhaOx9+fIo7ZHl6A
iWZVTzhxH564XxFdMnSk71dDppDlxCuot3vG9+42caTgb6BlZR1L5tmG6pGviYMw
NlvpNR9+QNj/IGO7miZs3TSvli4VjaSxjAw8qmvOoYtUV4TIPewiNxPFV/EFL6da
Mx21q3x10ELlF+909/sQ1RIX+TZtPRjJGLGML62pi2O9dghN6Bg1A1fRUG8ho35j
NnXi7BDz9GOTJGxDgILqsgbkxCN/sBP9Y2w+7W+doHvBZrSbDcQc/wKnFSQUHD7L
Lo0DhVndm3EPiKyN0QC98gP1GBozm2Y9XK3b5iViArhKpjYfYIPNPV9B/nrAEJMX
fq2fqLXS43eMsXsSA4J/Sgn4h2s4u61MlWLalKLMYEdI1zEQ8CFvSQsOr11QWIL5
H2d438IDjNIdBmo1DgnVc6Z8tbwq/FY2Yw1gbGR5R9FRr5pDRC+ojMTqNAy+Mi54
k7IJFmSzQfJywmOVFEltYV9JuLGOr2bd+UuLt3RHTlmmb22Zcn6hcweoe0GL9dLq
GVgrERSW0PjchXMBbHYGjjqkxvn92cLZrjlgYEh07m+gqcxnMQ2sTCZ3QZ68Sg3k
WcwrFp+miynkQ7rE0VFZXcsyde4r7zYOX45Z675IWyT0EFBceg6QXd5wY/OY/KYG
bJkq4n3ICb/GOU1xk3+xTKNiUQ/Zla2H1fr00IvYhyh1fjo4yy9sCR0P7VMFA1H6
0F1Nf8PLFF/MYzhd7Mv12Nfkm2Able+jEovqr2ZZBHdlakwOTPcUtLK2s22inLMA
47vv4uFcWDJZ4is9z4B6qvdGml6ViS6/eNbQGfwcTlxM2B6drzk86LIwbdmwCZFD
dQgXkidyzGI7DN51EeBNHb1r6ISN11AKI8OZmO/y8ysM0juz1TX9NLhCcNirKERD
+DNbyWGeCPugFYVybiEFLVpySHIr4CMKh1G82Nt1LFtbeDeP8m3wHyuKLTGlKtfq
NxZ1Jly09VfUbF8a90Gax32BcifD+smi57YtuimYpfa8xAQ62znGiaI3MNxzAXo4
5CvRBYbC2OIrt6aucZiX3gU8bYFNKMItbv3c2yUAAyMQ7De4YKzsYuQjGloU9MtE
BsB2VLHD41yTC249AY9YdF78MmjAwFjBhSqPv3l3N1WqEzpqG/3TELyLAFSieFCm
TC/5Mrtu6OI+AONK03nstlN4Mp/3d3FBgxpLVJZiwxOcGaxlMRcobWkGf3CZuIj/
37V1w10a83MKWKqFz0pJ40rrxm1oqSNra0oMzg035Ayz6l9QUeSN//oXvQkMv4FM
MPEt+6A3ioEQsL1suX5N2Obrzksy3M3sNXzrdGs8pJbA5y4tw7ih4nOnZqpvYzeL
/5dKNHbbt2rK0peE1m3+Vm9e2Q68DarcUnHX6gMDaGnrklApRPaY55/Fer04uLt8
dZ5iMoOL6cMXawj7kyR2BUjK3gKE0HZmmVX/ZL6ml1jwyAYtSLUfuOYbBYhS8OjU
jFFB2jtGMOIBkTYR7PK+/phk+HUY47cFrhnzt1SyQReGURlVpKj+zAGUxTROBP0W
8zNh8TpVlc+eHQ8un7q+z0uBJJqVyxTQlf8AWKRg7tSviUDNywjfn4t/RrY7FCne
EXh+zdVySugapHYwKqJXaj9PoWVrpqnESLHBDyX/m0RhwUnR4KsKcR+RKRqgfFGY
KtIXHFsrncLQBFVR+99GU36ml103gdnmqpa2NDQ+2LQA1m65UjsL8gg/7i8676+9
SnJf6iO20RfAahn/Kh5sXvcKzzg7gz1XQKraoB1ZhE0M3Bw1EuPxUIzDjud83VDK
BU3Sa71g+dO0BNOJPmLui9uiMnZQpmpOGMM6CMptFGEyKaaTfap7sovz6JZpGrPO
c5jR4oR8EZhrfbHSx4ukxx6osMR67vjX++xNYN6s1EiQaI8Fpq633G0kH7KxWFVA
rD17kBekE7VZInC+BWP27BK+XlUoOOETAdjvZCdd+HN7kBkue2HdgdycjNt1sFMQ
2/ek87osbWdzuv0Av6y6pirZBoTZh064qRkcvR6E52uMJDTiPb8W9dk4y5FU8TME
WC1X2vdfjSa4zWAgtwfO9D3axYRxRgqXT3Ad9AucRH5/zMT3FW6eDiN2PN0Jbr4c
PCiUGBdhor1pInazOrdhm4o1inQ+V8fmvy5ivDzcz8rqW+dBxPCp6n423B1zmv8U
Gb3bN3sCeC81Ir7FDPADYefDeqpFnIGSFdgzYdbLebPsZo1kdYYy6EL+6X+CQUiK
PAXVY5WfDMeWZkOdtksZL5UAcd/zY2qSTyn06v8dvVbuXMXoOenOb6a6bGljOSuj
jeX4g/QcDixXmQZ8YZRgoZ0Kh9rrJL/akxE1U8vh205dDPpsqylE1CjWJBPyrRvm
Ukp1e9tmQ8m3nLLv5llXQx4l9P3n+3SXizG9jm/gQnH502/zF4WBX2l5pvfI1kem
QOptKhhpUxhbiA4W7hAHfQRJKH20QJeyh7Yljn1XOVnWN3HXRanPfedTauodVLED
91KUIM1u+gaNtZ0hwrMkIazL0ep+UkkhIs7DoKSvdFrxl1xABET0RbpYAQpdZY9R
ONU3e86SEPHwurpJQSsEptgmpGG2IeMu+6tqowsxCdtVtDBNaiwYMn8AesEKpfFy
3CspaNsE+/Ec3ORwi8pCAFi/nP1+te6lFIOIgydBOOZoN50zTaJItSckyzxJGMmw
Gt3d2rDLLgu+64fyaIpxrIe82sMHJMyOcB22fSsEUbSeHc17H/vLZWjejbUYkn4A
KqI3ezEc+vZe4Nq2nU3tf6ctM4/wmByI1sLJ0tGYm5tQfR0E5t7ucqen1uwPmzwW
wop3W9N5X0f6qKfdwx4tndDvlYwVtbNA8U+F3ut+O8jhgCLEH0xcdjC3xZKvYB9t
OsaqPH0YWhfj8wTTDAwy8ijbBJ6Zxac7jWGE3FtSAtiw855CqsIPq22iBAl0QM//
a3VIfOqTd01HJqHOyWGM1JqwhepuzWe9kHYQGLCD5QaocMHFv8Q/T1liQRYhu3iY
FhiZ0b69Yj94TpvHpokFFOaZPybw61DimlNLTFhm5Eub+uQdjka9+rd5+/KyQPYI
QoMWD5nWntyccTWs55rMAu5aKefNjwxVXNccn7u5z2M3k/mNv7ErREDODxvGJgx/
YeNoPDpmm4mTLkSrpYOWgzO0qS3Ef0EbRk1C+axD0h1GILGSQ6qklRUc7fvGN7XL
MrriEoIiEFwa9jxzUHWj/9+eXaBgE2dH/vRqdv5XWrziVfiyUZiGpplaSk199du+
f653qUzCIA12WjGMAWfAVGxqacfLg/CD042j0wYUloR/L4HaDXPFIa5UDSdWJ2Ct
DSpxCALdruTHI9ZKKy5maKF1Iq2/xt+SZvYwQluTIpwOmMXhmyZ2AlrkUWKG+zeY
jwQlVGyZcscUVVmIKzutGcasBlQ+pOC4XzIhlDjcRsN+sOzVRdtJ6HETT3HuXqAr
ycFFk4jWb4+pB/e05mrvD+AcWlIl+/nXGl8S14zFIUoX7yoFPezXV4a5kh7qYzV8
fOaks9cHW0FFgtUrjqejNzQ6ISUzAHd5lopz3ALA8eE7vILGK9v2GWlNvXZGtRVl
hCxdivmvD4KGSHDFhenk4HD56azJRgMSp+a7bXP7YRSXl6Ol69siRvDWIIm82SLG
TdnAYcAPcmIN0VQshYqbBR4PwEJn8Du6DRYVBtYzuhqJ3FrJBpPIqe1AbqjdH/Tt
TGnZRJ6DOhMOEypV5vo1lYHRpNC/1+91o/MrpxeMcycGmXD8zphqUjwedVB46L4T
iAkWJ1Q1KtILHUuAdgkq2tET2h1KweodEI9+P4NTibvCm5lwOZU2XuwzmoUh1GiU
OrL5DtTLiEQ2hZFjjsRLHEBlLJVrj31aXmVotJIVb8M6omHG3kV9Vyh95IE1vncG
Sciz5tHh7sKgnvm2Xgck23CLQ4ofYuOgagEoKQZXdpzxtIxNXn9iWJP/dSQI4WjY
LMBcCB+uddtauJume4dAxDITQ+LFqNaerihbrsAAPmtsfmC7cj7uUKetd0yJEYTT
NONdB1ctKDSiHsxhupldjka0/1UiTDwGIU+kGH23XNLwch5cWzghX4JTyJIBKjjN
GgdyVBVK+UYbup+HvkAky7v1//kRWKbkqn4pUsR4I4um4IuYdUTpqN5/IMfI+/Fd
AAXvwTqZTqMGEf705tnv0YZSu7KLepvS4B5fqaCtOzVTCFJIjVtYrlY0b90hAwY5
3Pa54D2tz5Tzjr+fHDNTydrFYpNKAJwkyioIyOxa3HYXDITkiqf+LI/wYSnmr1dl
qoyPl8uABEoUa+DbAK+YGNIdhdTAQ+UXz8SUK7bH34GKI/PEyyj3D4SQfWlW4e5g
mBIETnE7MX524RQ/CrIyjmmtSpL4VONDTp85ZM33EMcH+m1Y0UkpCIXdEbI+jTEJ
E3Pk3VsjcD3AxF8K0/CXrRu1g+QHnxBex8lEeOCGXT1NRgIAisL7uF/viSqAdVpn
KaV5G6w9Nugze5fNM9FfsSby82TTbJs6+B8PSwqj7UFLS5KqCPv5wx6YyNQl473Z
UZZ90et2bs+ztd5MAoqT8iDQU0ObJA6FgNLFgdWPLDuDYSpHAq7wfCVK73wCQP8X
Z0s/SR/YzBsgxJb7hm8xiiD0bCkuqbcaYlXiQvu3wAvSGmcNC2qOYkErxNmY+esd
8o8mu8wGXI6NjEmBXJjL5yLi408vZ8mFds7SgvZsvbASvzwqk2PD4r84x2Mp2gkZ
+svc8BtYAYoQJh7gffLhXAgoye5EnReHbftcWepqWEqUZfhfoM5qtT/k5Nb96vIx
6paKpftY0n40CiK1l/FIgRIc8YzeM6i9u/l0aXU5Y6KxXoW/uccF2O44O7p8feJ9
slJLFvLcZ/L7wQvqcVwc9xbnrsMXwWAlaaAkkZlk62weB0+Drx8TTHTQa3PMKW1Z
mpxJflwwMEW9HOWWuwMrxBxrENdE7VA8k9Ikz9hpk8Ez0SgqT5LZXlMIfExMBlIJ
yshfC/NYvweUjxs73dly/f44qel2YW6YG6Nj9atb1EY+ft2+e5AnLQZDMcs2gdxE
1hXbphymEbPZp33wRlfUCACk3/mS95Sh8tzXf9LqZn+9EtUsBgncsqv8LJBeH5vn
8ScJ1KgD3D/t+ltA8x0wTd3wBK4kTXqIuQIgKiyH96/R6bz8POOODiQ+LolpbWdi
5PyTKDt8FCdw8Pu/YgPnJqh0b/9XYuhShmL3g+9z4VN+yMoVSHMa6LQMVkBpzcPU
boizBMLQjeF2ZmMtCdARCWQVn0MpZzp8wTFm2P5NKPiA7BBOHr4aFyPfZ4pcfZqo
+vSh872Z0HUxPStO5xE+HmlAVlkHRlBWxQXvN20caKpa2RJAEHHEeDCBjOwUd53n
grvLfo/G+fTWOl/qaK2ao3BPG2kXNlGXrt1Hg+rQyv+hLBVPq+GSDziShDMvUbzg
xwOb9gjbFkvYYV4b6b899SOdl5NLVwwmg/S3F7i+Ud62BOBEecdzJjbIOATPR4HN
K1fCtudoyYdzFciD0vHL5QwnivH16VM9cGmA5bt43CKY0H37kuZPQnf4HdYEr3fY
j3YtE8/419dvmEv4SVMOpxFRnSxz67D2dIFKKcnHE//cp6UxejlJgkClzIAxerRQ
uOXjzAlektBaEoLJ5jao2IRd1SgE2pNYK+M1u25OH+syGnhPEn5jTV5rUcN+0mIK
TpQLS/IqXauEoNlnuSXEpohEInDqFvzX7H5X1/eBDGAFo3ISlcaB3y72IERRC760
UsTS1/LaoPYKKL83h6zWFgNwajAb4bIjzuvKFmNmrt/0AS88YbNbJVa2V8iDMMuX
x0rBduFYHgJ93qAPxWEuJYDVmTsLVNMsVZ7gDvEofktL5VikCYvw0QUa+ruZ3UcL
daAZ4b0W/OB7rny/3Lf8U+VYLj5tHkznbUkSV0FLfL9DM1IvbOFhEXjtGy94KeW4
bpI/OLXpK6fc0tGurqEXtI7qeDJh8+VadQC+g/Xn3lAitMTys6tLowBkVcdsDJxj
wEP01cVQ5YF3tdDACDDlbRP2pSB+GCuY9qbLl/KCAdZ8Oz9HYJu9tnca/g5KgxFo
sUZPdYWgKe3HoiCohnURxSv4keLL58HXiRSAnnnNrgOFNTCJ7ZJn/daQK4cfkjxj
yU6xwH+D0SSJZMl0xIuK5pKm2VLhPkGrPVJdQvMSoITt5mlr70odZXoKjC8tvvfl
4YJiMYNzuLLXpoaTrzuEED6KNDJpOl3dDNJBH6Mi5s42zeeyuWZBOXw9p7LKYpLv
UQqAdyr4BrWXasVCsdP8Yrq5a7HE/x077t3H0RAiXYuzJZnl18GleG2kWIppW1Ur
pyObXFeQaPro4EX+2n3L7e2Jqxl05lJDb0O4TfSZnLq/xXb+kmQR9QPHMBnN7S5+
WkhiZU8PDMvqtEIdehOIEoxY95fDhzCiWJkhwJNQZCqFFX9TK9W7D3tryQWhYLzR
gri34l+yKibpym69PSQ0axaPE26Rt3f5+qnrLB9cQ4cwmxYDUoPxixQ/K27GSS1k
ddlaNZWisf/zUS1AO81CGTUTeG2xKgQE/FJu9CZh3xJMwdEd7ARB4UzjUrnK0s0p
q3+YhXBTjLH18XZ3vS3CHnBSIoFgwL58B9xGIZnN+S+2SpMRy3wx2ugqo8X4PDXz
F2JZJpy+rCa3xW3aN81lxMSJ+L3Dyubr9xn985om2PkUb5TXUSB52x4vBiL2xBKo
LuHjIJhFmhhOifA1V0pE4fL3Tud+NhBiXOYBNK82Vu797TEzklake8kJgXFDFNwN
TcK8fZ0xvstolHKFdfC2OJlmIud6j7D0q5QsnBVMBRAPRFKp0tpYMPvoXSKwY3B1
4+j9Tlzd8KVOM1lUm5Dy20nEZaH+z6O4NBBD3RZOhpmAMPoxsopnelaFdbdvelRP
m/Rodiw0NE5p0hDlUIXK8/oJykjduCz0NuzF2+HGgwDbDo3OeHHDW+8a3IMgm2x1
UnPzZ99wTgcEjPbFCdDpoRDdAmsterPtzLv8YQfZmfzpw6Z16AGlgJAoW1YZ+hYO
n9U8UHOJRC4Z2u0Itme5htl6qyQldwCs+J7QeDmGueBi/yRHpNJkhWwH6qYaFZCL
LXlAL+b3XSMyR/MNptKhQ3hOEyO5kRHtIjRZ2T1afk+GqSTfAfTqUXOQ4nWHUdaL
vmlzFHucYmeSjuoBem5kV2XZ8Kd74uaswaZk93KF5E/Zf2SjCcEmPCje8e+TiJyr
7qWLEEFMzpiOZhVLaXrnspEnIWoJRUDF0uA6/AjSnx4FoR/liXj4hlb3RMghD5Ug
Vb88HU2jpJ9CXM9T7X4/3E8aVaUY4mgkoOP22JiPuahUHuCUgSHLEX097Las6xkD
WaW/D5MVeLQ7L0dDUS190/UCe9P25Bocw37nG8FX+c07mxA0/8mtIeQ7cHw8nzvA
2SGdkP6fAd9WHDvw9Mjh8LAat7GiaYpsbZXpP3dTBow+tedZpHbLzllSORC7OB9x
6vp9AhSOZN7CPWZ2BNfikQ7Tz21xIVV26hN9q3R2AWN1ih27glHYA4S4+yf56gts
PwMQg5yuU7PyVUE3yIttBOAEC9gFV04orgHjlyXdwhWGVGKInolfhJNGjA6S4s3j
YLP53P/MxcXiewhaWJeTT/yYuwVGtiUIOMhHgzAPAIx32jeETlIncBuhObFHgJKt
dp/MpXam5YlGa3wxxpyiVzDhvf8LXzvNkYB4TOkREwSMXecvKQqXiNYvMPkA8lYY
6ijeuHuOc0EdHtZO6xpZJjokP7P9weMI6QOsjUL2kOFEEY6b83HJ6mRQd/o6Dy3E
Zk/ck36EqiVsevpIeBOh4GXo/1qO5Mm8L8z5SWjRWNXy6XJtHYMu0+/Zn2EPo0lg
0nDCjRl405Q6mVo8hqH070v1aEJDRkmIXcw5jZ8ya2QqcHblTBJGHeTI15X+lmkM
acTOZ9PFktAAwt51AgMeLVB8nl2vd0tB0GSwTLSwUfxbG4j9wo2erBKZPX/2dPGz
X9J7mmzs6cI3QIk2zKNSxKBvpcMWTv3GF/6y4jJp9bqHmNuhHUhqNGkZrVN3lEdB
Riabn7qh8MSVJeeopLKTvwBTp0prPEJwMX2dExc2CZaMJOvXguTmr/wyCUbvY4o/
Gctq0F95GySFTVcwPdf/wZ3XDg0gftGaBraTXegEmbL77mc2lSEpwaBuUvRr+Idc
zWiidC/nejHnCNcktRNNye9bqoPW3C1Wv+P35uGtVcPD665HeB/MUU3Y3ggYKJlh
ldwHgaOeK+b9qPGKLSdDW0R+HkEjgWDXRrNh3oEywq3TTnGaw1V3AWJmnpzNL47M
2yzey6FLxinwNm/B0uDsMezRxDzcz1JY4I54IphdJ0ghL5Zt3mqJhc5p3QkCWMib
V/bXlVkpKq+59/xes1KbU/wGt6FajvPkcLYQLJlT1GD9o41IlgR4LXsQ7nNPCZB0
2r4666FSQ86Xa7py4Me0ak7nBdL+ip8tzhKZ0syHcOQuDIWopYkDqglfl3eyl78W
NTd3Ob1OVCET7xlQMrQ+IToPWI91QY0NYCsApQJtXdlYijVLaoRP02En08ahY6Ia
4jFWh78iUKoEpCuedyof684tcAARUH+JRPlGeb0Ex03flOrSO56dfr7XJfCTiRXH
/BCFZmCryPq1J7n0H9OTuyw+iKM2xCHYWqOx+Yw1rE2kF0JgxN00vsK5KColsP68
f46jn0sSRmEsQJISJu9ZqzasDCNz+l/Kl4hLasbuH1wHOEZ0LAshrqindlGy45df
gEDzj81IQ2Wa1PP1sX1wIr3LAYC9APEe2E47UCdg9+Gl3tWdfsYCOQ8fBCiMG/o0
I6/9Ew7Pxv1w25DYfShiyNFVvC5XnJDaN1u8Mqx/jXmGstzZLy7eX5IE2cypdWXz
sZDyUgEWi5flX42B2+yChctKSJ+LXQc9pvhfN/5lb95AEIAsMuNKhN07K3kS8HS9
JWp783SYlGur5UeiTtq5be1uW70uXq7atMuDEGvWusO7JCqOgDUm9dOO9oFWC9zw
qELJzcDvd3jp08sWAVM2Avl8RfYcIIUM5IVQe4/fsSvM8cavKvWFEzVKnKMXnpjY
b2LWygL9srWBVbCO3wHBv0jpTdJJcmj4jZ4WpGOZg/Ei4dtNZ1tiimm0ctiRq5AA
3jMf+9sqnDxaaLpE/Q2lt7LcVtEx9hSxZCTiYMCgCthz+asuf0Dh4yvrLgF+mMxq
4Z1s7CmDdfu5djzJCRjFXcjjop/PMG4SBVvSjASUyQJkirs5aEcqzir9R6HPMkrg
lrmM771V0Cb0gBCQ6zCr/lnOayBMzcGBgGsIim6GqBRgDg+HXaWmKzpN/VfrFBP+
B9eZWdlqAqgSeVNi8+w+HiAzIhBlCKQU4IYWDH5Nvtnqp7RWAq2cc0ar+lDHfkNh
iwAlABxqQRktWDYytCMBaB6b7pbp2qrpt/nngSbWHi3uMimvD7+p6a7rEsVgD10g
xcZpqGInJRIY6iqShumcJpskpsgSyBQhvEVyS0QIz0Wlgwvy1H1tGXU39QKyl92J
vHNKRsLAjYQpFpTFH3gmz40DPHKeUGanQd1epnHV2nGP5VbZFbARmN/AoZjl0z9I
+WYXioPNRScpCpvk/VSfOHK/5szDmxX0HlUtzmSJHZ/O+JTIV4Pt6ugEYpbCGMec
NmyCcmEksbv4FGj5TWJebCVUirHvCwWJRc/wUH52G5A4IKeEmBxOZmvm2PHCHqLt
R2zLrznqKoA1QwP6FsG5n3IDnlDmyRVQUpgveLsi1eGd2PpkjxPFtaOKRpB3PaH6
StoFX1b6irdX6y5ndY/I2/MSLnSkQ9ELDfKN+RKC4Q5PG1lLuEwR5OIovaZkWEWW
+l3EQd2ODD5EaHPNdx3M3Lsm6vMvYFu+YGlh7wDt2whs/tiwb7too3KU+5Dr1qxy
/zoBRGEoP/+oUbjjAG3wv29F1kD6iI+P6fj9JFd9F2JQHFnFX0BLlFgpy+1yFAnn
8Kv+W/4jva/h6H53g3i/bLkZ3c7RvIyuhd4bB1VZ2HUT0vkbzz3tGRAVTs+0cNKS
E+Rz4tklZ7JWJyDZItmnDRZbuISCtkXZBU3iQPwXEKgr8kO2lx2hi8ySTWYBqu+i
SS2AchHVgQi6WJw72Pv904r7Vp3eLUHo1dICUjId1vZjKj0tV7uUN0HaphpFnbqg
eX9Biy1rY/cjMcZaZtdLijwOEP4rPJGOJRKKiSUhV9al3rzn2BtXzbe8GfVG+dSi
jKHvWKNF1IrX51xElGpIdh56KVKr2YcUSObNq+18okS0ZgbNhJDC3lqxOXeNJIef
Gz4Z6HBK6uyL6e3iSMS092i28uHEJ7bK0GBaxQvu/vB25lNlNcwT+6wpf2+mfx/0
AfQM72AKTOZ6TN25VMjNQSrPdBm7sUZuYtt1b+dAl6ZMbjb5jckG5JYr2S/099DY
BsWdqDKWnBL+jt0uvhBGmOB5jhKXKDyBPwV/YJUwc+PCxoBd3aFvHa1ENj9UejY3
ThDWcwjTXw/RZfvJoYqJpThRf9CgCQTnleXNlx3+o/rKqUF8hszlmO9c5D6bNVZt
qM8Ffv2wkdeUsqs8VCNg7m+lOHgbQR+0mdmIoWknNZJxIeY6VmWg1bRdI8iA87et
Cfk14XAbXPQZOIkPX0s2UnADajlY7YuEl7/C6Nxd8NhcRc8HCRkXuNxhqwfbrVBw
ibVqb1+r2BaqnTvPTd6hyqyvsMS8h0vSGyHC6oaHRlGbONSQ+i4kr+42hFl0h5gL
vmnaalb63LK/I8ctgXCHUXqcJCIMYgLvYpoYJbmR0fsOXofWiFKo9BOR7Jg9cpGh
i+f1/VQyNzkv71e5yLT+BcfFaMLzcp6NuRmiOGI2wqyTagfSyQp4b7gEZ/WaLe8S
tyqF16oy5IWpvueZIML6jZjx/6CFj4/GwFSMpY83deqnQ+OPGT9rk/Sots6D1xJ8
O0GC7x2ypKthu/vZwv8FQ+IFhUZpAmauVSc/PQZFQ6TvV06/B9Lab8g/+3KKSUUe
NefFv3EntzTuImmOff1uD9UaFHz9nPjhoojPFKRGC67Z12G/PJgecME1mmM/1TNq
qniz0AUMSaX2Vt8sc0LYaL+z5f2I4GfS5FQmsR2BmDeQ5R4xYQhqNF1VL29Eg1W6
mZAqPj5enmMrBvLKCtsqtDbrAwssWiCk1soImBuT2zU/ImR9vOOxIDvv1B9tQ5UA
WiU1WTAx515op3ni5TzM/sSqOlk8yIq3sDiYgxh8PL+FbDxpjyxluvey2Xc1IQr3
RYAji8VzMUy2L0DlP++DkzRYbqWycMeenqlMnS62w7W+sj12+g9DEyPAU6OPLVAL
k+vvWqepOxSmyr7RG7ulvU9hmXXHMn8xgEq+hXBpYXPnfnEstvuGNax0ZEvrOZzH
bA0H7fzCg210a7kbBAvel2r1TodwzN3NaAnKyJdDIDXEeXtGPqMopddu+X2hA3Jj
RcJ31IFYwA5Y3t4cijTNVnLMlZ/cvibDYHuCRztekIDG7Sm+DUuv437fuPnf36Ps
itkHB3uaz60gKvvG8Sb+gXq9wDWf2zcRS2YGVaQmZYAP7Qsd5jjlkYF5KAwCwVYO
SpM2qTvh6peV99ZD18Hh4pSI8rC2Ccu+OwaWktONCiYiGzaqZRDTGWdDngKZISpL
ny2Z6+ZyfSSqUBosKmpQzxGcdn8nwqOgMBEasNUa1p/odEbEAd73MEcXc67HXwJt
4zk11nCXKzeuwyM4V9OAuAtSl6XULok1dg/Mk190LPsmlLKmGcA5cDDTV7oHXqUm
sTtbixVD/OxYBAWTY7Wxk7DKbsr0jHhQMTTboeF2pf20ORO8Lwl3rtnG4xxMljjq
T3pa/gloNbfRQRcTGtbhxn/fxq2VpcwN8w7xnhS9FBvKotxvB7XI4pi3oqM+Qorr
QMm7GcjtZMCDrWDpVgd2oPpsdnz6WFltwYUPhs1C5THnu/10htp9jaZCF8mvL72t
Kl7iybqX4WYePX2b8vzSdPyg8DjOZXmrB768gj0o5PsBtGpnFgcExhAl60r6yuB1
rXuThpfmGAZoFolAyoHphy40t1dYDFGpNqlyQx4PrYQQaaWCZ/ELdUTpQZVITKvs
F0JvDr0M8i5CZH9omy4+A6hsmAyQ4H8xxE/yp8KPCnY3RGczwyf8pD8Grq2YuVLp
nZ3PBOxlZm2VfUqbp9rOSrtjIQcjYP/t7OAZUGR8aMCRNL+Ko6vp4257Hu9U6HSg
L692ya34NgRe2g/Aby9Uca2lCJzwNNgXrWbpD7yTdSyJ4ldWdnIDFhB2ptFw1ohQ
cl/qILfXFEifGbTxuPwBhheceJXCCAbWTe8P0Aq1db2kJDWSh0Cunbm/LaTa3obJ
Mbhqr38rjNvHtC2rWVtDU5pn+qGXIczo2x77+inhDhg+hAe3j+8KhzxvH3rTtiKj
hMUA6e1OzTemULgE7jGnq9ylPxYOYKm2tmNXuOJGpG9mZCsNdyGCOvUQwooGD3o/
/KUUZC0kuavtFCj7VdHdU6sthspHokDmNMRgViE5fZ9FX1d4lZTXBWHcZZu3JwO1
e/fvJukpI4wQ/gccSqSnSM0jg4LnLBUryu40tB7HP8AQ027Y+ek31k+JJtpCilxd
R3/Snayo2+pJBGXPp/+WcvXa39/nYXgf7kqUD7VRFuH//M6ZvMs7wImL544fZln/
G91AqtA28JgU8ieie911KTJY+TGlk1X4pVxwzQMZ/NhePP57Mh4m/FzlzwYyGJgI
+4KTCp31U71le7083kOLLPgeVQlAZn0HdUcEQHTjjEN5pUmNfPrGmbliUBq9b0fr
SBQlJTJVCE9uwTldMyTYbZPPW8Qbq8JctEmmMMo5kjq1sfi9zEvDzUND4kBOcG+9
4SlZf+hQf3pr5+CORsTlQ56cU9TD3n3wFEnGPh/tVX3z4VpKhD8irgQjOJdTnYHr
SMY1Sbem6DrdInFs/ZqrrsMK1J+Ztp+Oo6U/LfUtGAeDC8xQ68EnycGmp5NkEANI
s1DovH7WOPHR7LqRPRgi9sTQgBOc8qtBecBQLWg/MDzo38gChXOwruVBtZ+DBd9J
tFu4lniXpijC/uSzSWWOXAXGm1gteEks3X8uU9E8B7Rn7Gqw16otzWyWMTipmHZe
+tP0Fmh32UlGmUyU6vsssDliYQ+7R7n7BhhlWGaey8GfOhTx/ksIfSnw4GS76K0X
mKU4bqSw8fkPuDHn244t5GVMqLfq07AjYhG+DdEoZ4sZtUExL7oXBeCDgLBkdrz7
iZSebsa0i9TBsd31U+kZtckY8XSj6QMbznFBO3AkDDJqeB8D8HTt194YQlNuI2Gm
joCyc4c1E2lE7wMwDQzgcBc/q6kC8rrZuu8mFhf1M22zQbiYK49+dyHos4Ml0RK7
4ikddwkb75TzgmjYXA1dapnbmKlV2gU4wxOycs0hfnIA2xYqCG2+glbdBRWKL5gh
seb2Jf0z17Y/93423O8n8QAJVotlMGZgMpcAZOVRLWBTTgqb1jB2sX8JxaGZfzgC
zmLHnD0dmIh7NZ7yo0Ae9eYSL1d71iW+3InIyZ/8vDEhbAY7otPcMOHh0792f74l
kOHqj7KVWbyrsF+LiJABapDZbSFx0bkTZKtyUHJTKLQFTrcCv9GECmPgutkFt/o/
OC8p5KZUZr6roYIoJOnbkYCSNREhzGGlZ4KLbvBNRm+KRreTjXXPW7VSr5rm6RPH
AzDJL1cXYyNn2U0btqNXLR6VXovxzl4o9cYjyJpWED3NIlCOp+7XOD+aC+6exMA8
haCM14EIoTZwtf9SgAQK/X/clv5w63DMTrjTGKoZEi6631P79ZZtJ6oQPqr7+PLD
+Biiidlwce8LL4R2cU6SwxoN0qJKd6pNxR7sTkuwj/0UXqO2VDtNPxKjPrxwdGYo
V/2hERomPwhHKUJ11C1FFvHK9MCjuVAUqScWMuspUwXZvV3IUdRov1VDfM1FeBZU
2O65wR7tDlgOD5KrPgfRIZMwrs7sWkYfPrTOP4GKBgOTOTFSLwXNYuPY+0isMWbz
r3kwpOt+e9r+ItufsbplD89g9JtTXuwOe8vJJsjcx4x73b8itsN68PHUaOtcIKGr
2TXRqRGLAnkRvj5bdqL7/Vxyt6cMwUNzim8RWcXOFFhq/zZaT5oYNjPtNKfhJ6/l
Kq4dj5SYxKpp9HA1hk6XpeosKOTCBi86Bp/I2wRTUAGRCjDm7qkEjhjhHnsIsuGl
Dr6ry8S2UebsltryclXvxkjYepatu7Ua+/8P9mYEfV6R83KSHNSRgT+qh7ZjX4B6
OlzWrwNiAxKFhvy3iSYr53fDtjPnhNKRW8blxknqSDD9M4uGgxbHefuhr2VCmFmt
KuB6pf5Y7mzSKtFwKToYcJG4pGyaf+tJHN5eLyIgB+kG0Bmn8BA8x7Lv2lqaM5jP
WGz+93zDC+6mONitE4I5/iLQXa4m8XT1Yx7Hfxs4iiuUB7nkB+mdehWiT0eIssWt
8CG8gmOwT6A5ze39EFaqZ3aSSDP8KIx0O3TkUxVv5XvmxzVHTpbZ2zakK2MnoCZK
MOuZdKbUPgfB2yEd1KTyP1m63CNauQUwOYkVf5TGMyeu09dUbCSAvZ67UFpjMl+h
fVzYTGXEhE7JGcx4XldkP9bEcd16fVCvs77IC+9n81p6/NWfB3eXDLbmYhUwI7HE
rETRFEJvHte5XzXWszWg1uLIUaCAZKx/oViPyPD14WESut3ZWfZ4jUpEHAQIHbJZ
0UkMQLp/bnlHIJdbsTUxMdx3WXJAQn2qlLw1vWR2Q9eCebtbzpjDOUtpiFy2d67Y
FzkUPMq1F43I4wa0VVcRlyAv8+KYgAh05KHGdgTUGDcyc9f97wMqFdXbr5CutKXh
a7fdeAVyMRwqIyONrnRRv8gqTx1HhBlM0gRI8AL483O9rGj5qrN9F/fG6y+794YS
iyzaMs4MRPGluJROq8g8OZQfDXsKHlcVQHrtUVe1mKdasSxRrPWsGfboHKlexzG7
Qw1L0kAuwmYb8zs3GRMted0pasHAqrtTH0vbsRQdJJXfojnNMMPy5IbJo9Q9q84s
NiCZk0l8FJ9vTaS0iZnZWhXoOa09XgMV6KtcHSOFp5puiKbR78dRMMWChzjPjez3
NnrROPv9NPMjNJoAhfMlJwcz4ttkkn1JHFdVe1GJ17wngeLyv/0IttbAB3rccoSn
WrlEt9yzdY7H/UkPtMKS8aInY6mq2u2qQh3T6HKLBzKKqKz8dHtjQnZ1uZTfg28K
BoBXdxIdhTNgrBeRv9MMKu3RNMOcllEwu9yFwWeS0XA/YYKsWLEBTVB1hxjMDpb0
s8zCMACcAf8zpuWzr8wQtmLyuOEdUswnXcf5sCx/MSJ601MBwsRHDqgxGOGeCWcm
KVIx/V/1ABWPDa4s1NUS7speGEkrNCEb/Z8fHkYz7F1Jo/5RlKET2PGU8bz+3HMd
pZFsw6SSgqKx4SBmO8FpKAlng3YMavqIpFY1oIW+Yfo9yMG6h6MRilquKMP9IS3q
EDDXVP0a6Lcu0hE7yHVtPaRzfAZAcu9QkJyv1Av0qrB4/bRrm7oN/vnNrMPQo54C
pivx/ESFTbu9qmB0d0rTA3cXKWjfwgO97fLUJaL+ELZ94LdQQ2ZDH0nN0vciOBu8
AQR0DiCAJoJ+S6KgdQFC/pyc4youaAdEd1F46hA7p4sMsFk+LMYdV8Zf48xLFYT3
lhxWE+WYkXFBmgBlOHhX4rfirGlxRUP6CqaDgYVYVl8VTvsqdUyJHyYMMZZ6ho0y
OFCp9SmD4ALXVZH/GLBVUrzKnfs36eprBxRfSoDhrYpFssvfAkWDRbHIGo5/0hOK
H+DeqDPthxd9Spga9b7+7zlxU9rGYoSZ8U3KPyMNB7Z45Np2znD92NUREEuTR6PE
W+2U3KvslgeYRSZNDWXtcJXHInPyCG0kQuGvJpYQWm46tS+bTuTvGznQy0+h5JTy
YtFpsRNkseIa+6VZew7f7fWhGRuIDdE2fw4usnN7weu43bweqlbNQIG1OGibZEQC
VrcKUm6MemTPIBMP8xdcIrIqS1xr/GtX3C+Qnha9Ny0+oyp0+wobEq1ZGCTncyfs
5NYizc7hQBNWx2OgcuOPT09qIKLWh/9DfHUB1m0yBOGYJ866nxZrkV/6nL0f+deQ
zTUs3EGb0Q2WwtJfPBtj1F1vOzHkAeaC1tn39y55Lf65qJ6x9si3PtVGqfzmcZr+
TH5QUBllugkMMBaH/2y8IhQLsXc/fyXm6VoSks8h+9Yidfvjn2YHF/MrLbfsvgtW
muezeBngM+oEKcjF+++FmOy4pQPlhdRnuuc7FmP688TE25wKIfY3TCVUdOKpYMhc
WAxMlatjFrxSRgxCa/+fnxnTyubTNCBu1p6CSrLZj3ofO6AtoFZh3YunUwGphuRi
QtyDuQsaZNggk+PH2Ral4m5D0iBozjKk+S42Lj7eg0ZvGDOGSceYeVCIBytJRYWo
V8gD4DjeZFH4bFXSGBUWQHUKCf3aJsJFlyzK1lWFZ1Rm5NTz/8TQYKumfItMONuN
C0fmdv3ORLbzmntDs33OjtYmnxo7TRQCKIDRCdGYzio5zasgrTMGegviSNeBEJoX
EvjouDMyO3bCgPDU1BJlq5SQdGfmg2935ac8dNJK6bCrw21k+tHHOBepnCnS85tN
1eviRhhbMXjjTw0ptk4Wx2EmpmGOJwHKD/+PWHCF9Ef0B6ECc7pyNVlTWMe4yJ+S
qZJ5C1FLOfvSxzVOt+elz6cSFsasSG5qPZBCO63EZ67qul+FMT8LJyyk+55WIszw
oJJCFW2mu/cOSsqnmMFBsBgNoZPPAFeT73U3f8vqXT6Dmzwc318OSiMUXvZoSCxs
ZDTEO4vBtHzyrkn3/kTOeIHpJM1Js5XZ17FbrYY5b8BMikH5DW2bV2fOUKmZtZn8
ZJGJXJaQF9YFuDLqG3qvT7h9W9tVbyDGyOYeJMK5XMWjappJLerfh/+UYwEeWytF
C3WW+xXFxwqrsL8lmNCWztzt/2GykR2SVkQrL2WLK32MrYpenduMM5oEG3wjREsy
BtySNDjD1oLBkaOkS2b9P4GNMPlD10PShhu/tuu0u0g7mNp/nV5SBU8+R+Y/dgDO
95lo6yZwq6JNjUSAj1RDK7aboWSsl6xFPINE0LX4nth3v+u0W2T86gS8EobpgKHu
qcwmEGBHmtaaoNGG0WpTJDMT9ZVKDjR6dISnn+Jazz67F6hxQ7kJNAx1jYeKdvgW
is4QNIDMhHd6BEBoYcI/yvO59qdjQtidRW5k1aAqe53oum4LP4ipR4Rswu8X7BOQ
kp+nMoYT9Zi3BqEwO/08VDH1Uq/4szeBYmG6erokKSLSOSFgRUs9Z9hGi9NEq3Kq
/t2kioFckqaVqUhNQY9TlGjKUkeLS8jMZ7AeNWU7l8zPLzSPIDDvKO5MIF9VGItj
W6KRHc4F0JK7AS8kKUVMRd0zId523yOBG0U7LwMnM7/1mvLG4O7uEAjKZga3x8NJ
HUEIAmmRidbGb+z/oVdbZiw5lBW3IuB/i+o2qrkFjVuU9AEtL9F+utIkIt11fIYi
3mr+Zhaeh7uWnXYCAP/C0REdzO0yg5SkUKJ0DoBRFG5RRQP/ZUzS9QmHOfDixrfr
n/XZXicFc/54p8TKvjxkJbfOKMzk+8QZQbQnhGTSFJCWBNMVR53R791DJ5A6PW0N
smN+X2kY+MWgU4foeDMAWdS0bAPqUvfudew3mEDPrU5V6ibLwi5LDaRtuYR6fMnM
feb9SPizbC6VaTUMAY2/NK3aJdtvR9bBjE1vM2LvlhhwG0qO0II0536oIXyTJK5u
vXl1eLJBnYeqlKBLInXgS1d0NrpK+bWRqWIFCGTh4MSNAV1dsIshMkifg8VUkPo+
lNvzUJbhs9eMo+XxGK4m0u1ajR5Ia1SDxbMIJyILHJZRTSJqhL/QM7OzAsjHo4Hf
9biN9zkGkkh+dvn4K5Xp4XsdqEViPRhHwB5XgNYge95WzckfOiLATFQ+DTFMI/LN
Mfhiht3p5l5gFrAuUpCL/EM4hSDvzsDXUNQ+xWkk4LZotwTewAxmfd7yopPaEXYg
XL9TqyHIekSLAn5OvkoqngZk6S+WQEQW6N710V8k0SNP+pEzIEVpH/80CI5/l7AF
VbQZlnNO947JrJxZJvb/MUobop0RzD+yBUX8cFNiJ6f2hKxPFnBVrYPZtxkoXs2Z
LD9AhlJW62yA4AIBu/5tiEonRzh3EM3o1Fvwcsypfm7HljM4rwwRCQtBa+t1hzt1
B1Eq+56w7iYJYzhHQEKsXOrBJjD5bsPf2/jJeI/xC8kgcLzaJgjIyUpaThw2+ye2
q0VSKrwiVriXwtaMBHQuGr5ZcVGDwEcoJQkvRbw4pli2luDBpBK7vfq5Dti21fy8
iczzgw13nowLC4BDXGqa1lvRn45ssQOCVP1kIrbGLbpl3qQeqUTkz3/VyGDovtl9
osDnOeeNMWlZaasrFX2USsfdX/OzdJRsPGXka0qPAqLBMu637qDRs+lHIEiJLC/y
tnLTUMJZCOCZ43hv+/EJyhA49SWYDxcKKabSBs5Y2/b8iQq0H69ZO+JpC74czlaw
i/7/atSjnWOKA/UZiV8r1gNiSvE31VCNIlNBoHm8VpkDvcMGVFOlz6ez/Y6L1eQQ
LtcqUrssT9i1kzcJU91FhdaSkMA5BfXmyrHhS7p54OKvb6ROa5XqMfhbJ2jlOgxN
oC+lFdgKU3S/eAwVHgsNgoO8XcCtO323WxbCs4wI7NNd10GRoNTzdWdDfdjU/QW2
5W2Xkc/hab1MruK7wWhBC6HyPJLPFWw5gg19U4UgPGvtmXvMvM+6rKOdr9LDDEaG
9palWaRhjgbB9AQn+rSlAvlHkvp/ORRaV+jI0cAcYDU0tQ1hruuTIzP6MkRlSOGN
hjjyHxDK7ttvev7c/aaE2Hs5DqMYEB3Py7ojMJ6X7Hql+LB/UjYKIIRirI5uP0Nb
/WXvcFa+nod4RWLSdub1zK+tF0cRnAwGlA4zHSUo4g5iSe0jFsDz6lwCpysMrWYr
OOvoeLaxNV4F1zo6WjD1rF0WkJrN2RgP5x9O6gro1NddXhmG4gFEUFhrVEkvtwF5
rYNBoWxKqWtBMwDCl5TsGzcTraVtp1cJQVEXaFnV3QatP0aD5uyP+d3QRVsZgixk
iy8PTAPEIFUuQm4IaGAITid91gbCDAkY8tN7tlUyBjBbedk1rx3IX8kwRs6rD1Mr
mt0g1gFSQ1kijaQDgFizo8XVu/8lw0Sol99RvjKR8CKgVdSDMwagstHVzcs3n7ey
r9cZvXvkVe5y1t/IbMFYEcorPEIWjyou47U2Dq8StObSneD6CPsVMZrWtrvvzafa
SbmegCcXgCuvn+0e6SX+Y0bJ9sqYin7Tn5rscd3NxO6aA+jPT63lR5b07qKKXAxT
4+zEYoVO9VLTvpMdBY8o5PVGRVyW8zCUSIG2HcOK/cltS4pPu6NrjRIlSiJnuVRR
CVJ++qFWejDjPhTEIrYQcv+0o7ZJPkDfppr6xTyjHphXtzN4irLajL8oFIn+OaUv
i8gSsOtNjk+In7Lrm2uvY+2Dsrd/TigO+w4xEmDfnrrysNGnV2ZA6nurT/WiUXnw
pStvAZ9l0NBb+BjAmKmStGqYPDihHSd0K7BnawEo0o4WUR5KfmTqoyEDZKmfYtoj
bmXyzWlPu2dW1LOBvXji4+VdySHax8DqrpamduTVYx00alrlW84Sht4/s5EmD/PR
Qu3zpgDnnarUKHy/yz2wdF0FXhHbbsDSPd/Qe7u6vSHUDV7K7tNqw/ryEzcoXiUu
71IsdQiXqnLcey8KUtNG8CfxMPb+VO0+fFmIZjsrsq/n5QPS9mHCet+n846tWFSy
ipXbfVxWYRDtzqOlyYvXbtHA5CDE34/XVwKHjxPYtiMtAUbNmM9SKOS8Ev7tlD9z
tjGkPeBSefWzTq56GEHStcvPqHoC3JH+Ql8q/N/aSDjL6rcXTkGKYj72XyOC33eH
IP3DUCzMovW4u577vaZEmxE5KYmq6u0axY+sOQDrgWSLqLyQ7BfTS/EKWRYa0C1T
qAt0QUsekKxF5IAMO4F4ip7AY+zzrKymHSR5gzaEajKg2U/8yshZ9Z35sW3t/feL
7WOu0TGs1VqZzmxVZ9OXrwtbH6aeJhWlTMirdUNl2ZVfc+niXNr+j0XoLkhE836L
1C6hbvWJjFH0+uVo60ivGPKWDlgwqNHR4j+hx5AF/5ElTfC4AYTf2u0pRim2GJIT
YcqAFjNw2odT86GBpHhV9jtHCAs8MBYRJY291J5GjzVv7hrDVMJyf0eCCN/Hx9nT
hxg2tWKmRERV6OgHC2IFQw9njQdIyS35KbVmkIZcQ9FcNbDV54O0ZsBsAw9p82ka
9POv/AAZsZ0SyxmVftJ+m0CAB59Bv8Vr6f4FaV2eWYtvRZEG2/w/PysOhXkAWGB9
AcrHOukK2IctqXKOlY7ZSH+PlMDwWzt/bmlA3Fj/nBKJomXHl/qCdCeOLg9AXXcS
LUwdunyR5/aitdRDRxXNt9ARCMa4Dco7MbiXZapnN+RrLQvyzYVqK2mx7D8fxha8
BzKgW/oVhTuB+dJo7IQwQdAGxlVDJXmf78F73juZSFGxPhNiSt/GN0WGed9iPy5Y
xrKc4RwDb9sxtZcnR2woIZ1uXcyV56fxnsswrZrEdVxzYsLwvO9hcw6lau0TYgwb
ODgNZLCHut4DEKVmZDrX7Dxihl4heNqgPwOiucCYItK+ok0cCIKN5uJFHx/8i9C3
NspgPp2EIfQQKJHPqXAKtPp31pHjsFb/3PfoHNMxhE2e0BPyP2SkhL94ZAksN1yU
rsiTzjBaZ7Bs1Lk1lWqF970GPCz61+s6/DHiknCyrrcuVuYq3bfhIaKTpXWbmj2c
BLtGz+BSRxX7RnrA9Cp+bES8BLNidi7ZAxKV+1n6G6hVUKro6H0YZKFghXxNLFwy
ShR3ItFizAxdr24ftQ/ZmX3I+6yPZk45JCwueLdbQnsk1LI+MhgPeIlZLd4VdOqF
U6sTp+wYNIf+ZJ23vifcq15j1KOyT9TNyfw0SJNb6VO6SzyavLfqlynuxk4VBDzS
PV7ivopP91rVT2oq8GfOzhhuRmpogJ9jT1uDVjyTgZ0MpDX0cGR0P5QcJ95Yqcl6
TgxvKPKGMVFjLk8KV4ZLML9Z7sG638YnqpLMHI2LCTgIxikjHdz0zY1l0exX5nFi
/NVYwlh8AZpJ11CdVNqF7cahiaKHeCNxu7CN3HdNmgk6r8EAOxi5JkVdTomS6VV8
69xQp1vJJX+sIxc3xddGWEJBk2QC+vRlGBacMrpGjKnImcEP8p0K0758r89GjTSr
6TtgRlX2d/7Zb7mLjc0altVV7EUZv41juWX8h6gFVb6OoW8i+rk3Ru1El/PqqI5o
iZF/i5W2A0f19b8UBbAGYs8R6UFOdUt+1oLNH7iMyWGkCkE/f+/csYpckKI6JBc3
A8oOm086A/ZSawxaceLH8GSscj9iPHiRDnQ72UspmUHbiuB/Wr7v1xjrDKEmRe+a
B0lvjB76Pi2wIfrsK/4XhAXkIi9HDKG9plvz3aYC/MKqKSBABT/CI46YMT5xYkqo
x9+TLcQgygIVO/xTC0UgFzz857fBibUJyk3S3GhEgXzQFBOuoN2/oykGPjbd3HHA
rOKqFa+jg4UzhBx9j90a/Q/Rr0VsOFcICzHxafI1vJofjF0ofSXnuMUOkjWMfTJv
CR79gi+Yr1nIdfuOyWyoN3b7XbJiXWBM7Vt6C873IkKTzcEmhlNhCpoFK1R+tm4h
NBp6GBTmBkNWHBMMd1hQzLYn0/uoTnu9wKIOLjf0PPPv0hj0qTuHsTFzNGzYW9DL
Aoca5+E/XeKhIkLf0C8GMfY0kLkrnZX6v8e1gkam0h8YCA0gxH0g8Lb7r6Rm6bMO
Z7IZ6J3xdqQySQxMK8RCL/+K12EfF2qlyG9+HakliMYvPA9m/uU7q98Lvdm/BPYD
QQP+AdfMOob2IL1plO9/HG0f4fwndFnwFXkW1lyKIfJ6Lf0ZQNXYMKnf9DF+EDPZ
UHrHJPz53NeAYfzhOTyGl6nt0f7JdRDBSmF4MWS0AxSAw7x8UVsYxSXyVv6jlVK2
I4IsiSLZIkFnwcqjas+7kshfJXkedN6QEriprH4YNeg1hMvb9KjE2EVp2DIl8csw
D2fxsATj6lUzblkh8+CWgEEE7x3DlpEafDfUsFXwN+AyRJAxxaCZykGkSgxVl8yN
R9QcytCHUhoiAZkEsL04Z5SLs9wnC/wrxgr7VKrht29f5bMfxla1+5fIX75ckpsb
FtDaxrZcSLopcj8dXYWt0pl6erVFnXDLJ0nIdsxkChoelwWjBH0ibs/sST7ghBIm
hAI1hDaK4bfFrUhZWZ5xGJoEwf4IgWvrzmydBXKQKmknLkpcqQsnxHjIGkHy1Nd4
UJSDKOZouqizqmR01tUwHrw/mO61kG2EeBzTb0mmmDYja5ZRqSoOYpD9D6OYDtTE
T2dYyh1Uy1XC8vDWpwpbMlHOh0cAU2nQpgAxymjmNQSjahhjeDKSIuHfSTJGRlUI
0IrrfDUJHmXQEr2hyWbpJSAeNeNn0yjtACafx6SWG21Ud/y3riKS4Iexd3qNM+pc
bdw9yUl/a7M/QtS2sVIng4gR1s8BK4KjKEIcp1bT/pazCB561HxhUWJgUTX/9we9
hkgNm0LiB/s8RG5TcCZeb7uhV2M9sB3Lqn1LI+cOw4d+F/t1AojK0zlaDKBLTuir
jjmna5yXs3oAoCUONEwD63ZyEYPSmr2tiVDC+GeKrHd4UGjcQRGU0577tSbpX7An
W9g7pvbZXqP+BUh1LZyOJxqYQD9fYNFYAi79xxSfN8bPswUdv3ojuuCVT69KgfjI
GT+DRdQjNKk6wbi3/r1BnHo+aousnl9UQgcNxOUPUhe/oKNBeDJSoXbg69lb4Cgp
BdVl4sNVgAlFZSWN3qtm77YuA12hbMPuwrN9ZpRzq8qTrBsz6Gb0mICeTiA1LPIb
y7CFbqe9ZKzaFdsz2CP3h+65A7H+Jo5fuDUwea1UZiHoXGOrv4IjaucOXvxTt+NJ
wXkmZ8sPckzuWYTw0VpAuPrYj0QQOthnNKhc81u7fZFfFHw/SREHxC0U+Nx3N+KU
GPrSa/0XVLGHcnfFHTVkTQofANv8VSpu/bMEd+qg3Mu9742TRq7LsZL6pc0iQr/u
SWi2SqPvm3FH0okJQYvuEJz+UiLisWUccIolYt4uEKZta05keu9RqvpVMcbx4usl
pDjkcdznPYP3hcxBbmSpHp8ml6oOZ34Z4VEgUuoS2ry76hhqWZoDVb0lfj698FE9
Jvs+6NXExX9z3FMwhiEhwfeCSf/nfNOfJa3mhVrVRA4XE4UmvpNoM7ukS+lv5vts
nVSDWJkQ1hUso5shSBiKoWtPzhHLiQFFxs7Zkg9PdWembtrHI3Q/rTC92IUNSpgu
UuF8EHDrMTLMDdZozuzW028Fwi+U8SIAHTQ7y8Wv2AT56ALz2hstLjUscfThaSaH
3s+Vwd32Qnla8jScgGInNmi3HbcW6gAIH7w5tdVRWW0YEgu5rQ7a6JSaW2A5YPd2
FqsYCrP67k2wRRbpnlyxFQLlipbuJNSBGG1XRhr2x2nwZNlXk3PMkzwSX4YNV/nk
uT/zNbI9433EF2x9EqMAcFzjTh3sgMstyJ03VLZ1vm3IGY9h0brIDBmmA88MJxI7
qftkH8N+gtXDsxGnD/bh/TDaJebgJLQUk9rBI4krEpQ8mYlfE8BRU/OCsepm2Ko3
jS1poJDJEM2b1F6RKUzrwlX/NobIGQ/xxyPkCGZMfCTPurRCHFLbIgD2ahj04Ymx
GN2iFYLNBIw0gueHHam9WI3/PdvI5kBDcVoNBb1cEwpunilF0VPPY2cAVNokI8NT
N7b5MJtED10tFWVF+tdVhbB39Rc2+lt/a38RY7GGfqHi4jxAt9pyI2L8qeGl2cow
wGj511Ecz3aT+aZCc1BJJknUiZQyNGZKqHmch8Hxf7rtepvGF+cdqsI+KRRC09Mv
vaUQ30ara+KC50CJCRKjk3OpKWlncEPlnfYRt9J6bskdIlsJwqW2j9FPd0CbZL23
yV/N/GRsFsIdVBWC2f1CjzOJDesXKinS2afrvJ3rrfyAxmEeQYomMuXoJ4Wc40Ab
d+Xuhk0gi5RO4bOmtNdo71TqR59IabOdvYTJRifVzXNuGZ17GVnb9N9H0rA/bwFQ
T0kbecOzjcIX4FPVh6XfQt+zRm2N6SnuGLr2sHLE+YEFOZjFJ9K+PIYm3YL/DL/Z
D33+cKPQEde50n+8/6zsfDfCTcC5BooptKvEtWhnyx6VJz4zwowBwWYX6gyb6fVi
uR78n+HTkC9W4moNGzg/fcsZ7Xyxm3KuQqoRuEBUJC0VectHWJX8XRYCQTAMLzWS
U6Pjp8BYBWChXtkEJ/tTP6LJG5+nSW5yA+eFrW+tH9njWyYHXFHoaoL9vf8Q5kpL
sPrkjffPh0Y7CUlbM67YizAHCBHPjV/H5+fnb01NI3sgVFIQhJCBLRE8SOu/4yRw
47ii95T9TZQ0P0OXpUg+lBGcQojJVIKGbuSnyl3GkT7ObhbutXyNcv2D4/4CVefx
Ovmiaq070oZuu+PLdmF8JitBTffQYlunl2IhSDicc+hRM9dTqF4NVaxWLSRj31bu
XmYjnGQ7hifl4hbnOQQPgRkgEjNfLu2SL+qeUiL8VkTQzw2M19j5nYBYdWfAb5uF
SYPwLmjYMVY5WOKL+CZdJX9+MrRTIZa5HZGNS0dKNJVFUFxhRh9V0Uc4RdHSV1fA
xWFaaAUkSNdP6mMWCvOzrQrXK6y76rKEGnACb/Oh1n9fD2a2IKorb7xjFDOfbFpW
9ogGoicKMRnfAr5Rov9tUdxuFaz8wIBFAt434S+eJHg5TSW4CUh92+ZYlELbWLBd
ufoBViMapN6VJGOXBT6f3RohJiNfUZODVk91rnRnCjSD6f9gu867y2Q1K8iHIhvx
1EUjw/nwPQsH1aenF7ZBKI8ElFklLuqDN+xDEn4RkC7KKY8dOJRefO+sUN3kRHjo
AhXzzHLYAOsir5juVdM+QHXvfBS8GYvuwi7XibGjzwOKv13EkTPxmpuDQ4EKlJpR
qFGNEpl7G+YqG1nNxAIczWE2oQaLIMG/n9Zw/0e7iaNIpRUIH9nFmGc4gS2Z6O4c
tF/+SAjHniVwiIf1lu5Mt5sff49l+yTuNatUw0yRL56Y1PcrbWkvobrx6l5nBmx3
LHTNNsywToplV5XHMe1vsKTUbtgrntKQzLxezEI4CujsQzADduMkHG+gvv6kd7yo
WbtqeF+S42pGy3aqa4krbPlxBiCMBpocHSRd1iOFGnvD0SooDytYdadHeGbyApsl
S7TaIigv4iDjP4Ufs9gwqcr62ZwAA2SzRHry81hbreMdZUQkHo2evbx2vSMjd6EQ
nvti1MkAMvlmMXzEAp7SHuW99Ljx3c74aWXhDwEWIiwxp4yFlPxNb26FKXZN7dOa
0fiODdLwtSl0m8M99Hw95PEe6e77JmejrTfPhnGR4J5JLqcddWg2wu6bwAVubnWv
7Q2lcMrm3Ay7+mAEgcqeXsXSymtbN+BuE4+t+oaJnpNzdKf4mgeINMhdQKWn9EMu
1YgekAENEBYd/ExEVyoJ3zRjcOgKp+ypGeuLv+fHIF+iXV9wucnb4eONSYWcnmd9
444YWK3VHoijgV80Fk1LSf0UTafEtJPwkjjs4CSyiuCaVjo+41QGqckpZyun8HHt
nX1SLulYlv6tGVQO7pekwgY8M9nWw2V/xS5/9Put9eSB1htcoNJLeyFMSAq70x2o
5qQWrt/VJNhXN+WcFi5Zbpv4efY6M04CZRV9WyxKql245dnr5ZSTXj3+v6VIjUOc
E/H9HQ/soianTrEHuL0kbqu/HaOta3w9yYytJ559QHQdCabI2MdIIzIBIpZaqK6/
Nq6kgbeIC4siD31TKPI8ALHbK9psJBGMfu6muillEGvMdv4398xhhzu8tm86YinY
iLUmq4Ti6y7KjAH+W7pR233cSUksEex+a6VHd8qmaxxe4Xz0BBeMhgZkVRGMJ4Rp
K4zrIqvHwhBlovWVqPItNsG2Mn+LIjUv71irtCq3GmmzvRFi3MkxnT9o9e2pcc7R
fqBHQb1ptzMk0qGc7nKNagenKbV2hWFBoFM1cZek2lzOuT+bSkpTDais+weexyT/
/ODgMbxqczpK6siPQRW/sYTty7WjF9IZ2nAEkD0a/BbHawMBR4l+U5KvVB8XHKGf
P7dL3ya8Uqqf/EhC1zxtjzJPDnrMD7NTEUQ1o61BdTNPyE+OqPw2HiARQubuDU5s
L7PNIOGQpgrPwNXsTZowakTEEKSEfVGiizaciTfaTTzvorvUXQ+gfcqgMp/s2kNG
GITxELoMML6RQ4Ed2U0S313tdgXEXarplttnCp2ZlRoMWr8ABIQCtG7+2AuURhQK
f6MG65efebvh5rAUjqfRVhFeR/3zrc83Vr3WYU9Fvm8b1N5JgaEy9+Rwo59RXxpb
bIiBNWuCZpvDjHeaczPsc9UqGKgG+IGsN+RbuPtdBdpAHXwTf7CX/HwXvJYd5wRr
+ZagbgDIpvLQ7eRinjBOmd3nc1N18FtP6qVoF9wDIF5ew1qwrE24shAAnDwKdT/Q
xuhvXHucjP5fQogAmi8Qm20G/VykGSZPBxcio/aH1lLE2eVAuElT+weJLrGWpMuF
pYeCqAZNpXoKjCFzXMlO8sK1CnfmFka4ey41FCNCHo/TSL9JGwLc5Jk9xw3JI8il
DJrnkBfF6odsqFSt+PcM9RpdJGfObvY1MCP/gAKaKruNT2LCMDdKPQ2C6vGF4wBP
XwnJj+G2H8tEJer64g+0g4U3OMHsM1BDo78vn/F10Lh8uo1KkcbSEwOISQkTDQ9A
UIP9EJlmwF6xUM7IHNDqbX9XVxhECTiVvUPLXLEvsV87XRJ9RB/RFwthqnEEvJ0f
QR8LovdgY9mMU9DEcADSjEgxloYbxp4u5dbUhnQRVPi9/FHXwB7jWiy1CqALw4sL
Wphl4IfNlzgA6+Nip21AHCttZ9Y7+MUufoFxIF1Z4D3XYS/siGQoawSH/CfQKNTv
tbsAy5ZJ0GrUxPr55xgXc/DeEOGh/hvgYrwEPIiefE1CaED57IFbftWAcwHlO1t0
CPun4atifa0R1r1L3np34FQzpmxhnpqaVzqwHKSAzGQZcz2B7idJrJagK87rzvZJ
820a1x6CLCeqsUfUSxGQL4X7Pzh0lfVrQa1ZrXivO4y5UrNUMod3OTF8aDzCDcgZ
5+5AKNe/Tw0NmP9IVpWTNb20QV8/Y64vT/JYButWMUMOFYGnzs2UBflQE2JIk2x8
q3A1tEz5bMfF+t409j+Hv2TuCi9VGrDq+ymQPhqa6R4Xn5gOAV3qUYBG53ohtnWf
bmGr9vV2P3s3ypeW1h+PI6ddxG6CRZdSgEILDj9c+EyvXxIjWoBJVs4QRHhudz5A
7ouStN8R+vDoeKWOV72fIgMIy0heKrmdn73k32RDQ4Nhr852mjtHbeeXvI82MYo0
A5p7dVV8wsF0ye5wmC5+cXlQ0LpyLjwApVHKFLBO9273lkIaqdR6TBablUCUnuY7
+Xo2J/dHY9NiXmOHEhkxiXgt0+GBIRIYtzMTtq2tKcCvf+Y+ImGtU8xAEW5Y/RXp
U1M8IWFbzCc1MDRf+HnQ4UjuL0Kk36ODa7qsU6V+N9sBJg5BD6svtfLqU1QRstCH
kQmDHs3UMKx+PCV78KfcuzCiLUH12l6dWsMLykIjO1C75Mk+WzrdQ+F0JVEQX8Ik
34+wnZcZ/qg9Lh8H9ydd1RUoLTYbWQPPyv+d6ZDxUB4vARFwgKAoGDFwq2xt1APn
WMTfDs+R3/zLU6ikv8315jW1Ip0pCL+y0LD1W9bZsELEjRLjBzmP1aQGZ7xwxjsc
Tg7bNgMUKVTCLTtIAkpUZRGSkbn1tuk1o2yYDblYoiQEhLIsev7F3nVIAgheJbRj
FCvYWO8738ULLypHlfxPfqb9EAANKVsJpwnZrAxYKxuTwChEQsxt4YbnSKA787O9
xm1fuGYpMvqj1IR5mq6a9jZgMvXKFRbPQ0ag6URcI2IdjsFWVDf2EE5fraDk5ktt
oNylsXf14Gt9JTFX6JK5I7fD+pQ22Gy1c1YIZjGWXaszJMuoSQhKuEnNQy9rKaSB
Rr1WWfRhVShj+RfUFUsA0oom8FrvSUkVGVl9T47u6GdOk67BIKdNGaC7D3L1HQCh
Dz9Fq/T4L+n19s4hQvgy0q6qovhYnzKxZWZ6rwbr9gW/rG8gq3U/x90fBy7uz50W
pC75B/IOeu96bDPQaASCp6/aSlz15wcFt8/q+JFwtiBfiuEu14mEtW+1YtsFsPa0
60W3KvWn9HpmlGMehUGjSWISFLxNrcuscCF5y31YiViTpYLTOtsYd5KCaBnvHN/7
7hnzA+/e/4i0bXN4tQKNDpFHZWjNAiIgZ5YU0wan5ZeZdkuHxerliA7VRUT90S2e
av1NRKK5yhCnS9oZHqpdCvDD4554KPq+TO4eDYqpv8D0rnAfmYvvL9mckGeWYo0M
4lxH9c3VDNwFPQZ4/OeD9D26M3nGq08yBzondwF/YdSotIaau7n5GLTexUwT1yJD
feydmzHzC4KosZ1Mi3nydjgYNIOZdwXvowYQQI2liPhTds2fEnjJD6Rsx1uS9iiD
E3b2QcxP1Pm4nz/qLU7+pr6qCRtzVwA86u13EfGue+DPc+/S4u3zBy+MngFxQf7s
ampe1EKteQXtIfHJ6yRA8JSsHAJ8naoLiShSfqJBd2VJVh+Qj/pRCCUaGQ0TsaAq
kATYymJo81A2jvIWdyiT0ov4O72D88reIGiybwv3Mnw1B409k+0J+d3ssTDtysid
nr4nt/HbkNBiD8XEhpmDYg3aQ0WIXIoEUovEzgkFTlTHXF7xpCQo5HdXs3Lxzvgs
S0j+m397ZhIUfq7utkh+iM63/ennyDvop1TaRgbwMzbk0g7/J10QTj33X9aq5LOI
bLGv0rW79d2ChrNE058Ooicb2e4S76mJ9rrI474SdL6Ql7RAWZ8Y2xzx5y+Dxmf2
K+MdgmzrHuK0UE3g+wwpNa+sHkg2zzET/+Dojlp8t3xdeDmGx5VVrukGj42iflO2
ltzRKIiLVH3vv34VAvbQa8ZoRtYLm27lqW7jJiph36xsdrkTDoLOY6BpS+MibaF2
hNAYYAp5XRCJG78HfkAc4/afnI7JIm+RQs+pLGad3ac9B9ireyB/Nyne/zj1cIho
q3ai0tkduwx1oBTyH43wVpSEVZ+pcAcuJFaWBOYaCa2dbHAkr06pyvYnpZzfKDJM
hagAW8nlleESHMBiKfFu9sjgxc6vXc8wSBZ9XRORY9cWdPBxETcpFDHhVjSFrHKM
p1N7xsqx6RnYC+NPv24k5FIHpx2e4kvdd1lE+M7EsyiqmFtMhgzUzF2fU4bW8UxV
QPHVyJAfBL2vGCPKQIx+aH2MpphX9scEnu83IqXOOGyXlB6H7zSY1LMX9GrN/Dr/
j6MzClCioTAnfnFUQ21qZLH5mtNG/1zPeG/UuwSLffipyoGLeeH7J19Lz+FyMKy9
2BmSAnFz5G6ULX0jFk+u0FjJVAxQ42jj86MImw2TJws6IIAKGTrig0vHRpkjx18m
nTLRVt72zShjtgIlWHu8CjuPMvHHZViByLixxIuZEu8HruEnS/PUb8jhUnsAbymW
+0jHteFRHYpd5G3uogNxCkxQl5DGzEQFUaDACm4Yo6j06R6D31tBgKKlJfjPxuAM
DunDWm8Zyajj4XI0T8kS4mAGobk7guwnPu2LcWnx8b9qvem2qHyBgRt6yUs5Snc5
6YT0d14Tyny4YYHxJRmNqIkO1sDuc8WZ1Mv4640RPa3oAorAT8uSiu7LxT4U8KXC
KFVhMIKy0oHJOUF96YeM0XzMuu+pXvJhMnTyLXmjIPVigNdKxEQpKSeeq0VKzrh8
m9JIWdTvaR+CMj712Vwv58FjufEBZvzI6NwMtLAcmK9Ix8pWA4OILAVYGOa75L2Q
25MSE6DTFxqxHzcgsNR3o36bf4LcmjXBqhnK16qMcxlG30bT2sEmM1sSQD1vjDt2
pJGqcrO3eDEcr6CFNO8np2w3ybrcfbFb1cHnD5SMWc4IGIRk4PiV1xWMtEuPhMVv
U/q5M7aTzt2feCICjYLZ9yWjfcTXPwahfOXmSkadU7bmM5MLy0djVeBMeUc6w9DH
hAvjxCwZrwA+hCS8I30mvVD6LLFBF++WGmySqSAWx6o04Z3uJBbuccwPFFNvWdIn
bkD33ZYQv5G67zhR7YtuT3lF24GHxAVxKAoQnDBT931xGVSBCMfjpH0W4vbjcXSv
P33xq/aJW0zSpg5B6xz9uV7JK+cFfsmjlhT7gchcH4N+J4lk5yWSW+kHZDShMQc0
SbAUKSriQ3cK9yjQ6265q8NbgCRQKBMRi9RSb4R97DWc7V8dEKE0Bm8/mzGhYWxe
Fc/wQ2bVOzFik8mecblzTR3kbXeWDGpeAR8dxUAVom9PFM5LoTIjzhpLYWY9A9nr
6HIl4zXvB/HE68SMgZQKzllWXsG0yjyQNPoXNzzBQ5QPYtlNV7dXttCAYgcmUUn1
BejOoB9Fv3wCKuqyo/MlzIHQVSPa8UqGgumD4qv6UtA9fBDZIrB0bEwSuKrHpLks
4FzNSCaI2LB+SS6jn+E5dNCJkrAr4Rd8R7okHO70PBGLEhpQtXfm3mb+M82LcIDw
wqHYQE1V+5zLipgJLugNKriapegiozHxo5EZ2M//Y+O9/hVRnHoviHij96f1gGnN
jXC4ABlLllp5AgbkdsY1JSe7wlIagM6rSKpq96yDOETV1cQry7bPkkRFxUJvwVun
DkuGWPjfr0ZOrsahgBlGKP2m7r3rGL1IGnW7GLxWL6pqajRpfSB3Hf09gwwVm+X7
hK0PIpRJUAW/KmnQi7/uRg7NtKVGwwG+EyC4pGeKf90a/G3N3MPfUJEjLUBNd+Hf
W+TXTwU+ft+kXnm8XInT2uYJOZqYOkToj+awt+wOw4kxloROUr4aldINUlfEHxx5
qcRYByXmB4B4tn4e8SCLlrIwfHuwXqQvclVf+IbD+MG9bw7jgBFYyVaMuRHS7hlW
xE/fEccTyTq3aznWUs/6qebJBju1Xq1hO1h8TwX44ZZhxDmiACVSFnXr1aevIDK5
8e5fc9AigCMCNjzh9vOwwpO1fh3m48TYC8tJvreCcW989HN2jqVsYZvWtXvmswFW
6Aw0HsJkzJLaPQ5nKSwRjc35ZC6jQJWPByGT2NtDRhcmLekXH1xPkUgkkX9NIu2K
h2nWXK2ePV5nFyxEV9KRIplpiyNMgGpqTt5K+P2XGKp56Dbtf/M0hztP8hClC0+V
Sp/eqEgZDosFL0G5KO8Vxal7CfC6oZIexbtb6XDRsLtZ9ob8a+uAuLPDT+QWDTsj
B2gDYNc+UMBOnK+7Ikt53YeOajSbhlSGdf+pAhEqJ41/DEM9z3UQ+ANgBiYlxqo7
qOyOkKn+OquNhG22McIQR+Awzs1u3B7i2VhH3peMi5fJzTmSFf1vmzZfS8b4k7nY
hmA8tNPZkHODxb1QZWxdAdPmjuuzEq6IW7J/Phz6Omjim1fustpFqV5v/CZJTtOi
1fwbCcqYjRXM7XKdXUauD/Cj2JcEGfNSd2WfYfesGAAa8j9TR1tnjFnsmIloTh+N
QKoveqX4stlp20oH4HN6iyWzTfXejogsvRHvMm0p2SfUMlHEYg4l5Jv2ZDoeRNgn
03ignPerPE6fsmepWh22sC2U9CfccJIdn+NlIQnYm5tNA+66sMpDy4dgxWsT9iPr
AMXQ5FAkdzib80bk3zIiS4kMHpMP0pD3sKEr9XIwpoY37itnoOflyWMR46T+zItJ
6+fmQOZ6hL0an29VP7kPHsVbQ97gyagz1aduKPsOauBv3lOvkZ9xEvLjbGUATYQD
7eTM07h4CDg/2kBPGc4y/633MeXOvSFexImW+5hwjZoMwoPRQSqrWAiokHNhR10E
Q02IPic6ACrEnQxa/PBadDJ/tJZYWqSC9DGgxjuerzHDvO2qr2DG7AAvXihWKyc+
F+/Z1T/hWQBtE+d5Fsmc7RBAoJmQLeI+Vbn/RR3n+Y2JbUnBpgtFv0uQYq7t/OIv
/1reoA1MMLbZVj+Tyqg4MnsS0SAIFjRNXQqWmgB0W0d3FcyiPQjo0dzTe3cqcgOV
D5jxU7hw3Nu+A03Leg2FFDAYvF/J7PYPXt2vuQaVWFzPMJGjQN2VwSudUbBkNoCT
8wlmhcrGD0by+FRn3iPuPz5X7KNeqbiRuXu8DvwKlDE3AKQDorPA7Ml4hHX9ogNP
XoLdr9H5Z2zg/p95GSo9LtaMJ/LNnVCJa+ANuLgFe0C4g9A71tWfa9K5ZbedFACS
DTdWUI/vc1DLKvqoLAb9wCrAI+oA8jKXMfIjga5w1hmfa+oq9ltSadLWzHpiX4S0
oUvyghz3RkjhPp3KlewL1B8+Ybz0BNNtDy/QFF5gzGo7zLvlRLnwXN1OwqIl92u2
VOfS6r4CB6JlYA7yRSzpgFza4IEIkpGd7a34eS+lusl+rGY2GsHO0Wm/M8cXdQeq
Z3u+bNoBnGF/fzRQ+mirlUXoSowLATbH3MB7HDisxR23yRQqKQ5LXWhoMGiqCnLt
xu9LXSj7Bj/hrkxjTdGm8rkEsUIEkCw8vHVLWc1+2SZV3jTiOGMTRNm/pALfvhMO
XVnP8aEUkySacR5r9Q/v3tqpfcxJ+GNMdZpWkKZPKQAoQRjZcFMCB+Q2L0mgwtUI
hpn2Mb1gKVbVHJXV3T7KF9qphMepo9baXP1oUKVbzm+hpMv/EBzKNXlIqdp8vB8k
XzxIugtCQ20HG6nGb07afd0sdZotUV/3TnFBaPVamnjhoQeEfLat/RpiwcYQoN1u
z13n3IskEyo/KSww0+uI1MqxnhDQO/znJ24ocbtmauazW8ZDLCo7qmbUzUAZK4c9
J+83lkvuJiVYHfhqGeeSJdXL9dhnrNP6NBjXCeaD6TyorNJ/KMtqJhk+OORA2kYA
K7eHxy5ctI39GlQfyQIPQ3EgE2e8qOnMcL5187c02sTM2gEUERDmB3Y8Zl0r5boe
YefCwqFralE1czlB3USh9GMitLcKL6qCclIa4maAArz+887fX6L6N0iegEACqZLb
GvV0AlxDtCDJB7v7Nbaxx7JQLhlp+zKQ+5+pzrQL9KTp3Q51xo6h3bAV2NAzsQHu
xMrOYchK40QAaSZxsrCj18kaYsJUmAHrRTOeemyPUGWF2tVmnFud7JCuzW9GaaP6
dTR+ETFe6inmUySiqNU05tbzYdSVtYneKyAo0IqKAo+JHwoRAW8ec4BsscxTQorX
UQgotCkvdWylI5p6i4d0fRVQkdTLGqG2WHca7pNx2OgvOFOO118kAVd/i178KC8+
UEw8NjH/8+rEalmF1sjwBVbQ/DtoAklnKREfpMJZ/5tlqzNr9OFiiL5RDojkNwAc
k0rX1rXiQf+SRMhD1XoHzR+FiwHLt/35sHLKRfKlbgyCHj7u3GzMxEk9vs/IIW6L
B/osjvq3VxT9pfMINlYc9ULbQyXFZeBIhtHnOQvIwlvqth8eiTbbIHyWY17k13B/
eejVo3fPCN45NedUO6GbRuTVMVHswQWApSPoSGM24ShRwpMfNdtudYKMxYUXaiEa
5jFfWNdQ8+HdsZh+KBKapEKrzbqCnw9kJM8mdwepjcPDU6fGaD8KKVS6GEPutLny
DHWf62M5ekrLhXtvIe80axvKjC+WOBl4R9Nki0r3yHozHJYmNhHBJx/CtwLj8NUI
G7sirRY/UJrm5m2RdmxzxJUc6Cmwj6APGX9i5BwM7Ygr/zaW3a6pw+UTbUxXr7c5
D9Iaz40p7eumuQAPuCkDp8gvrcGLvaQ6j+m8ChyKYH1W3uOi6aN+LwvuIk++o32b
JLwl9CoZT5VPo9t+HwyfjYeqV3SU8y/rBYkYzU3WTwlzyxXle+r0EQ/X6czMYNgz
dI+Dl8NO3Rtyncr78HZ4CtpIElVUO55TEualyheAbBZTLZDoun5c9A32VdHLpOSa
IUocDGITYRAQTjlZvMNnt4X9QeO2jxUpMbvDKftYxACvXnqtLNqN14XrcaWsdoEy
q3La6GPbHKBZhqetJNFgyF1imn3lMnKb9CldIkkmvlOZhigMnAVgWWhUYi6wAHLQ
TaMH95KPCsQXtgLBhpTY5wi2oW2JqwqT1X37gTerT8KL9xZ2qhDcqN6tcu9Ej8b6
aqeZsJ4fkxte48DV4+AJsAIZHzI+tXUMvP+8VQnIJRLneSF479wepefV3IZs86Yo
dqLfFiNg5c4wsgMScOMavM6LJhYqlzIpZ6WQkKJJx/mFMsyd4HnOrv8mgn16/cgl
Gg2f4YBnkYf2arUr7kS/QbSnf6uYMnHBg4L6tXg00yDXU6asnPABj2nr85QDmDAA
tYNF6yhHJXs6HRStZMtm7ndG++nu7TnSYFlFI0sDTYm/WCccwxDJrmLZBsSSwco6
ONHXtmTshnchIxWXu6kWBCNCwqG5V0tLqRHM86IiePsX4kWYao9CIAw80eNr5Q4d
r9AglOq+2uaCItryKGM7wBuy5SoqXXhKY58NPLYYpr8nUFbXD3C5+cuIiItpWlUk
axbTJ9dYrae+HwZ1XkVvLHZr9Fnw2msad35lgEjO8bJHsIBob1VqYDwcmpMByq9J
KVF2lbJV2rO5eexDM8kP/VcSo+8CcbB54bmJrC7AsXtHKQxH217kxGSVza1Bw5LA
bPDCQw5EdTJoTzNvGle1LuH9HdbnXXK8D1WdF3K+a8fAhXn1gEv+SVeWX4b7H+f+
fscpQ752lspnOzfJUl8Q/rvAAxi4pOLfTYQhNsDLUoZujXjleSAgdo0soV2sXK7k
O4L34nLnNMXu4Q8MiyF/7pUAYe9mdpK6ZHhMs8uGc8P0SfI6JCtAawuWONYaACid
5AKPZ2t/EeTwTUEDFmPduBiwA+669+qF+hOzdC1By1YhU/zoQ7KOJBsuwLD6qoGE
WnhRujkyq96sjdip79lpp9YZ59T5fj/Gp8WM4iKwRCwZzqSV+PAYxc+fUF6lSGVh
TMvvRnEVt8PfWLB1ZzfNAgYPVKNhCfQ8GxPRmeBN2NDbmcyNAZrTNu44QClLSkL3
R5vLwgHiROlrGr6EEcptsafWel0er5zOofFybGNhh3i6dgU6/trcrtmTRDCCDJT4
ouhOiTYfD5UTpYALktche2KFgOIidOd3qlJ87+lkkpZqGPWtx1RXa7n6vGSBlYh1
9CjQPJgxHYNM19f8DMVV/5hXK9oXZiD1iZT8Z2TyVWa3FrXYvWJnh1BXhVWFcelN
ksz7OcIyWFKGqLWNDfUrAjLErVigEs4VYBvtcDX6LcHuLNSvSpubjbd1xyCzS+fN
B/GbwAskL2FoYRZQkcKoxA6PqCCmgTPH1Cles7DdlTl3U+B1YJYGi6EqQFR+IFRE
czchwOT9edTz+nBW0rgNtpfxnMXf7z12HBr0A3QGiwY7etkahiJgn1+yWTolyYll
nhtP2u9VIkNHb3Jztv+NvkOF8iKdh/UbnmCkY5kG3/8I8vVyxDxnfXFp5eDz7RU3
lsu7GcU+dbNmujY/9PsMnOnfAfUODWoqDK+G9k436aVc3W/6ZOaiY8OEpZ6fOPeP
gZJR2+JCdMOdtmVHdOhr1hL+pLiESnybDA6QQpeuTjUCWVvJ+mv4Uc+pKMzMQdHK
nsDX6q6SihS13DC+Em3F/Am1qLi0PrfxvX1YgVpefZJ9YEY9ytQmHQu7a78e5dhG
P7wEyAAkBaaGin7olmHIMG/Ee1XV4sNPwofCfJnIvwvwVldWRU8mSa7tJ9Q9NLAJ
R3DX5cP2ywKAwXWmEolMMuQI2puSrl1blNd3BGCWdzCGJ+FYwMicv3QddKwGl/Mp
8cNM2jC7SikWbwLDn6qFvKDtGRVyi3Ron0SPehdlBs39xdUHKz6AONm/Bwdmw1qp
EXmCSlAYJxVPXxJWSfAKXu++laX4TYXXcDnR+MmBQ7Llwk2wnLMb1+4nDT5/F7hf
xX3/xQe08DQeBA1AMNJRxAF8VE6W7vQGmEsCfgIBDBbbn5/jWn+0ZkS2iCCRis/b
fA+pEb11BCDXWA4QDmiOerDyiv59U9PadC9NE0IdIRCSUWllP/hvwQTNrbtUAsZ2
Gb3Dcu8Wriy20sjC/UCzZ0ih2TbX9JMW1n2zVRqo7i/XYkvXDx3vjXVjQC6fSTYj
ewbsuJeNViv/cG4tG3RjlMLHV4UBBC8EtuzfZzrzl6vWp74xTDqsaE/qT7eB/o/b
pZ+AHMJ+oSHApg+Drk9a7dv50fKyb+Tlj23XL3Dplycil0oU9QgNVze3XVTINTp3
55IA78u2whem6B40jKK85INtHhBH9gXUNQ8f42Odeg1e6mTGskHDd/d7BmfFY3O1
iH9U9BVRm2GnEWLpfACDlej3lsmwsuNvlb+WrdyfRCNxxrWK+HVBOV83kvwypnaN
dCTzvXySF9Amd6kK4mpNlMcckJBh0OBgFONoza7UKhstDpVmYesbdDcb+XY/grMe
Bs0Tspehq0Uf4k0IpsL8CEvQCsIs7UvEr0vv95tIN/CaBFMIbLM0vsc+d+b+h4Ou
Uy7xx6JjTZij+qRVVX1TaPBqNYaD3cIULcSbf/cmOBEhVTegdbkfjdMdStkdDE0A
mnyPHx2oXEIH5YlcMFTXd877RiUiOIeET2MP5dh0v8IxdA7XLcfPX9CwCj8HzHZc
fcm9GtQMLAgY7sSoVmOjQ8xIUbjj+hJmNqnTDbRSrAdOj6/1dRp6UiHu3KKrtLJV
AVNsgdffbsqKSznZJjiE7kQKuEE2IaA0AxYpljQvM5/EjWJjMrCAEYjjB6wRLrJc
Eh+8Ka9BjhymyEhHcLZ1RnkaMfgpjUF8oJy3pTS4F2ILcgyopm1tTKszLyjVbTvy
IpEjDLySAbtzA0/SzthAYq9G7L0R09PKTzA+GUh46BzyzsVXO2x+ym5G1WcsfiWD
GoBdkiFMHtETHVXDaYoO02Eq+XdCxidUDQQjAEUx/Jj94P9Kw+w5NidSbpI2dy8X
1+zYM7vgd6uBY7kRTk810gJwLxPJ8HSVa9+Z8a+x1l7nmM/ql/z/psy8mP6zQEhX
QzSkiXwVBnTLaa8aH6/agpjZqOLGITPa45gMclM+1R92ILSLAhmxh7kiYlHteWAF
+goLwxQms139P+EvcozQRWcFGch7eKfIVeSRWNVWyW9wGNlx9IDwruryfJtoGols
vQFe0/RZHL3hWy2LET2vRAZVBRIYDOaibtAxRX8L17nz3Rz772AWyayZ/sfoQ2U1
zn1R/09KFTne9rpZKCAh6tPaO8oXUaMxe55ukH/tGhryQPHpgXN3x983QdEPGnTu
yW8lkGeQjawIyIMo2zR7UnSUiwsmib/Jzqx2t0i503CLbn8pNQO9MCS87boV5xtu
6tZV0+cEdJMgZ3GKgRS56rC9xpOKkQAUH+Rez856INpdMTKjerXz0NUXGV8MLuwX
Xwr4DPK1A9/bchTog2g8tc6y2cemV61Wl1tqHtcO+qQg3fkwOgM01ljuxzrYPcBl
ti0c1iRqsfode7IZFQqRYzlcigqgGFOPZJNRmw1UMrwdktyZWtiUYoMDjN7HAVqu
ahXzCM9ZcDDNE33w9FCbYJAbKDaLuuAEg/7WkHqMEKbMaVSV1HxrytCjByzfYDke
+JZg9knW4oMJjFhj2KN4vlZSJspN4CN2U6mdD5+bfzFIHDQJQ+ijuWUziNZcHCQD
NajPwHLsfeWRxJtX7tqu0mxKWwwfwU+pXVAp9S74Prt2v84NprcNfiJ7Y9Zj2aPI
MLYUU0j0g2fVMlYoQqzoFP5UFRowW3TpU3BZm3PHXUgPZrPxFPa5zLBeHmJGSKcU
PW+y7CrXShwLnXi0Y6BM7lw9Pj6nmXkMrgRC3vfxzvQ0gmfJCe9CpX30UUoRCcxe
mFQUKQ3epgnFw7qnJxP6p26kULpKvHj5wGRpns95rxIOenYKHwEZShkzel9MSqGi
oGzMQMxB9MoOO9hGhbkgEsI944Cjga1BfCHHMl9cZv1jHzaNCf+rFXDpsYNAaZQj
h41C3Jv+jiiImn0ejjTpGESyZPrxqdL+FCi/pdBCGE14qkOITEzxisTrQFdHkMAB
ApDj779iNmWuiilpLl6loYs96KKz2mBr/j0lx/Ob6dkMnxBNJPL59X/A+rkpUpf6
ITFNAi4jItu6iTnV2G9vSG7JSwDOzTPHtJo77Y1g/bi7n70LFDqn77EumYFFUZRz
Dx419LtmWdELUJT0gs5evHlhucewbZjfs59QdDAL8iYXTK4y9Z13in878CtEpaQT
XAcheoDbP3sPVAj93iXizB7kklqkM2HaiMJ8/O5HfAEbDfXH1td77kCiO3w/8DKv
VcIQDmYrIdeXiPuge9ToVC7qYIrwvkxoK58aK+7t6I0DbguMOvPbvVgpXZErNlf/
x8ETNlTKAoJPDHtSLsiDdic9nNO0cWyl+ETPBnaaZlOnDA66YAHvtFr/aPQCM6dd
pOJSAsURw8nOdhTp8k+eP7EJAbQNAPgGR55j4MpRvIqdNDqZ6VYS5KjponNRMDON
AXZFbny+npL+aPtL/H7KrQYQBKzPWbRzZhlwOnCz81kL72azQ7kxAGQQtq9CxONu
zd2DNsPXrT8th3wBGlFTLca3NYV2lBlfcVHSEfWdqtSzOemyYXT19wEnpp40oq5j
GXwJHEQzUb1STFeAVqJ1pEuzmC12JmC8ccqH6hcHh0nJ2Ge45zlbXmu73LEI5BTO
6ZKAFeuHqZDBgPpk/CB/aoVZ8FiGT9WOOnp0TKtJ3CctbBtHgXpXn2WGLnAjpCNL
eI8kp7M0js734RjdnQWGXP19b6p1HfjWEeyuLK/M6m63AR4oukWBvfWeZiO9+XhD
az4tcF3YgrlTgr/qvXojUlFtZ9KsuWPu7LFQFvcmrdUSoakN55Zx3zPKwGTZfXmB
bAkJs96Jn1V+ZPDMd0JjYe7HUzrmNQZL1pX6IyoB642VmCqlENsCNwtlduqwdQS5
WzpRj2oazQ5eVGcOC+YpvERqavCF0wNZgqNVOQKB+eHagDHHRg/oos/P0b12x3Qw
RSA6zEtHz5/X/HNJ8Coa8uT1PoWwTn7mFFrx0Dyj58T82iJ1UgjkZerFQeEwJkhU
DvG2X+xv2dk+cFrG9s0T0nM+EE0m57Agd32LNmS5PSLSaB1WwUTvIDS1b/yEfMLp
7o/dfU9EVRjaoeH+MMQ5DR6jBMnDzrYDQI1T+0UKWnNnunU3Ei3DVy+YLpJx52LI
7qNE0snMN2n8V9k0HusR3kHUPHLOtdxmF8wQp75g0vmpSxlo9SShLT877dfAyHkK
c0hf8oETK6lNKgMD9bBVuRkYkqhqBasRbLd/LOe0kDtXO5Ot3Se+4Nde4IDOn3UV
Gfms8ULF341E5MXA0rCvBvytUeQEQFWKQXhZpJHe/x7TY5iu/RW1gaZbj+xzQd+w
IEwylaAxxW9zEh92uY/2GlNk5ZZ+3jezkLDQdq5HnT6h0CgMg1+J68gLhEWvH3G4
v/i5qjff+awvKVIi7VMkX8Xw0v9xbyWguw3PIWEbsh8oC1qOATsh0w0FdLFGhPcH
ABw9LzaJu6hZW1xg8mCjcPpXdVwgt3o+P6UguK+1CqTVyyyhT8WEbWnHLRCsvKrI
7KmFk+QGiOVx5JJS22tk4nRk4M5y9+oBfIuSek9bApO+TwKkOfoP+YiEPnOf4l4L
h33AXxeHDOpAQhq6G6UEfUcoNSYb5jFDKW5jAydgEKmIWmzZ9Iu/fxLGNE0VBUFL
RPp27ROZ+DtRArIFTEx3G6oztU9/RGrUqEA5rRj5Bqn7wXjYWwoO5A0Abda9ly/7
qiLBMsFI+sSOB4RBO/2nROFeSbvywrH0KwL0XmcDRCRrFerbV2VJ4+hLqoo1bJQ1
+THOc9N1E8vECj3VfQu+cnnS+HOsFZ9PHFcHZrrKFH7HaubDwnvMBT1/kkqWTWTe
Q2Z+V3T5chGX25ejKRv63rDkK/Km90BJiE9lpGCj8yW4PLLFO95psBAIchgmjMu0
dN26xKXY8ALebk0kEz6FhigfRjR5E6FWQdULlP3vL6/RVqSjHTC1PpObsOO//bib
DlhpeRAkSmDMgqwn93Tr7rPfWq4amOIreakRreM3szHe5nQJGjnRLu2nW4d074O0
5qpW1lKZt7ruOpimAK6bSasQbpsSSF4xppGiRgJblySEPxwOHixeiFYspFyA0+NR
e+ydxQHDlCOgC5fr7/1eGyNLZUQqkyNyMOILXtL0Ri6GQL4wsrMeXAFlSj04yapI
glq1HKcioVjEjmluIhNF/idIagtE+Y+uBBcHknXs9hYr8N3C7wZvCgOWT9N9+DZO
pt4j+Fw7ChH0cedk2MaoNNePnd1jAlN/MHF4IMgyTt7pIL4vpRUombmPAlGjq7ST
077bm6sa8vCFpox5mFFhIYTp+ieuSlPBa1544ZqdWevhJu6AjKCmKcbRx8gHU1I8
TeYnXUjJntkeJ4dzdXEWWfr6+5iNAiaEBIZptxWg/8JjALlcP0bpSulnwyYF/YBM
JS55xXDxSUigQ059BkLj8z+cKMxCJ0MeFkLqTESy0oLx4xWL+ebFr0hQUMuUUimL
RmDUFeVs1PGLqHCtxpXBc9Q9znVJjXfAJ+OO8s0gbaNDMVnd+UPdvbOJjj9t79+f
6FwDCDcsTyyHN01YzcrKcaugu/H5h0tJ5O1wI6M4aVTDZfI8u4BCph9Ataow91zK
liw4bzBCItBAZTa85LHHEctjBxhk9vzh2uyIKrG/xcxWQOABwaG5/XhDXN6EicVp
ewxftCkyOCWrJvLAiT8ZEQmWSb0BxPk8IkVbu2RQvd7lxGmihgM+Mn/kvMx6rRwJ
moxdNWvMdYISG7jm58gP2z2mQD2N2WeA6gabaOa5Jb4a6xZJJHZyeu9zy0ACh5WO
PnqK2LU2iArMBQENo6g4nxCFXyzso83YUXMm733O59kuWafwDMiXhaV/9M0oOS5F
hgtALmCb0TflcuAeA+vem4IEHBzvxDN2DIbOutXTwx4EGn/2ZF1zwV5cPrNjlRra
dbkAeaOOZ8gv4AUobEgX9ZrljNYDp3BzLdch7+XLt/Lu6Ppl9uD8paFwaxWH3a8e
0C9BnyVqROR6FrLaq3ytNI+QnGStBTO6+fwechwoHkdqagNaHqQsKnJEFt5XBL+1
WqCmlAHx7yeld0MPc5tq+pD9QNFP0yqlYMujS9mb3C5Pvxac57MglAC6lZwx92Bj
ZQ03dqIvsdg8r+DfYHZI06guYkK66QxDkhHE69oAvvExC6NNcrOznajpGx2ryrGk
swCjEMZnEmEIYbqT8s7JbfO87uV36M5/u/5AB1RRhQ1mSFOuBvVcSvV3kTjYdjdg
WbZM9w9pe1IM1h5ya+ZZvE0lPvapVOvjKH9G3kUZbP93RvNnqhjEsWPEemAo8b9C
z555KzuQVdlvo7EY5TmZxQuUZ1RA1Gdvo+UAuhUv2ahMEKy4OACts1yW7C7EmST7
LIhX3BQPvmPoPbMPDrOqZOg8YK8d1FBXpIqf411BQyVlPAJwCCSYqCHblZg3Pz4B
Bf1XpRPYNbQ7MAyjR0nB1MRJsLjr63kRT3w+xypz0Jm+x1BH4ff0D6tLX9i6oATo
LmFZ8aGfuH5dmxWBYOmT+EN/LZYwqhaVCSri19cPQK6SQ/HQEIIC9s7HFrXLcsbX
QMzZS281JK6ZIox4Tal+IhRQALbSokUmINXgus+Q5a3AitJS79lqdggDGw9zuMIX
eJYFCOt2M4hGKoT2RVRY/vHFH3n7f+VFiOBGXamyUP1ifOFqXawVOpys7DcrQVB9
smErlNDyCMivGNpdB3zG9jb1FzmQ1R8o5C7tmrQs0HnLQ1OrvU06+K8NFM3hXDPe
8eFuL6geLEyRxjK1mTCClaKg2iUdkktN8IX/J6hhARwVQe/aUHmyleFgmN34ApMc
o8w2e11g4fy6Tq9ROwe1a4HsyKekayg7gkkDrNHGuakgnUXsOETyrATIdyzpcx8W
gSxux3YmZgxUsTlaUgQv/WA+3vN6/j5cPK7PsJJehufctaBb0uOtZiFwPDcoHzIf
wH3ACkz8OT5HV3Y4jL5wFncUDmOxEMoI+7VFqHbNFCPpvczYswWmDFSWVlnSOFQs
6YPXip4pdJvQDEOM84YfAGzxz2dOGHCtqExvG7n9yqGGztDyKDin5hrEzbdjNg7r
mtJwaC3uvnrRe4uKO8/Kc7wp77sTTqUl0wTYX74hLrzNlWmP9ZXzXRqvl3DQNDkh
wSAZCCA0Qatl43ZkbmJuuajrCpA30Ra8iG7fDgGaSB8hd/S2g0SuwwwMM5OS4JOI
KR0nApNmfy7+xF4p/NlonIBXrZGvPeyebZZKwvt5Y3GMUd/6bkY18ApJUpFZ1Rqe
lBqGx8JJeedfB5Z7XLMrmh0Ja8LKKZ2db/3w6YNDyd1VsUFMBptqjQNRSYe38icl
KPoj4veC9jX2zrvdfLjLYsoXKPVIgbt0OYKijfZ7nGDSb047PeejKdqP+ZjHDXKv
VFS3KDgtwOt4h6oNMJU4RcZgzi/qoeOvi2HyWPcjeQqaneqPP6Ub244jYL8ljyJ7
d+MwtTUh6FOMXzF5mQVbZES2SETCmrX+QWdO8AJaC+G0v0weadrkw1gM0UQvMV1A
aJ4aLkdyiOrjkpeU112ylXAwyanbUhyDdIpeNxV8hh+uwEXaXt4cRwqGmLBPBn8m
JJm/VTtFY8xY5dZ4s+jZt0RE7MIknVuT1VDicdpR6k8GE5QKChIZRBZ8781rudvE
QSt88poYdLbWjKKFr6Sn/1me2YKWy6LVFGw08BCZTSXRqa6TLKcR7EJILQhaazqf
bi5lsO5E4GR0dUnduJIUbnTWBswRJMReEeVugr0la8AyXM+IKiexOU/b60hS1cRC
kUM2LSMGh7T7c5x0biOddWLtbHr1P4bPkBQKtM8J/g9noPFr59dKW21+QOvOqSdU
+NispHhC+8/kXixtELksRNyOjLDPuZC/NNXqR63MmWVGKZ5aKZnRvw8Pan/DygTz
FprpzuGgxCcoLOt3ZJTowAZZGvp9UKGdQw5CmtYBeOVGAm4/VgsAnJEtCXKHhGIb
YFJBiWw3Cy46PyKS1gGxhqe86vo+4V0OJHbtB4p7b/OWuQ2i/8AsW21a4GSNL1jA
UVRUrwBxEb3Q4GzFZPNxq+hj3wHnL1frnpoHkgSW2yEFtcMsa5mcc1g3HBLLXrsk
R7/YZaYQg8fJPbhwiPvOXtd3A9nmsg9V95TspxQcLFvlm3QmcjbpqYH6Jj+GQZ+w
D3OFNEykjMlKD8KwiGtRcIGRMKOEQOWwKmhlyiinOvYq7GNcPvXsfyijul661iE5
NfIctdZYFvMrXCoa3AmBzOZu+jKjN9lWB2S0NvZgQ82UdG3RFd0g21dfYVCnkmXb
l4970FNqyhTqkHdnI5RkcIXlzDNNziIeCRl4caPq1ryDG4h432O/ZnJ00w7F6fQ/
SWDGUlAzPTLn4vQo0U0NsS9iStpMdIevp4fCNerP1vMhiqZNOZG3uY/uElazGS0b
Jn774j9Lq/b4fLR1/CUsQMsZgXVa0zIKZv1SRqUL8N/wGTSg+ETu4koTIRGq22nz
GzzYBsc3u9fV2nUPZdFWXT4NQ4GX0keeRp7zCEnDbUUBHpF3r6gynOTv6DSi3VtL
l/WIrW+AO/ZDRu54Y86B7vcNG6DOM1At9w/2vHyXzN6EeZGCR26Tqnv3GP2k0mN2
DzQ3mheFVOIvDTjmF4VkOpq1lLuIyNOKuFprOMIMJ0bcN06HJ6Ge4/eAZh8Uy4+d
pP5fX9p1z435PB0nhD8oqXttB185AGatF6WZeoHtSoiCGcXTe/B9wIQm+Ip9F6RM
ZOsGDjSSRjdIhiwe2uSzsR74Jezz2AdrFk3N+34xuDFwVifO+rVNyaXLVHjT2bsm
mefiGsjwFRXjLwWUMSYrGWOYTIj0OR94VEiCaTN7FDXGQ01UvTvQxk9vYKaYueQf
P3ffCsa4ozJDGZo92Qq4vYcUA7xfBzJOKX47lLTwEfO5ARF+DXpaDvzp0uDnQM2d
ntMj/M1jd0I8PLwQJU4tempxnN/N7ex5g9avwend0nbIi/aySxUke2RNuZunw1pO
h92OJq5gLataGKjp/+ZfGyz3sUjmGTP4QDTKbJIxr/KGpS1oSIMvQqoVweRKHH7p
FHVU5Pu9kQEOoNy+qTHHaPT2Lqfiy27Ds7R9vi3Trr19xhmxESBWfYjFBOH3mvHA
Fwj4b3Jcv/ixnn4onWJOWxTYIEGRujsRwu63nVLTAeKtRYrpgIChVsy+HAdwVM7t
GxbAhEJfYDIcXYmwAJxPQnse9JWpruRmNzQD4xIg9QzvV7140Z7cINF08lTntsuq
RwaoVjrkdX0XnJrF0ofEVMI9jCxbTyLBdvc/8J7pzE91nTeO56fQbtyezArx1aE4
WyXUCOX1Rd69RJqSGssWt4dSYz5ToFxi+oCE2dOMNxcrpv1ncAo1R0/zFL75G7ie
gPeJAnyVS75ZdBKHeSgxnYAS5eq2WvT4vwfa5ohPwAdUm2hHLxKqdST1ippexx0u
F0ZhPCOHsj3WBxYtjD7I42TEtY1XstDL6/M5Ra7tFaab8JcwxECwOBKD7H4Sn3oD
Xs3Z1tuc+3kJPWCyS2mO56JQZXHVGq2mdmW/EKFrjJjtLX4gxt9XbIf26ncZplpq
GbNNMGa/3/+2wApifFmRzZyRchxSYenMFlsnMn1ykn5PEkYFWzFuZQiumxDCsJQo
TFURHDHjs60bcJg9jfiLcA9qxADL61VhTpFeQqZmiu3wJG3ogEL3O1D1QN05YaL1
TCiAzA9d67Ak3c2blyUD1rylyIZVm45El6C7Su7h0xdDrbB8g6F1GYZM17YddWij
AlhdMazUDQPgn6ESUQ/q8uyfYekwlUuangQHweBtjokLs09IbVpe91Ks9ZbqSxQJ
S15IqWroU2y/CS/iKTfBXDlV2P9ADXHwSd81wpVeQujENxlvwZofp4acOC2JGLp5
8O3SCrNjsDuTD987GfOJffNav8AwaV+fZgJi8RcI+tHIfazhSCLDct4jOGL1ybG6
I9tvVK0dGyjEJ/xr/z4++QHg7AJcqTWaFLBisaL7biaD/Q+j+TjerJZ+7ocQ9l75
l+aM7oRm0tiebXEC+tjReSTyyyO7Yf40aZtlGeT/MCE2RyreczkOW9e/IhgZOJc1
KHc1fVPx/P+wLlsFIPzdvQyF9CoX/ph4wwD7Pb/nTTrXA9OFZoa34oE7GB9WWepM
rbEcOwdWsrMOJYNjdOZLWsK8mwMUXbZ1O3kY7VsfjFPojWrf7/UpgoXFPQKGJxnP
68T2Ea4MVhQ9kk9i1htGT+HfZU64JjyOiGpt/+ctRyU12EIsQaXAl3CNS93mDgD5
j50pHDdKAeAzet+JAZq7HjW72UnjypgjTzPsQcI/5Dh2VnZIwtYYA3shXCiu0eK+
fbmQejZ9B5SEHq3qU3rSz+t8QHaRjxOZ1F63xOifgCRJfdwh3jD5tAzg1W1ZFQzG
Q+8ROLv9m70+gsEXGFaNpI/8Qq/D2ytiGOYyguOWGi6NystBR8lgopWrb5JKihpa
xpUNoCWaaLrflSOi5L79v4Ky+yoNFSy36z8lXCj33/nDwO4pBejBNA5GXt3XqUhd
m/ZJGjgu3blo4Rg8VtwlUPuVILpWG4fN9EGOGSTfelgv/cDiB4QGLxrbKxe1hMEv
41vW00+rmDeGSooCI3EeJzHSMo+YUm4bdjJDSHg6EOZYRVTLavBrpNHp5lfx1ufN
H8HuFrs1GGDuDJFpx5qLiC/A8AEgm2tfRvX7rIDgyiG+rS/2XP0HfxyRp5/7IuZf
qFWMr5BTzOW6GWcTJKv5mx5aUOXvv7pMo8aXjZRqfGduYdVShiGoS90gTtr4Etvz
/dJLGQTsglyTpjSXAC0yWH9uaA5M92VhjTb1kKjdt7WkVAFot6J9Q0kbX5Y3Q4l0
gUeojlmud61LoRFns+m8YX9UoSy2J+EuRN+1itx5hc322vUWjsDBwRs/NPzjmEve
7uRly/HD/I81Ndrvx9mOagzoajw8x3Q0DSXPdlfsyxIos93/noLN4hXrrrr1UWk5
RhmFeHkiszJt6mB4IHq7woj76y4LRvvv7wUvfpdQiAeamlj/pOK/oEk3WkvM4jXO
lkvSY6f3yE+EmJVsoCeaHtg2oPf2UvG8C5zV1qY/HJzdS6HXEiY4zfvJHNjk4UGR
3doMJnv/rVWiuj+CJW6gLGlTqOdKQkN+OKTuMWx0hnzWr/6ry1yxDJIdIfP/E5NQ
IJcCQzsTM6H5ncMTd/iacjEAD7wbJZHAmNI3VugaK1MxoCMNyfV4QMAjE5+J4wVi
+KhegSdoYRF449R0dX5wUozThWSlNbLYAnYMth4g3SBXvUCzUy7diDd2cgzASZR4
JUF7NBKSjugxgl8U/87e8RWoiyidjvlS6F8DnmFXp2hjgm5TWQ3O23BMsx8mvacq
dzq2RRL/TEU2TVfAYBlhhBXD2RW1vhQnSJ+Ri9Qz48CTi+/nSHclQ9eigzgpE4Ko
MhEuydOB9mgLoHIsWivFR3Zogz5r1o71QGJmCWdYwJ/MtWlb0RQJXimDzBqJBjR8
DrksAmu0SrbbpBslCJo448MSVSQhZypWIzTMfocgMrVne94DkzPoEl8Khr7ZlNdM
xbiZ8lOVlxn2yGYoF8U3noGXuyMmzdvR1UdP+P3np9EKQH3IN9tti+NX+bOhwWGi
qpNPmhzjwtX5gJEh1z8+mSM87IUIeG7qZ7DpjVK2l7JiMnLxfgVf3KnfRZvhsyIa
rKxd0Y+w+E/HIAfBf6LhNbPWPd/ZHjwz/muVafMrsS0Msp0v86hoGKcmTOg7UGZl
mrd8S/kQALsPxN7ud293dEPR7U+UQlyb6QIy9QFEx62Sl+j0ptne78nKmok375Ks
W+LJC0OEaRi3L5evoc8Pe3g1z4lLa4eIEJX3nspP0zvAXUfEB3m3q5T4a7tkq5h4
JtqhimemKT8OZUAI5h/Ew3gRLTecGR9jKogoKrRcAT5GK15vw/zZ3j3Bcwyy1wSc
xbyHahXgDpQGyyV738fMnAKcUimgWk7EncHIpxVxexu6z+xgs6diQAeQ5p5ety20
2i+PxqvXsPxuyx12OATxv+gcCwAL4IPR4/O584cqZ9o8E1FDX9GEGsHHKQzcuSeT
No8eeTMj5Q8CF2G4Yb2XNgIlkOTJrjnDfBtgUrx1jeLuhdux3RbmRN9vsuA+Mq8D
AeTRM/xAxlwuHrTOengOB8VwTM8f7XMI6z1luU7afaRXITbfCty75YAJ5H68lSmA
G80S37yrw71m1azxvU5i3OwX8PmQ25xxApdQAFW82vC3Zo5xZbnyQVAY/8x/sIEx
fwgYRg76yTiSW1Kft2A0kCVuctXr+yZk3izEWDSGwl+yrKBGftgnS9XIzm3Y4Egb
HjYHftEcu19uNL+Ni5lPN77MQs6/hG9m7czCNHQlWIr9ncyYauGU2TlaE77Hto9p
ZzgPKrOdUbKUf4ExZhPfCmv+uKMu/dwqcDRi7PEK8SysA6bvGat53/ECiuvLj6+R
47c/xCvv5F9ToPtjtcpKbkndtNKCb/KGtXKMPAymk646zk7HsZcIz7h0F1BAZ4mg
SmrHuKerAg1CQaVNKqIii4zUeB8QCm39ml6EQht0fZ5LHRpELcO+Fb1y3I1TLRCt
R1u/i5OOQLQsitgifzR41+MHzvw3oF2+EVtjVu3ehBtPrc6MH+WDO5gPj20UyU8A
TzkRWaIvV1RP0rG2z1TSyr6hHqn1FVsOSdcK/+xQq2xykDtadSbB+7srtQEy6Apl
ssYCQRDCw8gsYuK65CAo2eN9eCfEegr8+af2J5D0SYiUMrOMXtuCx945h63t7F4b
II9yQprsiKbFJ7yYjyXAXLqFxzibiexhlr5hBj0UD5iihhmaIWmAUDB74sNJUd1G
4gVCAvUtgjQSf8IJ6LGXJu7yYhNKCqYeXb8ulkLJMjdOKLhf7Hd/SIp3Y44g3m4j
J+io352rd4B38PZFAfbcQ2Xg77Bl/7r8qAJrjb5a8YzRrRgk8G96LduK8eXHi1C2
vbvpM/GrvNLoJqhpExJdLQ7M5htyG6MVLiGR/aP+h3tI4PwlKCmqeKSoLlsukP7i
fRld0WWPrX4gJUTeR4DPc5OFyYFeTpsHz7TaQFbj1ous7eOqbWdGr15rrUNWFcLL
74dPMeW1WrhyAah7wfxg2+sDWIhiDK2jeegb7ALUIayks7La0jdgEo+2x27uVteB
fgSGbNdJ232EDBaudZXUh2GsJp58TFByS0kw82POK6y8N8Ji8xuWeUbQ/oTlEv9o
BFzyyP1V10vN309oBcUaVqItC7jcXL5CCdUUtHJJAT0e8b4jJiS9cEh7GWjmmJkS
7lVfi6LMz5zSPmIMaw0AZhqlEi+aQ7LUcYleCEecxwo3AU3fJ7myjC7dKi3eV50y
+qdb1+/AZleR2rJe0eS/TSRjenFlVY9txqysAbD4vrJCG7Uao6cEsSVD5t0WMbAb
h6Im1YUN3qpnzIwvvtexs5XLoQbQC0pO1DJp6LPBDDJOzIITiifESsY7GV0DfvNI
Lu38Fg0QS7lp9UQY8vd3iClXyzaI/utPupb5IN44yYcwA7dG2pI48tt8Nf4r3Ki6
+web0DzHjtjsk4o4r4WnAJcE1ryfnWJagjQ4YBxzVFD+wD8L4KPnzm+iBnckA2Fv
WxejacJrnUdo9ZegqQTqez6WiMnLzHVY+M1DIecRXk7ORRguC5NjSw/mkdfmBYPs
ijgjwI45p3oP3fFmvQKmF6MRRF01ev/OxCh42Hen38MgV/H5MUqZNwFLgzoh8GeT
badH56s6pzJSNpE8SGMLByZ17n9L5ePv+fm1exyIVlaZTEb8agZPaJlxtnCHtY2g
59tX7A7c78igpnnkQPqDMkVhEs6o1p5CProAWFLT+A8DGdchX3f+inD6pANr03gm
9fdQeKpieR5bONJUeYpLHsewd4VMUoNQVtD4HxIr7W0Xs/F3IzOHPOj9HBWc4idw
syWm4IwrDBWZLY1He7mMG5qGnKwLscB+ekrSBvVBwVJ8wcOcdE+BIY+FrwIjsa35
aa9G6ruR9bhpa9izWas+HVhsJ8NmH/9UvTTB8Jx05U8Wsa+CvDtmROA340l6v9iG
DWU8rqe7+tTWiodD/cCRu6eKeSJ033eMwg4dJZXx+4WDnHqBb6bFENgK5XHACXoY
7YmZLoUXjLm6+9caQFYgK/LIl3sk/leGfDdoORC0UyqG3nZ5AGYHsU9xArD1pPnT
KbJxYX/irwOTarLUVQzsHouzGrmWoWUgQh1PmuZ49avnJh65Fbb3LmEJPC/F55uU
A14uLnfa43DDb51maUz5V9ljT1r8qSGrMMeNRZzf8yRCTP0QYaGVthIXn+prSyc7
ePgSk8h89xjHnrx70pIxHt/5n7MPFM3JTKVlhkIBLG750vSxCW+Ll+pf9RrEYWHl
ybq2hTLDCgC9ZQRwIkFzBBPwKLoW3tJiznjDvBWEmYYZhQju4da+oBq/sdgqIPir
EamjtnTU+DjZ5P3mzkvQQ3ho3kINsZ8p+9FMpBNu2SgULQf/4ymV3Cg/Nyp4f2ch
7v85eKI7U+fAcZoEUG+JkEZcT+EqXWxKagzSRkiBmIOqyH4UtMbWzRJ/1ezhg5Xw
PdghHLNIccek4Sl9mgZmnaCmo/r/hfuTPYG/xZxAJyzTqOywSl+nDgy/QylMAwwx
H+fGt5bKA5taAaNRZ90s95SptdL7hfCfYQdqXHZWjDDS+KsHpjNXCvinHVbRe14N
jVYt+OXpoTvnGDBOYGnJQf6Wicm1c4BZ+GJoWzDp9UaAEnkjPAnwFO5oW4Wy8e22
g3d7l3NH9+MaYKkXBPcFRDHMP3/NtN2OMg0pFOnXAAMBHWexmSGP1U68PVCrsZWB
gYQW75pT8FYi1LoQzp8I7lJqazd2DehuUMQtp7Rf+VespXvuT7N9uS3KKWrB99Kh
+jc+agzRzffDlnRw2p4YgsJ39mot/FqdUZn+lnTxkc1nGnf84hbyFZO9h+aLrHtU
e8tL6ozAGqMqFeEA+Akc11BVMxzvD3GZigsTzGlQQhkIcQWJEWwhJrIYGAPmD0dN
s5WBw2XxoTFnHcRJHnT0FdLcBeyoh/1mkXZST/65Ho124IpwRrD0IUu/Beanf5yO
Hj2O47ZP8Kq5yM1yVMG+0pZbchNegD6hWcTmcReGCnmeGoWKcf5Sj3WEwrjPbGPe
sWs/s/KbQaV+WP+CMTV3i0GveSSvHBe3Kg8nDQ7Uit2oiGU4BcDfDAIPXwTyB6ug
TKTUA+sjs+Mn27w3DHYuyTUffBFa5iel8e2RlhlyXAotPITj1NvAr82atmfsu/S4
TSrxChnEuVT66a/pGEgrXUcK6ur+Luhqe2rHdxaCGZzNN2iuHwtTWTKyj9qTCh+L
j9etz8RnMv7RqKXqsM/31oHZDkxVmIIb/IIynTn+pa3VR6NS8mcmw9qCX6cSVMqz
9Hy26p/ddr+neLHqqCV4wXayKV6dnMwi53KCKRuKjoERbHv+RNsoyGR9pyA+I78B
aL5REpl7a7lb6enOCaUBvMvIVnalCkXNgjuoL1fDlIO3rcRbBRX5jFZ4BKR4/yW+
8x4LPyWcHN0sCugqu+WbE7VWOQusyaKHX2Vmt/PdzC3skiYazijcnEzLN067kw+R
htdhpaEHz/Qe48IDVDl3SvmWr0vsKOwmAl4igEkSVfkWpu03pSy/kaLBMP26fFqZ
K2zRS2itvfnubzYSzeDCJPCWiivUAPufMT8M3OtGnHB3OKZIxskJKkCQUJr1IFdS
zIzZTq8ympThGknvEZjR16XXVJZAG1z+bl6shp3TLZA49iV4+Na4HR4FcHuqo6nW
eOHZRyu/F2ZeldWuYR+1m0FdFVna4MxGbyEajqnU25Xcy9Epiks1Fog/Q/UHTeIk
Jdn4rS8onXomJbsLy4U1N90dKJxfsAeUe4JzLIh+1ok0V3ncqa+C2e8OXvlAuEJh
LFBhcRCM4TGwZa4mfPZLAyaMro2X6jrWA7VxRa/MQnF4vnyjpgWltjY/MCeEBmMH
SmZ/kAufTjLF814Vrb2iy+GHiDzXJ28nsqosjIwVb1+/COGSZX7Jj6anJB0G0GNh
oECI3/9KnDea2oa/X0YbvhUFr57jyeeVCR1OQvQOwrWjbOfEy57lAbJKkFlB0KKV
odSBeHIVn5zTGjTsZcPuvatIQUAps29E3o9wFibYjqksbwXkYjh2RW4npKIv3UyB
F7dznTSxbYw0mJF4DCqOAVYXLujwOlX/JpI3o7hsYPvtLh2Z++5KZ38UNwGR0Xgn
C/husTwzqrl1JLWJ++d7qjg3C+Wqrfev3WFhhLRnJnLp3QNtSQ7+viV+lrFnSzMF
i/gVbSm79Qz7hSvSFscDtxcsWo7hUFs5k/COo+aqEDGgO4mYnJ3G24oA22JzGi8b
TJdOW8lTVFKasB70s8CA/RWJ2mgeSnsSpMkZ8/HK0YChYndFusWn63uaP+w8uZmH
CCiHrr0K3pqfjRfcIROB8DHgzS5SPvDlO4aGMbG+LlHfou+BSbz/xTrPPvDVqkDG
O4S439ufY5TeMqqtYIzUekIW59hOMBtrpC3g1ATNXFR+n9pBzx3H/uS7ww/jlXL/
oBunWBwnZ0r5rdtUKQPvGl8Z9SN8SPzpPFPMitQmRznqWr6mMQ5vcTeKQpoEFenq
P0/+F4zZPRYTC1nr62C8tJyvDpdvj9erKusaB7PKOLJ7f6gFalWMB0wxxdh4fLsV
6ROPv5/2OtwJJyVRgCA6/tjEhI2MEOnQtrx0GWVFcNZwvNkzPHKHEwKUr3FsLPgM
O6xRKXmXNmzo9X3UCWd1iXhcjpeBsh14Je/Cid0sSoMFhItr+maRGMD4socvL521
732VxRsRbL4jFXRrMKbxPUqt1E87HvrRmH9cihEbz5KoeAscOQQvcrL7VMDwD/Pu
PwvgT8EBuWXmfCp1b6M59yqMljytvVrlMJpuzhzlcUAjMnRjilu2WyH8YrGCy/p2
Eqq3Lr5l7LJrCofPBzFjzmFpBXxidCQal0ulCeC47FaQOj8yw2IWvKkLK1Y38F11
hfLXJPFmE6QXXzhRk7brMWj4TBONlJ3Z4Vi+Ia3Fvbxo9sa1cjtxVpitZYKcuq5r
nEFV9c1dbiJNXgTkCfWzGjIBjMbizIjwLJTCiKF44A5OyAvXlv7QtUA61ACKHfNC
XRQ/gNlyhyUTWXbd8MBlWrYL2xsvQUe8PyfXUB1kcUVVp7YrBRpz0WlFgAfdpfSX
x+t5l7y6SrZsPasP3ICuD3nbqreJZH/XbEWu+7UFt+DxRvcYZRo5fupj34FYswNq
3ZvM8dorh+KKcz8Q4CW8zvBtdEzOC3hj6lKfqtmbNarKFqj8jJclkYQCh+jGuq9P
7ggah8KkqygymdFItCNz1kvupyUrJ0cP/M2wNZdrlnDkI+14fESFnlrANp6aoyu1
8vIKzr3LbchXlj44S3xFPcNAxihyaUgjawO+hog5DfyDFnKUpznuNtNBe/zGG2JK
BszU1ynVP+u1KfGmhtz6TLDTEb71QsK0YwkDwBmqCKpuPcsVBM/BuGpOUANVqArK
4hecTNTI/8Kkb9DkCPNloxWqrlpHB7gomtgL7RhS571qji1z0vfY/iXHUTNz9a+j
G9DYylpeYwU8WdpmBYZLG6E7p6qgrsuQeiNh3NBRVXrw6JKnLCKSwzE52MmonRua
ZvjSVYZd/aXTmApAox66bcsf96rQAFIp+TJRiFqG7KgvjORbNThrmeaWhnbiY0wR
A5fV/5x+niHmrJ6F15F103mkqvIQQtJGuQhVUusjWqoS0i8NgON7+a3Sqircks2z
tMBTHA4PKJqIfDFdC+5cL+BlyuEHu0PrYnZvuUuvqyl9VVglFmMxbN6nmCNpS+Dc
pvKb961xgfSgGPfgBPoLNK36zJONj69Qm3ocUTdHt5JyR0jkQr4FMkYQtp43uD2g
ASVZstBPuvBHSKOAcqG1y2C4ibqI3ftPGthuzf9FyG1Bu+vkhBRkTFIjWv6iSnLN
MzOfh/fxkln4HilGPt3RwYyMNqShXplMfDZhKxhBfEjOWlSlal5U/926hMnkO7Bw
qYH0AeOHnbpj8NTZd4HQsLJfcVFqiaNuggZClbZZrHj5semeGvrqkYm34NHGt4/Q
jbSEaZyK+ct3IHXQhW1ELQ2rw8sXt/Zbs54BvI6Cpu9tN7TuCmlINJjmECBdHMt5
czxJw1qDp1eGlpPUDKMtZQfNtSpeLBpDi6eFxbym+wfDrLfaQPvZvdtl8cSOTPOF
N6sfCay/Le1VRjoqMAcxzsaPLifaqyDEIJ5en1+cli9i9u3BAam8e8LNvOAFny4F
fKLYhfezrBZKBBjqY6XSAqSM+XfF1bfUn25LCwXqEsIrXTtcuLLqmKUI89AHB7Fo
FYU4SRTNWtinU1I6d0mLECql69uxKbCIO9fD3PnNEZ2xmyI1Mlfg4wbLqWHxbGxC
G5wbprAaJctfxQ1EYDHPNpC5txAbXwo1XIEp1XfXHDfqRhbPeHC3rY6E6SunVepv
sefeePgpBB8c07RPXRHViaIOxYnWNQAC2V25APqiAXa2nnnFaXi01ZZEQVsAWtb9
DmIeY2BJmycn+g5QvabWN0A/NgIIOGa81xMZd3x/MG53hMlcUh8r9CbSeYBPipOM
a5wfoHsaP2wdrHyA+s0JqeII51BB5sml13WwW0FD3A4sYeDyGZ/I7KFIEWsIH0Sx
AfOEGLTVbJxCxlP8DFwVxThr7Agmmc3ta74KmyxLbhMDb8a7+Y25HWX6zEr80fXT
g49cfvRDOdy01D8mFBQNtzETdjQlHCp1pR8RtpatY8ZE19t/MBF9WBsGuudaa9rS
k5Hghggn1IQdOeC1AUO5IPhVHFmdBd1lMpTob3ufk+RBA9KCNg9yDx1WnyZoFscs
X4901zxp05ZhPiFaf+z57ODkAnnudkCfFUfGZ40RNPo13ZJcdsumPAeW9smlDzSc
dZFQrvxUVOJMPspNFRa3mT03RacM2/48kk+Vj3yhDhf5WnW06szkumz8x3r5WBux
64N1bfJZf53DihOJgotTplmXEY4Mtaogddgi5UD0weP+hKNIGLdKEv20MP4/y6dx
k6MEoWr43TyzWkvH1DcPU+Q6PUi9pf3nr8mLTK8wAyWFgWxyO6KproeFWJzxUg2i
aJ3bkk87ke3+hz+kj8U2DULF4nMa3M6fRya3nN9CjFUYQNcOaXpLOzjHb/YNaQ0u
43058IfkGJCkowejhDzX9u5wL1bmd93KNJL3fq3at7uiBw2I+rcCU3Xn1mcZIcXT
KfewzHSMjeRMd8Icfm6RYHWuVebjfrw86PuLCh5QxRkTa1mKTOzT5dIJoNfu9/Yp
KnXaqf5EYMymbuHamfjRQEeSPEK8q6LYYo3hyE//g5ZfRUdOSuHr/EAnlrhTchEs
Rb06QSPZvZA1MwgQVUBATzkomVX2XhCoiktQFm8/R+sMDG10Hgpd3YTv9fBdjJYk
FxZ3cIySByDlrzX1Hm+T3XmC9gH3DHPPHv8q56Nvg0Ks+lJW5A26L92fuDuaoJsB
uMrQOK9eF7dCFBau0YXKNxBU3jbeyj5KKvArxOz8K8rwLWoRYwOn+E55sao4X0X0
lWzkGKWdUVfESZzYx4uDOL878UWRavl2ONFCP3kG9SfPS9u9sdzKJuFGlM5MXakG
93eDYv17RutESoAoGA/DIRjFZxQIjEGqVR5YicRd5M9uYhrOBcmH6wU0hZIBBMqf
MGNTOAaUMIAI1VtVjN+/rFXvvzpPSLVrP2fage1Kz6+K1uO0TlZ1zUnqksEBNPWE
gCiS9WdetE3kYtiT0eHJXcVP90O/oUepSag2PSzK46iMfZ8RY6UsuJIsdX8g7GBD
+ecIgJj/OkoSNuKM0r5WuPZofs0v1+eHTXNoqAVxhu1N/TgIMKlkkiSk9J2hKAuE
ys93nyqotgXny11icGxJZ7CkWFNNlnmxYik9hTeCkKmJK5sUhVk3IENBLvAuKrkC
Qh2Trwb66jKP7iqqTub8mK37rgXEP4sUc95PrIqz+IE69XgrlWvbl2kugtMXFREn
dRZ688662DMcjAHQ7TvRCvxgrr6oRWKTNSbitOJfqDJu4oSLJHwyVRjgmueIQJOY
oRHZAGINr0pKBYp4J/Qg7PjRiUeUKghLmo7ycK7k2PkLTomMc/KSiHTGbqXC0ve6
SR9B1z2ok3CGP59ZuWqeSJ7ueBrO1b9P6+td3ggH4fphBfVgEcXy3HZtU4P4aUbr
joHKI197QOfyI88LOZA7zd4F007BFXwYBqAnI9AFlLB3ftHwR9qLGxztjTr0/JHW
r5Jpgd337K4nZgqPmwo5ZdrcGY+1Ng3Iwh98c87X87NZojXw2Lv6Z5YjYHKE0AE9
LWOsMF9B+eYHrnbCnGgT27D/wmyVL65mMQ62Qnw2WSUWrbo9MfZHYjnbKA+6Ak9G
4/7UnDORceAuWhLFUppIGl6lCa0UIhjqQzX6vrmDvjmri59AsePX3LAjLVVExgPm
gptU062ElsTW36uFKvROrlABJuNWXmDmDmloyijtr2VVpBX2ME4MyP0BNtH8Qm3K
MfEHJIa22/mXtrGQ+XMhKn7YjP9WxxlPFHJWMlYIo111R7F5CrFFFyZKVkp/6+rf
g5ep1MA4KmzycgHf3TVKrju03VHbnqOL3wh6fd60ytZSuDYSbRQc/9SlcJZB7/58
2UH25HDzFgvEhlVKRX9sXFsBhQIHW9UdvTFxgn8FIvvORkzacDSl3FshXlQpfdPW
3IbnvfQU7T7d0xr8Uh4ZdGmysLwfcr/+lOk+93bPN7IPohY6dKBF6o894qiRUfva
JFWIPDvzQMGQ63bUe5tIDi36Bl1UNs3GDur3Vp1U8UizlmK9+sgonFJijYex8e76
+HNMxBSnPmdHwEremoikUQLZ+E4jow9WbcFAsgzhciST/qZtRCIrEF65MfodzQE/
F6Uj6BFeokLZxs/c/wQCJeP5Gd5u0rHow/HkKrnvyhBBJLl98qy/uUegY8ap7+SF
sOszKgYkfwxmNqSKXQrlbKdc7DQxO5/JsobEzgYTC3AR7h7bralTLg8BaY/VjdPh
y5I9ENC+BcwYlBl0cOuJoqwyQHkWRIo+RtGrvBWzYIH4wYucvGUhiCKVvDQxG9OB
RsbKla1DbwcnfFAgtBSfAf+31VM4pGg+k/Lv/preAUldNEuh7fV/fee+5gAXzdwa
UVhrN77Kfg2f2T3UEmBOu9/YJuEFlIkHb155j8eyA7hPbARZp8k4QAntZFbBejxv
v6snMPnCeylQOGJb/pZ5Kq/Doz1mb+LgxgACV0oB+d1KLMSMYaKlTVmJteaIllA3
nHYcie2l6Yf0bVmY5CUtXDeIv4JlXlabQc8AYRjeFn7gPE7RFGrdQm4HWOKyJOW0
GUOGlxq+g69Td2eY599Ubuks0gKAeZdE3jc3DXNL/BkKpX2RBECr89KXlwOXeB0h
SDHoozN6R59l5VeNTcPQDTZTTfnK0ysTZgwKH222IAabL9eIF33au8vwsqxj+j8n
lO6IeSHRlOHcWqNHRwYT6WTnf4+JYME1w5yEcstBg09jEpIWw2NIgUHivbsDIOff
QweFqoG6qbYP96PdwoT4rXlDJUWkA47qWWiPZNQl6vH3rHUwlTXI0P3saBPmF3dd
kx/ZidDzdcLG2YJKrViJe+dc7aztrKAJShWj7lio+KqASEKZAI3kBQm0jjyC2PoS
zlHYKKIybLOjfxE6dRCysLiWNqY4W18/nz+HbDauR/cjifRaDyH5ao7k1tBXCV7Y
AMdiFqT4PGW5ymb7/826N7uWsaHv9Khz1GVvoVmqFISdCZm14XrrefsS1S7svae0
cz17e7MIfR8kLPuhqrlRBRIpfJ8MgHrnFeGcRhgZuXk/1BbVjXkqHAlypaikY22Y
JbYpTl5JFEPvFMfR6BGbECeW0adWqH8dV91P9cvS2bJi8c7ZlVuXhK82lH+X/Fko
6LY4ctSE7kJL6NszM+aNOYDe7rw04PfX3i3U+NiQYOvpOBdZpeCg+2BAY8iJdLu7
wD8FjBI39dGSjlha2VDOalKMW04eUhRMC2IQysWkbk95/ZxvxiD2MNsESMtjtvx/
MnoInwn186mi+2HYOIOvH3lXFmcW+LcQKJt8mHs2LzkozIGlCQs7zwnG/3E8yK5G
hllq7snLClTaGwODJb+1ngb1qS4AeCiaA+6T8boCyY6RbZTyaer/9U3bUvnytES6
rmoWuICtEmcrt5ywUfwJrSFFZSH7OqYlglJ4D9T6VgsWyOEXyVXoPR9IG/wO2I8I
p+mjrYuk4OQNN9WTaRkIvVq5cQxwsNy7IMgjJmlFdO1wBpskc89pwZWJ6Nv/ohXb
+xDYUJnT0PhZFE9+Timjnlai9k3dLsuAs+rjKrCBmz6/iqbISlfAv2ljhdxgPTnh
Ys0CknrsOO3cSVcEOxOG7ojvsI6bdXL0xPrU6lDZpHkpUbtqUg5bOelQUWLYoo8U
2J7Cdh8ibQvzw+aka6obkzBaZLC8PY22M2Um9PMAh+o=
`protect END_PROTECTED