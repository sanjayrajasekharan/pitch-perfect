-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
UYurLFnriQ6QC7jyWO+fQDP3jiYfSIdaLDGG5pIRtjEhhvyUWP49hwSFjFRm6qXZ
W2HDPBG/7qZeXpQ6ZP1lAeVo/g1/6kLG8xdGUHUus+qUj/p162njC3TkBC4Eztts
am689CkeRf9wf/9MIvh7+WoL7FFHdm3ZpMoooGS80Hk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 111845)

`protect DATA_BLOCK
eqFaveVzgAUBsqm2rjWHK1I8WD4VXlRxxeEMQj2/xEW98SVlLLbW7Pl0CPlxEvVf
8Bm7PVSZ0iMosMC7H3GOw1B7W5p8dc/3++78irlpgzTfctzFaEIjjMDNHjp2O5ZJ
cPunv+2MnMjrUT6Om5Y3Zrx5Xt+6v8xBSmja9gT5gmpU1H39YZzn/e5PM+kSUpry
m6TUpuJNBj6vhubhmaMN0w8TiumngKjHtsh7/36e3h01DQFiMhD1vos+qSRYy63Z
SxiqsDLouNppP545hbLgcXTRVlUrKgY5alnk2506TjxQM7eNroUQDarx340g19Hg
syz3GClGkXRk2PcWX2Bnw9cdRAgqZcXV+88yiYXX+eHViuR/eKPBD/0Dslb2FHQ0
FqeQLYjLBeWtLUYeghe2F//tvT2d1S1L5pUyQiNtRADD6uGexYnKhaNmGysOOP6l
BHABk+vAjQc7R8RjLmq7gRZloL84o+q6Vvs/WITqe9FtZChKxsVtNOIrAnZryB9Q
diIOI3fyngqJEJyEwzl+ZqghMl4RK/MC9lY+f3BKu3+kAN2kEqwVvPT2mR7CKH2Z
JSWcWfxGl8ow5/BKRz2Lp99zec4ehji+iPjLBA2xrQ1xwOw/wh9sp8TCt9i74CGN
vYPGHSeY3Sm57jPHUARuhrDyUK6FEWCIgqRag+UxK5O9meLATpsWAjaJ5NtAd8Lr
Fp4CHBdSp79WD7hGLRDJcC6DObVO6H9uXL7G6GFNHMRcmMjOjx2WAlNYH09qyTOU
difPjK8Uqo+drUEldTFuCUgTgQkbthw+F8MzqdqiAx8dL6x9eU0B3ZhD2Uys/dlm
RI0mRUyVfqDVjFCXZ5uYgE2AYK67Cyd0QIoDkdcQj27pOfXtq6IJgjhDRAZDhfWV
45btneVhfxVhSAQw9z4yt09FMAZe8JZ6mOW7xqr/Suu+aoaMtRQS/5Ck766DDq81
Mu3t8jTLaZml/CgL5P2l/DsC/3/g0Kncd+erz6+oqqnUGeTEysCl8B6bkT4we4OV
1hJ4GDX6O+Rsr3NOfs+MLdsZWdniR9KAAWDzR9CGXUzDxtB8XDW1yKa/xYXPu945
nLeZ70npS4rgS9sxD4odt6BTqaZJAv9c7KkT475YI07rpQ6D3dnsQEhna1tGGdNO
mE/Lle/K+uFGsEovqL+EmwJUnTyn71+Fa0gPVx5UDNl5yEWn6+eDmFCYkop8TFZM
4830Ca6QHuwVGIyGGuFKlAn90DDFJS4moAq+2jIWdorHQ4mBXKEwY79UwFOWmGYX
CUYxYOqzuS1+DgJvlGQC1YUVSzTVnFsX9fJ/GFkUo+kzETD2VHxLQ3cUYrX8jXw4
q9zscvs76Knrcj4uTZJ6WcqT3AavlT6Gpdd0CDQUD7XuimaiKQSxIXGC+ilJ75eP
0SW0v8CMTs3VVa7jJpBCZdlHiTcU1NokjvS2om7XERP7GBAAuK6lDbLvtx9P3xyz
gDbdaG6fJCfMn6+TYlo90GWNzGJB0tdukILP0XNNp1904nJ2vYnOz3ab8SvzTgIj
fsWh6j8n3UH4UqLhKbMlODB0WBtNVy9kzul5U9+N56mbuhcNVOXEmioT8mRU51St
RpxNfRhmK9W9cCIw+l84RpFzwhWCeWSk91lTyraWidmmldXzM1qa4siKsL4HQiR2
YZENL4qJrw4jpbogqfaSyB/Q9xE1RvXEgwGJM1VATXgMe+sQ9bgVpnqBbdXcng2f
uw8GeHPFuy5rSIaHkbfBnKVFj4QTvAeRmvfSKynOVquWcPFsTZGBNUSXYBF4e9ZV
v2hxwW6OcKs1Gn5EezfsnaRjKgTB4qlnH0ndZxfpBkQaTn79hA7ImIUuUq+15BZ5
/Wf9j8pqCFLqEyHX2XHvLIefpj81XJv68lBD6ha7dgGnoFtW7B7/+rKKRflCQqVJ
v5krlSbOvIVgbDORg91snn7aAkAqFYTNr79/qQdxFU7VBzYsWX0Gt1XfC5WTKZxl
Dr6LebT/iPb0kANHrjbpAWDabJuT2XWu6U5wjVPOyLq2MKqgFwOTARqNC+cEF5mm
a/NemZkoj6/LVDn4wlNxCH2UfWEqHrMTGpucRJGq80V8LrEY9AFCZwG4qtwXX8HT
cLtjmS620nLAihbFEWzGKE442WoEErpAVVCxcsxDACI2kJRKUMAH2iQ1pbVrSZyw
cwY0vp5pK5HUEr/QqWH6nrS5VsyKZQL9sChliuRAY4JpK/EGoM9vIFHPOpT45m7i
V/nZAkURLd75UvQXZO/Abj/gX3+ZeEBTJdMh/fS2Q8Z7Vadutx42Hgc4O3tZ9nE+
E4olfo7/BGseP2q00GakWZJgnekJkmdX5gONYXUZVAXZJE6lvtoHfLqm7tzH00Z8
S1FZPCv+JD75+fIqigH3GItBN7L4cPyWnmYT1sBV9R/oB/uwK8EP6RXIP2GBlqTM
9GtJhgI0S9ZRT6dduR1R1LmZTvmxdAJOVMc1/U0+PekMpAh3fC7GWTi79CVEmzrC
7OR5NhSEgcjVxJm8dEwMyJtVK2a8b/TqBRq1JLvQ7bh+oTa2yT3FNrkjWN0Xyrj9
fkb7PWLUZ0NK1pRXdrAlovK6iRBLUvr32+sBAAbJFQ7kAYi7C7Ye4M5ldxPd4zVz
vS8gUsUkpJevilD+1otmY9k+GB3tcCP6lYKl53JdiYVE3V9iAIw96kKMnz0J0YIw
t9g7fiI5XfkNr8IZVyOUzNb9MEiVsq+mNLVfVALInDzVf27EM7EzpUqPG2HJ1GHm
WUhVKoVZ+wLtrph98zqOgID9XmBqT5BT0eA1AGS5l3tWZZ3H64aD1bP5DCOg6EQ9
+yRMdd4IQcZbRQgPkRz86dNRsM+JbnNpr4xr/Q6wKy5r9XyfXvP2lO0zj3KXT3LA
C02Bw4HnVoW35CbRnuebmcv3jxe9tTBYUX0vKXsGs+vm9wuNEAaCPRsBNB0UiFvI
gYwI1+fskyLp0/uueNLBGCedkH27djtwspCFve9NYTOWhXvZzwgDGwijNKCOAEXf
C37/sziJjEkXzyKJXXfdB+kyWghVAHquTX7DFZt7cYtLQS1FUpG3AR0tZEom6ctR
WY1OzKbcTo8ilWtjnseunSPJtrYc+GtMy20HRBMc+sc7fTYZ7irajQ6mAPDvtOo0
dRxcm/nKwjFRIZ0eG0zLW15l1dzmrsyRAoVBQVvKhPqvOBuAjl4UwJ2FJv1RUqRj
Xi69f/jW8+39SMHZX/Wn5TpWySWX10OH+vtuSB4vznPy5jBS8Xz1fAfC++hjnh9U
ZYnpYo8+osRxNDeQYiAu/N+vZpuHUP0w6zckudCH7GE51Z4VisP2YWLBty8y5FYA
bBj0axPg3IEHZ0Cu6qYXKQT6mqMfR6g/4as9mVj/Q4XHW61zNDCcyaS70u03oDg+
4irjV1LytvadO2Hzbs1FFx66qz9PEOXENziJX2tjn9kuGytkoYDvtG3UNZ8qaXNT
t2Vc2O0jIjjUHF7WjS5LaUl6w5QfR8eTYsDeEmNcmfyh1RH/A+itl/k6mVRSbCcy
MH5T9BIk7Bm9/SXubxSaogQ8VuVnk5lNrz52AeJepkRZM1nlLSnTNGqAOuB4g+Kh
FuX0bxVcV1wPgJ6nd3I9TStU1mH7c/XjFG/q9koWjsLyUyKo8lMqWWW+LoZ3IKp8
ecc7StId/GmH4Rw5PJ1PpXgjychFZvHHGXyHEM7pyIJGzefvT+aEvoqmifmBPejB
/2Zvoqi9OQUq7mEgA3bvi1NmXRQaQBhzwurgv5B49rGvIWbFAt8lDTWsf5v2pv65
llz3m+oKPNM+rpNbH03oXiX9mbIg/94oo/M85+MDK2rIS0yLPCGri7x5J0SezBjv
DUwYJpmF/cD5P/x+zM2wnffCGbWe7YhTnOk14uNeXmJweXlSK9t6TynRVrqmnfJw
u0g2UwLE0EehYUrdyUzruLmfQQRGXXSeGaM3JMWtkL8koRlKGrmZvJqZgJSxZsZF
GQ2d1Owtkx8NLT13QzuGuuCMZuH609U173K9vOOogMmwQW9XSnzfZP2EIJbvd27Z
tp/UJesrsbEVVkIiNSM9H/cqwWQwc6aERpsc/w8IJqd2mf4/HoCSuwGBzG4oEPrJ
mVZ5yQMNzSTlHIWpPCVcIKnuF+qaQjWzm+undPmxWrhDZuWM5hGFqvbY3PJMDmw4
R6p2x9snUAiwVDhImUbqs455ISzogW0Aj05m/sgQv8qZcem1mTY3eQyZNW/qLvyg
g6T+fqssGdNNnD4MwqCHFcXIU3BqWYiyvMBpLeyqYd2+dBez62ospF2qIlNaGoE2
vGJRppUjVcFUvHR9YU7XgIWGcyOouo+1oAwPYWWy8wORiTla5imPig0Vh+1nwxRe
BXSuX1smf1ZhYRwFzdc9JmYAIDxo1LzQPuRMNXplUHX6dy5dj82MYMhhooJQDIxO
DYCaaTM9awomZjkQoEbgTatquT2pzlL1hAuMinT8rRkiTCmvQQWbNZ1MPEg1fQVg
wqas6EVhdkQVDIg6Cvyew8gmQnWvTk4CxAmJxrA2r7IxrXIf6JdoFjtZaU0B4Obh
8SRlY9xEJOi08VRjkNCXjOxFkmseFKHUaAPa806hp8Xo1hFJ/x+uRuVhwTltI/d3
CCz+FmXI+dAbN8jZim3w59PmtM1ttRL1376of+EPoKS1guFTmp3IBJY82NuofOPb
bCEweTHpuK09CUU1ewb2KtndRPHgxR3uJilZMb8BjD0p0x7dhHfLusEgkKpzxCUB
kaevtKk2K4HVjRhLEfGlnQhkr0EQyGHCvxI3Odd1dqI5O1exTObWM1wh3qPEAxdp
h1K8W/Vr6ROEQZroihp6JOHij6B0ENKLJbbExIx6b7v+MSferQLpkRxi390B6W0w
/rmeWo3wqVuQCo4x3RJDWhcVZYbQoj44l+JNb4w7BpL+DozZbic7ls3y5NNTxUsl
pGybvz6CjFRhvkV8Opdtv4EI04JDtkIRDspbroHZ/u1b9Ub5M28oPrJmBHrB4O+O
3KUmVbA6FYlT+XZJf0PjA9WCYRP660hyNwGVdq5+cMrJAMGw1tQ4cpR4sB9BQHLg
4ilc1Qo/lr1kPbDv7xMQvJOIm0jkOiIk8mUPurEIvOhZiddv9R20dVCMWPDbDuxn
Gy/KNKE3QdOtBYx4mhUX0cloa9P9LhYuJLYUYNyXn/Snc49uD5DJ0zTJJ1VMB0Rw
FFFqhOuGblPv+YZ7evdS4pX0MnZt46rhuW0iYWJKALW7L+konpOP7QAMLxQoGA0g
ZryS2Ey3G/RRaJlOK7oRSMiU63QusjfSRBIsXSggXGkkJNzbeN7peIElQJkxw8Lj
i2mUrBiA0dpQFpgmJjLIAfIinRVVU/uZtqU+unSnxqglhdce1SKHrUpcKj6UQsqD
gVtBFefyDQoJPkeaoQFISFdusuUccpkMwflnUrAVkV9HjDUcuHQSN0Yeiprm6+Qj
YgUgSHYx+DyKtdvVypQWdWeU6r9KaoldJuZ0Xz/HB93Zfw5gZ5vimOrMlksQc37u
r+eRdnkm8DDfFaX3/rpkIk2soxf4lX2rYeHnlE1pCDEHdqb4tWDsHlZt1wxZsbQp
1fLQKsTzdiDvleUg6mrn7YVptps2+klHKF3xF3xpHWg4GvgAjW9kXS18tIfHA+7i
pG5/xbBm+aNW1g/ar6EatCoIOKAYFZn4UpYeOor26hZXxhIjCWyscGq1IX+NgVPx
d/K+189b7Zt7dy2Bn3kb0kA0n9sqyv37x+T1DiWal/XxFyEpxYbx3gk1X1KFjMKM
Ji+U7Dor5h7c3flW3v5TFP9qBe2414HAI/RZQJpR7I77g+O5/lkb45dGjPJ2oOUc
WL6ixCWa5osU8KxicyVVKq4PMPrOmM9LjLxoHwS72mYaYTe/9q7vdTYcw0VegevJ
VbUPJb9jKygBe0KZvCipyVAeFhBWNZFA/uzFlsSOg4airfRTF5xgVn+nqV75yH9P
07yucTt/TkHs2m04Nc2/j8fmQq25/2lJW11rVTWLrG7hnKrP8UvyuXJ8lV2+fh36
It+/mrD1RowzY/wtchzQ4lc6Wt97Cr//SNHMm60iez7xkCCcm/knqUtxKK9msf/L
e6hOfGfnpd2H+HZAHvfRiSvKKprUA+qxmOL5/bu1M9SYXc6jOwn2HRZrA5uIc1DO
h348ft7PMi8lKVuQpJ96LaioEckzHgODJdcYN44lJZdFQ5AUAsa1dG8glmt10R2a
+jy8tKBs6r0Lt4gERGt+lME2UcJCkgq9DsQMODZ3UiHwU1hPBy6bFQ6ukmjgHsgh
z3/zyHG2jMOyma1vv+hJ1UyWWink/k8hWIQyc++NWWy+NpD05gQmYSL1cT7pz4gn
itfagxavDRaFGaQ4Nif+7r8aVD+h3r0vGu7Gfn4z/ZZw+5+ZxdxoGdo453Jpr2lE
g8E6RcK7S0VuyGQqhlYKggr76KdYDefTOFbaE/US3JBlRMbDwOJNIRdKRiBvus32
XgvxMbKCsHPxrEXjNk0yNSLrY4VgNnTOCH9KxzqrBTdRRhR0IVfbIDN5i+dRjBoY
PKLSQXfLkbfvnE4elFM0Gd4EGbIA1rgAvH1UfWt0Ge4MJGWO2qQj8OE2Cf62wV1z
3f2YrTHrjyBlJekK7FJiSyTe5hQsincL2c95UKC57bS05NKcMZjaD6+CCOtHmg3p
fbu5tIi3ECC4jZ26j/TQtz8R+6mdBowTj75iQr9SBPwUUFokZ/H8DUaj6mHXZYQG
nwnyMz17wGSqcm4C+7J5z3U4Wi73UnC+EijCVmbxNLcjj4YUPdg9UhtxZrL+kZuT
Kjy1hph00Y29en7U14CbIlWW17oKGTFed1Ajz51QvSmPbxn6TcIGaHec5Udf+6iB
1wSGmECEnhgvI4LnSLLWdjyMsgri6rrZ4u99PkvVdFyvrQvROCZynLctTgRrs/Vx
MFF6exhc+Kgp6cLnaVRJEyM27pc9Y81/fw9iW21K89eaboDcT922ItPIrlTEsYxB
Zsx7P/tUAwLXpqATqpqzy84Qu8QXVFqxUDPqWss7AkCJlnXl+4ccEixs+ffHte2P
fGAZaC5DO6n4RveJsaDYxvO7KayPlwUNxammbBTWk3EpVoWaqRDjIYcATft5pHO8
qTOXwgju9K2bAKGalfU1ESJ6/5KRXbA84QPCmg11wx9EINdRGnRpleULg/GsEvTJ
52GAMwvWZABcYuPltByJ3IVZ5cLpPUMqG5cfx06jTQnul+OmjtnciXnU0EO50J6H
chZxZJkfVPU0nBmuR6UjjJk0KAZtrCjfSNATcsoOV6D61D4ohZd5cyQr2MG7jxXV
JkFBJTu0EXVgwd5uz1BLPVBUkyubaoiMlwgumOhD+JLjIETdIN1q73Ywhd52S2mi
0vgSsnv2k88FQ08urFqksvXco/HF68R76vHccRUe8ATz18kUxKpX+Q4GOgnUK5Oo
m5VShusIBxYfzQ+1nrQW/X2Zkx6q2aH+LtE7nsJecZMc4MMIf4cM8EfYYnzMR3A4
bHygJ/PJ7Hc2iq8cMmYDuLM9AJ0NAkvHgqY8Cvjcck+/okX06HlOpO4WBr2C+Lf8
o7eY1eA3fdlD0/4kvKZGwXkZ8577XkOgbcwSHOzju7xsVv4ii9BSGkrXvu6ojYnc
KaqrbPFhLuq8vXIEyOCQL3HsLt1YNCxmYp4l6+YKgSVRh9ly/2MVwA1pw2nhcv+S
RQ2CpK8KGusBPgW+rfu6dT7xTGdKq0eU9XFfQYd3ERt3+jkXv6qaIB/7ztxUT0EX
Ti7qxCcwxcPhKeomqdv/pJ8saATQvFuNyVqQAC2qnLPgd7AXepkcltjofaJPFdDj
UEt9JayB8QpgeZGB/Pat6l+nmR7sRQ4qcsNmMXDXszq/cm43klx6UcyGP6Kj+9Z/
wBQkjrTOH/G+rKFxM8y3jEIrE4mvNg0MoG9KhdglaEzxHH+hWZcbG4k3gDnP66Av
0mE69TkLb2Uh7kVoaekS87w6Wp7NYid3LKOtcXPcwBv3bdk4nURYaUwqHqIFFlM1
vdxBMImSkckNVYc5bzxvYeGpIT93+jfZij8Y/9nS08cD2535bICCyhgIyzUHkbOQ
z5aPq4rlHaSX1EoiWWzy4HRvdfUqZtvBrGpyfyEVX8J9nUZNRLCz8wHPtsB1TUai
0ytL/PucC3JMkLqUQVoiD8Qx5QLlmINCmhAZ7LEzm+SR70NBwt2guMRvymvTFAGJ
UyCkIpvCwUQivxiVaz6ZyOL6JKYskKHY/3jtNpUUByiviqIbf/y9SsbpvH5ffDwR
IVa50gmeysBHrbIpfDoVJgfzkV93qxLchAdgHr2tceOoS6FQbPTyZOl2fRh/xb0a
cll3JJhFHhth6+YYG/NY+0FcOyp0FI9iivGi/VL5lol+NeOP8aqCUUgL6CXzVS3L
w5TVkdZm8PTGIY1qJicU+kANORgLbegVtQe56/6bu3TmfMHe0+WRNPpHT5ei8wNy
JNf0Z2ep8QMqv/Yw0n1Dy0wtAOpyjhyah76GX+oGJsaxttPTP+5xvkIDGqa25j53
rGSrvshWoFK8zAQQvrS2LnnPsFjRhUueothjIryxCQmtfss0AeiyRCxuJsRK87jh
pJv3bO8/yMuNIYaCzN35zE50LlLe5OmA/N/hSPw24YonFMRSVVegqEJaPlBb6Lc1
ZqCCO/jtWDkzUuRhELdBnOcT2ND5/kHP3y6h0EcVyxB9Lr4CxE8ebKUvIimu080M
SzcuaitYkT+PghAGTiSDznQWDHqwQnqySCyP/4clHK9vRM74OScLZKq9Dk9SvwLW
btOlBmGly1VYuJUHfCAkUBow5MRHX1+QhCVsccF/UhEj0mvJaxLq24n2vApI2L89
HOiGl6xhvqcMcWVS+By/zkZjgidBmWDSA7Qd/gn/Z9eHvM6qoH0sUVO1IxVULmdb
02nmugMiO0u0mGgXIyhA1tC/JfVcOSyFJvX0B9Vc8iBZvaKiv4zttHaHZm4zAo7n
ptxcAYmC07Glpi68kMs+Xl5lN2zNtm3GdYGbQjdbZv09lBbNlqoBVLqnclKDhXye
5Qb6uTLKqYgJtXGoZapnSDGeJiQP4AhdLHTkn8AN3+KM4xD3Gt1g8onKbIezgWHS
+CENYS8C3H4DZcoxxBCFFMdmbbRrn0+W1zryC3XnCTYd8D6DoD+0DdEFzeKFo2gF
w9nPcN7ayrRy6sFF6OldqOYbBSceWkgx/B7L8u3KEJOD9nRyDsyWaxb9hcdfkBU6
B7/ctvW+I/80LZW3Ao5iq7i6Wmmo0RaIBtXJTSRr5sOb1PDHTmavEDEa4DU4JeQl
dBcIlghLO9z1mzCe8pvxX2xfL+9S9I0ljyroivPbF0gfIoJhuP+8CHlv9hCQBrzr
Ury0D/KjW+NIg8wBGllhxxMZKKIjCWwEBCsfgrr6AOSRj4FH50SaELOfDWQipAMB
RsAO+sDY7Zc14rmO/uvxT0SmKWBvBUW3/V23NcJDzLURBPdJ8EHhfCWnX8Fsu92j
HWurc68/7sUYcddjRIfMF5ToXLC+C8LJSJvbh6MJDqiEbhWJKNj1AHkDQmpfc3x8
QSofCzX/t9XgtI2GWJZ30mO7WJOz66Ii2oURNnGeHIdPGjwOBBFxFlbK+GMQ1tHI
w8G7xE/R9aolO2r0KOqSHED5ZehtK0uqGeYazsJ+vjmzGFesLiWA/I66P4/Tj9AK
tYiZ/K3bgI3xT/2YLDNHsZEYOWkDWVAUSdziZLBdS5nUrsdusE3EAVTRdNKio8rT
2uUMT9yEoODXRsED4hucPfFswve2yLgr6BIqO6z+AMBiyFNKWb5/1zJhHfnUL4Bs
nHgLxBBZRIDLZ/n57b2PEP3yCPdinE6NLUTsyZHUJkAKf6EJRlULskTT2Y9XuzGv
P7M/zC6g6Cyx4cI6+hpF/Frz4PQOWhPyGUx6XSMrv74O9kqTkeUrfMJxfQFZZ7Se
ATJ1t6hk5s9qEv+OU9hfEU/rOPnXGCCP3Es4VU4GYUF9bEe43DDrLm6y5idKOe6r
q5SaEwHhdo55Ke5HpCIt9BaqMddQMXOFzWsgJhFsNwpL4BryEXt7ZHlEvon96rlt
S8I4C2Jf/vzgYPQQTDzTaczkB6eLJzrJrZzqEotbNesIPog8i1roVe5K0zGLSPrI
wD+qvr9xey8EJSwaV8eIffIi9+lfpbXPEGLz5njiL7y2+B5Q4CB4O3KAhgNVrhY9
Fnv6XCH+jMR8iR34UfapJOwyuliAg9Mbl3m7rLfqKQ++97JjClEQYB816Bq7NlIQ
eNED5BYgK13ANVHmBrh2KLQVfXLzJjdoXM9K2iEtqbDQscewoNcHMKysBmzj9irr
7s5lr2GuhFA4kCw4hWpnF/XSs0FyKxKcRR1+Em8q7FMbVcay7AWtWk52e3WkAC5x
VkCpbJDBesV/wiIKwfDFlEf2r/Y0/S7LLYFG+2xdIiBUpkHd5x4973zzSkYahmhV
j4J8OiyEcwLC0asSEgbDXyOgljZtQiEsXQCWhyO7y22kSA9Qh4tLQYB8ZAa4x8K/
e5Exv3hxDPiB2Dn2FV76D25pucSZhEYqpTa2CruH/05yWAG3xLNh0kGKsijrSkFI
dda8+uMfoljVF9oey5jLxIJUU17Wjol2WyIT2oAD7/YF5vr6IsUDaTyQksOOzd/N
J8aoU7/ED8Ck5s5slLleCH9ERSgGj9X5MhWocG1v8dJ8eD9yv1SMftoGQlsmF8zt
QIHCv6svugYdbPtnYuV/HVMcyOH+qJiXnQqisBhT0UrkCYaL3BoP00BtjhkP6xO9
l/AHRcLxF2b3WkzxUEVKVi7OOpzk6G7CxqffOT0xa7vC6sWr8hag9xwtDCCUR0xn
sr4kEZhVUp8hzmhmfUagWIf4v67FLuD95zT4KWtchti7Dciee24B1x+5+s6/vmUK
8PuTWlWLfjduduCLVM5etgs+rnSrSCQfWGEYqGRwy37CJNfJ4RyQS48SUlyBIOU1
okmmA6vWwRMo196F5bH0qgzo5gr4KpoAxJkP+oDc6T0/TxPelByWWJxnucbv2EXi
vf8CWwUEj0F2NMxjRzwBliu6Eqd1Q84X2UcJO/gpUHfAYJGycolRcTCx6bT5LeCi
ZEIn+AWMXLBVyPtRcVUT/yGA2GPN1zBGNv+MkkoGMqkQI7uwDiX2LF9VifupE3CD
fpy3Uv4o4E7cwOmEZ8UiqWm8l1zWZrwXfyZdKfJQkh7y4oUve+WavsG6+NRScPwK
dPOOcJ+S4SHQq3A+huAojns1XuVqVfq31HEXLgRNTWh/54lxZxbgzvHOftlh/K23
Xy4FmWhuUYczoyAwHkbwt7kWYDWEHPmv9ylVzBtTmUcTe+ejv231pMCFjsSS3Qgr
MNshjJtbjMlacqnJnbvdbsANk5DFg57BVVry/a8EpgyQsrlQsSYFZ8e0Y7LKAMRH
LgAScmR7/GMO9VNTbAVNoN2ISJqhTQtX4blvGI1R471X8dkR7nYlXxOaNE0HWZRC
Z6VMgAVxzAQ2xIZH0e1+qi+ZwrL1sIQuELJI3hNXErEbwPfbvf00Dk/q2RxA5Kc9
IyKaOOG7yfnH7LyHyZ96HsGPHEYrsgWww/ho6RkDHedlU3oYqxPm1JQzO1jnGmv0
ClFugWzkVWZzG+ZkvFWIx3DJZiH48qeWFgMiW95nnh0nFZCSTmPC0GhygFla9sdC
ieyExzAzJBO5VIej7IgZ9OeT7DP5sabj3ZjewGHUpxRa/R1P+RQP1BfqzJXaYk6A
N1YaFzGQjIvCuoWCZoo/XQXWvu+PooD+XguQ4+ss/qApBt/ceT1lLUU9FcJf4CmV
pUVvFz9kCEdLw/NZkTyBkhYmhl2zqgKK5nhGh0OcvjvtKxxkh9bursuMHln4s1T+
adfUGEUMME5UBcN0Ebl/G5jmREQGyS39tZjzOwyZPMnOtl5LkvpCkSn+f3UIFUcq
pr8I00bnnODK61NRNkX5bBwRAFz1Nb+o1I+hhZfxJFuAXo40BMlIT4hy+AgfulQG
dV4VEyiEewCIy+JzHi9ysTIxmn8wWorH91I+KYnCCIhwzOqIGvk7N7HFBeRp7YWP
/iLvqiKIsYyTB2yefoSPgcAUHeivl0FMLpZPghaTs9NeVXcd9bvvMR5Wygi4Df7L
+Ifv81IyXojj6sqHu7hclDfB178s3tpcH4xjbaadmOPhaCo6ibYMWB2SfDRlMRMk
4Cr+XWQjxhXuxnyOrjgFzNjB2eJKWMdrIj1knXzEfUtzOeAC+/XgiDCNxsRUWVhN
K73cT7Kkj607JXJ2XSxbBp7mq6JTwn7bgBKEmRbvbvs+s2I0NEiPoNTHgGegHYoB
D8hSBxRAm+YmDBSm9goTca7tHBPK5Kb5A/5ZodlwHH0BoV8fOavB78iWI6jYhnK5
4WwIHolC1sq7K+AW9MddjEQZrxFgW1ha0MEkVpcKyK/nWtCpWSAMG1eGQPbx5d+O
7MsSyVN+yQXqUfgwgkHp5BU6Wk0xp+Iu8lwKScYnqZ5foMOe1PogNO45TW7qunhg
W4XBNAZwzgnfRUUR8+y3gAHAqpN7i2WXxIJK70dqd+fzUMjq5TQbQnmBeaoauWFB
kkZk37cP5rXiX9WEsUsiYWwPsPSQU4tsZDF9IeG/sFymv9BLhTkph7eyvIJ4W7cL
SP1GZqWRV72iojc48t48HIvc7+NnvTl3zpkYpQJIc2yymXwPSBZyESVuQnCUDcbb
0UK8bnLijSyLpcvFwKj+3EAKXIBL4ABNVx7L2hewbazRRAUCYeKDc+YOrR3sXIIl
6a09UQYy3Au9M7g+K7/tauNggN0XtuLgqj7z//GfJauTiCubQXKeklvWelKjpBde
QyYyE15rGe04S+e5bYxD0JssuQJQOCkLV/9VVUgEr+pC/4iGuz/VNvJly5Inv/Vk
9H7SQ3+TScKchwRJpfA9XiPU9alcJrAbzAa+YiZcafkg+NFng0CFenChR5NaBWRv
oaS5KS+wq54oQSNdpC19T5A2WmlfDKu6N6aWe5PpfaZFWdZzh9GCbYX5CNyiMYpz
HKkWM5UZleGODTzV/MlvVmns9l4jirrPuvN+9m7U76UF7GNCZR44O5M7i+uqHuxg
yIyt0EV/bbpH5ai6e7OqYgHqj76lcmlXaMHWRh2c9Zj6EZpLLGSzdU+wQeewsiPB
NKshy5wYDTXFrXGku7LOAq8oWck42vakJlnJ5NtaEY9v+5Aq4VnIONQvsll25Slp
dOkgQqgypNEkjYhgzyGJjfXuoV2gPp+pROBQ41G0/6L+zqK8d7IduCGzW4HDF+ru
ynbMOI42qrKVpuCBvNMUf1rrRvZHKJstvqcFoGy8AmNR9+VqKGIu/iRQda/MGNhy
/H5mU7APE23K2CtLLGK0vYa2ZUroCkzPR4l1syZi0uoRy5m+6dWD1XFuc1snFowf
PYePMHJRCeKYhS23co2ZHpRYubZ2vfQtTt07zZIc9e19tojxJK4gfET9PAuKs9x5
JSxpUuwO6d23kFMF+c0Ca+XJiBExrSVAqyIzoa3QZ9tIdyqYQvkDNC3AMO+2Rr/x
JIUU2bQ6M+cTtumhDbpibYzGEnDvxyW3yMlfzK+qrztBaN565cfrAN4GSF4onjHm
HmOH6a5woprfcictZtpnaEx7eMBvvMVMir/bF8AP4KJwMP6tBslFrH5kgY/NvUp0
iquOj0u8s9eUR/rZcu7escUlSWRNOkk324qd4fRxwA8e+dKEyh31xOoOXh2IdsZ4
0EmyYJbdDzBU+cG7zxzKInCUgvgR6ckjN9r/B85LnVVCvYQBmfCfpD9/v2QhG4zN
JEU/HHtbASduJbisv3g7ypfVFdQ8auoacFH4B2UqTSFxWtFSzm3RjsI7rhw9JYOM
Wc07sQ/fCyMUy7kXQ85iVMVIe27d8DzdzgUmH3rgCzzPAWp2y1/Yx1p21N+GGl62
9kBHJg7UgKHEbgAO8BzggcY/LffxZUDfOTUpIVfYv2O5uj5aaQP5hshhQaSwZ+sa
Kxf2YoQA7yeeKpjdcYNDPmVAGuGTwCxNVf4yk7fFSNdHVeyKLOnAjdBmUWENjlLG
WDQ38AJeIKrNKW1+MBcCgfs1kircLDEUSW/AsBDbyouDva7SRYZa6QkTTHV+Yar2
b1+6JdrTi+CkfMnjFVApZ4obokELWj2NDw/V8LIZedawZakzgX/sjCtrXG/Jr6D4
CV+ZQPyb+j8H/s37dTFWcUdreTaLpcT/BIJgyu19fv0djRQLkqzkrDGKB86OL/oe
tTlprqOuZXEsO7dNtKyDEszfN3YmgroZNJnQIX0uBCYOsk4+nhv3YpXDlenwuSE0
HYZjPC3lu24Ki28SsV7tnXYV7wTX/jRX1dEDtwHd0/93pzMe9zZSQyFDnUPquUfi
Svwqj38SyFCm2jmrpt/TUcWSadXOFgVhyVgOrME8CiV/F+kABxUtqaB9Cz0bxcWv
XkGQ5TBc0T2cubuQ+8x9AcQhK2UKyEQmFT0/F0kA6fKW+pxTXsaNJWaZU4t1nnV0
hdrpGdrJibIw/CtlQNE+2btiJvxirHI0DYt2ZngGh7kr3b0bdec1bAnfKkg7QPV1
B3EnXW7KIl1Ju9rp22Fdy2Ic+gVQN8991E8S7sZhKpYBfW3vBKi5g728iEB2An9/
KCaVbaCH1+i+pNsdhIdtYR8eRdWpxdiFueJ3hEex1a9h/qtmr9ZdM006Fe5sfrhL
Cef5sC6OelWuq5A06yLb4M7rCSRBgQDmAlViiCpyUzKlU7B3rKOn58Clp/WQtIyn
TnrbuksH/bMx0BeykWS+FzYce+KyBo8k6QwC5iKWGmmmFc387Q1pF0pOj5i94KCT
85DlevRXmidRtF/uSDhNipGT54BrZZHM71e7mVjSNfOkVQ/BPp9H7fZ/xkyXmYAh
huSJfx74KOOGbMo19J65o4/+AlScWOU5j/BQtRuCAGGwp1U2/PLaXJZpO7w2zH0r
Y3NDZ8Uc8CkKIpJ4NmIj127GWc1jTa8xRHZdby/sDHQcRM0c+tIG+45MCpYiaOJa
mrYgX2NGC64N/Rej+WgTN46fJQll2oBMOMXMn2rCCszCMBHgbgKcTRaxM2ZK3QbW
cJM21SWKlynIjAfDJMukW7gx9pFEXFziikExViR0vScwnKyCAb3P/CYEEIohKZBz
WwPlc56Ai0NXoL2Jsrvav11n96Butkmb8pC4xtmHTqInZgGm2IGVGCuFKadRtpJ2
Z1sfC3C7HdO283nh+isHuXVr76ZjAhJmzOutAdXF1NpJ6o1P1pGMopulSzHG9CiC
xSsji2qmaj5DFoXYv7PEAIUahtlOYRf0oTlIHl0ZyYnB/Pw/Abq3HHzEDbYzINH0
EmxDwFpelizFda1qPcrXIaBqXucTKh+MMPEw5VQF2lC5M9LY4NwLbmjp+cxVuTd3
JbsFh8Gz2WsVpqXRoXxDEKw6LRBsmvdEoMtUk+9omu++aTZqzyEPkJDj1HsLt2gM
sXSMJjg3gnvL/YBDOE5Hb2XOSHGtVfVsjtkgP6sKMQks8L1YriyB2xIz+3CxrEq4
tnvU3VKVOZJRHfTjC330G8THtG73yq3df1YouIwSkhdIQVxsdD85PqGZGK5MgeUj
RzvHOiG58rXm57yQAE8jgUOI8ipjfUT3XUOKqDwsruG5q16dM66HdcUs70woCwL/
OlYbqZoAr4CrmfQGZlJp8khM5jPeG6l3TvzEc2RuGgpyXAT3MXQhT3sN/j36dlps
KSLtgE1FqZ7H7f+C/gOOFkpbVbci2jkPcz5MpsaQV6S7BmLHaUk/YKvoODnx6Mde
DyT80Ka+fVudoAvrHPW6ucbZTwFm+YyYyzGHzwbGMqg+1IvGBfjOtc21h4wcvPUS
k1L972X9ZheCs14xu47Yjs9iShsnJpwtbXKcJR7CAwcuStJhqTkdj/vHU/LrZNJ+
TTqMSrmuAXsX1SFY/xABiI7AVCKUn6QFzA3I5kXWJtALwnzyxNhBF6zPcrdOpvZu
4YRaZIE9TEgSKMK1gAA0H956AMZF3xUhQHJll0jxQzCvVajQRh7T27rqAsXT6WRW
CdVHSYxle1ORj6RJB8HDVznRza6EikUrFNvaglEWEVURrhUc+Fz27bfLsiEJNtbl
ej9tWB3MikVp3QH6vfeOJSWDwIU/HO+wk24JNaeSDiR/Ej4AMJPMOTntYtg+AxiH
LTZ8joXmER47admHAxEl4brZEggQjTQIRv0tZfmlWR/B/09QW5aZLTF3v9COW+B2
uZEV7HmnJ1t/YWDP8RXLNdYotodQhyj0KNrfz369MpO/4OaZZPFVuNg2KJMMIRmb
5w72v4XSImjywbel4SSOlQ+YVmjNM4a3FzA9DGoWT0sWqYU0ou88WGQAN3wCdSpS
kD4Ivv+Q0YqpwLN13T1c2SA9l3lD9OkXh5lrWZ7sWZrZu40E5BA5psV9HMXH4Q2J
Bo0XcESL/9XbaobRsPs0hvXaFW8CTC9DKoihjs/4Z8m2uy1OCiabqA8QAhCjUGJQ
4dIhakF4LQ//s97EbBql3nHZuXxqWppWCowA3GJcPGejSsof50dZUADVm9KP9knU
39ogHIb83jn0rQPvzKI0v46HQlu+NuTBw9fJ1efwLdhnjHCQ7IJb0wrBN68VWWRw
I35alb2Z65RPO239F7EBXAs+JEFlNcr5ebTpc/LYKe9AKF1VY8MnYkOOFLfDKoFj
Jbl+AGNBSn3T0TJ43Lrkg++S7Wcu0jJOI/dpsvwRVyqUVcf9bD3/SRSnzxzZiLl5
RES7IzUfN0cmbZg1lA2O87XaBeDJ9Dw/3oypbeEimKz1r47qBM/cLLxsw1LpyKC3
gw0nUtBOIM4A4W9YlMBlU4zrawBBFaJIWGW7HcPtdaGcbIIMqZOI5TlXec3uFjwz
AkTezd3mes9qm0254ZR9bh59V2XlmBU9vorYCI+uHeR29LidgIOrCgh03bqg7yOy
5xAWFFJGlMSbnzzqEkpfm4kv3gsw3FOt3zFApxLKPuO29bxvAMdRUCdK14s0BAnm
IoPW4DX10mqzWq9UdI/NAejnhE3JFvEkGWwxrFCLo1Qa+f5Y9tc5YDwbYG1l674m
gFdgajgXCVIZ8tStrsoU5gOMMbGopcM+/aWjrOjiEK3wgHWDROBbJwuv9xS1urt+
nm/TpeUBIBQxBCkO8N6HnCiRo2DXNBN1T865T8iYOp13hfKNapqqbf+lKTI0S8Ln
hWhxYDpulUpDEasb9JoKSXWLptk7A1VcBFid0dFoNRoq2rHi2/qlrcEL+DCilunx
CrkpVJaRpe+B6TxaS3QjyOVn0EI5ypGe/K2FY7tqfrDUDAPX4w9j/IaUYs/uFTAK
+dpw53qyQbndnlYnLEzRMepc9TwHFADCRKeiJMhphEPAsWRe19sAQtX87PYylzLg
JvCECjY5ol7C0pVAMMR8d8NAH6dYrCRpFx1ItpYIjUNOe8HH1ZCUemPR5RjnO+rh
l74tCVenHrOHRseXUQr9m1MiUb/PfhPGksoz/FNq3OEsgXBzbVmHrf3t+c4n205R
o1oSnHlVxwZlqmRRvgj/Kqo2YvbnUQiubx/LO2jWsgCZPXbszSW/HfIWURQse0TM
ZL44XmKUHXlHnOD0LiR9g3dBUV8xYtdcqSSgGqtXaRDNrGfxkqhSrnMIcrxtWktG
z+TgDWpm12y3uxHsPK0Bh4ySkSlm108k9SXsnvYju/OBJvFnaBLpH0Oox7O6SW6/
18W/1mTEH4Kj+acEpKU10Iufrmp3YaA+GvSvJrefWtoDZcRnHLAZLZB77i55ngAN
rVDkloy4lFUrwOa6uTJc2u9aZRcLy80WW53x5LulTIlfeW4Hkf5qTQsDdZbsgWyg
BaYBSNdOSEjpD/qL2U0wAPlmhV0t88Y34GNJPPVxqaJ38dp6xoVKxkWX9V7Bb6hX
8x3j3xE4FDB5Nb5RhDubUSWKHTUYAkwkX1PMjKB0owxTu7E7YkzbSx7Y9nFDibAO
9EorMfQVH1Az858P1b7Mb1XeL6f6CQIEYZMkVzrtwyHEj3QgVCozssnUKBZSpmHX
QknBUHZ3/vUZHPfbX1kplDcazYsxDm7oQOdEqP8AQtXkzDPS2XSCps5X3AlNCrs4
K5oTzDIPOawy1StwcXTr7HVYAf39sTtr4xgsybqEYuh9jWRJVkptzKAlEvXpJAxG
ZD1TAzyUCiAsePQi2MbLAhXqymQPYbkK2b9UyjA3YNacU37mEfzZAGF91yIeHDto
ObndBqsIL/r2RjuhrGQfOmYfAJ3bVjcpIdZBNsJ0e/KhpcpaJerXOACNt46B70P6
HzgPlA6zKV/Acb1gzjg57j73Sh+OXwt7JKVooweYtKZe/QZisQ3GqxOMwbH5Zeh1
6+RWJ0XKHps9LyT+03JMFxbJwm+JT6u0C2pdpz8hYhQKbaQ7eG36rqubUid6O/aA
mcMlDVL9ftX9Obk4ew2GrsTbewnT7QclsyOK1dV8sGOch983KoZLwaPbANW/0M+6
Xpg5Jce8/KNzMXlaAro7l3nM29AmRyRg+Je87qZsYgPHKFzhccn1vf44xuqgtkVL
d+FQWliYp355lGVB4TVDvgMLRlcD09/v2Wq3QNoudE5zDxC5FVq/JCv/Q1WpBQPS
osnxxma8KqG7WEkVZ/rPs88K0jEuHzIGDdkbV7ujjnqsiCSWASfpKcN6bXbSLQrh
3ZLSKzwcfYTEG20dnUfp884nY8jY8sdLlORP6N2B243AS/5tjnmvPMwQy3bOLV4o
EBh9IRooUElhPiIt2JPyO/5pf7BgBFt/5m4Y61T9WuX/A38Nn0/7//zx12E9bd4U
8QihNq4gravcBGKYxHNQbb4lFHWVezs1g9QfxHOXlo6rXkcqUm9cADkZoFJgXPIr
Fngwt/uhCiXvauPmhb2EXyLdKC/EtIuaplTxYjuKxJ9iFGP+WYAh3Qp00U+9GQT+
cvaJ0fIm3RUWPROqR8iNP8igoP7kCEKfFp1lP49+VIc2aQcmP10irXUAV0jGZfSH
/JBQFVLIVfasPInLTum7oe2OfER0yAsM/rywDaPaQ6mvzFpMA0MAEAtGGeQ5qxkN
MbviA5XQlIMCA2NDkAB4OG8UT4W8aZKcrkj+tvSpM4cus88YlGNPrNechXR+OKa1
cbKauGYjdLyw1U/x1/ZGn0ZAR6KMXl3j0zPirt7lT8I7gxSQT4A5f75XFSzLgxh9
vX1DNlNkJTF2rXPMJOQg4R9QaTPS7UChXXFOzvLonhA4XiDzC2WEWahNJ/ZzCGGt
q/LUc6LHK0ZG35oNRrwCn6Kv9dd6tzr2ka5V60NuYk6UxK8J+sW0ia+QZZXwmNb9
iOriVy7xaM6iFB4WWwWmw4ZGbPIMP1BY1Tw11X9uaC72njHTBiMkzpsSkE12tnTK
wJNzZjoplJ9Z3V/wBnYGwvoYlmgeutnwIx/XQpGCZ9X/Em3u0Q/LBhmxwiIYt1S3
xWm/2AQB8m7ja6T1mi5E4QHlD+rp4n8QTs4xVLgUzm7T6QIrQ8e1oROgzTxYUFqG
8ey8dM4mmHHf3ad2LFDrUPM4bcMJU+cKWBenYFqftb7kZmX4xxeQuH+8vcP5HAqx
ts2X2nbSqLY9B4W3UjfuUMSTD3zqAShgdk5zU2HPZogamVx+aiQxC/N4fiiALS1/
0S4KulQj9dEWtsDAPwjbC2J3kFDBUHo4HNwXmonrLkLCrtjxS0z4fKPiHoBesY/6
XmHT8lappZQmURPgeAnop2ceSZ8Ix4J61cYdo0k21v3w4XZ9PfdwF5J3zNZml8e4
AANQh7ISwnr3tWdhatIveM4FTs0NUlEi/yxI1jqtZ3wYgA3fPCzR9BkHFtr+mzo/
imXu/h6tTQ/Argcse/QWRiOEnD2eNcaaaZpE5dmw9OQTWZvsf3zvQOPx2khH8AEg
QfLaKUE8qTbpEwgTqEZF+xMpOjTFdwGgGTdrK5GhyGenCeGhpIPkSQSBXFqqAcNU
MdswIQWSl01sig9i9CbvAR+QNV3YL4fW79G4dBuEnxcCxs3Ec5XsJNS4qSFvSUsT
QXb+OCQMYNvhY7lql05vsLtbFIaGzcJEmrKf+6ITjRQrAY/gAnSW5pctbpI7m1VD
Lmh8mVt2NY29Nek5b55Bhs+nybOd9dhMudiD37VlB8NMHL1N64pNbC79UNvvLTsO
C5By5deK7aFdGSSvhGs0ZZf/15x5Q2b9prQ3HsLvQa0DAMmW2WanyVdmdZ2eftLd
wIEWmDgcGCWQTtJtgzS5b+viH4gBdnOiSbd7DTtN6OfwvRkJqKcoQC5R86SqJoHL
TfajA3uMQk07gC2YP1py0u4ZtlP9WlOhRScg2lcHejuNuROg8fStZnEBKX4smnp+
uo+x/wPQgm6OYQqajmo2HFJAOtlr9W9wt3SiYkVfTKLAD84GLO5+LjbvEm9XP4oa
naQZkDeacSOGJFmTKm+hZiIfr3ynGrFRpkv2DKVPW/xX8cR43+KjKKqOCap4sHLV
Q1iFnRsf/0r4KvGpLny2rcZinB7tHaX6128IPB+9AruGXcFJ1xX2g229dsg5XQdZ
TzmZPfByWzZVrR+HBS/SZf7rHS6L/K2j+0f/YfUhiQsDrPhdjmFE53upJ2afgl75
Uv5H5FncxqbGGR6yUfP+QsVM6XBZOYnDBOhAXwiCtcfCFYnaY/7opw3LP2YrREz3
FL4/KlHSRshgPjZSFQKCoup5LLyLV8wVPOHtx/tyojzimqHdJgQ3Qb+lr5qxQJ84
AumIMdaU9RfvFgoF4D6D8oBxQlpW1QUfZcAXLRrkQxeVb+BwGMXp0wSkINOxrj5L
aRwVFLs3Fqd65rAz4hGL/qImeC/RVeEE36dVvdXyFy7RNq3w6bq1ENugtPmvxuAC
y96nvP95R52nFvTGR1F3QeQZAp4RUq9NeIe+PEdh4ZQNhJKsvMzhUSDxhOKFxgpH
fsQMGHqxuka9kjtREJkDQEaU6Hddvdo1cYnmhlpp8RHxJxVQ4jFuCqWsVv/JE5BE
6jag0eZpV27hcwYMIsDbF+ZqZ69o4S5x/xHNPQ2tLaVQkVpu74jAVyu9Iu2QJfj8
oG3JkkxcWq1Z5866YfZ4Wx6TTWcyDe3aITaoaIAYWHfw+FWeruC7pBuTiGtGGr1T
x6tG3RnhRLPF5sogKsUqk1fA54DBm7kxf0SNPMynv07JsfQcsof42hXfg29lXzuz
VxEGWkpRep0m2yO9XuJlqy/248lo2V2RRKXKInUmQPexdzPqCnzBKeBxB29/kq2O
Zs1Sa/4uBYIPhUUQTLt3jpI+J9IMmGp50Kt8TL00l1Sa/QE/tGXYpwv10SMypSZM
4/ajY/8Depr1zNlBwUYaWZEUQ4AygrZCWLOCstwLoQs7Kes38zJg9T4MuW21k79M
tlH8teNhvt3FwUolR2vKC2edREGbZtbA/1QDzxckMjmkprsxfLV/dWtJ6s8MnLSi
igwpWLQvRBIGYliY26JMUafeievbjfhAXST3n6AswvtiBMe/qw9gH+TPvF0S1FC8
G8fJb9KvNdX5MNO/9vK+AmKx8NzaBnkzPZZUHT9gfUKCzoqa3Y1YZV8FNwr8Fhfo
wjZPd7INLX/G0aXXcMBF2ZARDXiJ7JwULTjbK1NlMowNrFRgwhXLLL+5gscbruAH
Ow9C2qeeR88ucCjNSP8vkuoMV6K/AmqA1YgbVDbZWQ+S9hSyCJ2M4RLHoS2e71Vj
+EVr35SFsRxiZyVQZrqv+4ja1v1SfiQSMvQSnEuICBH+u6rTvihzaFoML5GPZS/B
IEBPi2ozqCgQEAXs57hWphdhvPv8hX+pNsZiDJN3AkQABOp3o30gLGofxeWx36F4
MHmSF3heRqws5gHn48zG6OWZjPpXPa7Jfcc11plpCcARBD+g0CAkO55iCnQyDJrr
gJ7vGx+6b593xB1tgBHh4oZQHh5rxggWTWV9W0Shi4PqF7WJZwrxAamno5xX03qL
YVYZGjH5kOBh3BZ148fv6ou4BHEev+cAUIex+GJvuWswpzzQtt3o8pjTajxVGGYG
XPTMmVOy5gklKjejtlh0HazG38G4UZ5jK5YGm5ej3uTtl9+J4rFhco1gRPooV1FF
9YRwk3JR/iYJvR83SRjRSl5npLpurSqJ34t0Khvg0AEHbAn6QoxhurW+TDpF/8M4
1fxGhYI7f8cgyBlnprHqPEnXa5zmq9lTxsvxM+e+vOEtwyv2CyzPaMjgaVnYk9kc
E5CKzUzrgzzDoKPGU4jvLEYW/AOGx9dUGo3UPIcm6mr0fEWAhuGyMCQU9h6wR/s0
eBgUWQvnDIPzuaLsKcGaeW4k3FTMjrFy9MyBy858lQwrWow4APCrs5M48628kwbu
8fbfQCE3mkpho7eeNCk5EzsUNwweirJq/gG/PTGNDhImUR8l+1HjRu0nG3dKvMU4
1WNCRHjcb3va862jxdqNnejrZtZBnqq157MbjXMNtL6t9StSaeC27t1X1Cm7KElF
BMw3k0HLNBudHM5PXPh0UbqMAyDzdaDei11BnexQkwzaLe20T64MvMhveBQObnlH
GT6ptqFMmNKKrT09Mkc7hsxFmzvDrj8JbXHelH9WZ6OX355cd91Z9Or5HR0Sea+l
iXMjwb7oIVbyQk7JxtyklUew7VFoZ6OPd0DSQdj+0QKQRxZUZR2Q6tisntOpOuEM
IdJ53Bqh9ZuI5lDY09+BCicrl30TfVoo4nzfX5Bz5K8CG8D49OpQ9rO7d1FJdCrs
hYDLQCbhlN/L6QRG6RC0rNMfgeOrIOwsQCfoGIfDTT+TqX2PTw1IfUjyixeVxzEZ
Yj6TuULnJcHGK5u8evRTkLlYjRyxGmknTv08Jm/v7O9Q5CmhfwOOODi1U5rOkuHR
5wVKyzJO+dXOt4HuYLjlirmdgp1MkEDCVfKBktnJw3pmSxKYr4APujdZvp0vxwX+
s+n2l4ex8HyfSu3JWCwWcIdvy9EgmYS+5ozJ/WZgUJsD3JYzvHZapx6e1AMdEIcR
Af14GE42PCGWrP32ZrBGQzLoIBweazB5xuf/a0+Gjaxsl1LhMgniAlLYf8tcDcLv
ImRkq1YsCqpMkWnfdtA7RYw3R876A12hdqjTAQqWGwLmOoD65vJFIMWSOC9STohz
QU3NZTsCw7AYn6ZQZKRNQ12bTPhQWEHrCHdbLPhRutRvMxL5gZvLje1T2H/ShG/D
xxgCDXRNuVnn2JYEVvq7oOn4XRsVsKHtk9GhfWvd+1taIIdHM4uW2iJpo8m6d1CJ
oxtW0R6EdORU2bH62mS2hLfhUNCKesqgOcK/hLdqnPXGj2oJYNP+QinmryKHkbNa
x8B28wMfIVLGSZfnm5VK+IufzZ05daVrOzTMgns7KXzqnV8p2IwgffQxIa3+LZEm
zv5eMisbO+NUxxTIyC+O26C+wMLgz5hZnXSUjmNYccVkd4gKflC4m1Z/30S2Xndj
/XVssnrPFaOzSjxB6lCcnhbUfVTLwVrQEfXSvrmRkTXMcuXW2PShnGYX61wNGHk2
fuMA2mr0Q0RqY8PgMvngX1glVcUb1MxBezWN3w2nMe75J7IAFUd154zJt/KjgExO
g6fFw5WrlqkuGfjCspdRMBi+h3ARXUbDRSEVvxvT4Qwg9hBK6pT+I+Q63keToV/q
yFBM7SioP+sN4Im7zuxVsoDM1U1H32fwxKisZgvlHGiitVki8110EOWGZywt93Wb
lnlUOAtG65hlvGuApNMtCv2rUGCM5N7R/WWn5v3qc5oDwSsFzUTOgGpwVIUiUrNJ
2MrI/z0CjmcE1rn7BSiCuu9E5Q/AaI6od+GfN2cP22+EdwqQiAemvq4hOijcxRHj
AMp1UjsrUurcqNOapysoGHHMNtI/DMvSi/HPns+C2/NM0fqo2vwOt8l7rx2W33+C
C/QpCF0+uEgcv/sdxLJmrzBF/Kl7mFCJ9IPqXwWl3+G/hc2SY4VIy6021nkmgLgW
4A5TS+LAUeWIilcLOgvv86afzS074tB3r4j6cAaLz6hw6e5PUrUXrqrBPUYVb0Ao
O9mKUyYS1jda6RD5mJhWAl7ND0zKbZeCOGrdUS1q2Or8CDH9LYhLLT38oPwWMGv6
EsJLQbiLXEn6QzVWNEUryrXe4GjBmfQ6vRVZrKnm08cZ3dIQ8VIxmDOCYHtDsu2J
S2lq+YmEzXC8sVMx+hAjCMyCIZdgMY1Dx8ClvjaHwRYx3kTu1fgv8iuWC6k7y87L
5yjK1RTVDDTfqhK9SDWo2CkeCeV3KchjtXGRUgpadrIbbCunc61VV4FhlGJVEoha
c7AObKz0FpgetvTqE2YP7yiVwCRUOx5GyysP4G7KRJqO3gaV/cbrGwKYB4L6nVsC
smqUK+0T6AJhQ1SDCPNpIXe1ixD/KAkjDk6UH+va4Z28lTv2dFNu/HLKodVNg7Cd
79lMPbe+Sp07Z3T9q2kzZD9haP/iz68fLb+ekdScHThnqhciweyAVB9RXgljvBbe
Z0X/osmoLs2c+9sLgYeclpjcqpOAoqsDqky8uK6ES/yDpkQmf6piIweqMHtws14b
4heBXIbf/cwkmNfEfMuAEwqhQ+hLlFy/Msh0NKbiuNc8FQ2+XQFCIt1TkXjcwcMe
CgdG9teu4rRRyGwHQpV1iZSL9tktvc8m+OmOGGPXwNpi9btbAYwwTEQT7UP6AIc4
acrfBJCWnFG9g8rsvwYt/YFSgfx3+afXghbARvLU3mAv4ykQsGx+2iKwoHHA8gg0
byQbSdKwejpDwD4h3Ony3cPySRPfBjUiYF+d1vntIPxniuatlyMcXe59kZv90257
jPmi6nCTTRKM6HntNzVp5+04Hx/4WeH0jGJyOgqmJrB3AYM4UBVO77TDdm/mVSYq
z2DORnv2kjQ12/c+bCKObkKdoFN0Z//CWvRyBRaIqXFGdsf2Tmog4MRmIY4iLSjc
1hRZY1VwPjeigrzKXSnXgETtGV+Mny4gA82ysvQTUorCzM+YOpMBYaKGTMIaxBJc
9uECW3ke/ToXmNerlErLE7gedVhenxJovEr6pJa404N4RWd6bUWH08zU4lhaLGwI
gNheyzXJ+Oqk4FVjBPgs+2Cm/A6LujybckJhJMgk2nlLFv7zBkIyLB6muct2k4kF
AtRPVxf6ap8HnT2ZzwUmGZnQu1suytzTMdSn944C3MFvIZypSAjlG8Rw490xRlXT
oZwgcND8oo/xqkh0tpN6jl1gINJDdYbfnK67jv/OTOni37nohIgVKHFatkppgL6c
R6hdwtFYBOKmhDFypc2pCZXvRwrGuz4SKlZHCUf8DYARmg8+CueYo5BKvMy0b9ZC
4K1JxZpQBbA1SPClOa9ii93guzG7EdIiavcQx5233RFqs29mel8iEaFQqsEs8ljp
8Rc8VBe3YVjvodgDFHmYU00/F4jXYlaTFRTMcqjLYa9MHMFFOsK7zzEeds6e3aPZ
VyeEjjIDZ+8xF1gD3V8OOlUsZAhJmYmUYLFsq10hhJ8W+M2oo82eK6d29noepHAT
g0y0vJtMGdGyI2r5IrgvGACdTYS+uxjwO8w90gcA/uwWNn67L2H+Lo+dfx4tJNbC
u2CE4/v8BUjBF4phAQYoTsgp2f1ablxsqZV6EMIwsjXZGOU12rzMbt2/qzMmj3mR
ue/jj+K+/FRWjp9zY3vFG8dZ8P9N7J+E/2lASdHSn13Uly1JI6MkITpU4TFrjFvv
csTVFMZUEkt+gk0Mn3LODrG58AbFTPiqO9+zi7bomopa0ZG8w+l4c+wwG0ckBWhP
vTXgkeOi+CPdttLJsYdyfUajbY9T/EKqOqQ5R1OGkKDlRio2nLhzwlvIIlXT6fJB
ARLsHwzudZ554/oS7mpuKI4QiV0pHXG/ozCcGOC48BlbNd9HNoQcF05CWY6gfJXn
NMJYMTl8IMY36Rw4NCGEsS5yp7cvNOV5Lr9HinWr4CqQRTePkOB6lVqA/+WbJ+m7
JnCt8vJU4I0Y53J/n8JIaOSegzBla+irg6p2lcciqDRL5EQcKiru4OmcFle0ZC7t
IjSU2JvyKnJYn6EnqouaYyBd16TsDqivme7+0fy8klpEr74aW/4bs7L/3i6uLCal
UecuUNojzVnrIOjkrhGeLjfRtXfR6IMUsgUaa76hjzu4ZXFNkoNCfZE3zO7MycMU
SpDyWgozSWJS/wpYaoeVRo7GOIDKuArqsv8CmSBkGB9AH3tnLoYcW59xdLZRK9Ke
LOp/TjbuH+bgCF6Kyn+ZEGNwLYxaPb/SS5KyEuVKBalBquauc9UqxDewln9Yi0FN
djJWyFgH1dNNd8sy3RD9ztF7wbGgomvnr4316B+RXl6xOoWePW4iofzdk1IzI7p8
YjQ1IJzMy1M5WrrLAT1yst03B8ohWQ444dWuBOY4T0wKSwd9BfvWmYzJv8j9AX9g
/Chsvy6kS6m5oHd0z6QFQqicQhPgqlC+OGMjBTJz5ZSwEa2tfNho9cWwXnQWc8hw
fR0kUd+l8BhgmRTH0oMVOC69NxzBzdN5ezSXhmVyFRCy1vUaVZTUS/OUb0V99a1X
/hEX8lpwC8iobrjpGJP7QB9zQbbLewRqdyhMQsO2tmCRuew8DfnkOJKCx5uX4gZu
IeZN2ZpeG7bbWggMaEoYoY1m1sAB3z0ghEFQU4A/YG6LolxYOfJ+iSBfcUkHhc4e
lyYJiUKcughulbLTy6ukJjJ/nZ2pUT7snxTVZpnaup86QjuQXwrT7U2IXYPleKDH
2iNoih1/QmauH631iSpp+uDfxp7PCxMBihV2YpNE+0whlHxoeI/BdniqG9QB/VWR
GDvekmFSFAJfT+xK6LZnKTZvmNwf163XK7xOR4D89/8Mg9iwJZm1Qlmhbs8ye+cx
rtBus5aLhEamnZZbpvxJPnWjWiQP2ZBTZJwTDoqlqH+SuXf7ZFF+uJCzgE/63W1A
uOW1zKXiUrlo/da4Hx8I6UIj+X/jNMnaCKZzgbZJA3ZWk++48HEb5nZwyv4N0UpG
81YzL1UQvNTn8IZxkJiuOAcy2B8ZmQrmxsQli/a33NXqA6iJh+NKnvabDyLX5oK8
ft9uKwL/Q56Nec7JYsUMzzn+iQtpdEKukTqC3rGytNHIOvtqjZaCuPgCK9+tu5KH
Y5B++Cox8Ny9yXUxPsjBTd7ssCCYAtq5vk984Ajco2o9Wlid4kNRlw+fxydeUJsf
3lnsQw2FNVjkxz195Ud4ZKZy+LOmmynwb8H5+eLqpli5ZCudmmAtztHlqgo95/3D
5G751d/qGUa7DAHkhWFez/sR+oKRGtdssbZgc+CdRDMOxryDzCGpkUc66EbZ9wtC
OudfifxgxBCgld89gR9COY//F6+imcUO4xLKxYZoTbKK/uUm5N9PH4xTWaYSaR86
JKxi9Du0DIp+VXjCsByQPqDXSx/rDFlw4+wrYZXFE2ASK2SdPs23qg0QITB9otW0
IpGxEut8CRQ5Msw1l0g3YPh9ofRZ06X+QAdg0PLXJgCSLgKE7a0NOi+9y3FhPUlB
NFPYuVv6L9dsJ3TFa6ASV4AyqOeR8Osaqzod3WlL/HW9dPRFjVdkwBRq3uVM5qJG
ccyuYt8dPIKjjKbysOSpZM7C+e0ujFc6m5cU1oBx3RDPf//p6Imi9lpCIabk/k5x
pDXpSMKga1OhOyHQzAor++uDo6xPHjh3SZ+Rg+Sy6f5f0eKm1GrpSTjDqSDIhHwF
KJUuV/pVaJXTNHV/jPnsFKzojevqf1QSzlw486Qr1UgHIvLh7tXaOupl9DW+nZuB
RNCH2lNtXKjj3HRkU+mJ4MvEBABHQ31rTnzjNJE2/7IcfCPqPgxAi88Iq1O1fT1u
Ow9Ws4t2jydhjN3FjF4/NRFxSr9Q88IYZTgCOZ2jJwHbDcKowt4wcPizrpJv6r4K
Bar7NVdmVxxHJrOKJJ8GKZIdJyVdngt+xP2vzynktFmar0lwD44aFYOxq3GVFXsS
X1qc/nrGfATdOwsXKa8t70VrqddrQGhEJPv1iyVHL1YfZUJ+egSE81RosFR37WSB
YxFhlY4egndQVqLz/1+rYZoptJNzRaQxhotZuFvpV5OrkZ5k/tGl16JrAXAZLMuW
UHzQgR0cucubyh7xEx3hsHR6vCLAcLP3slcCFoEDcwhFp9AJCZ44gKtTt+5awg7E
5NgdQ20vkPHgrue/FkpTqbVXNaD6MeBwjjd+7fh4ebIMj1vpiRXr4jgEEEOY69mg
PzrEllAp9/7sdxqOSeoxK/reDKU2zLzok2EwuOAhrJGDRdhc5TXMt8KTaMFFN3Kg
sew6mo6hneMFuvbKpCr+a5FSVZQsjuUBuh+DsVPQssjrrkUY0PEdK7j2gINFWSES
tuzK/07xhII4ge8mu1dhQIG0EkJKROkGOBxv1p+NYo2JQ2u30hEHxpSlLzbLutAf
iwAgee/l65s3UWAfSSLAUj9ow7GkPMEAz8Vae5RC8eQgnqTSekNihe7hMFU+/XYy
lW9uK37CF2g/ttuYq/INxLiI5vaRTc8B61Dy+6AyyFQXmhblvX05yJCzIpf1c3Te
rTwUHJAgdudSQVxe2igb6173x7YOiwjVhKzaEZ7g4xXO8ZWCMHO6n/Xs/FzwfVvd
DHCSFCCOuM05e/yl7HgqKQMdMHcPE5TdhAFkAjydPqt7p3aJQFcfc9PE+4mHp/Hv
7+4+orM0WpgdBnKtDfVcPRISwCySDX1doXeo0Odmy7T9g07O0P7lEdMbDVcGtjip
WNQhoKIfZLZIhPbRZKnfVonxolgC/pTwrxEQNP3edhJ5nDkoDMrP/oELwyM6nDWP
Bb+gE1Jhb6CWLc9wXAwprN6rmZeZLKGhEg5Kt43kgtozyRnT1Qaus9YBJSBjH2Rf
+LtyuLffxf97Yz8YCqB8todnL1NhV8RXTBfAf6KT/2SNgj/3etEcUweXZ/9mCJCU
yiRkC57etc0c1o8lWV5/xDL1fBx7NSXaUrwn7V8+lk266lZ6e8oVYtEq/9XZMIof
q+MD1OX6Zot9T6pda9Tgc8vJq2dRcOgxzyCjK2H1KeXX2lVfyy/ZJI0QTnT6eojy
rfVRhfbEjAXUw1EtCPwrjPLL33d/ng5MI3wrcNY6XpXSADUMZHJeDrPFFJFlfiAS
PIdPtusBxeLv/MpnrChANPdq/7RegZFX1BoLeUy8E7qtJYfCUHGeyApK9CJtu1mf
O/WHWWZbG7As9HieUu6A2Lw8Ebo6B6XUnewyUtYhrxNvIzkwUrmv21nv2rvYUHex
9SThLU9A/7gQ+vs9GDELItsi6WSUqugCInHjhmKTgwkiJRpGKn7/6x47U3fuBJ7K
VAF4PIn09xYdGHwkK0Il64YbZlE1Ya3GQ8ZNiN4OROLnkcHLWwtC1zxOD1CPjjxC
J3hKK3tWzJhto4s73+MNEvaFJTw7XyfUyt9fiPxAuahZdGTSczv7/GjXIth+Edxd
UwoRyeV4NobkePQ0EsQYeZBCHui50XprLCTT3JOemAfJlVEePCINsXWvIVMfIGZU
GPcDTvjl7r50s/IAXMlkyB6m/P70R5xKp5H57DO/OZ3QSyZBGws1bq9tcVi8ikSF
9HmLCMwFLoj415RXqJk0HDlObxoGtV8hK3JWUD1bYOn8473mLO8cfZyNeliiqrve
Yc7HLQxUWwp4r01fZ83p1D+EPQCNedp/6mLsRY20Mp26NO6IuNpD2yUMyirfT6Na
px2mhb9Izc0EWx88NzxZJ/78Z+ENSGe92MPFOZjZ6Os74SyvljL8UD7Pd4NPAmzA
78SoxtJXt5161/oDR8/ZQBXTdoFQUgQ+qNHE6ezMeQ9B1KdIJ1V84V3opnnT1oHM
PW7pWLLs1c7ZjctyBKQQ2UZAKu8n0NjCU/5aBLBkhwidqfLkh6r3PsgMI/iowr2b
+O+zHXa2Yj1IAa8LL3CZWok6YHPq/nmxssLzz8S/RfiZf+nJEC04FtdOdoplvQca
OsYreQbnD03M2gZTMC/wzElhPn8Z6uLdHdR56x0KEzoR7DW65dXJ8ABTPHDM6wak
+WiHEIQ80ALl1M0lWxKZauuoZ0dnOK2q/RVT53kFRPuJ3cErri5oi7bO5RcK8wGV
a1tF5VXQ5ZsyyAIRhJ2j7mbglb7HAllVftaj0sHCKis2vqcEz/OTLqOuA09SM3Or
q0kjagWOS1MCuTHViu9LhbhUsLffzZCv/5YclxQpObGtpSmi2P5kMB8Y6tn7Q0GU
LMHgKwU2+Y3PAv0eNmvexFqUrLJQ8s2yWZDJI7dZAq0T2q22xhkBb22/Y+bnZAcN
McAM1Mj8sas68w9erhpx3l742jFZGbhXkxR5VwA9Fuf5a/btDf9fagZvO96CAAv3
JDoicsi7pNSj9qb9k2qjon0EeP/E87I9CJ2aJ40nXCPuJBhiLaAAtsL2+8m14+AY
vXAhP1agTry+IeiukR13GKijD0aoKE/craqPiPOdDWoSnBVyw/RBcMo+oQLmUyUH
sFqnlS3dayyjAx4PQcgAIpYSuq5hMY87bR9H/M6oMzlVh2Acpm9LJP4EqjLH8HIm
YiU4hA/yddCfd87rBEZurh1gGAG5icqfxzERcBEMt82D8S8i0skBKHwvZtZUIJyI
zGKD3xrySozcY+EP7brx1eE0N4rMcY0xgO8iGkc3x4/dQX+foK+PczrLLLQWBLjg
i6YPSvQl+acHUgMHcR87ZxkYBvhlO19QHgExDvBkC/0UNumxfRX5c+fbE/BGIFns
4W1StP9atq5P1bzQPSYwWbFT6Yztn/CWAVHtN2l3lRa+eE/wshdjaodQ8csqI4Tq
KNzGpGEvdOx1aqHLn5CGOsKgvgNM0q5q/SspgvyEwLTHFq0cOcHdVMqtkQVQuh/2
qLW71gdv/PZ5919Mj8lSk9QiBS5Up69uBR5sdlNKoIpsiwxqGK+4paCYYnEpslFq
5J5aT5w+KUjtQaZ8gqeuuWCv1YriaxIWrDpxdt3gi6Y5Jk+x28nEUv0uMYcvfbho
v5twdy6huBq63MZDgeFLirL6g40WRDkFgMFMpjjKRNN6tqExskfT9FyjAqueWoBc
mQ7yPcM90az71O/9sVZjvjHqcAFd65KanOdIHpbM1DgGFAJQCbsc7dHqjC03Ee79
l7YwG2CVIGum6qlsg32nEKxhk+3WUHkKrV4uwNWOd/301PkKmyOOUhH/VlWpE06b
haoKA/FOdnZwHJEYG3tNf6YJ9pRmfMH8PO6rjcU/myBWLP+ugaMap8gdgwqwsll/
xhLWkHtm7lxhGTQ6zoKfXUAVqSUgtuGQS9WVKwUv534fPh5cE3PHS79uvh8S8Vsc
zWkqT9huXjUnJUOLtRQP9uBSwYxamQ+MyaY4yDEXAtKlVmRIH4P20NrFBmz8U2sl
+rqws6v2xZXdIpv5TRfzWbkEVg9T5nnRv29NTlf5wjhl9RDD8ZWktquRDgfMGWE7
UxQpvBoxPPsyA+tDx0cqpntshN9gjlscNVubhEGsE1SS4Hm+Fl/YrXt/Wa6vRz1l
DG6/bSdKg8Icbh987E8macbcnNU+DovDZKwRBCO5uYkJnR1Johjr5QfJ9xkLXLBF
p5Eou3iDar2hts50UPF+GLC8/E6nGDXl2xa/cBK1+WgcQEFRYFdlWbEioXJRRe6m
YS03zSFZuxssgew9nOF7kbg78q2vGD6yP5l3P3jHoxCaoC+IPGM7i6156SXcW2Rz
bPXtZVtvNr/b0lOPONd8jaXt5yX4E8oTaAn+cX5p40wRkFkaiXygczBSEjtEpRw6
cY8RWCZftSeEYAXDh6nq+of+9iNzXc8UkLoMFpUXqopiwkpey5OJhL/XtkNeO4AK
szfaIS3KoKJYldcnXHO/4HjBa19Zu3gYlGS667QDf3ZNw7tH2Hhx6vhRKJDciZXf
6ocONGnwidstvAuBK0A/GpvOS0DCV2fpONNOp8fc7VHZty59dw/tjQ/Zd6sG27qC
rOsG29B1c9vWvVTMjvfmzt4XsKRF7h1RDFv2+X1bZFd1hqiSM9YMmCppa3eOLFew
4hNHm6/inH9dXq/zW9U0NrQ/+bJ/WpGNAHv/EwVWqrK4lbU7XWv9b3auh8nZErFS
E2MKiv/HC4T/aAicnfy8G1xn+Sa9FM9BfQplMmROHWt23Nv2T+zF2sirjRelVPqK
p435cWWLDYwTmgu0oNt89C/WJ5QCC5M3eK7tm04OCJgZFXr22nkFqK6QKPUIn8j5
XDpg/KzdcF5azIz6Vzf3UX5ONv+ArBWE+XcKRefGDIHVjiWlGncEJ8FqNGIYzpfu
qPjw9ggT7S0l+TB9sEr8sMoMg49iF6zArSjedUfZjY+zQFP15fihjhf76dJJyDBw
sOBKI2r3F9CHUYTW2YlveceDzNseGsBFMZDYaPBfpdLzwZzPHN5+B8f92vCpSMst
OJZuFosbmOvL7EQsGqjr1nPDjKVvhFX55HPWAb+rD4X+Mzt84lnp10Qb+GnGOYcJ
cMNeYCghDSeDwmJCAOo33GJxty3/3oi/vUxIiiPq/BcWxC8Vh0Mw2x95PTgC32LW
hPrc3Q6v2ndvuA4lJHtoi6b8UMZ/BXJQP8uYzwkSsqq1r7Lj0bm5IcVJeIyYRN14
yyLyme5lGh8pnRO3SJPY7bzDTFbGaotSGCbOCPk64ua1TD6hZFgzUsrKTBGxdX4d
ffPQ5bihPvXzDPN//GHLgpW/jGJG0XNjwrJR1eXu7wdt/pjsHuaCOMc41s1kExb7
ZJlMIo9EWiG+oQz1E28Mxy8PzChvkH9cQZIkCSp2WZdkmotRVf5CHRNlpI4Nn/43
MOmrAqh2So4X3MsWgkYFdqitbyHnJIZazR206N/iKFSIaniC0c8TU+rN6um/8VUz
8arEXYlnMA6L2swd8jCSkGPB5Z0Gqngxg1HB6LmXiLC4Fb32ylrcwJkRwEvJzZ/x
pi8YAFKZXy3G7mlChx1Vc0dewoHXIgcBUNPIluKathvmtNAusp6WDbJRACTdGqK+
HwPn4lRVaT/aACTDbjvoyvYQlt4rCJMiAnI1EjY5P0kE1bR2UrXK8PAx2vtQoDBl
ecloxFEZlOOMqmF1/PQvc/EZxfhEL8h6b6WGw/lAEvxLGjJAUnNJG8170Vf8pVv1
IJz7AZO6vUxzE+Ot2U5Qe/XX1vs3ej7+Zm7e7crGq+Didkz6RqKaJbMmx2BxZBaZ
fYMahRI2ypsCEqENot3uzKuxVGCwuzCVxtgCn+NIIg9q4I5pKQVagj8XEH/7/r2z
Qg4jK4UY5NB9DAHqtvErkWMY1cXXFpsoxugGNXI0TAUSI7UojHq0V8YyAfudOJzK
uhf5oRe0tfrjHg1AOI304h24Mm/SP73ukOgHnLkfUMVyH26PmLcIeBFueQ9LWYCe
B8+5VkjUHKOAIjrN5q/mEXdC9BcSUf4Py5fZmijFSZyr5423eTifiw6V5JTjDCsl
D71lFLYEtOuxbFW/siyIAc/sTi1liVxWSuGCufrrU1zsSiKaB2P7zaKfQoJIUYhP
ruh7hbO0jmdvD9SwAKXS2VNEjntmxw4Mu05MmW+L9h5T6W+1RJmIunZPykBpDP4B
hqzYelf7MyhWCsfTmwBK5czt+NNVWP3xa7pTOx3Yc1tNafJHJjgzly415Z/qD82s
l4SJ73rxTQvorBsKNaqnT/JfX9iseNzNPxAnZo1LlgS04/11Odx8owHkzNljA8aV
y0GDdNA63K1ZxXB5OHG6ZMsuxTupW2X+uKbyG+LStOPXUCqG9i589v3/qGOA9eeG
7m7n5VG704g0KN/tt2aMzXhjFSYJ7O13MNBlmF7QPpD+FNX/6YlAF/14burFQiot
apGK97dkOMxi/utvKB2qmEuqJrsSTE3+/ETX5khEuiRHZhJLUK951GvIiqiTFKeI
+FyPIpVPIB7aAgCsdJCJCYH9CpKDbahqjXPSfF8J1ncNDAUikz6bO5siOLtXqfUe
jls/zvZEHLCMsqRmdMMAT8w4QFhqTCeuJR/Vdjk6X6VtAVvbV8CZO+ovFQ6uwSsc
pB8LprrWIFEBGyOp1vKsL7y8+BWCQetmAocaNUjAcqwK5VBeGKGEF2l5EFs7Q4Z3
daVibW2dQvG4gIlMEpazFUbs9vIPAc39HUIP+nkgLtFwSmPBOyAkcUCWW1mNL0KG
3VfsUI1HmA7i7zX7FyN6WG+px2kGezIWmcoLU/K4Kx5YNuk+9IR4v7UP21r7FZeI
ZjCNTEuZgHXSOVbvRmVdUYdfQaTlTNBR3PDxBQbfEZGPMs5ZCcS2MC030YC0pmcx
2q8U+pECFS2G4M6vu7Kc3WAgFnP+MsVe1turVyI3tJeOUiZVcaUVTXrAsd63AZeP
WslrPNvSKsohJ87WCFXtnnL4tIKE6880rIOrJHFYC6dFUH7S0OJYqxEgcgj3NVH+
PX4FroB+0PbSWX1QjevGrd1Y2SwJ4z7MkrGI/KOj2qPtsQk9ZMDyctQZFiGdibL8
ajDR8wJHPl3tkrWPPKhbFWksTEnXXmEkR+ZzWpbxt3Cv4A+hBNZ2gN88L+uIPhHJ
6GoMn7NNjZUOOfRohiksZA/cOzRFhT2LUxtj2sSvDQagKtaf/z+pQUgvJdE2c2e1
z6FVvYJ+BYncm0AJEKbWIFvY1UyorLe7Lkk5RvDvQaQuZpbWSEafzJcrcEMXSR6v
Fl0QmNrhD/R/Q9NOxdWF8O28HwizyAlK/m8M3PctFW1+dKvejUssH0vZHnsrAgSz
D6WXMBsN+Nh9TG8VvLFj5eI9mYk6NemW8OuE+LHww9S6VsjOlu9uhdZxA7C8UepG
xwBT+O/1w2Yrg6XV563bysGT1EjlWGeX9XbE25UIezBwRIjEEZAOMOcTX2TtQlXs
bm0rachqjTpUyGapntkpiXrPcGWuKea8v11cqDZm2QfjcFHU8chTSCwAlYMuibaz
vxEgQGbMqDcV54wozxBd7mEVG1xSyDdg5D8x6RmS9g5lkvLAzicBqy/5TDM+i+al
4nJU7n+AGtR0O8n6PRybCzOukSzBnJJRya/xP+djIT+OCcaXYWVF5qPRnnuvTtzv
oMjXW3z0jzQe5ryCLJKj9H2kMLgwRZR2p/2AZKw/wb212ls+X8aB0A3HeyLsv3FI
2+E2KLtq34ISAz8N+fI2xQNzjfrgBbyFfhTlC/s7BtPVEllwTw3J2cg5BUkpGH4v
jWkZ8gbSsgpCZ4mlxV9g39grXyBnSYOIhFf+mYLL0lXbnNzGztMkBe+nMngQCg/L
VOaG2UGNb1b3oot7OGuR/rL80gUUc4Y+b/YnjqX6t2UbndPSvbxuxrYo9BJPZRpX
WjjT8fPjtJ2fMJRMRExCsRWx/+lJnFCO8Gk54rIaURBwrTp8ktpWNePNeVK4MijM
czyg4bBHWqFjP5j8Vaq4mtBfivLpSA4k5+bn3Y7komXqD0hcspT98TQ8a8jYEB71
a/7PuQOixtIU0l4pvTGBcqzDYREuLo97faum2wVsi7ciOmyY1tDsgKRIJhER32AX
wcz+iE3eKZvAi4SQC0jChEQqn5qAiUGi68a4aouWG27ONcayLd4ma9Z+4zLhwJQ0
RFUt8E6OvTNMxQ2eFj/xK/xO2kKCpQuUbeRcO+G8gU1m3l3onPLYf+VPc8YTUU+Z
0MXodp/OUwo6i0aRbw52IqafvQVx5gp+LUsrmsPDdhC/8Y3pKkeBLxU7Ddl5drUk
CxlNx+eAbh+xffox2VjzVHjGGypr/pTyuJTsVRxQorl0II6zbAfjCT6bIMEm7vnp
xbM2+6DpO+yxjzxhWR2SZ3Yb31CAwBiDOUUyjStUIupgCS4KkosYqEt259PWu6aQ
pTWnDyB6cFwBeU9beUg2jXx0HCQI3uOxtgk42Bc6DTQuJEHsoW6gQjROGtLDIEUz
xLPyYsX4/OTOwtynqKl2WU5zEWNMtGk50Zrfefw/X8ckYre30VZS0jtwtmT+S5kN
vdl58KXzGCF6fdMr554MJ3AHRPEqermCDM5eitrCpGmm9fZ9HVgoS0BLQxv/ULRS
K5hG0Vhr6/hpYHIvWSgZHfkcfmiEWsOAQWjt+5MiNrMLmE7jL++q67+Md+9y/3JO
WpAyrkafQj5ttm50j+BxZ6Wjr67RYhleSiebo243BT/gWExpoZAVMDtVVb9Tq08u
CurKn6KACB3vhjG2Dz7EkZLOxGxVZLBDA/bluniJYyu3ZGNcHh5A72Dc3FcPONu7
oq3ceWLIobQCZl1tLf1Cjex4/6hzvw9Bcy+584onFb0ztR2tP6munTM4mR4MndOo
42nsOAmsXpKac64OCevIm4vBYACA6+9IumLms43JKkdaOtoB8lzdQ6uXiogQ4seB
5ws1/LETG9JDcnA2QhV6JlLyHjyraq47gp0lGD1YrnwpsvuhYY4BgYfsZI4Ae6Xu
mU0EnAUK303BKSRUcnytVhYm6po62/psc4JzruZWsTRKWAiqHRs5C3X24/LHtLW4
Af2u8O9yc/fHV2b5/Lb3CYdkQBXk7jP3xnh9hkcLY3iVtsUPT1TZAZFjjOYljec7
t7Qrkeg8TDYHcTeIwUc73ft9f78SkNjWnb4BylZMdsXeXgRw/9cGlTlIXa7Qy86T
33YT9gegt2h1CDl5KPj8a3aLjeacJR+DyPd/LU/ur/JnXPEllpcR25lb7QzYptKc
bMLgrIg74AUUFHe8iMwePDCUtMoeVnhNW42tYPv8+3cwDJpYJeW90QlnfINkGWPO
lyN0n12uD9mId3FVk23mROMNscUhJDkPCwpVDVng8ffZLeiACRBYSQg8Yez2qqxU
AxboEQgSeq+TchUtzJ4H+w3qStmEUPiNTHB90jo1tTRbx1t8ZGZ848OLmyYTaKMy
lErYHpU0i/oZppjjbY40SG/kiSh/HRL4CQ5yQ9gwoqx9oJXZfyBbT3kIiY3K1gDz
j4Svmrb3DUclWFcZ1Wz1l4nZeq5JpWoZrFQJ6DDRjemVGAJwjZWWOnIj287pEqUF
Lr5fe5tC+qoGtcPMkYLvYmAd0xALvE7lxoab9/ZapWLzC4zJ4wlwMywfmdGjG5fE
aYMdCKPA+YX30v0dZR/FoFivw9tBgGOrTFNv+KO4609Cy2/K8bqtj6iDvCTw94dG
rvZ3Vm0nmoWcLpvzONDYBfvxNB4xyahn9H4yZdnci32TqRwGVT6vjKg0JoG359r5
/TUpsMTGv9qdcWHT7OzaYti743bMIc4VWaS1Az87v7RwZpwakbaEJVxohlZUn5df
zxFaPp/Xm0VMbSdRFy6z1McaITFkF6tdBVQ4sqQDckN/EPoyOxj+WuMsWN40SRnh
JkRbBor3XKJl1E8OZ6uMflLqykb2j/5w8oPRuzU8NJYEeXFXiZD3DWBzw+aGUXIb
q2AUp9M3JJafF6PkIzj+oCtjsBJh1ABfnAO4lce1GP1F1ShgW2toStofh2obdxVT
jObZ+kIWRp30Xg09G2k0neYMD/cWA+kEPqXzb121pGfO6bWXHBJeqhsaGU8F24rL
MybbrXC6Zf1ObU1wBMgZKa31hGd3d4uwAdfejrVDI/nvSGP+THejVwCfAqTXYho2
J9jGZTUtFopN3ts3J4n3quQmpprj8OPzRmsjf+uVti9QdhXFRT84SPlZQ5Vaf1sk
B8RB3WMw9xkYxRKSdn1ZaLaShdT1HRRgAIkdQtZPxoG6Q7sDbV1fUGFlw0PROJbV
kkM0MOWPEdhaMxmaH/p6L/pWn6YVsdqUQvffuzNlxsmJPw/Wn2jJR4Af4wWV3Lo6
D+Kwho5sKpTsv9BNlkgACbmhcVDvygz91uX2O3MPnOwKGuLtxS7m4nZZ5ypk6gAv
p9Fo5exaARc1c63NH6UMJjM0owQx1JZ0NB52R4BY5+OXfc5PJNe15Hm0cg+Mza6d
8gLDtGDU2CYyHSH03spXuHlzwD3HqZ0fLmRtM+7YWGdnoDDzdLirBKqmBiFFKcVz
e8WjXjYlJa91cYvLIRFfpjQAlddrIdEm5U7FYRAxsHBHVFmEc1OD+pYtDVfoc3b6
y2JVz5wazU40GiGds4C67BHaICv0sFwmc2umXs18QNVDE9TXoYAhUoym68poFg0v
bPLYWqrNFdkPt0nfeFc85og1baAz4vKfJk4j/yEdSWM/01W111AxzwSqq4DR+rcx
ahftGTWprPtq93B+nAZ8yrwWriAtiZeu36WegeJC98qsOmygoJuuVLMRqNwqAa6d
WZfKXDJppU6uJihic0jt5eUTozjbOPu2NJF8zTzohI0fvipxYOhz+UHmbAA+8Tno
Skt7i4GemsKA/kFpJ5RIKOMCMCxgbZ3QNWMl+rY6u/HgMZOLiAsZNb3oao3c2Q4a
yP44XmJ2UbhG5PmwT9KTcvU7A0WPu7AznPbhN9+orSinEWSuMB4PlGQ0Yzjb/73s
I3HTAhhpgiZ+f1k+Khg7AWXFA8v5w3J4ZJ+PKz+bPRs3QLea584N/0Si8KttCO3f
AlGwxIjg6gmCJ/OJsaPifDbnqUvaMwUQJmAUVECyh72CvBlsdRPgREkNXYiM0sR2
NtKaBOlHFU0828XNUUAqWcwEPTnrrXCqx81Uot5CgP4Io3qbswmFgzH5jx4tc34M
/Yty7CWDG/KaO/9C+Osq8Bnx7Gg9rI7r4ofkQbmnNvD/VqUekW6u83aD3ygNradq
g90Awr47HDfrjNYHPHV49r7rAdLwaM8AW1lLIEcUMqX7RIXBYUQ+4uGX0ow4BJaF
N6VmkPyVhwDFFxdjDpxnQ8bMdMK4Xk0AJenJTwo9d9Dslgq3GoBor6gIEwisEbEd
IQAS73VO6vChPFq02y3/pJ2aar6IPtUElxr5LPPYgc8h1z4bhPF12JM9wElgsBHR
o+Zd70bL/sD0JaPWqWo57s7RdHsxwPTGrVXWHMvS1Zw9EYp/N8wdjBdZPZf5D9Hy
P3I2zSeV6B7JbFczBxmdD8Jo6z4Ak6e0Z4486Cd92HJ+VXcMaBOL06BEpZNmfSGU
H9Ukqto8N0k7XnhBawqlxD1uxRX8QyHTbok1W0WOOAZsREpbVtmG0ChzewRfIpD3
t5DmHnzRrF8xFPf6Nj82zeHQjLVVad3zUkOsAlYDbELvHT5FCfeKzoDVsYlRff5z
L7ouhrBLHuyIvnGocHpYMipeFrIoCg5aQB1ou2uNeYNbFgDh8XBDl4dUo1x8815Z
LoIXGQzWQBK4uPA4vFlu3Z9MCKhijzA7NAUhsRvzg7acH1nzYUGbhLNsN/XmdGDF
4hvwMp2n7MMYQ+FrWteaCWNa8is48HbEQILcO4B4PLztEf4XvbO9okw8VzZGScAn
LICksty2YdRAr5GAnbMCSOUfCk65zOr5kJSnBEcKfmkRr62QDe2kIIhkUE4naptG
irhhH6/HwAHuvbz2SXfm0qhEXPOtxyH1g3q/VgvzeiUb/mCWY3R6I4ahXFNzQyvl
WDj0hbJj/Ddiqe8igGX6hOvLG3SISaTlB8rlcS0UFFu1c9R4OWd0D95mDqDdkeeW
aSVdhhWbFnMEozkbDelEbEiRQMmYauqL6J++5Isbc3lOxLW6/fhaHTa/ym9Jm16/
wnaNuqwIFUigkVD8LqVIB4Ha/txfvEnyF7oIn5etyz1csIWR+xegLZ0H1zLhi6k6
HfT+AterZYttiBecaxl9zhugW58FqDJ7FueIZWzJQjC8lv41pbkVfS0C/wFWlZet
mERJiZui3tNsUDqaheuSU9VY3NBXkOKhYNBkM8kDYi3VjPWCjtNFcAXCOeqAJRXU
lmy7oQeFxiZQ9v6NeUs9CATifaRmNQWWc4XUncnRvoWtrWi5BCQ70IQ3farTptop
r43/IdCT8mlUGsTDZQ3duIW813B2FFe3Lr1FgZlHXH22Dk7oh2KmdzISyhfUKwsc
Cu4H7GgAeT+GZfnUdKASQrzZNUxvgP/vbTDGYx3BoLh9anFYDpI1o9XVLXigua4M
DCfQjsLNY3PIEqx7bNyNXyJ3xGIWKSi4w8wE+AyAqYyeLmkaAouxWlPnLiwoa+Si
JGUgIhMEbx0SZxbS1SoDcNxK/iUH2wzU8zUB9nEZjNyck3zXZoINWzM9RFQRJCfl
oTttpd1+Zd9oaNsfOOBuwO/1l/DXQq3cElUO87+VFDH930l3svAJ3vQQ/SThgSky
M/aOsCPbHqJxSnr95kZSFi392SXgPcNZB3Q1LZFjlqI2OY9V4aG/hHmxCnhDXExM
58mVIU2QhhXmQXydS4eUU0p4UUNJsFWEngrVmP/7KN268plf8Ox6iBs9FVSnaDwt
ITMwZuSMB/QL/YnmfesNFSMyr0tEux4q22a+8xZS4xhQcTr31Kf8xUZ5U3a7H/Tm
LUYApwxtcwF8WZ2Q9eLqxpWkxyPjWE+qUqjW/t+D+YufZyiFfRlAVetEQoHMrRJz
Yfpzx6379r7Nplo1CJzNyAJHjpO33fgAkkrL3XT7nPrbuw8dqmuulopcxW4BPciZ
B8lheiblKBIxMZtS6p4KtGaMWxD2qLkAFeG2thhOHP/Fd6aiEmGwimjF2culmm4k
VWi8XS2wl12QMzn2W4PKZEDRYank4kPPW03FyQ30zkHFC3XVH0Rbmv0i1hQdUR4j
Dj/Q6q5TWIENzMduNOIjIqCGVBYQ6DXpYP8YrnLXd6fGr96HMB7w3qpV+mv5/eev
uxeGidHV5WK3uI+rQNB5Xyiinr2ADa2p46zqEHr0NSzP1DpXbJlpzHgTeV34+ISz
WjtuJriLGci9jEU+L7JVkehGGkqceWoAhL/923PpFlijnzUhuyGaZC/xqvSLXEC9
woXcRgyRZFqqFLKiHB1iO6AUBu6SjYm3mjlfFuoK9FHVN2nXkIlz6UwiMcSOGQw3
De2tC4tXGmPW/caI6ylFAtm2YSkvqzv3tEZcwl3i5DT4oCdxdyHJgVsbeu/5Kq/q
9Pmr090Ls6ZV1raeITzok4/QApzeLvWCFXF1LpadgChFLxXV3xwOTHELyLmCcj5+
uLSMJpCHzczUbQ+V/Qm0JiY3b8EEIwauobWV3pXyfnFaceJuwhTs4PeEF9Yy9khe
qNbawX6FHA1ULbTUjKFITmNZtX8jvGwJ1St7u7ihzQCH73bZqoM5W4Hum8mpPedw
JphNusqWCEAIFjxx3qQK1ymkkpCTiyEX1vRbIg/5KraQuo6akk96AD3eio00/Zhr
4/97sM3+OHNTVdCRYMp4ZtnliEakRku7RLpTFN8NXr6ahm8z4n4BrVxj/31d3JJc
GxfOdzVKgNqgLTD+TFQ5+cK7RnESu8wEXmwo80YK8d54N7JZdmJLITwlLVyGyB5z
mVWEEuwSOg59gqaTuCddJ/wj4mZbyVyNJxt7KDgExUwbM0MKgMSc27iSGSY6i/pg
PMoGnqg+RF9m2KI/OXpiJBhzkERc0J9Tdsm3+c3Wb2szzs4XGBlY7mFN8a10AtuU
hLdB1IOZ1J+sxAw7xGmpr4ugWWNwRgqrRAN3lu3QijkRtknp0OO7IU/EofJtR0VX
ObiIpS3o3Qril8p+RNlkZDi3feYdhnb02J+AjXQDB4b1MeMhw6ROB1cuSlivznXZ
R0QM7qKiWh9fRP5pdIkyFzjONizn6P65kdaRyqsjcWDKRSWl+fNS+CpulvHRaDgh
MFQ91ai2WzMXPOBq5Aj2W2PG67hKBM1bDzJMsTJx620BXPRK/0/67o7EgBbkEvxi
kuJu+9WfsQi0d/at1D93gjS7RAt+af1tmlDFsDZCxS7BtZTliQQk/FM7Pldc85Dj
SSo8g6UVmATf+/3bG050dJE04GiFqkTLHPHBinL9HxQcv47BZUzXATfGkTXzwvwg
Lb5ox8vLEPMMVcAegXmCmJuqXh52IGzHjnMNCb4EKInE0V9Ty5/QLbTGMPey/3Us
v4qOrLVa4dE3nIvwLK1Oa0bm51/pOUccMgnA9kuwDXdnxviX+u/IN7YppTzBCE/5
CNWRPZj8eFaUV0MRy9sEbzkdd3W/L99H1pUXnxd1Cw+J6fe+R0u7CRCdAkPAixRE
piOMLAIVcdp2YKM2km0ba76AFRFs8pwZbQaUGlRWsLoUCAo3GEMNjbQ7uMEZbIGr
3k5iXmbmdlUGO4sTRZEphf9SJK3/mUF270Bxjsj+vIkHeFv3cNNyql+kDchB6CZV
8djkr81H6lDowLAQ5EV1KnF28fCySbjB6Oe3c/TvFHyu2NiazdWplXvRaWwrY0Iz
d9I8du1JGv4ImTT6ieF/7bH8V+ZfdpgzglyCwXDkFK1pq0vbwhjbdM8jI0M6b3ph
8DLQC81uNOrF1cxRgiVleaQNdxFk1HrYaiSFLuig6h5gL7BEHRVcOjZiL9VgDOJ1
dNGjKSlJWvSkRLu/RFzPkhzEdViboIYFelCQ9TWrVA0gIKeGMY9TqwR1LbJbiwua
DMYD7Aa1u9/+ZXFcQYXuJOmHTUEPSlzzGrGoQTJ3pdfC/XZk5GVhPVC+HT8YnjkJ
em5Hmrp+aDTCqMdAH8CN0G9mFYN1UqhFcpvYvJ5prfZ3RTgTvUqFjNAmZWWI5lmM
5YO9La285y22AjJ4bu99qxQ2G2/BbIphxT1qwumg3scFMu6ySib5FBWRy2KvY7xn
bkE7QNcheWQ/LUnmlvzGA7TGNWZht+kFP+RXSwpaWAoM9Pe6UqnemUlgHWg71Y8x
5VExNHagsL6X+pTl8Yw6snIfCSKPwq75L4yOdtZPVrUZJXXHnV8amp+BG+A7Cr/T
dI3pYXWrmjYhiKask5fiUaSdTUxEcThq8RHR2CJ9tBCLx7bCQQdCte6166SOUkXk
FBhhTzWZIFwELP3eQfiaXOUC96iOCn0akyHTnKmweGSUq1FiE7+1OmLbKt6ArT3F
jxsdwsjHVctIde2MMh/AEUiVZObE0n9zi3b9b1QyzG09Jz7UXvUpYWMSDhUyfp68
wZps/scVEbVKnZe0wvIykoih2gxrky1c+MSdQGCrXI7emkQICowxfRyaDu5JgKsI
cqc5H3ulHErHDnABJhFUpuCuexRabtXwoLrfjUqPzeHSJjaTZikzhC5i9AjUPSjq
vaP43zxaBqbzzusRd3BDO4wwx/v7BkKe03xrd4CDjdYPqWEQ+cCv52FfgjbqUYMW
3cvEIzc7xZeXOJNKHzePU+pvnzNZXEx1kqg84/B+l24RbX59PGxcUNKQT8L3HSoT
D+VyrGYByp054OcFJceARzuNvXRToHFAXoO9qkVjvVLyr6YY5ckX5wTWKRsJYB6G
/+TgjG5+9XEc6+3f4QmNNigdIZZPjwPthBDuAUG7UdmOIPV4LnW/59EFf0DBLykj
m1Emxo5cOlz1BK4ywPXWgUpt9kkLxEaAu73EWSiLIzhHo9n9dzATqHbaL2OlUA2g
lmPguOpWPvhP8HcF9SU4SbF3NbdVv3v/HdkntA449I3PPHx+jJ32tiwDjmcW6X0R
2KWkYj8GsdSO0ce5XP8AG2bFIP/agzJU3LrV5eqGu9DlR4IYGCtMdxiNLLjJaFG8
R9PpAazB2r6uEll5Vd/YJbSZDX22jJdn0vyFkNMEiPB/iv96fOTuIJVvAFuRkbu7
ZSfkokVBCDPZp8kOLdfsQtP33idO9tlcIq15v9ujBxXJ3QR0Sq+vRcP6egvu5kAS
JY9pbkCVHzG28/Jb6CJHcSJd1xaKD4vAPNeksXLmd3DX3cQP5B93Cb62cs9pSN0C
aVawJ6W363RYiosGs/s97GRhiDGxT/RAhM+WYp3ufZFs9dV3DcLRWWc4kvo6OxRu
1I03ANCO/JJoFCwgc8t9k8qAZ5WKjmpZyonQatfi5cBAe1zhlnDkiLRSgn68urIA
85hjXAMY1pGMea/rNdvkg7C0mifyoEjfFoXifVfuKxzJswjwE+bdIkHOxhhMhgvC
o+zCC4+UG4bhfaIS5RxX1K+6LGWBaS0RIaBfigwPnMcj0LPx/b0uaTjNo8txVarz
Z8fGh9Gd4muEPx7JA/BeNocxy67d0xBghPOn4BkcyCu0Kd1JHZbesv4q1xoYcka6
NZTufjwtmaQlrinw2t8MWFHHLRp85jfC2RcTHWBCttfcF0Eet/sNcF0EYmloHNiG
DY8paGfM1RS72fQNMSLjH401ZFfN2bqWl6ZGQU961YWHRNxuLog4/29Q+Mxv2bFE
fm2jOAMxA7FU3vnvydgwzczHk/pwu5HA9mLrt0Bx8lzZKpewxqyXAYWZ01kd0mmU
EObpFPXtQ40puGiLegauoytgTTdhvefZ693oCxrBokOhFw9Svf7JXLkLdH7YYtD4
M+IScp7SgHH5xS90HqpTNi7ypavmoIxXcBb2F9r3CbI25azhQonYzuWEsuwxpgDX
cGzxniHAimSggOHKzt1RE53BQSQo5Nf90cZ5bU9tpmOXbJMOfsZKEU4vA5t9ZwdH
4U1Ku5rvHH5siX/ApwU1bivBjcwvANDZSjoGkGn4qRCixhW3fCnchC/pNn6P17mh
e7a7DrChmEMWGjLyXw2X3TNlNNS3i6Pu2iu8bi6C3LvmDCmlPX0k3UDoi3VUDTBR
K3qTIqy6Yac4e42lJOyuZbNk5w6oNcDzx/T6DYkoWCAGi/agiXKNsNYDpvJYZREe
ltdZ7Cfdi09SYX19prunuBfe427RpssBKevj/aLFeSVnH1y/EEXs5pLmWC7hEaz/
Hkl7EBbKar+QjuwLzznMT6poo5xRjkn3v51hyJmsYaZeEQIDU584Zo9Fu+27+BiU
YcV4DyIpYLEHmSnfYk0Y4g0OycN3jwmLahmAbIzc5HLHlgmZLXGjhgyeZ4dRRibK
B6gc4mPouZQtFVHU7DOtlzgjJa4mP+B3sPfCSDhd/clFZ6cQQvUJVazdPG25NzyW
wpKaDHY96naKtLahuGCLrRXG11fzPiOnXpK9F0pS/XtGjXZbMWLrV2bkponMeEZh
isABZGyvwozH5ffNe2K3wjvO7mv1C8F8Q/YHbVGBkpXOXXqFGcbCSuECApw6ai4N
XFeIaLiWTNPg3GJksPE6mGp01kMhNmzvSmy8Rxua3GVmJTrRypEYGBkav93dXM0v
k3ofeANaAemlmBd8FhUmLrhjRuAAch+PkyLvEunshwgoAzfKLbd742Ty+DPqROcm
Qzwoy1Ja/aUMcKljMMsvD1aKHNgli4M4hy1TL6lA/PPLKXwW8rf7vmf0iGBZTu5J
eR6ApGejCVmcv5/vD4kjMtj2YuWnM7hq1p3ilk/Cd2+0UMWdD+goe4By365MU6uS
EclyYjGVHz9VX7KGA0bKpukQTjLpd8OEMzCDw7nifhgY+9Ql3CiMZoxm1jduZd9P
ufsOgTpcoo3QtwrZSgzYgi0zs8qb8OHn+dDlgE0vPrmOdRf6NY+R1ZukVesZD2SP
bg8J4dkYqnRFCxfnnFtwmDIERzAOG+RwsvjQZ9oXTi++yk8+yX9AvsakYged0Jmh
ew8/+/GVVddBakGl+T4R37xPcc/f5EAAho21CTjks/XDZTgLsJLG+3EAdiOH6ZlF
tSEE0bXR7xhepOGY68WP54drB706iunR7LnKjHxUcv/tiIIjLR+sjCasIieKJs0f
ZFjZDAslJ9K0NXWxMLiMYoJmSSTk/8pQlVLvNxH6wneBMNY7Gsqc+j1ABO2T250v
GLiolnEyWffM4f7KFXlKBrJqdef+hRstt5rDb53udxsnTkzN5hwxpVADXz/L1mNR
G1OM3srnFHpw0ZzDgPX4VmmOOnKQLsBwLn0h+pZ8bXHv6nhsW/pgytNgjxkR64wL
LZ5KT3OxOAwdZNMX8iwYr5GdEe+4BOOSttYfZIY0tTWQyTP1mDbNSBJOzUlZ9rAs
B8HYfATUV8ZnyBtd4mG95CqDLve7i/QCxBMNcEBTMsH1fl2p2PV8OV8wR9zO3hC3
ykZ1u+s3DfK8n4GgHdeFGV/T9l78qbkxxdCp4+RdHpVMBOWZNFfYSXktoHYGgJE5
xzGuQ08p9famuy0AZvm7InrNSvGbxkOWO0OA679b8NUvcQBCS2nB4KbdKZdzg3Os
4CJP0Q3mHvXh4JAqb+p3vVgO8oSbg7ELI0WRlDvGccL/eV00hbL4xTXOuwrp0l70
vPxQiwZfNC3wLL2Wwr+AUhq1DdYmyIq4EOwyr4PKePlMp1/6NPj6F9tNJaShS2jB
Ja1+sgMQlGkPoPErjzFGpw+Ea9/bsNIFUxuw7QEwTZXBsOBMZZqLfWCxPZzlSl4J
EoXonx95mxx5Une3pn2Iz9SBkAaF4ptumJv4OoqgWSBwGkCX8sTj+0BAnU4HBU2b
manxqPcrvKKqyzJ9d8Bx+MFTOSjpeiwKZ4p9DHSinCHmfTguF0o9muzjh6UYTrO5
2gQxIRhwY4RmGHQOgU/48AkdExR2CtAwYkFPhjDqmcqadRX8SafUTGnlWtlpczCF
/IUehkfad7rEeR5SophRTWLz0myHz8buahxxc7TPfSk7Cc+eseM+bv6yfPtg/wEp
nX8nK6qhPBqbCClLFW5Gr1H8IKnJSi15AL377T0ratRqh+LeG2HtVR7AVpGj9RKq
89MMe2DS219U0SSzsVm13Fpty/H/P+3heL7L2dhOBDouXzmSvKC3HkBwBxAm18ok
NtqGrYu6qQ1eAPnl0MaE1XA+VFYTQY9mXfnIFx81W4bKFTCSidrTuOR2IH9qae9v
/vMe4Ipw6OxgFCAeI03JbxTXXgHqSyCUH36aAVVA28XeANzMTCwJ07XcMJIeOfyS
QTDO20dYkkAclrzd1zupq0wCXWZfwN+7yOM0oLKbHEgyyh4pihXmHzMKodAp7obt
X/SAlInKTRFbpmTwFUnfQTIiyDEA5mvk257pZsxyiGDtZOxl28udvSgPZRv7wMMW
VCVu105MTmPeYBFK7jqA8X81JI1VkjEqifwnRWwzWmPhy+icclIWpPqsPXxpviBd
lRfKOw+NkyG8GBJRajEaq/0fQRVjSbdq640gEq2/PX+TxgM7VhwYbVIl0fjbZZTC
RaEwzU4JleZ0NtSboxGxY2AewJtpR5RnEdbeXfnPtZUfSi6sQ2zPkbgZU64kLR1v
goh/gcLKCY6Aqc7iHaC2ShDFzUKSIRVUge6UWo87JCjTyY9X1dbuvVvri5RNwZRc
oG15IETHBsPCDDIJuSlGoKw5a1i5dj6CfgLfXtImAN4Wx/NI72Vsd1R0IonWH38F
vW5SomotvvUw9Nx7FvvVyJLYN7+r9Gt47bHjkzQhs0Mzy8724pKF9QWIsgoWTGZQ
yp5JKe4HNNZZUCSV9bgoKx679mEntExBw8ctIoSY8frVTL/IT5Khxy8JKJeq846z
TOPOfYT05j9q6jEfOEDQvfCQGGNp6DwNMuNU4Vk8gWkaIrd7iedAEtlnzaAkfg/4
nGdFsLi/58wncwFZ2ktDgOMB45cngaITTJYaFp8vc+LA1RDv7UO5fl8ujIEswgkF
GzvAlFr6cP9O8P/HmIfmhTzlMf4FSj9/umFEHgeiJcPzmI0XbhP5sEFMINf1s10/
74eXWsKl4mqyCacanI8B+1orfGs4i/4wCXkq9uuxKW0Lp0vHw7dZ9NzmkbAZhumF
hukpXZiZmxVn98PNi23QJdfuc7M5+M/7QRCdxEeCUfmNIMQ2ubrRiKmx36A846H6
5ktoNu78IQLjjxiiIvmL156+sE91sh/ySU45Rrb6k5C6JQ5b79KpmSHf8NazqrMJ
97q7nicEl4r9cf3fYtyyXYj3E5VgCn6mucdMhni66XtuqY3gUDWZrqat8r2RzN5H
z4JjczbteaHd/URUjy/CQ9PPaV0+XLB/+AHMc0aHHpDqLmwHCVBdPTGLdkNeKSpm
DzG2tVSA5Z498ju3vGstrKpnPNZIlgQ1PMO1OD5XubdS2WeCGFkSSEtLmfnHWVyn
RcPaDW9zXKDCW+tfl9oGeJEJ5F/YS5O84vRLhrweHjnnB/LxwgbrihqiO6IdlFB4
HnZsaU2FSYvtZjnUiSRN5zFKkxW+NAycDXhNVbB67QZvytRPJVZC2qxipBNEIIx+
t0vGFi22QxOQPTAB6CPOE/0g7IVF2ANgYPa+oa6Su8kHTKaWLbZlcK6FwQLT9gfO
UGiXh32gd2A8n48MOoHGrZEahmGSXM7i+FXIYyl3fkG050aCGx83hXUrZtOlAo1e
DPi1EyolcypDsh9mwlsbFbOh46/4Ejw9aBEzcS6coNSW1bvrkgzViGMeEtkesDro
i3aE/v06jKz9f29AfEyolWF8FduS09iE6Ef7cWBb4WNP9nWgLl9+BPt+FUlFy+gw
33isBeJ49ouELR6cHF8MYLQXhhRi/IaeNV+7iueVVS3RnYFWZNc4vTX05XcEIZOy
W54b7rqPkyekaLHHKO3scxyXILrEyvyupG3yfUM+MCDWLOLU8Xc6bk2FmIdpFLbx
rs4BmCaxrUKI6+eMEdCB60bXM/vd0X/t+Da0f1r4QV+SwtNLtDnRlobqDJPY2Wir
DhNT9Xjm6ZMezZoMRxFDdgIetWaF893nlvbrUBPA87am5MgeVhT1oP/xx9BuyXzR
MM3kJNiUdKpyZWxmrHyEN93XzTDsb/+yvsxgeuQK8fo71YIJxqA0dfFqxXfBBN+H
uPzDSgotctQ7A+6/JhlQP6NkMg0CLlmWSBbc+tcOq91l4NhNAxFpTD3a41LJnEkM
YftR/ueWjJnShVS1uF7YNvSDl/mStsE1G4PphkYniWlIGdNhUAcZLK/Gg93Ob1Es
oTUdXf0cR3BBvmfzxy10cUxDi0CvFQt0Ra5qNXP4Z6tTl2I46/Rfopmb32zU5URJ
/7UP3oW+O29c5Nb78nu2Gk8bGlLeFLpT4okgu2Q97QFhCZLJk2EdGQZYG3etsKal
OxaJQLiJq2JWZTOgZNC+0Om86C2007SZU1bFBRCDux8ISgyNMATG1X2uQ2q6DpwM
rgRcL32BO+iOf9qCzk3oAGAfMZJRpVdUxLjHAVNsnnm/CXDa771hTMI1kbfgk/uo
EG5Camgmtfp+2bMkl+o+LWjA/Fcpm6ikk79dNl4OcsbmjxLp1iuPnppAOBmFZr2r
sYF51v7zH+AIZkmecBILVM8y42C/vgHgH2jmww2yS1QC+wabFqpni3u9TRIbPXBr
WTqV5wCzTG3RsduBa8Vx+gCws7EK/1fcZS9/cjZODk6uCBABcVfHjaaAb1wGSOw9
9cp7YyGDPyQNGV/i6rlYpoNJy1EV8JFniJNDHT7zwHj6csxCv7KhFGqhiLgz3P4F
Ve/cU975oR3/KuB3xa8EG4mjVbDGY2StsQNFh23WBkl6uKHRZ0ZQnt7zzI945TWZ
yvFlPo6Ps5kDE69XlEwx4WkfRho+RVsXDvb+JbQk0T8xzNMiqhJsOHx/Y+OCtGk5
GZFA2TOY2T4QObbxgsn0xjcfmBFoxmnFfiy3JdvadSeqx6RdqMfgQFF4jjo4JgEm
ZxQ7mlh6nB8+LHtV1GNWcqJ9ysIipW8uxiKg1j/ymrxOiNjiw0f4fhJtTKYPcRqE
xwMCaZEjhR34lT1QRuUmjzQ2llqSevffT/MQw3UgngusKMc78BaljFPdTdAp9cUB
aUhNKuN5m6/TlbLg0hmLBBRvPaUZ8lZl7j4+brqBZFMLekFQpiSaGoUDLfh7CdPf
z8oU1FS9KgmmEmXgY7nRlibFsY+YqWQVF2yJzijkakr8SX/mh8djylwSbbbHIaqS
+QAbOdvp4KsLqULMlTdIq7nQ2K3v7/qr1Z8cSiWGo1K9ug4PvPTUsATW/EM25kQT
yHHXqa6UaIupeCQMmJa1/AAzXuPKk5Dz6zMMFx49cC9G53IcerCjQVAVvEWmzg0M
ox20iG1aivZve0zupN07sqiNgUgInMjfPSTrikX4sYqXpgKqwiJxYYwxwBsR93Ta
KH0HS2GFYt0ygGpJ5Z1CnhxhSi0DcGrqE0/EIp2JE8wduYv5ZGg5GVP/CkoQlhDh
uka4WDWYZLN4aj02Yud/IsZwaXL6jsRCXHo1iZ+BEsa7hqCkix8fh/j8DU0SLMv1
MH63ajW2CfzdT1F7zgEqFbeq7xHvrYA3WPs0yr7An2pxEWyBKAGCM9xM01TCI4ct
cJqSuCG18E41YKRG5CwpwmBjxfh2Q4lA5ZbjIFPGiUknzQCrbigx8uI1hKV4nM3r
GFvJyjGM3tHQIQnIkJIYv5j5WzFsS3PlEYmh3sFKDFWl/E5KvdjDjJmXOiU5U7jB
MF3j122d1QlqsLZl/AO6zxB/oUolePCyjJi0/clyknIbhKCfx1aMkm/Lyphs86EG
hTaueRV0ba/jxlDGdWocm5DTh2frrqyBTkVjJP6fb3sKWuZqU9uau7PL5z9cSAhm
ueK6r7wCzKC3zjJtKY0v2C8fVGIhvsy+lM2CJId6ortWDdJq3Bm3xW5VaHDWbEip
6TueLSxIu3GhsDblmYMhQAcRzBL7iadh9aVh3nwANzNT09qvdyQOXaGpkoMDQeHl
y6wCLxHgYI4a0ZZ/zxONI5Vu/XXJy/OVAxbW/Ag2sulJPQwgB6+uKZ2y2dWMU97T
mO1wO5Iw37X7VB23QJnf1V/wO+5MSmOEDb3LBjvWf2BsRfy66k8Tdo2zBg+cKP6W
3Cn89tRex3dbFWEWrB9f+dtEqvLyuC/cpPE0xoe5xnC4Hd7eU8USxOar6KhvXxrg
r+HvAK/eGv6WbGs6HzDUJXEVq8FQxjas4FoK4KmS7R4edbhTubPjsKWhwBPABy+s
KV+BX5lNA1c/oI/9RdOu/Hd/h72Nxj6pmT89KzpzbGMj4wxUsNEyepXBzXY/P6nl
VGx92xAzXgQLkwNtLbVSXd8QLpesjgDZpsTtuXXna6V5dcUUdRke1y/kDRoxoZej
I+P5SAQJD0KP13qrPGHzlPQCfql/fwvsqMo20xs2AiCrDH+3fjvIVngwrFoAw3cb
eKicERzE85TLOeVFBMXfIV++lNFFhxw9Ag/LZFR3wWLE9N9Be3NVR/46CgrUTFKj
LOZ6Qj+4HOXTojZ+lCLbOzwuL/ClQFI07CFsF53cFEyyGVOX/zOtnwvuDraG1GaX
nH2jkR45OvpBEjix7WADUdYpcAjLZd75Xc742czH61CzdlmtowCIiZka5h5oV1Ld
PjmTbyOpDmVrT5zPePAhno022FWTAKLcAlLu1IxgA+xBHraIIfrTkp2fBhZMeWhQ
qPBasYs/fG5+UeT4JJTjnuhAo79eTKAsYKIWfIAKW6w7F7LWMKq+PG4VC5u6+4HF
Us2G51qsP2KaZd+5sGXcnNCcm6OnbmOVD37RylOeuXSOs5Tml+Xn3MT3XuzRvUjr
jgTUpTRSmZsPa29p4m7eaB4nIHT/955IsObp5iH11uqOTo57SLbRgoK8C16iuWDP
jY04AD51rMwLhN1L/1SCUfDlugezpsAmsf+vGFzsBRVicGsCGBUqucs/xJ8FWtpL
MZVc0lidAjtVFTPGEdiXTW//FqCyb3DpMts42ocdptOpbGB52dbg4OR4fL/6ilQs
hzwI+gknf3yT2uIbImFVvEa+r77MbJFUIKTHewbsfEeEvVsFKsB97XF/RuDjFAf/
7PuAD/KfsoS3J0gVptmF1zt3KEeqHOcx+HeafJ8T+7ACHBlzTj4KjYo4LmYGo+3q
/RbrnOgLw9a+kIg1Jpk1Jf2fzWSMl81SbnSRbIm7yZHRg5yk7TCKqGQT0q2p9ZhW
3OdyqwtNwtgIRLUv+Vn1dDKLVFylAF8fTmSWorGAMv9llFaHqB5Pslc1n0jETOB/
cIgOhz1MBrNZkYWawc2MVSM8lVCex7IoIcbabFuFhsmRoyDjcGHuFugXQaOuhLJc
wJydVA7acPOMPtBs5BK4kPIO7Y6HQCT0Bpz06tWEgwVxNpqLDvl0PdWQ2XsY/ra0
zRYB5dD5Ryu6ZURjMo4lDscM7TosvLkT53DCfP8K/WgmwfYF4WiSM7+vOj/EwXv9
n9Nw3sZw1y6rh+rxPlTpgReqoXXL9b4QKNohXTUF5ont/TDwgFds/GBaZI8PepAC
cY8pnvivwuhtso1V1GR+wU3GXwsUws011F20z9hau9Wg/S/7zEFhmjwSaCu/Xnf/
Ulr+7E1FTFLVW1OCLfjRRc70FE+mjgplW/yZUDtMdKJEOmQVbK5rCswrVJ1FA8Uw
Pyvo5HkMjdhFw9I6kkCNv7TqNv7xhFTSihHfssgkroWKWWryk8JFiRKMjufsVZ6K
JOaNgH68HMgx02hztUQrIR1CQO+MA4ain0D63tjBonS0u/77PcWtZkz+NRX5vD0b
f39h+nu9ncZ57KkeISTkTCS+aqTKdvBhbpuhCBFIWdqJGPhpeDaq8fwvF9hwlLyj
lbiYAXRIDFIygFlrjFukjA4fsDHr9tlvp67j3c4TQITiBA1bxdHvtxCZhYMEYwbm
avGh1kGpB8/A2zVErp7nspsPnSYAMerBIcZpnuW1tgAHy/r8n5CkYkciZzFvE2ww
hFGzzuR/AplXPiH/vL+losTu/OVJRCA5HsGFLJfL4e26sTO+Gy926qvN+S1IGk7W
OnXu/eyJB0WUh6Ifz6J8ef9o8ZAT+i9J0X7neWMB4bYZlJibChYIeUO3oTMkhzZF
hMFRuUQUJUGe7l4gNHT++W4gGE5UdZGwZzyltaGusbWohFJ2PVNYXsz1SWEBMb2A
US1+9MrzP6Im2aa6h1FhNJnBeYqTpnv0g/I2ttfuohGkUifWol2AL/g845m0xMaM
OxC1d9hni/FbLnDlLT2ie46ux75XzWNQvmKj25MYeexy4zBnFa3p5Em7R2mrldt0
UIk6K7NAIdCn478CoQIuqeP9XrkfPiGg3dy0JUftOhLU2lNC1Xwg4MMLZOv34fci
jWylD/tGUualUxMTEhvYnKr4BPJe0525bQd5qb2HGrh/naannnhMjqgoHXw82GtO
wCviPsztfqXe4Cx/Ny3vNp3cpnA9j+ARmEkc2aaYmyjuQpPX4cH0vF1v4yCpQ6so
6QcXEF+DKPI5tl51QwDrZUg3PSi6api7VuJoCopJdbdtEhlVmuQtyI3phEpVLK9Z
qZdMvHQNSHXwoFjuMVtGYm2y8p/tJ4mfrjDyQVUJxjPDWEUSbEKvnbGHunl/F8hm
c/0BikNlAb0By0BFnf+PmVnGjFwg+xJPukIAxmx3YnHZ7qmb8gAeUmmc1ddFGXx0
mhFa8LyOc7ydNiDvTqVhKyezAtD0ou7S/foHlmSGT81YYC95QLCD48wkmcqJqm4d
dR3+h8y7t7owHbemv/UkFIlpE4B/RfZcMvBRKnSOJTmDnfN1Zw8xCjna3RrcWHqi
znTZaD/gyJyl6GZ0i6DfIrDdF9yrm2e21ynJ9U4S8zrrrztC4Qjnga/RL85ZIyKI
svtrkv6KsXJyOnnSbcedRfvxAYtQaAJ7Myke8sSNLPISmfZZ+ao3VPauKOWZpKma
K2qGpS3LsXEdBL3mlH5rU2hoUZTWJRxFY4V59wWOoENgV4cMQp1ZsfIZpdPrZuMj
sEEL+F8g2kMpcNkPB2Zr46cHTPiWwSJvFi8vdcBa6dtFkMoyE4f8gyH6emfP1lWC
nKHgHUY/LP6FNmng3xmvdhTUs10o+ZZpf/lAH3o6jVXhqI9GPDxPTNjKSzuwPUIC
Kq6CAChcLcUVDgaWGYi+eDCAr6NJ2a32+71JFWzErf86JtVpltORuuCGv1uZBiU5
vc4+k8WbJudbUtk0Q4X7insC23+r9oUm+QFh+ktgUxJ0ATWG2Bu1UiH65XB7/bmb
HNjqmFaKwFbgXlDPWtL0oqSu/VXv6YpcJfsvoJOOKu1P8hVvnkblmaiO9w9HxI5G
GM5kgMao3m7DZtdutZWMLj/2A4dUA2IPTpnNIOtFbiCwDB4TkW+oHRT/t5Pn9dHf
w7zcSSGZJA0SxJIoRtC7oVLvSNwOHxeSYRv+ezZArc3zrXmNcFctPsBnaj/RU0Wo
EpxePHRzPBGxOiDMSqo4cZmdZXqSKjGnz2vTa7xV7kQZ0/wXPFRWvt/BnfH6dKoI
ZQusznJ1PUkdoumY4oE7JNPJXjarT2KpyQHMpzpatpRHIWzycNPOgKvZnbtvqNy0
TrvBOmAsU2Mh/P5dd+mHAMimXPLPXrgWfIwPhnB/w4AnwIWrQpJjtoYTj/7+iLaF
Scu6Eu6EPXRU3A+IRcZ7gtT2b5WGqtuMxFVbVaRR+h0f+JS7eh5ehN5rs7GMJXH7
05vl8wD1ptVIKeUgCixl5jAM0UG9U+Y/GajAhNQ2Uicq1Jxn2YHnHkxulegymSXo
ZhuqTOYII/1bz92rh7E3XdroIQ4LRyeR8A3p86iVIOw5swktvTTiilKmM2iSOVSD
+4/ImtRhOI8E5Dyl6d1wEl9LX8r5EUY7AzA2k+hlZd8a1NpH/kRcOC42HFKI54Ya
KMhBzE/0L8+ZNdRt72gdBXTbBHg4NY7OufrrgSztUiaRBz5O/vSLR5DcmJpDsIxB
xkdzdvrSkAgaRHLNJFMBN4XlXeaRGU4Y1SUNo0PW5De8Z+VKSW7ihk+YY5Qfq/Lw
LswaD9iG7vTKv+27vcHfsKOPQMuSXpLqOaHNM0Yuj5qfZ0VcZdAfiK7fYYyWWx9H
A94l474w9qTqwLBx1Qr/gn0Jw4RszdzqtHnelfXqDioER5cYrjJ4FpiqSzJ7BqWR
Dkbd9p0b7X0NpnokaL6cQy0LjsnSsQ2vWCWRsf6F6ICTaFS60KaI3v7w93U4BQky
zvakBSPrR6Kr6Rer1OD3OGb54uhf7QYMk3Zq6NUCpD5WjWSCcGWxFAdXBtPNq57C
t+fMydt2YD15vb3Qvs+vZJRq5cmiEECxgBO+XwL9ueIFDH5oQWcr0bc/OUPoYAuc
RIAWVPAgww6ado7XZEJiI1te81GAy3KMFjc0jN6MA6+tCih3NlcwPmQN3FyrRnk1
HAJHNuTqEiAquue7Sa57GFSgnG8oLRFnhEmJv9IrqJE+lZIIcBWSJcfsSDyrMxrq
ZIGyZxjL8uC6DKN9yUuv7nX32EJ/EYxnkFkU+78Hlq7Pmm29a8Ta+tiwToQ+Mr4c
mo4yTVWUpd6PVFiIGz+6i3da8MBnV8V/fIMZCeWJ//F9Q7sTVhBN9fbuV2SxzBtP
ANbF0hFLsPoQDGSJqdYc7zbpesfbiqkTure3F6yKr1IdGjq3bIsVsI0OcT29RtBX
rKVbJvWqGxiJUkq6i/pPIWm6IwjOhT1i60k4KxI0JEw/s2WRk/3d3Ju21l04LKXl
yJWvWR8k6RyQPYFYOdptDEceuWD1XXxfLGS6PS8M8JX11X9NoYqNSY7NupWb6jNX
675d2RapWE4cU4F/OW8nXGW5Sq/Z+NqlIm+aVwyUmHr2LQo11zr4Gn9JenpFnz2y
pWlrDaR4t9HWsUriYOtelIwtF7G8Bk9tt3chV7QsnTcRZpKaiU9PUL/RqD5UjZAt
hkUb4OUNFiIh6DtG80PkierEFxQEN2J9YlAml9FT3euML+dpYb5lviSXF9EEJ2AI
1M1rC7halzBTTtRJRsDztp5yIh76JgBn7GryFWdV2p/XYplXRtFCga67bsqjo0GK
r8Dc7hnikJOok6YQ7ZlxJWVy4Rai7UmuniYoNWBSH/FIJ3lRvI0bJF60BvXATzD8
NhfpgHw4dVF/TxBSzuOkAUSztMIc2TXQOOi3RyNMzbuk67LhtyFsOURFygH258ea
z2Tl1lkbhjV2tqHESsna04n+vsJn0YT2KAAMnmw88SPf9ISdFPjSvkDfADj91xeJ
P0Ke3eNJkgXEkweXAkK+GZ2Fl3fNKCjTtoGdb5yrj98EbBa7iILdCWT9eTS9xCbi
umVC3H97eXUJkDKD2/Wx9ad3rYHClNI+4c4yoeG7cugGW4rqOZH4PBu3Jvib+t6O
5YDm1SEQvdODIpGlIUHiBpOS41IU88D3S2a+kFQqmDg2dCxl3Vt0eBGrSi6gM7Pm
ONc0a0ZNA1GnFb2zRIr4DCRdXGOgHuOeyZIgwB536N4PKGTa/wvRA2AF7CP0J4cX
O7Ot/USNILSGXbWCMU9VhBF+buhYIVEXJf7+qkMMXv6fCNDzZFq4e9fn7ZtnxK9V
7M19HoMxoQqthFrzfSPIxVqaWHeIr7VQOeRlYtkcTJLus3n6+xBojiEEjzmk2mw+
f0udBgJNsf/IS0z9owotX78f8XnegB7C7FRPrNQ+Q6px9rtCitXc/IZoJEW7o19p
3Ax07VQvqSngjR48LCW/wr0JBMT23iyR0rky5cYFmRn2Pg4fF7D/+/13Qve1ky4U
tTpDB+i/s8VQMhLRPxSqzCdYQjQa2B8fv/ZEmllnFpZZy1RVFQJmM5OfMBUuZgFX
LbjVauE1HE8ZsmL9eMaUxAizGBrAZA757l9Tc7xNZBIlPAZ5AVNoF+scAdB8FwCx
nMkOOQrsKRTJMmFiRtj7BWoR+9CiEjGnmPLPHPsuqrhtnwa6mT3/KL9qn72+daJy
o05HAg1pm61lLu6lKVVGW0G4Q4JKn7ONZKK0fThg2wjpSA1OJTQ8ukjNux3pc/+J
8JcvjetudMsbeB9SwPt+9voBmLRFPby6+Hs8BqmUSQUiRE6gXjwUjJFEnP3WbjJQ
7V1RK1EeC7/HJqaEpjqng3W/VEp1UulQDQgAE2OJxDtuG4uCRh6G2JNy2HdwEYD+
EKnQ2FhwlzIT01eZEsuiMuwCrCJewgKxUbR3OWPaOFMumtJe+/InicQnHTFJKP6p
h8I4caYHggt+ehjATw9gwftIdlJZlXQF4mEar9xkFuzSrQnpPfv/bNMmhCgnPFVc
HtzvkNnXWgIEpT/zPNtzRO/VYoL3RQSh7bGiHFzAtZNRab7acpEw28K1VgyrkJQn
hMxOyjGrRbFeU56UQkRkfS1sKn7N+W2NhDPEHVLMVeZnqVZZtr4nvBswB/8VPxRW
V63uGueKBBbwQvW+MSU1+W55bDoCppyLp1WhrHG1SE/3gaVTirDSxpfGGcvJ+jnu
mhidSGP+ynsoBuAeIOpotAugAfBGJX3+RV36eydhCA03w4vUsfqTQky+tJvjxCzm
UuydV9RHK1fVDeW5rI3f0z0sqIe/EqJIIkrF70mbmcwwtDyWfrG0ZeeQOcdlNqZ5
xbXwMyxT2wpTIHEYMMi76p7FZerxf4aJnYVoW9Ceb8cLm8Ss+UrUoQgtbtflO+fN
KxFxAT1S3gR+/Y7YZ4f4O/Ph3d4FNZ+Rond6ypz2U2lyFxh6fAl3LD3J9xn5g27u
c1fpZRb0xNMLxUdswgwRPMy4yT80pygt+VpyCZJPo5208SQHLitE2nbvKzpTnRRE
5cuxhCk5urZgDxyK5L3EVz2E9UXpFDiw+wKR0V8FufR3wmPP7k+a3mUB5oF6PSPm
wTInlz6wO5MDLysJ8NFMU1V0DkW3oN/dCvBHXSG7lbnvOjANNAcunJ7QC1RtDBOt
F8pH2lr+wznCTaI6Ei8FEIJNV3zjWnwc4c7WnjA8KrxrDGh5WRmRTPRxKQhgoDsX
XQC/rc96U8Wr+aR50XCDY7Lby0JSEZaHhFsrJlZFV9MWkW3SkqYxHq+2PM63+S+j
37j6e3hpYzL9WHVHRTjWA8HzO7weUuVTdWD+Wd6CP0xhEUWX9X3swBxnjXwsOVcU
Q6XFmeuWraLoh4cLsAVlq14qmdURlFoONiXz1RhGnXHJGX44ILNqhk8nrM0V503X
/IdWlgw0w9urNZpPOZDzl6hroAqI0Dzigrx2U4b6pPnYQbuGizkJKp2XR/PNpWC1
Of5naMkl5y/lDtdVQAEOPXZ4LSqRV38ecsB9aYRP/9SiCBZY5AvcI5+rlIbFk6bp
qHs3iRrFhWbBFUR5KG1H4N1ktce9D+Pmz/IUvpOCyXF08Y5IxrYwi1JJ32r8vTPX
2BqNEXzImmVDqKj8PGxrifX0bi8lJogMTVw/V56xdYD+Iqff3VKh75ks2Yba5/zq
uDQHpmjR9Ivuk0FywxusTGZDBYj1UCnPe9n4xyPOXQX0DWiqE46Wf7zxkvRvGR0T
EY3CtyNgXzx01ncU1nMdCVjpZjCpl51gtaudX57BMY3VVPOekye/BMzAGG9MrMjS
fV4k8LRqDBT5aEjfqX4SDjNiB/JshKqhG+/+VFoBovE7MC2XpOLWI5Epka1GZGDM
sLE4/y6JqBLM7HeGWoGIIy5e02qJg3WxR87w3MqN4b8cL6FqAJplNk8nB0VQiEbL
hxS5Ec6sDZrtilHdFQvHyZYTG1b3de32eAXWJhkatbM+XWiuuIeDZmuG/6RO4h19
geQ3J88Dd8PhyEXtvYEWZ7mUkrzcC4kbduBV97uB2SF2PKrRWokHI2RpejmtcFb9
nxir/2YGkETC1iOzJJIQzNVmttlQPsubbGPAYd8YxW8dKAvlLFVIF7BEBgswgUhg
UERwPqCB/ncI7UZmZuHon+ziQLUT2EVa0FmLupBbELp2YcoiqbQAZYy/NMHCO39Z
L+VQhkuUvlJu05htPJU0GWhXMFSyiL+VtSqbVKpb3ijWj4gTn1ksoIpvsM9ABtgt
NRyYA/NPAu8qxcgbJmbZJy1JeOvMPKtazeOC5377d5jTRHjUPxGSuj1YjF2ZwXVI
Vn4pgmqLe8QIa6fudRj7WnaSF0JyYtCu5ZUcavRMVeFavFNWgtsI/OBhwa5gC+x1
FOTJJRCl252BXjyuyGMc2Pf9K12JhCaBhEy22299EcCcy4DVJXlK6h7YlTm0Y/Bv
TVoXGFLYdXXelqZzrcga9q9sGu1dFMRE1ZyuaoB0H+xEbaS98Fj9NF8avusp4th/
i8Wri4XDIicAO4mLdQGWN6iLFqATOnJSmSVURbq5/kmXOatJ1JUUTxeAVI7GNl5i
ifBTudDMlnb4ogwxokY0BKg6MojZleBQCvLS/AEMufZnP4RV7yeXKy+CD79RIpXy
LGHdYq1lAfEpZEenIcEhuMRlRxQ+d+/IbKZ9DN+mih/N9Jo2pbEFOBqDnyrg8J1j
HHUZERrZ6L4aO8RMzh8LOwUP56V3Jg0ICy/6cRVf9KESpzWFQoLKKcnfAHsFU5UT
v/Xb9Iz2eN/26rDISbgcum5dbY9+89v3O52DzxQaLzj8tPvgcdvyuohWv7Y8nu4k
h2L5vkocZnzrI3pJwMxyGSCx3fv0JYC5+v5iqg0Qkb7Pqg44iuV3paB5MADiJMh7
Xr7zxhLN+O0mTGim/VaahKpAndpa1eS0IciddZJVCQv/xImoLg8p6u7SDVVAXIpn
FxHnNnVs0Ig4YqHZHCHVt0gKMss8fqRb+vdfHEVAEwo1Sviv2KnyqnICZVS6aiqw
4nNxUuMqLoEiPhvKKEYANiKWMjCrwhVJmlbQBiB1rTSbkGoWgqrpHQD74pb8cLQX
tHY/pGnVS6l9+uM+NUbVQQoEYr7/ROEs7aIzYzUEFShzS/x0t31QeZ94Q681t1qo
8T9Gw6KJXEkyHWzmc7BBzt4RWt9I4eux8nxETLs8y9wkkQhD7e7dEQvH1v/iU2Xf
luIHlYBYY2g7ZxHXAgK3Iu5X2Lu6KjTLA3HVanZ4EZh8y6ONN5rTcg+9/msNtgX4
QbNUQQQFqNdTKw8oP3IJrNWi3Ywf/5hlIS2xOOAPdiSqShdXuddWTwYwQ/vI0qB/
yQqdA0In7f84/dot23o9Wgcc6FrzHtmLkd3Bt9Mwd0A33NtsJTUeApYjfqS4EtiX
wSxM/WnaCZSy3vhaBXffdQ2yYi1MNVnMZASyCFJlYl1A4llmlLZ/l6La8Aido/on
5CYklJcvTOTc71+fVuZxIqEw5pZsxIHeKV3rnWx6F/4ois7XfBQ/N1rRey0iiJ6k
jrrilUvdEYmp5IAwh3wrHOSMAz1TP7EPMV5TqsrS+WYjn575DtPA9MUPNgYAP0UW
Fq1rSVktmXNvK1uDNQTfI5fjaQ3iWRRxrWlQM4ijZVG/oQP2NfdYoQxqESEPCOTA
PuJQhwI1VM48HDiWZ2hWxjzXBRTyMGsFkbI09nf4oTyrShtLxNYPS8w48YeOM51P
tAv+qF85H2xz7VrEIyXPk2EHSW4ybNkRyzJZxYJdMtpV4MkFmlGyPf7FhHWay4Sg
gjQFki+3L2gXxkSk3rBs9hB8VmkuKwebIXpgH4KRVWBdsk40KFcialalWovV/BvD
SRua0TcxzK240OIOopeAUim19S8iAtVFH4Y6D7wy9IkjD9++deeQBJPmZ3q+Vg+D
sDVCYWNn+ZskSuJz3ofr1l7AOXTtiY7/JF2OFnOdYOPo7yv8OMrQLhH2tKOHHTUQ
Gryu3Ov2cgtCHSbTsCMsWAY/r6s6l5cKSALBGOPYOWkJ44fxtK+dQwot1Sk/f0+n
YhJtRIMBxfRDO8xQKY+WkTjVOqr8MiQUYHHKZWFmXs4iiMUFksl4+TcIIspyrM82
ZcSLZ3ihYQXRjBgxKxpnh0ck+E/E6HjAWltDZIAUKDXOlDW5e8zL6EmIlT9hL+pF
BumRVbGlyR+f0uAOAxsAMNQK3I9YaZJBen/d3AfOb+MFrRrAnXU1n+Bs42Whumle
Kf8eWTaNOCF2/no9tCC/vmxfZ08pIDhZZFe7/MKgWf6zwh2bntKLtT4AlXt4Qqvt
YHct7aqa1FFdLAWzO++o18zqa1tOo6CGvChxPXgX1yfN6MBZJzFeTRcspRDecDaC
wPqTtpP58A037t+zh/IRD2rFWGRAfaepoh0TomZJmFwLXN/ejKzTUVRX8TNvdEnH
znILzFgxiuAbFzw3ABlZWtw0N7YPKQh00neecZBn5VksSXOHISkwItQ1k/Y9fFDm
ZvL2hSJGTCUHNIk1ugD/VDq3DMre0b2zMoCUTDh6NuzSpH6C1wdK2rtGx9IDSiLl
9QzP4RYHoIgirzYr78UXCNU7JD2r526Cv4bQyJHCMISVZALIragjg1u27dC7B7yn
EbIYxIy7p6FXhIiWo12P+NA6ndrtSiTcPdB2y0moKcGlnE2EndjdBTIo/8nqp4jA
DICkiIEj7uDFp5J3F1Ziqwl4q2yN6H0ycTz1VmaralPRSQJRACbRZyVpL9e6PjBE
P+NSgS06Hwn4V5f+3bhQCdxN6lj6OVeK9NgATyIB/Ulmzbo38wc1lLPLrlQTgZTU
g4n+eZbV2cZadFNIK0CSmn5v3K1Appp8P1Z2RnHhS+6Mu7YzX26R1HhgfRDWiKsx
rtIiL9yG3fGrgYjTBTEqPwXxoowbg0MX19JokJWj9ERzEGwoT3o2zvkFwpaHhV/t
LUKI0Lq4PTktApO2sbrElg53RAadlG78imAweeM2Ly6crhOVdr/EcTniJwryAK6E
7GggJXt5eSsNspuJOlB/ogGe89cYdCZcqSuZ/bQXfOfZftyvPDNjRJLH6A/IQRL0
fwlm7c9t87TuekuKRWXBXKqmZMfaJNX3iSBWhvZJUSj3oFiwi9jujfMytm2TFIQX
cvPthxE2gyM5q0n35avizstLEixlmT1EIGijzkAbFSllunsFrvfxHl+KiRxqsDIv
SODXtviIui1WKqNaQz+TKBuUAzrSD3HYpAn7vgpz3q13BaNHVATBOFGv9QET9NaB
ORrn5Yqa/T7h3l5y/ang3SV6Hu/XvFgZnrHn5UYRv5arnr6mR6dylN3Cn6DUG+0Y
GVLx2mKmej2cRMggJ91iQDW8+k7SM++bnWUhENUGC96ToSwtJZfVE2PniUC0AMXo
6Cbb6QjaRXGP9s4ANMu0YgaB2haQi5eF9HUVfQI/hiQLnqq2UF7P1G4mzPyjKE5R
yiXrWthiuVnMzq2r0f0Q7ic8YVKE+tUgEAdUfEniBxjMxgTHMEwIpWYRX/Ygzzlj
RvRseo+XSNjOq1pMKOhHRE2ikTSDOtNg6DLagvINFeBLpod+L448Li+uKWNSVK06
TJd6BX3A3G1w6TYNxMhQ6MRU9AkZbwZIRLmC6q/axYpt82u/O+1iZ1Gd4w7o59k8
FZSyXM4HYbgSToyk/nw4Cl0S/K7MhufL8SbB8RD94yBYyjosOOl99qN7QD1nuuo3
1EwKPyJ85MJMgN64OaOFXy2JBdGrIVaQUfpejFwJHwCWBxXp2n48nUO82eSWTuDE
6ddn5DhF8+W5A4jR2x/ySdTMaDC+Uq4VgKX9WhoPZzc6sxNkCgqV+HKBOi5NGnEj
GV5ll3sUzTVGOiRyVBE6eZFvao05KNcn1vETgebal56umKMmg9bEP1rUAMRe/ZKV
+lDNd/bkUmviiZ1ziF+nFjobU3Skw6M1sSSANoqHzc1Ib1epm6nfrwc5sBfKfpQl
kZLD1y+xRiXOl9BNNJ0vMAFhmThbNKnd6xZK+VZbuirvRsr0Du5DUMQ83zui8hfG
dzHvDJp+YcqTfazpgsjEsgq/3Dk7Nl5iDtyhqyhwT3dkC9udCc4Gwi/bKgRUQ4gB
riiNAPB2hQybnamV2AKXNwpDbAxeM5iM6M5ApHO0IUavSaGofLXCqXVntdqgAl1M
SS3bHP1s49c1PKzxFn4YqtkxwA946MYYJjz05RQL9HjWs+IYWUho1vBK02d6fZch
0wvxNoNrXWBayljF3LLUicPtm5BxAc5tw4EZA74EiooovI64FQHpJDnGDkNHmPux
Jc5+jvlRLp+QL+5EbpnRE00TDEhaWL6N+nriDlS+U550MACcG7/EKYZFJpM+F2kz
FPtQD62Lpp1eMQSS0Zjc5Qw0dS0kHb+CYKqhWkHQn5hXJSn8lXe995YuJra2U3LJ
08Ldug1uqSIsV9gFCAFSwfP0y7nAbuVEuAQLSaEq5p5eYLmWQrHQ1WsG0sMUZHyO
sDTgLrju7GeJHQmp/70rLRuPLWQ0iZnRen+BKcx6RTfS1MnfKEnIp3nXKHDXn62B
61At4EMeOCdvXTKO/bN9poIiNiHqAbnR8TSAfED0203+i7Z1FEhrRHPz23Vqgrk0
oi6bK7YvaJJxvurkJ5Muaia/VN3r300awxNFMg5rqnPCXZLqqJhzF6JhiQinmauj
dV6mmSJYGXEl49A7rUGJTZVrrb+PIxKrumhCBbd6a2fLYo436Np9RYXnngfF2K3m
Yi9XzEW7HC1eeHT5ZbRb+Lf9VrJJcR6QXJOlFft1tSlh68zBLlRk3EKVTSJmUdnZ
YiT/lo3v1PIQ2yBoWrRM5yomp+73cATF6ziVCU0G7Qgf97G2CdL3CPkb9WA4JSXV
OPiYUlo2/4K9CAAoNd9G11CMOXWvnb1/feITpkpm1ijbrNkPE2yLukFPhvDB7BCg
bo1shD5W4udT2lkEsWVhMJwGxz+jQzkBP3bCLZErGKGAobHzR4i+TnkCR29UtaLn
C05FuUUxdg9z2e6Sl6DfOr9QFBgqcxmNb0Oa1QwxSstDwl8hO9+76bGaRvOotKIs
bl0J4UQvDlyrUX0HMx/ct3WrUIKdhscL/SO75g05810rDLZLxxRvbc+4xVLQrHcL
B0/z3cLlDTiYpDn+Chqcoqgybc2+6lOz+0pYUJO7fa3aJ+9Kt+PoUWDLI4YVZvdJ
E/v67Ty7Ud8W06s7Lc6X+YV2ylQ0tU4/Cu26XPkvNHZeXjGVlRyEj15XcbUZmwHB
VEi30cNVzKLbnBEDLonjeQGE1KencOqLaa9XghwiRkaVZL3jKGvwLGhuPeoozOSI
jR7hc/SNMJKVjPmSvl/lNW8OQZx02LcdMhFzcv0LsWNRDUfm3fcVmDOkAb+zVX/e
SnJ9ncM2NFEipsLne4FgumekAZG91H14nL3F2tBrAh3jNn0lhD8oq1es/y033aW2
N5jFMmEpHZMCNOdehqLGFcgIioajXYe2fVp48NhxCsmKMAeYinz3T2toTCPU8Nwt
aSW1sp/rh76UzLGDI2+hNTE+QcbTj4OjcB7Sgxc5tU6xxHfJXbn197O9wk9OGzFC
ZF60HAnZc2DwqZvvqYQhfpCWcXf3yULZtpTDoevgOlbvC+yOvlwsuuiW7q4gh7+J
AdibWtfscS7xhQ0sHn64c2l6ENC1s5RgTtTI7ycfs8sG/eHmeOdz/HPd2eDnMsY+
DVcs05PdGntkr0oWs0zE73raMV/W5zyp4IlHAIy7bG+PktlBgfUYf+qE0QLxH6Q5
uRl/8zwAn0VIqiGbImV+a8PU35hmpg6l0GrQGhunCcqUQ+YqHVs2aHYFOWH1xsqX
H4hLKcDs9RXlKOEMP972f0+tBOyMKBMKwpSIHBUvyuX8Bd+GXmoJP9vp3tSxCbG5
5vpWuJk3bMqahrIEHT25kOXj4EHvtq+Q8ivfXDawSxrWYtcpP0crAmKZuKUxkNN2
oqTJ34uWcaPXmAm49i8QgfPGiUcAgWdchssaLIZGnlh3WHSZHvhgEgV1/6Fs+Lsb
ycbHpef+pFkAcx4OBi49CzSjfqdydUxvDjzmfuFdaTG5Qhjd25Cs+wkfAunhYu5a
YAAdvVKqmD2B18norswUwpazr1hyeOoul70EehtJBQXR9vEUo9VL3T/uVHabsKST
haqVvup1y5AwOmcAtXGMZhlRtRf+iJg4AG/qoJOF+613ncKxFTyzO57m4WdRREUY
twcLNZYQ0YIRLS+eoDglPTD2OEhFqUW7Ivs444M8i3GalnljeQVE69W2l0uDXsuc
82D96FhxSs+CHwCexCEhwz9+MC5aYmmAWrinpWRsiu5Gx18zUggORrmwg1khIrHw
RUZFpl7QXPDhTJ1SXiiSLSJ7GfXgC/ob7lr2HKXKIR2fw9R12TirVVtx+mEA4kdG
tKh0HmwN+GB/6GOoOurF8Qfk6q29u5jE4hLZ5+eUn42ZG6gH/CHjVjlnSxGTdl48
ITUefMgcfX29GtcDwkrZN2UhcaTFRzYO+N1WbeVo2mKoH7TEl6C/YnkntaoM5444
KCQDKEPkrbPHZlxGmVF35OZRke7Us5NdqbUyLqU8M5Z6l9prHnI4uQzQlXf17umL
l3bKjHeuIwnDWSl40zJ3WomkfktpxDiy/CSLhx0YHqdXpEMBw/TQnWPQht44OJT0
AdiizPrC0X5PZWr9V0hX8kXE5l+eoWXoeYV0sN/rDIzz+occNGp9n2QPTWyCl+RS
z+ZDsvRQP8GTWpMgT+a7wrEY6hPMYikR/xGnO9k5z520v9yaKSqGoACOGZYCPuvM
x42YXcOXB9LN9yWyX/MzCvVSpGLpD+DZSoI+Dmog3PGxe7yQ8w/VlgjkSJp2QIn1
TWIsMuInrFLWnw79EWiSUspMbpbbBJgeY0HRMaD5o4ZSP4vbsXZMbASA78sV089l
UoPT1Cu58VZXVUvZKuEy3aMzJC99sEzcx9mH8VXfPQ9pVziCC8gu3GbLGDFtMxM9
vaqCA+JOjVrt49j8cmXSIU8WgGqCtlHDfdy/gpy6x3VTSuYjToK9oklh78tlJLDe
Lwlx4ZpXHMCuKdAHnZW0H+R3J/f3idH4p/uGOOSClFPII877V1iHKKG26zN7TnJH
7Izf6v0n8i1mvuBRE4bZt4bSMtn149i50MlMJGS48Aeg6oxg+RylnPgdcHbSuIYe
v5vwdR2Xma08MWIx7sm7KWjuwEFlqeN1V5Rp0FM0j9wzXz9xcQcuq8md96dZXpb0
sZviwIrUqjNGx0apete4ka7r5USq3ywgK5m3dR+IcRgmEv8Xg6idCip3xebvw/V2
pA6PwFK1Ja4xtsECZKIH9PtcuLIU/wZZFS3mYf/Z1SF/5MjDBgEfcSa60WAFz4pk
IgN9FFXqrw4yHsS0MyBO8QD1+SFfz/o+hXqKTtfeLzwnH9ckULsLqoMnBqZomOFh
68os7qQG+7qfaMcLJIyG0H5szmkZZ+poPqznFzviEM6PQCm1csqmmC36K61tzv3j
dvfu5jBsE0I7pQPr1rfZyTzVJXwHEaFVaPoOyTNht66N7pycu6Y/q14IBz4vtVz+
5/7X9zACwTvW0y6lCx+VGW/BgEAxEbBO/nsUamuPhQ76PXBa1/x0zXetGVIHXDZR
/kCCKPiOaJpEis3/JAdBCknaLNci7FO/AVpGnNPzoLHSTeluqRryzDAF4uSEI00M
TaW4zW0vA+1LQVdT4KENHBIXEQ4toNpI0cON2vQp3HtKRldB/jA3vFFzm29gc83C
b4bVYR6sX+45B/VzmNUTwAyPxdaANb0T4rGrSpIgKJGil4Yd2727H2X2g0GJMU4W
WlmEV9oN0yQP/QY54mF1nO5nkQ+EDy1FV9wt/5N9ibjHBFkrK0idxKiDGjpPsCN3
DuDiV7aL6QVf+sQTEErylwur8pn1iIOKhaFa2qFhrhm7lGfzQDIS4Kuf1cpp/WSB
aS8mGmC4X7UwOlnmoguCIQ92UFVKz132Kejp9uRdo3Sbfx/BLzbItds3yf4wlc6h
KykxZgpr9nN6U6Hm6hrtkldy2ZJWJ1AUvveQmlxEiSB9sdLdH2gJBTzImDL4wCGJ
kxfO/rXUFtjiR+nlb4cs1c21mDnTJLbiaID0+bUPReJ9vJf2NHlugMtvZdiDf0OL
cJRve1P2RryI1Py54Kpuvo5tAp20bZdrigbOwUb5gVakUdDRLbfnUN/VWy//fxSB
pQyHnDjMX3mR99VUGfiAIYhBpLKTebt4HDHGbgsal6XKmNpBS9ebqnUWshP1h2Qw
OpwuYjPNbryIQcag0vpw8piY/PO/dZVgszI3mnXRLIuv7HyBv3HJpd3PlGHce4mT
4/HH2uV//b1VJj6HV0LyuWcNC4tiAhVcqhyWSokiTAOvS5Dk1ReLDRQ/hoak2akQ
4zAGuHPM8jNcWwBKbVheufaY5dcDHHkRqq+QAvLemLzOdE39mMdxD0iEYgLwBHNu
l/xs/IhP/xqFj/GfYz4u+Uxyx5NKA2TyauEM9+9vF3MUJ6qSQ4RpXKs51R8XkyTM
TVGOuEurDOZsCLFx74dDuSZMMGHdymPlBmfN975lq+f6t0WfeeuRPzlb4Z1mjp1L
4l84pX7s7WrzRlDvtJbbsfrxo1gjGMmrZHI5sOZmts9Vy5E0czrluvqvZXin7in4
dmbzdmYa8MVkA/p5z3S69Yq/LjcE74pjBvHk4Eudb/HVsTUUvu3sEpakuMbkHKy9
rjlkl0p6ZMxtz8NNUUzVYKg0cztd8kQNby4cxTdmFc1dyZ6dmdy8KvCyQyfShjii
+pSeVCJk8poVXLGgD+uwOc3ljfIaSA4zGBU5uEsCS3uMqSCmHjlmYSBFVgwc0Sdf
+3f1kXS5gVIcekHdvL/3mRBdrFfPPsx/UP8/nhdWyHXrCF8eKqFLuqWyiH5UFSKE
YQtVTHBP3AvD2GIfySU+LzgamXLVmrx1umpDCl3pKfbY5u8fruVr4U7kWbgCcVyv
y4zyLLvvgWHSov2yswhdOySDcjs/eeWGCBZcABEuLlA4k12w/5Uslg+nyOpk4tTa
N6HDGwTrAj77x7Xo+/Tbi6N+98iFTmSvro8w5hE8A/i5SZPgBT07ojLe+QoNoG+q
FwGLm8/qI13LtNY5wwT8gSb3RskeGYEpJs1kgcgx7bVmlawJ87DKvjjLI7DcyFOR
ckhubq6nci2kwG0qdVE0ARGLHBpZ5B+F8YjH48VZcomugqVywh5FwIPi6lk4tNCp
6Ed+RFTg8/1lEHnzvGylmx1f9rhQG8zmVaEoETOk1yzTDyz7RgtBr0FV4n6Lxis6
HTvHkl0R03+NudEHvUcuP02wUZmpBhBpQO4ZzPN7xSchxfFtdaUlrPAqera7I7HP
PTFWN6is32nQ4gDWzaDDvzDSc9ad67VkHrHjwjoauvexk51kfW99eYYeotXdOS+W
hLb/sh48QRBct0FNBNGfbOURIKzdeoUuYagNjJGkP5hnzx8a2ACpNgjwTgNa6Pdz
OvrPW7Oh3TYjnvAlreIdbVy1d5QtuuzgIvd9I4bpFuVlqsWCwE0DrpDAPLu0VbfZ
Z/zjwikcLv9u1+yQQpKAkZ4TE+eo2dK+RZu4ebRPsbMuYvBxqC0K5DNtzngfgnLv
N7jIFVJH0aYNkOdOrEwBc8p0Hp4OY0jJJ2OwC64IBVICa52EMjlRQq/jR0BLK9Ew
HEtKOJCnRViI4ndr/tIrlG/ABmf6XYd42QfEexK9LcJtj4yOwFkwOCGtlTOKbAEZ
56GxpxyLrE1kWd9OT70J1iaX4LHSlcc1NWu4QtwHoEX/AUPye28RtMHxG2i2UZQO
0FJNTGM1SMnVThkzhpcvZXv8u4onPAjqDENfzs9m67QdPRXKPShlvUrVysMiki33
ASMjS8FGr+Gr/1qor4rsOsignot2SZ57pUl8u0BiK/pxApiAGsGPNavWPVBztulJ
3J1t95kQexohkkdsaQoeA6j13MrFCK0LgsTZOlevs36LxSC84umCDGWnV0egy5bW
GRhlYnBti2ZkrDWpUiCud4+v/NR9gJpdy1rtkAouiW/P/2LaMI57uTDm7vHQhUdh
34l7I/lFYBMqxWfUOHc9b6+AOPKheEZ0BfgTpyoFvJDFMUzU7ifGBu8+L2jxkBfR
9QAGkXvlRu6Mts9ggILnjzUdiMu5iB3WFezHsKGzLb/wL2T/rd/DA/qW4eXlTG9j
UECjItubMLPhN/og+7pJPpAhu19wqw6Gf4jLGEL0Ed2ppznfyVKd+0K8Mkktnf9N
g2ZUz0S5e2DPHRspsksAfsJ/YgHqw34gfjP6ZEkFgBBYDiOxI09HESC67ZAM2QDq
5J0l7w51XRJD7+IFPmAgSE/tftqSUrbgGQDxSsjj/KmrQJFV02mAvIMsVtCitDgK
eY/0p+/P5lZSPCNly7QTwEon3OgqzEu2tNslteA7WscNMOzLAOgU3CeapbeYoA+o
3Joyt2YZOLO9K6fZTpv5iJXwdjM5nBlpZCqODt5nEVNAt3UDIR0CMDQDc/t9FvhF
VIfb3RP27lGLyBG/4zl430/y/Ds1+Mt531poEv7YejpDxvud6u+/WqBge9a2qTfa
FsA2QFIzanSZLw+06ot17C78EbQCCVcO9LWrVy0Y12N+dNGVWJOyV2UWmGENset+
+Pc8fOw6lF1WH/BB3twn14h5EiWPVP4Mck6NW0ew7+Uw2eI/OcJuLuSyffUn4ZYB
F6UvkSXLdrZ0X7WQ4BA2ZaGXSzzQL+ABTXtbl7jLTIQ+uf3uKvyFto0oX3ZqZna+
uzgB7hqi3xAVrDHg5mC8yV7+Tc5HNZhl2dZLYYfgm5uUIlLup2F27Ilpbth7Y2jh
cyRaud+jUU2+XhlROtwXeCTQ6nZx1l5nDrXmUDzy9Zu7BRqQP5j2AS60zl59QbfB
iJQ0NGlMjAg22B+bV+sGEIMzGz+eY4j9TuMiO4Fyrlv8haE06Tjea9WCol28X8CB
rNixuOE2FmUK3h3MKbG0u1dHAeapubMaTlEALuCniIKISZmtZPGT1jVGf/4SC2JS
L+WH5wk2i+FGpDQBHPBY632Y9R64KfCo74Ai3j2l/fxARifHed+YVofjoUE2VErq
PIyqSLIlruXBubpSu5u9U1tXkemo9mhWSStKRQOC3IFYim2X5Md3b6hiZhKAth2V
TF16htxTbZhTsASzx7D5s6DbB+SOX3N4MhMAOwaoZJA2ayiaUBhOL75OGUnr2IIn
VzFN8Vxuj66ZlZgbs3gYSR9UIB2o+Pao8QPAkDs/2BH7L2eDu3jMkqIZfMlx7yvB
FUWNpIVtoy3daxqNDdm+gezwv0062Wo2zLGjvYNrtMHpfYIW17GrAerXSSExPq6E
oBhp+sk2wQ64uEk6qZONcYPs6RZ94dKaQN96h6EhZHg4aF9zxvt4aF+uFPY6GoRu
raALvmR9W2QqFMly1QTEeENKcy791K92fPIvArWg+PmnQ/hj5EZU9FuSBDgDWBZv
wQ24JkZKEwwpWuwpl6JGhqPVxh7z8LEvgm2S5j/Zke9gtiglJVMnrEH1rltbvqhV
guGvSr4oK6FMmtfkEGE4c1+fpcgO4LPQD9xsRFuPZKnHvnNnaXs+8TMDMr0B/Cda
lofWPqVabYE7Y9oETxOhlIjDuTL6fEGw10l6gEFeAE3hGbWTNjYbkiBHyOJ44n/v
TNr5B+fII3X5ZBFc7VOeUoS2jhwMn2bjnWjh4F9k8Do7dUCEI/DS5TCcHTtAqXRO
/x/c3rbmZuu5ydy978A/KoEoj88rtCVl5nkNZEGWhsvertBFTS3EToniPg+qobbj
7mQgrCFYcVi52dQAMrYKeYNc/3+KYL85Wme46KaXb/3ot1AEkIXcggsMD/VYzarC
J0Mk4dx9wTXbbkSiyy0k6oGQK0mm+mPUdt3mN34US1Ya4ADjg0esrES3feO3UKIx
a8QRCo/GM7lSDCGqGXbu5heW9DmZTKrQSWPt7c4U/s6JJPG1EmD9QBhFgmHMQ2Fg
81mNbKFHCCowA66NIQw6K38X05ZwsBfHa8BPYZfQPM45Z2rBaA/hisJkCTlO9xLG
OvaYvqIqVfj1z1PxBN37HgSC9c/+yZNK40TJYwQyhsP4sXwNzJnmMWVHqK06kGdx
7kaTrYj3OYfu5mzxfNCPalFLJ/PbxRDDg+TlGk1lGo4Qq+sJJdyQg8//dkO0/J0e
AFI6N67EmTUnRAiwC0N/xF4YaeUqgeK3w5EetGdYNb0QXkti+bDowJpuSXAo8vAT
d7/O1w07ECCVCGT7mG1SQ3FqMcEOw0izVMhgdK72A2XQvfVP5rydlSFjWRSCFArk
frE9gTXtGkX2A2XcRhJ+wkDHDasbKg4JF1uHxhjd5JpHtS/8DbNFPpaD9MPntiS3
3FlodAZxh7ZrsmeGLzFZL58UDWr2I5rpJS+z6ICdazHw1QxY8u7+oiqRinTthbYs
ehRLb8pMgG5gHqKEQqdIE7hIySd6liu7BEmLuFPjqOA6jeeSehTSD/ikeirBiuXY
qCT/F6eC5+prz//Okk6JqSIIbxdjdKVhN9cJRNHFS/AuZVY4ycB3KEhUCDgKQADS
rCpaZInOI/ycQcduA3xTTrGX5qz3TKPKGmLVL475iPcpeIiZpvb9jtgXgg6KRChz
grBPYvz9/BYH4+18hNHLr/buf8k1iADa5y87Yjug7nQgVrIiPRH53l9tEF4U56jb
BG6//eShiwpy7AkZzhjqvsaPxqVfNHQMkKZ//Hm7ZLVWnQrCFNOkV33IB/6/ycI8
N5EeBG9LsMf6DPljA4dRUoVyE5o/m6+C61qxgrTFrQnO+/K/KVzacMtgbR+QGp55
dAmzCluqkm3RGsV684JfoCYZvtX3uPOtFVbI8xzi+wNEQ9zSWEyATbGsOyVb+aac
xLmqT1mC4h76VAKHE4qskRl3ocwJsEoNx9gCN/LnwZ/Wp/WaAAj5I08ghRIAvnpP
UlhkBVdyJW8P0on0dtCT5EdhNlC6EGM+w+Ce61O3ZH2yzffsbbTJhY66VlR0fGqR
J97AP18SEWNH9+4gyhTiUf6UpXWpqtAZpA5J6YZ2nnGWG4cr8dmFrtop+8HFbtnc
FV+uDjoDhATLkpMa4yvmdUp1AkI7B6uA2U1mDqiWwBIQEnlXH8wnHPe2LvJbDNgU
jEhVwHYqL7uveww0jcst7gzQ62ypwmLiJ2h7KuE0Eu2OmNVJqIpXBsF4gGguzi8s
opnN3KXDTqejtP7pDaOd1UyjN7Hp7/SCwdaFejrU8CLmScLgxgW2Mo3FPXBPrXKM
i1U3mPo9JzNqauChO426VPF6FSagbJx7P7BYBhwMc7ivo2uZ07H9roAa+UC0oEpd
cmUWLdhO120GDNDtHWv8hAA65vygGHZaCZkqGx9yrtFvnzHq+LleARN/UtY89hVm
6MlDgvC6x4u6jX2nM85T8jtPpfVbmtff5B+sEfujSeDSD811pXfJcEG3duwALIgn
isuJ+7bTW4NL+wLLmalh0vYqFAahdlIzpR02sdM+/wx+RTF7283Ky0+WQubiFIBE
TF6mKyOcYJwP4qzgnILiemSD+vxbj9fgYTqDIpUWQX5h4MnYJU/ETFtoW44ii7kt
gt/bVSrf/GH/yu+FRIDD3YjiSY1cfsEv8BV5BXxj6RCHPesbEGHNSIHtu1F/b+xi
oC9UYEvzioJqVzUaI6mbvNB5XWdfGtsSvjzI4IJv4cdDqi/Gpt4fwgrHevcWuMQE
MZLppzs4OK1LvK3KzQQpgAl/htX7+IB5PXHMOAEt+kavXEWF5Z7mkztqNS/ARtQI
fJg/QmKeURMG3k1N5Y282YDk7nWJZHfblF22I09DhjmligwJE4xXPHpiQgUJzKVk
2PVMiXogFjdjzApFeJRy4vyBLGJap0+lmiWMODfy4y8jj3yNp92jXLKqgts+5+rw
WNv8L9rJoMPaWKGrRQIUmdgxP5BGkQWYJogKevIW1IoruQt003GYsgB5DMYd9B1X
B6tMz1G3y4fXBBd/kTq2gvSdlnMvDzBXlzDGtGjac0UJXr/FbWBIX5FgQaz0V9nn
zEoEibhd2T2xwoo6VwHE1RMngVEqM7ko1kSVBQKXx2Ofgz8F+xoutjpdjacFOlmh
KYxR15+hRy07iAdjniWcAniIRxKefndBQfH7SlJA1kL/iq9u8q9FezJJg4J1cqTK
OLwNsEJsPTxDx5zLgaYqopBek9e4G3ybCwkkngqzm+PVIq6wTsrH70b/R2QpQBIQ
nfEtBh9Xhf1MzqT/FnIr/KbGM7Wp1rJgfHPsJRfSGFmB0DDADJ7Po00zs4qPafVU
ZDZlOcP+pp8NgVhYDs2pjO1BcnsCg0ZYQ9hNWY8LGPq2luDN0sa7XOCNB52jHnHQ
/hyEZx+PqZnR2Jq+Dwc/a8g/6ox+EQs+kaO1NSMMORC6/BKy2PqhfcvUN9DSm4Hf
TaD+lQ/6DzLrrV64HUQaK48ogEokcM0MtTIk/klcf+5huBLdZEfrrueQevosRRYY
Iy08dkwzUm2NUYpErP9qYxnBtkSEVXXTCzHj9m4GI94RnHKmlMf3jYZppM37Lrop
YSFxsuA68FOFSKnjsKquOLBPW9yn02nZ8A8rpflRR2VMWdjiIkrAhBXXtUuGL1kf
R18Dxx/Sbijnr0R9EJcTvqsAh5syULAPjsi7fSP3BfFzq1dESTU87vKPwjPC+rWs
l5GghtyauqEeFtRs4t/EUxlNgpR/sIaBbLkJz4RN3WTSb1laK75aliNxZSGqrO+t
gqwhkJh8MkvkCWje4w25+TCzS0FFOr8dzIavWz+HObwxmmiXvCEu7pO6LBptVbU5
zVZqsxf0jwSiUbAWmz6X19jQ+rh5gZ251Xmuei+3F57nwv4lqXqFA7/0nsLF80fD
Py9kpSSDRVr4X5elszmoK0SOJOB0dZaBZIfjrB7YIfrFetoJIF+wNihsq5gO4HmL
UJdOhFqBRYYUHM6iA+M4qmuhownoUQ5Eby/QWi3JIsRLypU70As9MgDcD4XTAp2/
1IZ2bFby+tBYV/RupNMRmaJa+o9tCJx7c7V8QTRXJ5XS9/hBYuG8jUkjowEoxykX
dnsArW+rwSvPT03jc8/xLYUACz+KXcrA56UuSZZhN4kiKJGgrepbYMywOaVSW7Tg
QfWvuwmbqMRLNqJR2OhTQSdQ1F5ZPq6HirDa8+z9JGh9dB2wCGhWmgbCvkMDV/D2
G6RwJ7zFTYBA4fbPkg/z24k4Q1UsD5yZyplqhaAN/cCsaLW+yv4bgNsPgmzQJRPw
GcwGNO8e57DxI4QD/H0J2XbGhXO78Kia7vFLCJ3wMjGfm/fH5eLWsyVQveykozaz
zHPmkqFhB+Qv/MfBycTa59JA0qddDOIpRNmUx9N1ieHF5GTm+7XsgNsDW6Yr2o25
TeUwj6l/5PyBHjpc4UVUG10o/W32oR7GcwWdIEwDGYWeyDegWpoEgBwsFymz9sxI
N49rFiRyR9Ff61h/46f2UIiwys62FbuNkuYw5LohJSWflG1KtbuI7yjntCp9mWqn
nQ3M9wW+qxgWLnkRu8O3pZ1NJ0X0kR6brA0EWam4IeguWpqFZ6TM50H/xRmmU7SJ
WvJQREFRUNDQ71vW5VRbJvRR11ZcVKAvALBXLUFsSIm3Vno81s8U13aFNhHycclF
3G+pMZzQta7nYwnRVXnq3u0E7YHWXdlVk4+eFLeBE9tMjIS/nOhQhfo3WnlZDYR2
hU7xOlyXFpHYM2+Jr3a0R1GzVyg7Y3RBG9DOmVQbLlJDS3CF1/ssEm6fYPu9Ke7y
r9OKZJCFOxbO0oNql6JJbxUhBOEMu5Y4ay9Gn9p3hBtAUHJ07hfCmq6MCINMO6SW
3rdhioyejUDKGlUXw2b0/Mg1t4RONdXKRohkLwAI+se1xw9RDNdZNPr76IAxFbsu
gxXHxU+Ra0J9pSY8HuygevP2gA45NxikOu8sxOD1sDlqOlIO4wdcoG7OtgJSrCnl
vxz+6lgaW8ekjPjg992VdtSwZK7/V2ijjPTFb9JVCGanbRiGbYacalvC35qJ9hE4
49Qtp1LPz4ZFFpWWvuFeIm1G9fjO6wuEMPrJls9xiNeBQTdLyVswXyR2seQlVIeA
kJhc2kGKcRt1R+rScID4Luzhcuzj9SeawLtEMgBwb9E068ZzZESSYk2T1q73um9h
N0ky7ql1FYNMI6ONLLZEbxeKYImT+dVC+RoNyWG9/4GUSmRYJcnnqv0VGaNk9jcy
2c5peRHvZaeJeXk5ipQAWKKYeBDda8Qx9G+8mfhN4z8vbUdTQ5s3EWNGgjXlK8oh
2A71+y19rMWB0rjgVTWUh6tEqRh5RisvxZRELQT4V2880o+bAUNkwn/U0KJCtGhh
7vhyACsi6qe31S+xXfncSMItUOmtO0QYJCyZCK+alRJ61oiOTXuwx7A9L56RrveX
YB8AVY5HmliJjGkazek+bhbbeIvqqDcNpONwy43VGqp6kD5XqndfuLWxLUjxBnEg
pzHoKJQVmg1uYZXSq36T2NFbpHSyouh2+sb327ErVjJh3f2tfMgq1/tL5I51NwHx
7s9guA4FDP2pDllLOF46DIpCMBF7vBiPT6zb9Y9Eb1GcTzl+dkneTJraZpziHKD0
VUx193GNCaSJ929kU2b++e1PV0Q8p2mXABl3Nytlu8i8VYaCj7ZqsIo7OOzyL5A9
dIg1Sl8ldMAVV/G2UoI/MUaNQQxhIbtcSaLsjBYiWBAzv25CmmkQwKQdda+Xrtyy
4PhrzBuhejEOgO9+gxWrF2uJONiinFsGLxDejvELACVKXZRUGhhl1g8RJYT7Udk6
Ui/dNH8zDfF5+Gs8onkcfdaY9yDKQ64fVmZ5tqwRiOAnDe0APjGuaoOJ69rcyeMN
kXvsk1CbNqjkEl2SZpZF+6ks8fyGpHfKf3fvc5ro+W/og/Z1hkybe55RjUrWoNwB
tEJThCUv6qgfkdYJ9KuTxz+IghJ3J5Vs6BD3CRA9Ha/+FXB34b70LRURByQL+bs2
eNVLRZlmG5ogr5SvZR7XoRSqa70BrdNW4PBx5AQvK/SmsjJsOuDrBPUfNGCQg/fd
S6NZGcPxzXfUKPXA5ZBbyFPI3vfW/UzH3VzCEAl+ZBT9lZVYhVySqjNbB4WuHCmz
msIrGnTYYtA3G6XiFoEqfan72XwONCZrgX/dSsszWmCaxSO20Y40Va6RqNOLRJ7K
7qrqKahH2CRgqh8Qw8Rb4yiDuQ43DPRqs0KxvUzfqTMuwUW2Ckz+9vgc3D1rGRwO
EUXvJLL+qATyoeib+P3ButNGqzUgMqRnKgYcy301LX+EnUzvqQi7G+KQOxayB4nr
/dVbB42qFWc34e5ye01pyM9NzZClwVs1X6HSK6ZLBwoFMoPFVjPndZ6GFF3dRwRG
My4k0tSMVW9itDuwNTcU+p3LAMm9M2SO3K8tYkpCIKVisDf79OI1U6VGav9mIbfB
Vnv3ZxCH9SMZoQQk7zSZiIIGceLWcFuVgBoZl0EMtSRkZkTEVvNGukV9HsCvd3/g
AnV/rEplAGv5ymhkb6YqKYs2sGEguxLxOcFW43Aih/rLpBv3AtSE/eAEdN0SfauR
WkpBkbiRDxX+mXvUo0M/iI8QA72cDnZYIwahybQmNocrmm3Bl2zrwwf1b2U1l2d/
0HR8XgZNiGWl/BqhZzGR4jHqG5FydV6HFsQIc/aA9VRyMOPaROnhMvgIBbz5/nwc
FyYE1VCFsfFx9e1XI9eMhET9r8iYK0FrGOt2BMmpnXFrFvGTnhu1oQd8PcrqKnCn
ls7MASX9m+4Hx/KVaC/kUvfKcnDw+scDcJeE51u48R9MwBkrzfU44ipqVR3a6i22
0WSCgPxsGeaR1Bj7vh+BLvihKYSZ287tqhiqoEz1ExWM46smyiDB2ZErjYyLRK5b
DxAsCeAwYXa4YW6kzPQLWbfgRKVYcL6tdrcgXYdmurGKAO/F8CEgjgDQGim2aOi4
GFy/3gjMRU6cCbDb+az+tc4S8oPTEYP1zBTEd+LHYDef3ryWDRYSb+UKsy06ifHN
IGqTomRW3esGtfBq5cO8WGbkkv98/i1y+jQSQM5H4BUoayfU2XOI9Y1Oc330chqj
yieKLbeU2n7y4HijcAKR/PSOQU5wIr6qMxXlF1IVGn0El3zEM9lGsc0thUWufhWT
VRUn/0GFAbgmCQzsXHUI2P46G1xqvtFE2NpVV8oCA61yLWLhmj9PK/nLXDO3LdAd
tYf50P+uD9wo0eoOEeTBMvOks3vWLfsh8EYdTNZHxXvWAr8cYwLlmI3t+d4xH+L4
XdqyRiVtS9C/nzzikl0wzBMzog2JVJZA4APwTSF3+knq5zumI9JQKkQuaSxwpj/Q
0GAizt6T+btjlWT7cToWk+l0cfZzZQtXf2PkRazimZg9s9iHp0LWiWKTXTAyNlay
gTSNXGq+5oVBnlLSLwlYMkeZAp/8g75RlNS6g35q5Mt0otoiUGF9NLIanKi7jLsx
LHzVOBBtJ3zNvVMPkaXz4bbUnhr6Zkuvb/IKK4GCALaeoWGfiAzeRn+3OujhWFZK
pMaxaGszuvGm3XYcc30bRvrmmrr3Hqg3B22RWlZN8wqA2EIBlnUPtACIen8iteD0
T+sbF3a4nLoSC8LGmGIK7XGHICUyIlF9uRF7CcwFBHX25KjEkLBdm2+wCcuxFfS4
/TU8cgKqJmZXnzY/3ofUgn/khm34z7b8zViOGoIYfFVXLr5yz6KcaCPKUl/UkRId
KZ8Uiiin+niHMBoTgO6aaZ9jwn2nKGEXtsO4/oynUYvcW6NZMRtoksjhDLQaRIYe
+jnPh6FbbsiLVdiU/BMAU6R854Y1we6ZDUSJT6530PvbQAxM09HliBdu8gRSG4VC
8auZ73eryWoGBV4SYnHygpZnd1KBc5HZSi5Lt6Aaj9X6kjp64HsITGHB8bTdpNZU
5O/Lx9Q50t7+dCwpqPGKiTzVa0z9EiAdhEcbUrPK+mb2caC9blLqmIrFkCRl+LC9
rlPwrj7kpu7Y8HYcI+V1yMde26EuneLuDTzsSfmdg+7A8+QHzVbVNE2/x7BtRhZg
11DVGmHoOr4eOYE5X9JnINrsCJ4HJDKWXaDYadCX77K2ngADVWM5wb4MHMKHVUWk
nApcdBcjucdcKM/4SHoBxWJg5G6ybeFSNgcV4/6flPtCKtIHMuJt9nZBHrVPzUGT
aTz1iPFmQ7C9LsIeCdOHoHiGrQl9a1dVJgDUxBnzMCzBO2gcGtDGyK3hDCxzD77g
RXxVKxzSS0oyXTz+kRUYwsv0FVOzrh+8+dr/DFXP2V2K4IfuElTW2em/ztzYwuN/
07pE9BdGlh29LFzxxevxQn+1kbQ69h0vacJNHLet3sEC1bc0RpdQH66nnGYT6ArR
l3m0L8ai6QD+vnanPnaC25i31SatK3C9xSRNBaOkVmDj5Rw40OMNGQBUzma/V/7J
V3lUSXmNPLVmHvfvY+937XJ+G+yDxHxAC0f0ALa+/SIi/ukKCl9ForJutHweh4OL
Uz8rGsiBHLyX0g0/ucf0vgok/16dJqPuU0Bkm7qyc1jBQbiH89AxC3x4H6K3Tf3j
16CSj8X1ohqsnnsB1fa8qXhK0PYKgtLLH/1UL90zV8/3TTB/ZUX9yzNB7NCD3DsN
p5NRr9MOMoowq8009sspYInUnxgMWpykm1E3NgvR2IDhZSLjLM1JLWALyFi5eoJf
W8jsU4y/gG8qttRRfAKBhr9TvFSnjOyjfbC5s/E/92D3IYV8M038oyj25rho6kgU
nLt5mbr+OFE5BJxIIm/Kbw5cpmLSV/ROQJ2Q/UpfgTjjSjtJX2GQ8dY1MY3h5Vwi
tJLp5BBALnBaAfXd9TnYTjL0OPpvXPKsCcRfLPyeRDfqnVXzh7Z3OjMhsbOoQjz9
5bpM05TRldwsjhyTkj/a6ngfl4kKUByTGqtmmVloRQ4Xpmj0yKmXEPZe75e7Nryt
BYUZF/3egD+Hah5nlX3hLs0JLtNoR8EP7G0r0wF4fMjfn8pXdKJnIJ4ZB0D1N21l
O0NyRNXChOqu3rsWsqrbB36wpSpYfESCyLvEzJmNDJSk8AScUoOGPkY8wV7GiHJ+
tRv9UrnyFP0F/ajCJx8HmtEwDkEWwq7NFxJgYaRmmXV37Zpi3U9oy7Avy7Qztn+l
idleX4yCe23as3HaVWy/H7TPwWs0c0R+O6ATf3HLkeVUn/cUhJT2yonPpWAjGhBn
aXANF3Qx5Rq1hMDylAUyEzdQrmQTtiScKIZdMZKX38m1p14L0kcXhW5oRbRL37Qf
a2GUN/l+VktWUTnMoUJxdApar9IHhvP2MB607wJvoFPFim7JagpzMjVZIaAQPY/e
tr8YQqn9uhoPxU/+VGCzUVrve8K4dpxvwuuJ1U4FPU9iDsA8OtosRDktu1g12g+N
e4omIuAYAErxOyV9xrF32IDMQk7DmSiWx2/YPM4ai31fGYLAhxItVtasZ4f+caCr
txri/OxAwKxMAFMow1mWEnyUIdpApBCxkjtrPWxWaEhQ3CLyHD4UBUycVC3cEoH2
+Jkc+jSsNW3/gIqmAaLZ6RS2MMvejvoSI9wF4aZ97rnVt0/3gmMq/hsUcYGy+wL5
gKyIGuqwmNEyl1x7wxmwzjfFtDaHGMvcZsBSXVslGyCMNiJfiDkSASw473Tr0ZKW
rggBpKrMejQ+U3Fx6XS/bz4Dtg6HW/zZLLg9Wq51Dt6uWBulbU+cXihuK8NP3U+t
ERqTGKx6bSLl1JOqx6ajtwrTewFkkUC1lB6g42YfU9GKXwibIHwlyILM79eLItDH
FhPwV+TFjapPrARB+B92DfmLr/QyMSDF6MyJr60OWK8fG7s3PxOeTPhYcsZ2/Y4r
rNYC79hLKhzwzLL+w4DqPMdCZb8ms89sypdKQ14gK2ik0aXuqcdNV20ZCrI4ZFpO
K84YH5KyK32tGvXRGrMu4zz09pqm5rB2mjKy5Q+Wet89AwJmyx2mde8Y9DpWAGq6
iZIN7KrfBejwjOvaRnV6BuFaL+KwXIY5VPBazJ9CIzUPlmlw58imXXnwjMzLG3xt
1HKuKZFa29+owo8Wl89lszDeh45t2ErOOEl2cCFvFqoQxB76OZWfCv4HGnYnyPyh
D8Zdtx5N6EWT40LsYbeZquVxDwjdCf9FTnzvoHtrsDXFcEo2NGHuxsPwrLCdQC0+
SXdQqSwM0MjLPIMSs33CGnYEmtnYGNU2r0bV1Lg16gxBG6RzHNnLw/3nQzpeU1vo
IzcniXV507x109ZiReiuGsMTbcyy8SlvqysKjdILSKBuaLO8ro57FZ4KF5ANwoot
11s9EExQij9p0577lwQmY3Wh/1WS7k4C7SEE6599wfXDMM+Hd98rnNPfNpG34oEB
lFeI6/o7ZZzI7L4nbvyOUbQaZYYlf3ZdiaOAgYFrujCxmDqWwyI3gK3SmgEdUmHU
S/63ht5amGakXyqx7W2Rkn7Uz9aybLp2cNZSG+d1oFXDVICDT+g0T9I2AYHuwXI2
I5jeasD+MyEs/cuhgb6ol3wxo0s3JqT1IzgkfbxnaHq9bAm4Svsoe5v5+vdX1Ms8
dFn5/YV6I8arbpcGr/5zltqZcI8R5R0AjzWFGIJBmJtBXWK5gj33p+HSE//uPmBs
eHtwjeCG5SCrY+GQa15hURPXmZbT9NXV+RdQVV2NWXR6OpbM1oP2YDVHkIUGVuny
PcgMXU4SNiaTj6OFrTy7WxFE8ODd63e0wjpIku5CJoe55efqb9rENnjo4wsEeX/c
+ZuGNQn2dViFAymeBsIn0Kb/FMlyErNERJjG7fN7hGkKKFDU6w33asMmiWoySeGx
gR7is50H4VI8BTsQ79tunODU7G6U8AXTVxITKg0/9PM8lnUebLDICTLkcmjEuE6C
kZKeGaJ3KDRgVy5iyuE+EjinrIAYaoX5dkjQhtUUT/oAK7T0gR8B2Ki2CT4fgyQj
k8azCCh0er/hHnZYYMa1tsiKwSYuVnp2cKeMtETzSk3PGCju0vxf2DBS7OZasYb4
OJbRfcs6JRpsN7AQ4iJ2cDMrfOTzehtDQqMILr3oow+WYFqz6g7wJfer3pAylb3z
QNEdSvUchasevKFX9+z3UDBtPFZXGAluUGs4Kt0MZ5YPM7tF8DslW1nOPBtv5uv1
IItfSvyKjtRF1jzYiC7ZZ9MjLsxL86oxKQu8DMq+581iKjRflup/JzaAextu6BHe
ynb+wjYMvd+R1dipb/ZCgxtlCKkz74HGVwlrpIa6oG9bJFVBCqG8IrYwJ3k1+V5/
6VQ7Y6dFKOrQsPKL/3bJwQXTiLYfX1AeWvAaNM9aauXLAOrsaWv4QiluP5CGHz10
UqvkiuH/oVv6JN0FNe6l9aSAC4uanyGgoBssbUuwmQ+tsWKh0b6JdTGReYw7seeV
S8fCxNvnaJHqpbk690YZbe6aSZZdvDNnZpomQP/fde2K0iPkw4KDiESR5vXghkwS
nfpermgbLDHqig7OPPIdFIFtZ7Kv3SS0xZnagAt2vzOeibRRhYIVLPNUw2WPxd9m
UfHYxgafJKCO/+C6Qr2PB6g6XPrjraUCDt0VpI9UK6lQmJodkh7RSO52l5XokPrG
jzGPrm7LU7xkX8wtoDuJoR0ZqZsmqnJHc9ssPT1n6dMDS/K63rMP12sqxfYkcT6/
1yQwzQVKdV8AIZ5mwJTLfSB/tx13uyivMbPZBlKcXXu1+Hdl3nQC92yOroqcYN3D
qrE4R3hc7O4a197j1Og/rJysyzLUGC/rq3uM1n5pIPnVNEeMpF2QycBSDbhwTgPd
1u2P6hA9CDRgglGHmVKcMPlrOCaD/ppiSW2AAasAEfeCGxwpP1lRF9tfhaT9wHes
ZyADVtztm7zTSz9CK1GZ/tD8xV97UKljhAZ3FnjWorUjm93pD4g4bcLxZ9N5vokb
BMmjq8AFXJUtSlBc6NPTwrbIfO93FRHPerEIsttN2JUk7A0h366pShOiq7wRR/1Y
osjrlQK0dLSu3TjJU9n2EZWazT2c0Hbt4wxo4qvtasUQZp1x9b1sJ2P9pDL/lzdu
+aoCw/WCrBhSDzDbK+pUtWOoljMzFBceKlWbYiZwWCDCMihlOYWFr9zRqzdWKUcJ
QhNCYyOhZ3a0z+fYEDFHx/+N7HQ3P/2ZiTmf+FlmiJpECL1biFbnsSj2ZJAcOzmp
tZo054OQtmPC09TcZdXLIrRaqi4PbBurUAiTe5EckPEeoF+5t/ONQwaRcthXz2Rr
c4iiYQ3XMA/4d1n9Ayb+E1WivD+zp5TArziuz7XWUHvmYiDpuz3OTAWk84FZQZjl
r/uSzh6P/zqPTZiKvuU0ytctwd/ymMXb9kFdwiXGigzhfUjYRF0mK+cZFBtl+12b
20cWQH+njAa68J1/5VsHZskY5B3rsIqHIv6PrGNJl/9Jv4oHr/VzqyofahMRl7Iw
ZtbcrVZlP6iUDEFmpWl3Vs9rJCLUEiV/DbwFSzu6jHICqvQe9KTH7YBhobwOl1GV
wVBNYvQeaRvXGN66Iwd53bNjpHXM3IM+YJqeALYaX5vTQHF1KsztidExC3wsqObj
/PXowBw04pWGPl4gmL9BMNX1lPkLC2ltWRdZF4C2Ic78nBd1h9txk3v9zqj694fh
4/oDGwTaPg/k5ce9omL3bSsCIPGspjS1A+LbOWGS+Wad+SDrfhBBI6ACQLdUjQ+e
prFEP4nGCqK7YMiqiWhOrZAgJanuDrOqZyL/Vmm+IDyBNRRTFvQM6HpcCFDEQbx+
jq5JTFXavU1qr4OpvDFFAZPE5Kr/3jeViuLMSrWyPMDX/cskJlE9fjpr2AIF2W0j
wzDXrQrOZWxg8pQFROoVRivQmfr2xFoFrjvCGe2FMpcNM2frGP2qnP2P2M/lezJL
O1Mw3sCxckQVVOPgh4spfmMUrQ0/QrwvI7bJ8yTrSbQx3xrw1lOTKUYp8H+LQmz6
VI/Sjw2kXuQrFBlf1Hd9wFzc/V86B6qCIG/SDzNDtW/YBUITnZekfrXYX/W95o1V
OgScgVhpPMotOL1rwMR9rUUrP4eRKRY9xK7HOAF6dRAb3RGrb6QStC19jKLVQD97
bY+1cw+9i3BKr2m9S3PrRA914SjXdaH+dff2R8ac0MNIaYaoWWpPGwH3sPnfsNMt
j1rGtz/a2VwcmIp8p7JvEOjwGyzBTzxjLRh1qNQQM74AeqR5SJOBxKkZ2AKWc4Pt
YWkKnZAO7ePA/HnGyV2qwi04C/6eKpoBz+l13xKt1Oq3jY9Q2CojYtJtzXdPujHr
NMlxOOKd4BXa1qpsIxqw9HSUlwuPP/chUc+cTcWTmyVAOWysuiKrWOWD/kEEvdC7
O+M1xXCettpdZj9F0mFcA/q++UHxeL3NWuyPwkzfn1MSfstbmdsZWTXo/EtwvKr+
7eHJIUd3veyBD8kxM+BH1sVYmcHTT6gY08UzJgEWhauT4FY/pNq6JCLfKKB3rubY
5VfVMhNsdPfNSR5cFC3oBKgUYcKy6tZyaB81Ar4Djg8ChwtH1AT2E5pwJ4b+dyP0
bBlKjjxjD5LHlPLxLwPCfzL9/kfU+ag4zFRY2lrTj64U288Xo+ki/7DY4EE7ljvZ
a5YmpURxWPDsZVIYc7O+AeXluK1TQpXU+gCw7iwjaiZ5kimyuTMmo1fZ/j9TWzr2
PIkgkOfW/JII8UlGkevZ73nBzH9MPUemKOuoZjy54pI1MLhit35PVx0Xpp+aSQhe
HclF+OExizTcuH8wZ8cpXF5aRD9d+4InIvJ9JmH2ifIFou0OWb+n3dTjJ9vQVw+B
xbpGEjKeFYHSsHwkgnJa8LPHek0jqpN/rzfeDVC3+iW96FS5q0UGkQ0HIRGQFhBB
GRDQ/lN7RzFOhdkv1DdWNjvGwAkWL1fFN7/wgckGsVsJcLYaC2QzYVO9Rjk7TgZT
62J/05j491BjhgNk/O9yO6gQK5S+rPE4RAUbPJtywrj+g0edH09egWCd4uonTKyk
+oYaQnsCNM1G6UcelPGEYVgs5xlQtY2+7w+tJUnGTwZO0zToZAB5fk7F03BEoF1u
RewvADarz/9XJRy1aMthzi+6Ss1MlwN/6bbACV5LMWgHux+vQlsssvaw7KUB2U4z
JtsnAeX1KW9EF0AHLGITjrJiDDuHnmariyEkT33sfeOJyOPe0/CgXhy3fcwgzRjf
ys3e7xuX+z7YItTBeQ0I8cbqXqyecZHDK9PSYnA0mXvt0hRAnzUkYPyzNzZfJtv7
Lij2l4i8TMFMaqzjoawnQfChTxDTTbDJE8Wdy/rvcCpysLvYpIVFqFd2897ZLn7D
XqB7Q1J/PueX9rdDqlk5co0vnLTiiknULXR0iG+4AD91baF3GaBLXFXAvyxEV2qO
8C9gAH/8sP5agpP0JIlxaqTxUnDHRB3M2gxjK5viiAoDmwGS/u2tWneGly8T1mCs
whYEMI7Ee8KEmXRKLVRuy2HnRmDhVxcG37QqDCqJc0ME4lc9fHXNM4O8hG5j6Y99
okKthE5v0tXIvPLp1rs3KhBF70xfSEJmr537bEJdXyjm1KoAFsTcdNMh6H5Acyl2
9WsgsRxutXlQsga39krMUx2yBLEk5g74o2lN1+56YDkT83s0noDKsJa065XnUCt3
QcG0aOqZTSa3w4KqiCNGF9ADCIZ4PkznF3Fk2aeHKB1zbSr5nGpf6L4UcZBuCf1E
J6lDTcsOnvNxajJe5spL1xojyQDU5Hah9zRA4COJpDEF4b1kY0pGeYxCPUdmvYG2
XRStl9sxSh7wQSvA+bv8/XtuRI7GLQ/AG0XYuj57HTjZFPVW5xKha6T3K/GV5x5M
adGjh+r+Uh+KKflX8uTIZJFBWrIMmyyFLPFL1jQoZQb8oljbC2OU3L1XVf8JhrkR
u53avQFUKuIw8zRRUCN89yNzoKCqDUdD0E/9bKhcbMiQ/nzJLHRYZsEYphqodv8Z
h0Nt6rNh79eM1vaVoqyU4/h4lkTB/1LIogbjWJnSfWVHRtU67wa1PpTqKD/3i2Q5
Ub2ADSWX1UChEri4ATYH2SBFVBsUrKH/A63DWuIHfLIltwuyycIflEhKK0yTUC9c
4gIns6N/LDEDqre/ZsiBdNbmcUKTOFKWE48AIAgfY+0TD57r/dZgZiP1RcknVIpD
FeeAO8as7QYHBXahr08PTfNHOII0AHMwIe9VGsrrpDnfsYOWoRwyZtMn9gbrJhF5
godLzFpEkk53X6EoZtADgl2M2Tg5Zj7ojRePLKH8MBTlS/lEfEMvyt1TqiV4gB6L
NJg4+KJLfWvitUiTycpoNi5WMF+4nA5w1wYhG8//gppvDqJj5iSH8oySAUBcrR3I
zkfy6oCPas/knt3oDyHevX65/dqVGxCNYEjpb/osgzr5bek47Tqdc7AXQ78LQo3k
X1Glo0LzkO5Tfb+hyTi+4dFe0sufivl0S7L15Yyxt46jGavvRcqpqRHxPNWUiTFQ
zAxN6CkCSQWLsl9i/dOvf85xzFjiAtw4oOso8gSDgKzVK+yWKJdY3h0l1SL3tnFO
CMcnF/bAWE16y+ddb5j2dT3kmaxxEcb8EzuNIKRqZNjArkv2u2WtdNAA5Uf5uxTV
1gAnzWEHV64wA4Wg20BTN3E5MEO28i+eVIMUkHczVkG4Ig+66eywFvA7Qd7VxErN
V7Ruxjwb92PcHrou+bA81B7qGTXXVaK9AAgu+WdHWiiGtwYxbT8FOzhMMvbAbc1g
xgFbjIed3LHzG8DpGkTk+AnT7Q4zj5rYGtQL59lcRYZdQx8R78Hv3sMdlsiofRLR
oaKm/+oaOnUfBEXEJ/iW3+i732Ymf65ESwStOeflDIPfBHvxaS4S+170DxPHAfHD
qB5grnlBFMhtwOqIa84ArbEeGsvFHwgAmU8uT0og+u3/mmvBHUmmI200iQKxupOD
BakjfSqeCeG+yghMS9en5zC0thSsBU02tLvJJYMDxCiFMI/ZqUH5AZPaF9SBoPj2
QlDsQ4mtTc0Vzv9bU0u+kMDaH/O84c90skiN/S1+Fb6d1i3vjhPmAHR1WkIehal7
k11sW4WtqgYBCglUQsPU0oqAFqUMkmG2T5DsrUp1A8eCN8kcPIh6JrFhwcpO4SRw
+GUzyb5N53BjSLi/JcH/GeIWYt17SY+wI8qpMiBvAP7auG/C7TbRV6TTrafHD78s
TDxAw3qY2IFomi6W7XhLwboM2V6XnW5MQmFVl84wNUgb2dY51UEPVLTy85VKXPuM
rC1SZacoINRHUUwfEmomk9fcfGI+azrsoCFZhWH6gCPZl2z96j2SdaCU3vlEg6ik
dPFHSDq/kYMzxaysZ8o5em7Izf4PpJ6qzpLt0r3Yva/LCIBT8oAz08J6019R9SBI
c2doyBa/lse60tfCHqa3TAV1bpiykvaWHxcbpBtdHc0RZJQJtqiCXmyp4+tv/5S3
VfOKStmBdkvx/NBpaf7Bdhj4YjNknUUslNOrLB2t7Glq4/OvRXNYI7576QvuyDpw
aPMo/cZxpJkBEmlwf47jToXDI80lsFRe1Qh3Ciic+Hl9+4BTNArSJ6QsPqBSKvvF
jjB9WdaYL6VJp9UJo7KcLdkZnIZBqUfGggHqXh97oIlWUw+zeckxuhO0Fr45lEmn
pd+cYJtJIe8I7kUl5Rx5+v4+tMlTB3WsfCjtODSDvwTAS9faW/Wt42Cp8HGIxYwk
BL908V8RT6ulQXEwetvhTkL2b0Fey2kmpTp/u0QyV7HYZjhLqnGmf4Zzj/GFh6Gw
dOL193LK6O16lLScKmZuA7Sa+b/JRPZEVC4Gnuv0cdu/CXMhYtfkMCeMREk8MWmN
fhcFqQQ+6/vYSZwX4sq00/avwI0TNGH6eAaKK0J8gd9HqTolJZfsqp119XqF2dVz
pS2xNvNZfgwZkffcd2in812hPMPLECP7tumWxeWHfk17V9j3eciX+U/KKQJ9SXyv
0Tzfz/K2vSwsPK7kO4LyCjtePJhaYh3h1SuVxh7ESIsCihIg6m3rLxvVdSgtB6En
juM2wRjYaTcyy/hFA7gLN8e/6Ai+BjOurctRVAR3WNPcg2es4+/DPuAMExPdaQjW
NXDWDa8eml/MUchCAQF4fDoColeMHFUFhpBpjab5hPUb/QZEHKQJWx1OlnXvNz4n
tqldMz5H0dkpiwdrP9zEgYLLBco/wULBkblwaDxOmWEAopc/dcoOm2wKK33OxeC5
7yEVHYI4G9NKtAYRQMpDXz99Bk7xCU56OSk9Puxbtr3aki+y0GR9Mnj6k5uvnaJS
FiqwNWQfH1V5HtihmQpi7B5j2+oG6whkIXWVl6RtAOUhq5Dd0xq3a5ud4BVGH8eg
obBxakxJnZvHhzDHSGlm1hSz3T7HnPUzj/x/DvjPYnWM85h7PaGdSeP2O/82CyRr
6vy+JtvnZ9jwL71iBg33nNBqsSNNuRRhDK7CikojStQPN0tib06JZJxdFWHYorGv
uXJzC0K3cZi2fCT7fb0LS6lbvsu1d9CHDYz9JssV2PsVjuhLj4OIj9nUs9ibTnHk
NrfN5ZcenYyNHCy1wjxznu9/1gKG8odLT9KASEQNQKS/UyX9ZioiOqWwDpyt2OWI
JadAipCfkUfBkzEvsCaG7CRKY6+MFj8cG5TwbwYohHfd//zQTwM25JjSBkbsOW/c
5Y/vf+fNyFIg8hglen94SFA06ECtuzmUeo1wHwLmJaKUyXIAHQGjj49sZfT9jPYt
P+8pC9Md1zECMvVWQ8jBPmDx0xXZaNafM9fDAxdm4K70yCHBjiDkBG2nOnGPmN9f
kIdHX+dbOSFroiTRwhXqbZ1TYrCUvu50Yt9dJxwwapx3fV680xN+dTC/7iqLGCfi
OfXrsVtUyabp+VblwaUwb7OIsJ8pOEdjHnT1J93Z1ztaxJDgVsUnSxVOZxSyuu0Z
p8ZKBMHtfdZjcdooNo/KueJ6UvX5uEVmL6472DzDatlxv90NTeDYIlywdA9Ij4za
HYUeLDtzpLIbvXgJutgHRzBHgwTX2bus7nPAaOYyCa6Ov607fFo5/eLmw694PYwF
PXozQYzFi1d9xqSM0ngCOyNt4/1eFjSMEiuXBNQLN0KGe//CpVfxkBDGT/CQisnx
kunCJ/SyI+nSnji4w07gV/MrVKCH90pxA5NO3mBFw0G+3l0g3BjA8WOn+vs6B75E
4uP/rsMT2C9nNPwScUCGvbk7oaV7kRo+6vt47xCWf9DIpUhRSvE1osbbqbylFx23
1bkDwPZ1Lb+XtUgbFnRHgmErTIvB9coMRIu6OalBKN7PHAnahX14hbAwERPsdHSy
f7CvQMJ3AU1xMU2IbFv7h0nBH7WjVzPQLkZ8rLxUCQgwFz4Gv4VhPvV31cn8+ewT
iIqjeabgpxS7iSGs3UkfGzGRaE0+iDjzv4GndQnv+8rhFI0J0nAdAtAdf8Hx64Eh
2NR8dZbxM2LCcjb7gTxxxRaAoccYD1z2zh4Yu4/H6GGOolgx0Oe8QlkfsL9IDPln
8pQd9m6G9ihdJHBoIltDrFhQvFDTszu4Y+gQcC622RrKAoJJEEE+w9xCT6TsGclH
Ia/jNC+YyxdY3Zn9It+xEosm78GuTrKzrIbFHXFRHMZA3kbTOnjLqyuLFIAcimWK
3LZoav3fwc/K4gZP4P+06HbIeLOAvfnTTONIFxfYr8Yzz8NiL1QYTdk2gNTUfweZ
//hmn+PKvV2CbuRpDBpwO1tQ2u3lop2F7jiBq8ecr6xvgW2ptVq3F52H6dn9sD/7
KbhvEyPBOZKnbelJi35OT1++C4nv7nkFCwV9ou2rhdqHDZGDsTSdJd6m8qc/78Sc
pYaBL9prUwAuo8OV4FTsiH42tU7WQuEHlca3bYNdCgYWewaN2EF4hEvwxPea5ZTr
K9tJtabXrHZKn6w2ASjg/odofqJ3P94ArWAKoOfsQcb5EN7tVeOgUdvVswySBcYk
1t3ifDcRxTI3AG91UxKeVpSKmeN4W9chQwtrTmbnBC4YeDAHKAyWFb0e3T4lVYSU
cmEp2BPlAIOUbjaHI8gHyNwnHR989YkNnj8qoj/W/YdE1O2wbTH5kgl7kgzXSg+o
0AXhN26BW5c5jdmwXqZiLjkAQ2F+2wlbcHimxphp9a4HNl3YYqXpImYkrI3Cf5wz
T74dx6oBHid1rLYBvP7bprQvfnQdLMN7TKblOFxXpJl9N+8DRfrrrOKOhZbYxSk5
juYcXWC0PdrGUqBL44xfi8zMjD65zwsl/rVUho1M3hwOk3umMSwVsPxK1UoaFroM
h8/PScChmwM/NsEkrpHOXYcMRncS7pDV7QCInNsc0saSgdGcdO0JeK5KBycTyHDI
KEXFdmnTQKcLuNS/Tq8ZnhMLcnCPUl7j8DvJXkP4wozYrip1ejmWKB+aDmlC5U7n
qyj8MZvJOkTND5JEuoP6Bjgh48m6UBV4eVJpRDE1Np6qoVLi8NzFHCgeEi2MkQ0M
QkRZl+nr08+fbm3rWSGNlEiiNbRLm6XdAjdGf4iykN6zHgkhYFrNl6X7iBNoqRLU
vG37j/cYRXmDlJWx5lWgGYHF7p6BDt/vuuB9gNhTABHqcGwmsXehxpZurzfWJwmn
wyBqi7saIM5oT2i9UzTTRITi5/2/GEmCBs2Ka+fOaXnKqriocpCiSsIDvp/n91g7
Y2RUmdL5vlc/NHLKeXawlJG5CuTO5ZVk4j5wgokxHdwJonMqg7zPHF7Her3ZcSg+
y5sXaQwCKutpBCie/F25hChO7e2rMsCyRe+g1KYJVt5Ex+iwNoWNeJ5swJO9uTSQ
Vxlr147xsZDou/Fyn0Bx2TrjGPxJ8ssFzW/9m7TKuML7Zm8Pp6WOgL8gQ3gQudDu
WqkseMUQJ1a0DuTXGvIPrw+Txde+V0sevbQvHJ1NuQdSNu/zr6bU+WBLmYcAB0bH
tNMuHr9TUhnZ/V7GRpYJ3ntE32n65mT522QVSKvekTDOt2erGukZgxvHOjIvds3R
HdMyynGXwx3GVfGZBrxMhn/BvcLdLVw1SeJsqmDdpVoBDeA4rIfgNeEDZUfPfpNY
dfDBgGp0A+3cdP0QDdw/NtvTYCxK7z2OJ8i4jxFpyXJ+rWYLzfqOljQRyzbO7zJW
ENG3HeIR5L2Iqch/aWET4kMsN9ncJqf62BDgTKT4/fNku80K4LK9dfvgsHo678sy
0RupKw5YERqkvyP2DY7Lm67ztZdmcacYgh3GI2lSU5NG8l1v24e4A1JvEHWW7UqJ
UvHAJdtYQ5khLQ8SNx+VaJ7RHUIeJD0r2kdzqd9e2FvSbdL3Jof4QlPQ7GAS2S80
YNHKdsSN6f4cAvQgLWmXvIFze2p9itAcscr+89LjZ37GLbw5We3DiQGvkiSUOU5o
XzjvkMPu7w8NsMZ/VD6Gxu4pc/1JbewrmfHu99MxFVyLXo0PadRn4MWARIMHdIfn
wnY3NKHCoBSTfV/2wdc06K466EZ3StCwkruJZm27WzEVmhGTSb8+TbL03bRbm9B/
5kGrcnIOzmRMoW6w8oB6KBVfZMgySsQubgXZx/6V0Wd2f1eCf+3RNPkK+Hg5YvRc
PkguXanhWlbgMOXWyuTyD3EKB9/b3v1T1RoagoNMFMag/z0wCsUlbMSuV8SoZ2OM
10Ps2UPVpNqdjTiJSzLdQ1W52ZAcm51d6HYP5DAoNqOTrCpRr/v+GWz+UPpgB6mM
s/3RyOKYCTJtgHjJTKQTdWKWZ4zKezBNO8rfkRpVUWS9UcNaU53uHi+Dj+KjZq9h
8S0zRj/I1UtToxv8oF0hhpSJkDXEDVVuh5/QbSUB9o7Q4WMDxgGIKBy1V/crOfvZ
N/PNXysMhO2jmLzjpBW1585fdZYkTP525Mjz3wWq2/2pp8/GQUE22lceyKSbr5QV
3c3ZzccfbMhuxQutblHDgrnFDVZ1d+rr9h90m3hEW6t8lcVC3e4VLuTeEoJusiKu
yxmOGW7wHVYWCp8Zr00C8vpwoOXrhFhN3ZqN0xo6r2Oawk6A99sXbj2xRF1HhWk+
TktW822u2yTZLT1TAnG3ySOBq4cdr1uyYtTHSBxSI0k7aKyKNvVnjdCRcSv1IK8L
s5qfhBXxhQ6lZYgTq4E4adNLytsHq8blnbtYJv09tTm/sFiTCDyvtAc1rjMwLxww
HvF3G22XhVWmS3bvn5yQXUQV6rPCzbjh36BFqieY5CxNkfQoinzBm1ftL7gTzMYa
jdW6cFDnQ/gUSVWHh6WAhJNoqXNZFg0W+o4p5eeDdfCjb6k8JYoIYfkfk8EdoaKu
SkV2Ps3wXQUJyyzqB90EQuwn+4y94BnAe79u0KFED2wFQpe1gGZGYfk5zNpIuSS6
86T6PxVAB7itrulJM6MK1mvi50V9h8tq6J94O4UiBnvt1CRPsVnrQV8k7NhIyeUu
580tYwY9rpd+uacVdZIEAWRrYuWenX2ht2zlUzYGP8ZOA2haW3orXELUvELT6+LH
tdPra3BPWxL7yPa4oWRvRbrvsGY3ItOfgOroLkYTonTbDinGB03yFWmb3H3RS1xW
7hkRJlZSRfcSOgeE4VVCTbZsVP97VM1fWIUT5kxc8JSZVcYI1xuvuEfeLVhOcfCs
mhMzPMZVJxK6ZV/Dn4EB+4bEZbUSCKNmwZcytcEvI8wbqE73GwvRwXJ0/wyIq8KW
u8OiCRo5dnEg7erdjSyI2ZvgGLtDUVOAbJYssHyY4gUNdyTrR/8vOyWaDBifrvam
x00PjdhhRmlqo4J2qtGT6ez/yfoMIoPdNyYiPI0ypQDaAnYa1SQH6cmpQ4fNkpxP
m7gA2ht7Gq+ZMCaKR1w3uc5Yqvh+8vKEWlwR11YWn8UmCssLjacuX7GLpiaaqZGz
rUIvkgxHuV16+CfG3PdU+SMCqNe9pfHPrie0ZhuLZhmlvHVKzAnXQPx3aO552c78
yOYJvB5hYvSUyHIh12kg5voO3zvoQSIEYPz92NpMDFoCFfsItYQu8Qfo+PTgI7hH
/tcOarnu6TQNGokLiAAb4AK6haDuYeo6CNpCxZxbxmw28eivZlsVCaI8keAU7BLf
T+xjRYK6l0enioCr9VYuA9FLgM8lxRLphi5L8+2xGEMKDpdI6a4DSngJ6zw4WBNP
vklvJi1l2qzsHwvf1dm6+3BwCNtSCcw1GjNILFwrTGjeOHP7Lr7pmkUtcG6Auwyv
1f/wZg+Yzj/7aOt6a2mt1H75OdNOXftUAAVtplDSNZnQqe+GdP4KlFY6FFE+CiFj
HWkkaDyR6nmss61qDhrTDevlyFZSVfA9D4UWC017hWjgbLBvlnW2xI8ote7vG+IV
bVyYYo/e1EBuhC5jEsgyjyGwX5rJvUtQLhQ/c05hr+DWtFJSICegmAb9qxGVtoFC
OWznQqtZphdtwmnvIsZ7pWaSmpB5fwalSrkK70NijEiyQhhJqu0za7eQNuLnnr13
22bjjROUhpI3sHkz75Ebtf+3G/Al4TJBMYgIX6UPvJlJT5Qf7ErRiAC0enhvUfgf
V72NkQ13cMJob/us/15PC1jjePmUpdtBZaqFnyHro/vG86fFq/kTR3GgPS5s6mmF
wk/iqX4tZ1tshN8dOPnmAULV3Ivdni9QhrtOI1tAn/WwYiAIgtF6NiK1M1dXsONY
8eo6lIo1DFbCgx2U1OyEAxJ9GR33yU6e8cNKSm5dyGEh7419fXrXs+m8hW+GFyqX
QC9HCFsrpxs5dKA3DcOfpmk2vGjnya/qiWKifDlRcSkh9napK1BvJG37J08Gj+1Q
gESTPJQf9T2+9buaKcf/PwM/OrpOn6hQC+NiRxkp1A7gB7sBRuxbYuKRO8KEZry3
tjAsF2d7jY71LgIzmTwE7fKrI3D9mNied3hBRRUxxQMxyFE2HNEUTH9O3axqvwWf
AWUwuKCiA1yOSfjHVvz+MENfWbodTTvXKComJriHhIQlO8CdoIODiqVYIAsEsx/1
TThOEvbVTD1hjMeNBmye4Efi96TW/B9UaeMxlOpP40kS6wUvhJexMtajr95Yf98P
Dk2S/T0OuDVDB7ZFDP73JgEA8/2sAJS3EqhGwU0kfFgFvrrPD35HjuJ9q1Soxu9P
4M/4onHICSH9uaOJNBlI3jC0q5VzA/QXrPmUCQ0x+esEmPFbpOnv5k2gPu5RJVx9
AvM5LpiiP9qFMOVAxRWtjJZZ+hlcH2z9Dj3D2y55HaL+kb+vJV0rWuS9CbpSZJ1C
5g0ZfOYaR+Cz2/vHxo8IEbK0aZ6hwMgZ9cwSvaRkkzvkJ3N3M5hRZbc7YBdvbq21
trUu/i2Oyfgssi3gUJLVrwL9e3IFQqPHLA2IXIONbFDU3d+8qA4fyJ7h1eyqPEGl
/HeGEh47e/oyYOKI7iirKVMRH2B30IQsFFx8ZYr1r87LQnqB9Rl4YNOAD79nHLmr
ExFr/XMdYZ1EY5YWLatb/dLHxqGIG6QyO+jHJ+aWuLL71txOicMozo3j98eecSdf
qAPLshyci6cmZz+qF3l3CYhsv/LYcsCBM+R1c51IvQDb8M1JxcCuYE1jlJ8xaelB
dXhnnXfjBQ5bdEwwniDAbzOELYqjUViOFDAhOHgs9bj2eBCe/nidug1Ny3KaAiwu
qkLYWTgkCcGu31bdNiHBUVEqw8/FLm8n+3ofRBHCzdHNnnqkoeT+1zq13rORQvFM
eQ4W6P/jKR29RGebBeDSvkXfSnE8jtEzKRPP1jo3bEfKopWMllCm+elUEMnddRxV
bObtfkzjUc0qaBpOcyx/3U6EL4qqijdNBLfBhAIAfZLVlsdk/nuQr5BI03/jjDhc
kmMK4PPOi3oSCBsh/PNQ4GK1ovhY6Z5dBFMQATcjviGjjluypEH7TFMB0ZCNVLhl
CQ8xG1HfsLPFCo3coxFmkAqH+HEktJLVWDcouoLfr7+ibXAI7dcptSdVoB0On2+F
P6ZZZZGDJknPRXRCYrcu3dQ/YVubrU3TSy77y2eGqLnt+iE3gzlGj3+0N6GyhSIH
yQ4DGBpRonLhui29gz0wrIxGvvCn+KHmbSbmR1XF45bF/0d8vZc2DAiFVBruuDP2
K+rdWZErr4z+L1TKE7Mq5tERfywUHa59j8Xf30akTP/x+p5Nfr6JV34+jPLhqjm5
ptjaXO9YOoQrNBnDd9KL88DCwu3eUPDZoQ56i010fJriGsV87YXbwscwjKUq1tzS
NonqoYzD66kCYMyRURxzJAE1wbrpAFQFuS7P9kM2orUK6ZBhWpXUflsxCTpwLKDI
U/5NTMxAL/E8SoNkM1aK3E1eHngerkt9vBE84eKZvAZkXLW3gZnL6XINU1NT2nYh
BZb3Le5V4XNqZgiHtNoHJdDucMgdZdih3IUKH5Fz065l/3RInTl3WkIh4FOMQtAC
Y9JIWrLIZVctYGw0zHTx8zdgrqCGiSuhTTGcGDTmIXfE4ygLt4OZlBNI6YGQnbna
zqhOiClO6ctlmslWK2MA3vHwIXUnxVBAPsVyltd75pJUiytCXTpxt0EwFBLiO2XX
rDmJI69a9pgpEtYokP9xnqG0r99PYVXjth6SAUN3yPqTnx329m6vw4J/BYFeiLQh
aVG4KVK2xuX7+8V6mQ5nE5UpmNMUoAUB8vUejDZDQEiJhlDxPWfHCc4BVpEoVsm8
FsvThcTpiw0QYT0Jad9C2ZJaE34eY/KpHPjuGi9vQRQJZpP326JJPg9infIt6nCC
ZRshEiFNBYxgyhxxXbcMyCLL6NXlpPMTbLQg3wLYaYnlVr/fRv8vdfujd7S0lBsp
B9evdcy4D/j9FGBLWoazyxvzeea31oXta7VO4GKBUO8vQdDXuNfEUSXO7PCO9MOt
jpY2silXoK/XVQyexoGNiC+QXw7i01qZvJuXDm42F9okvVhZizpwV/kkDneMt39k
bBvZlRxP9yUCekNbP3mm0VI8fiVm7Pv2H1HDBYThuRJcvOAhBxiN5ix/FPVPD87m
tzsuekLOOea+ywPFUfAtCsTDimLrzyYNblR5/WK7VPLnJGjquMjEBnMb/BWcmn4w
MHHbwGC/I+CqDXlXTKSIuL7XtOo7tJSEoiFRPAbmt+sus35mZzDf8gK1RWI0e2CD
RgabAM5j7ffX9uE9o0oz5HkOPw2gMPR1hdTiJesQ/FZv942fxoHaKi27MqvEa/Jj
vbUWKNVmfVKXfKLVhZkfLhrlMtkhTN8bmr7K2MIO82gt73sRz8DrlwCF2BTIR3ih
bI1iybpNSHCb9EwZp4p1q+hwJAuR6qLX2yyIOxccSnKl7a7bn+pRAR+XmXekkhT6
vWIzTBI0x1hulJtSpFjjy0mqwuKNGptIrH/8waZ3ET8BHAzfK2bhY3mAdM8IE6va
LBLedRkDZ6Hj9WnHVGdpSI5R7Z3zF7nMMVACWzpiiQcx5du19d1ZnySYSAgHha9I
Lye7m6lTC3FDJk10tUyN5eWSK0f7r4OSHkfSvDOVEcoM2HMjhFRBYi8fGnuGzHmm
Qva4tnZ79WHVeZZdfYRONUDUCq6Qz1lAGJH0f4qlp5TXEmHn4QHb/LvGWHo9ERjO
Wkp6eNzkK5uJirqKEgQGwFQDISW/oalIleosGOZtdsZTFUL+K26JHp/vNj/PbNaA
cBGuQe0PI53xtwiV9a5AkRUZpua9hhhNt63P7osaDCAmyKA59MME+JwtuA54uMJm
CJsruwZEzzXb2mtzEcV+/+1zj766EM3IugUDhD1tf6zkzNQsqlAIzgSjQDue58a1
vaJYLHjMZw/2dBBOaFseQnydmWNV2JY+rXtDILZG0O4oIgdzcK+7Xu4Op3u6EIut
PayTCHLLy9yXRWqVoE2Cg9wNsYQmMlzSItK5ujxBbl8xzStEqvAeEm8iKpM/nfqv
+rcocTStUaM6Hpd/RiMyAyxILAKYeJO3fPCc/luDM2qM+R+Yg2CgyYk0babcSSPk
k/yudTO+gS4S8NdlMKT/fDIzFHekEd17ZFqzxTVYjwFKkJqYczyfUIZyVQ3+tSiw
2l3bFZ/SIcd1OIdA3ib1f4vO/wXhF3ombkm0byd4a/uPxvjcjP4IEKvqVcbxiHH7
RxGog7z/iD5rjzkHaCc54AyDcH0jAS/Ge9genS1O2t89XhN+ZtGd8QIhzMniAo+3
zgeuL4tK6ZwhWoVKcjH9M529PwogthIEXyK+slNT/e0qGmaA/pImncNotG4aFh+B
VpBoTnDEBh+d4nY9ncZQViSCoT0iXaBpRyh4g+JkjMB+OAfKPvil/aNu8feT7g+e
DzD1doBVIgALre4NssYUGhYu55mkZuZF562QNOv7UENYuOJjxnnW5LcCXENzFXGI
kD2Iah+B5LdCNNLKkJTUruIIiJ8orQpVZwWixyEwQA5+EGlN9AypQ+RHCDmO5ccw
yOOXCOEw+aS3WFMrTEzZhn4KT+U5T1T+/tP/kzknuNDMdVDvGTeulZ6Gxcj8KsoL
NaV7u1KCrxjtLj2rF9UjA4B5T26XUscStzKtYb9PYE7Y3RIxHAzlJYVLN2fZaCiI
npUlSFW/Sms2O216rkzvhFOsm9BxJ4jdngvtUArSmtvRbJ583KzKbD555wqxpuJk
hMsYxPVv3XMuBSTi4wjqRgrAoolO/UkhS2Nfc6fgXG5aer5s0B9var0CaNQW7hka
LQjPviwWKYBPrUR4V0uJPr8fAIPjLA+8TKTYs4MDBSum36Ky0wddOtE0JPyZAfXl
/UYKgvoN+7eP2PKFIxVqJ198VXhsjTMzDGPO292hBMXtxYL2k7fzQqx9y5iWXAyO
31gskXiispp/M66ag3UtoQF455j/a3ubYWJ42YUHmJoAiyZL4PnnTuv6mw5cIFm9
WX8Q9vD6Jf5h+8yzrTOp6F86K4F8+6OwtEH7jKClLdZKQTHQorkqW8uz2bkmn2N6
AIZLN7/24BmifpaekPgU77xz/xUCdK0QgYGx+GcK0ZbUiQvxjLUngAiqpEa/u0Sb
Fw1NLEP9RgF+FiPTn4TKJojqdFkUrY566vGaCopw3RHIytQoB7YadTNZeA4tKHJq
FPQnK1U/DMWp3v24hfKoQDV/a7lDjDI0xbquGkN0vqQJHAnv47nS2/6u8Z5ibvUd
/Pqxr7Um0HrjpdRIXEdd4Z3gms3oeO9ZH0b3e7m+WjsLKP/t+DxR35I94rt00ftd
DGxgg2mKxh+UhfNEuuE8DDbCs5juPfCOFnRWJXnQZsmzp5gIg113EzwozxMxjAwb
YmtmImXGX/s2ErgE4MYk4FhsRFzrNX2FEfXD/JUN1iAsWmfKeF4TBzZFRb8ZJmiZ
gGzukuk/ftiTK1z1gUIvOjhjCDSMXpoT96m1XjsChzzeWDUcx1XeADnE/w/WCfpt
+8N4pmBNnhjyVuUQZlkznbw1zTyJxdxbeysDljTYvyByjtHWCi9NO1yrcP01Djrk
Nbp1PerwGBfFc3eRMRy2ZFI97Hcb/3zYHCz3jMENDrFLJsZ5HcB0OShUmbVg8xuo
s8kXlLiBsPQypiSV4bNOkbvA0oDb4Sa2xFs69pwGvb8aecD8Bn2gfJtYjU9/z4gB
f3ixaRiX9ludRi+WBgdUoyvx80tuBra0sFuvojJ36wXhPWTHDc7bPuJkc01QXZHg
Uock+aq75JE8yK1yt7TFg+vpJzKedFT1cuFdIcm+CO9+jyj/L1gBbXzfiVIZcRgi
xIyGzo3F1c8IzQooC78LxJZ8vx7wf/lx994FQwzks1l4B5a/oDyv8mQuN1yqlaIR
SWT/9lWMJjYpd9HyVKnWCmySHosAZZYw9z+pyGEL5KqIxqUEVogZfsBApII3xMt8
rI/IADEas6q5Jmq7mQcLtifOksNbpOuvxQFxuKtXPswKzmrIBK06yatv0z71cdq7
dsaTXqq5lMzltMZPOKYoswML7/kA/efGFPnsSei03SM8r2jU9HxmDXWzvltRrPql
KVggwY7oGjTkKmNHdJu7fOkVu+x3EH9ogRwf36KpPW8sHtK6JUzEi6roZ5STxOPx
mbz4UCMPKm0tvZgRN3A1kFnKnAijli8HBSkwabRg2kW6QzCXOe58W37UnuTeDhQ3
Cn5GlpRJ/Z1tbRoeMplLtJ22ZzyOPYK5+9Sbz2EEK+7bYcDxi2qftP4eht4stxwk
n+NB9+892XGL2EuDnG6kHG5xJScNYjTrtaavwB4IfL5rGq02znfKt6LMERVskWjk
GZSFkGCtO18+zaBHUhJ6lg82hLPhd62+7kIdYk0/yHx/yEYaZ+sTQhx6BmmdkTjL
UuwpeyM7dNXGUcSHt0ZiepyizqBj+S6ZH4jyrjFWi8PZbEkYg3O78jvzyhPsEQH7
7h8vf7TAoIuWLaSefzyNaPqbIOD81411P87NG6z1+BcjS6/w4UNkAmDfJ35JUYE4
jaTX9Tx08iMhEr0LWh1HwLrLNTBdiCOJ3xx6IU61n86zKJN3EBkG2QG8O8HJn5D5
/SPMEYmkjQVSir+cxQ05O79iEM0uTsBgD9kxRbuv39okAx67eXtaKH4jGjaRcmB6
ULXMZYmhAM6MOUVgRdUlatiqpVVVYzdP7ij80977b0FK72LRGLIRN9DhBnArkwnV
Ls5bDlstwXCk5tc/8YsbxdDrtIAJxQs8A2tby2uW1YuyR0X2Sh9i0WINQqF1cBE7
9Ta7sag9Vtp4s9Ok+aBLhPZDrDXCJ/XpWVemvex12YgrMDQWiI0gxiemNDJ3LHvJ
w1xvUFVzgdjOF7DyskFRdvcMny+6iju2fHexZKizTPrACP50V8UB65gIoy0HnIeN
KVsLAVHahmMSnAZYdpIidiNIgo88Vt3nscflxLjiKJRY/4sBt9+lsOhgaV9i8TEi
VXFPY66l5xz1lb1nUmE7vVVO/Himr35gx9ibM3qFBr8hbJc83WbpaChy9N59fYx2
8Jk2jiegboBVQpwO4ZB8PBAV/QVKHDeo8TAiuJmnql0IRHJ4HDBz1vJ46ZaPKkx+
OP1WPXpVBjeKoIGrTVnftLVi81XP3H2Ntmd1GH5gECtqmsMIKOZ5JxLlHvMsZrYN
t5mrogWwHEk2RGNtky5xrGu39kR2YDlUbq9JikiipnU9IQ34u20+e2CauEyFyN5W
AXYQt1axtj0xuUCskSRTvSy4Z19gA0DusrNZSQdCtZ1MqyqnMXe0ZQPp/jNjj56A
uu2jRve/INa6x3IvpogrhU02BCi0afXHlKuLseQoh709CtcyQWSiYQ3aEn7ejnko
FgsP+dvDH3ijygNduzwFIPOSqNJ6EB5Ayh3S/dhrx6qv0DLkAG6L1cRDYw1Btdwg
LtPPRc3inyMxeduECp/qagBEkdTf6bPuvdFg2JpFsv+RbU+4Z79LV4B1Izk3+Xjd
QU7QKsadnSZrjxeILxudfp41DDtTrOoXdKD6lM6oM3Vd/PE1wdAwFzZndpo5HVQw
F1+86LbPN33AfvoQve/jyff2PO3Hlh3FPD7NB4CFhjnBnCbcF47cMJnt5eSLNQPA
lK+t4tYIb1tu+pF7mw8cl5TFBXDmKp10oiXhh38E1V7myIGm+BB89+MryRRjQtam
+tTZP4vSEdiZvNKmUlvxT3i816L5xVRhkgwxys6l6t/K21y6uhGX/GnDsvSA8RBJ
LlFQxJNzrqIKFc38QXZjMEkDywu+qjLbOJHB4awbjNVb4czPknzqm0qjWGOarnJb
KdnsPfvtjNAtVkKWZH+5OFz4RayEWSkMZqnrl+acE3hSUhTDlV66o8eZSWO5Yp1Q
lH6DpSSnM8gWBQD1+P8foUZhrrCanXNlGNbbjzM7ZRMH1TH3p2GJABkt64Dh7cnH
qR1MTVIWbLNyH8YvXL6Wp5pUsRhHxJRBQ6tP3yVbsZVKLh1YcSQq2LLmeEKlwaNP
Za9rjPLwYlmn3l9zEnkiDHsXzxNDtqtMiN0p/F3xpIPmfzulVcowFjkSY7aPF1ka
z+/io4NtcZJ8TVRgBtql4IwSsliXgHLmGalGC36Z8KuHUmcBav/ImhDPXPCgtxuX
YyiLgmH+KSke6rqL/Ou9YHgoTxrEVk6jwJEsnaBZbZ2FWrJ5CJlRKysuKk1WQVPD
KzLR9KyMLFiOufPDYbyL9Ea9GlYC0m/P1RIhPz7iCqdnV+l2M6rxTxkIdsAhKpHV
VaNbBT11PMzm+FPW4v4jB0wgJoKWSmPRyq0/Y/tW/YeXEJbg73wmue2Lf+ys4/Gy
/6HGF8t2zUur+GgukTMeEYGI3bPk58Y9J66Aiyo+Fa4sZ6yQuQBhnI5LPwVErRQK
PZL2yisjjTY7Xxj+97e5fTpw0I5KWQVIl7QFCXRS+Ip5G9c1ybTgTjTQTJYn5m8C
9CJBmjFe6r0UGA9TR0DTsk0Iouu6mvE5zyTaUORNScWa7Nnt+FQ5+s6RAWU49tsW
4sfYGEkN/Lr/ye1LUYH+58+JWZM4Jgxhu1HzUbN8ED+BGEmTKryViIIXDvbKsGB9
pjoO5eIDEqDAyn/v8G+71nc26UP0gDeUC5O2roux58rZG/pDpwnaa14zZBdx7Xih
CqZAD83cLJ9skK9ABcDXtRDZ2u4S8i8OEi6fn3YrqwekJIf1R8OglUdBm7LgjzmO
QUecZUkWBIsBRLYNUeT1EEF5jcb/HaJA1Qqfd6Oc/MUjc9L6Mon3c+8K8HzLNeDW
7qY+VokWeRKUSDn2nBPoWqdDUj64G9c58jPZncmgHgQ/OPsskvzJEsetsIDg7ocz
u++59S5Vkny1NVlkpoNMQAIb7WDUqlZqidx8ybtInQxVZEJkPQKF8xCE1v1QB0Ud
wLpmR1qTQuCVAmWXh/26C7yIc/egJIeuuGBV9z+XY8z8dCOwQC9xaninEXq+WF/t
vzgk4DLTdGMB/14UvVVvQaD4nM2in2Jy+rUBIATXxl4oUXYVzn0c04Ytxy9e1Eey
tsUgHkTyi4GzKSaPQHKrf1xu4nQvr5hcx0291lA0x+LtDvFtRZk1xKb6rpP+S+mp
xoeOg6jBfyXEpyINlZf03GHUm3mbi30r/Ofhuu97018u+eKAoQ2P+l+LgFFNViuw
HZz8gkM/B4zDmccBOsuad8GL6RJPtimmd2uh++mbJskxC4vnygWrydzjSdQwqECd
UVGUr4Se/4sPnT9FqUutCOHu6L0MnxYPNPbQa0leWzTiaUjThDv6mYwpvMgnA8Nr
ZDdea1fxx+JDoLaUTwilmWe8jrCtx43b8mzBxmBw7LRXKrpYpUg2/Yp5LmtBJHKn
PjG8fnMNKde6cMP62aQiFrHFX7qIRmwrqTAaFkTQbzSZHgLjR1q//TnSgpWJeKzR
KBLJTnzGU8mRpJp1C+FDTbvEMbAfCyQWofiYv0s7TLSr0IC07L7LhNjPOv6JFuqx
a2rwx9LuLUv4/SMagOVV5co/Au/Cdu9Elna1MubXosbnIZWW06qWS2YEZgTx2+ZC
Pgw602KSKYykS6wVNEbPRgBUY0gZynKciBjzcacOOh3pCzrbjdNRgC2bT9kyIVdg
P8321+TwstoNfKQu8cYRhdaR0J/GxaZGHWoBoRnGeK699jHw7PupFfOciJ8Vm0c4
peytZVLzjEpNFvN9pPWyB0IAtWaz4tQsN9IF0bz0TbTI1qKHlVNnYk7g9lfl4Yu/
nT49lr4zsNf9a6+FgHB2vpYFMwVu4JWsBOvgwrqlCp5U2iwloJw0qLvmRcuFsIEu
L2Lj9BWF1mswVlHwPrDHcuV0TI3N0h97wHd8SMRC+Rq1vqP5S+UyWPQJ2twyI/fb
3/P0qI/4refj+BbC1RmluH9W/fJfG20cVxa/F1x7jPTbtGZqRbi1x8MASXGtKSc3
hHTdu8ybo2wwZXtIer8gzetTbTbI4O7mxfA+2xER1/znnLP3aJeskg6+i+04RXTB
8dFXt9KKtcWvKTx1m4XNTFaQw3Rkar8yHosNL0d1/tm3iAvwLAkUiMwmihVEJpia
4xfub5yg3ia7AnRY7NB87TrfHtMmN/wpyYdPMU3HsnglGg+4D70nzcloTUezOXTc
WjxzjYk8ixhhNAynaigL3eVNvndR0+mufLe78nsOMB5lYRfd7UO9N6TrOj77TmcO
hvsr1adr2u6wHbjEP26tWMrHFRK/f2Vz39zjZLHnmQthi/YU1yr6c3bCOJ82OHCX
rqhxOAwgDCH0qSvLgn1Qd8t+N3mt8F6jvWcnaYvvWA00y2RLo1hpd6q8UdFK895s
Dd1UBe1aLCH09GopBmPGB871V6lU+OwZaP+l3eGdx0ngjQEVzWVonU+7ctBvleog
JOe9GK7NZyo8ZP4Sv964PR/dCgfuBVAHZRlVu4OGys6GLWR34Raua9W6IPl83aRQ
c2UwP2z4fovDraTx5w6oUhie9J2RzraKgCap5ILgrBTgg0HpBgrlvMRwoi08E5rR
akr8JQPaLVOWoHjlP5KDB+ZcK6Sjgoi9sR8QA5axy0w0dHLF5g3BIVLCFGWjMdkY
uU+UOOn/8x6sSkFUZ3aiGx9Pmxfzm7UfoTjL9a8kdeK0/v2NaePXiN6adUWEozOp
Bo11c87lxxgxF0ws+9mxSsAFFCZRctYRJRRXK9Bz6/KybLbVcUqCf+vpf637hP5H
59lS7H1J1rdtmhz8AtB/UGbqhjMT0PWjMFzb2W86o5sAGKrprJxvXbxbVSZWVUtJ
Jyk1HENjOSAThrVSl/j5i0xPthC+35G3yKHIWX9tWucktSQvbnRxboJD90w6YCHJ
3k9kRQveb+trKwvWGT/Jm4HJlVeTSC896lv9e+KOGBLS1fRNtIdL2YC0dddlcgr5
bDSz11qDs3eHaGj312DFQdIqb82zSWQ1aVXRSoAIjARJ8OUOmyGAVdn9w9/VklWB
roferg+iCgt65YLfAZ8FT7gYG3cDW8DqMDT1yl/Rbofsn83mvjKogFcjLJxyWdnk
LRwdfCWX0L0GxnVlMGp7IsKeObQfrK2/rcRm8I/hwk5QOEVv/AosdRxdsbKzJQGV
NN5n23SkBc3sE/RMIlPDY/d6RYvqgCkL5S03b+M0vyK4T7VJ44WyPylOmKU4d2Rg
L0ocvwHft8IX/tPrsRb4kQrcFCph7HCkjKRgzMChrCz/gikwNLQXeexapEMpF6Xl
ITl4DWNv5bHdJKarB0upvco9w8vYDLz221yI1dVqIlJqqmGNmXco31sAIUnzl5hV
iOk8NKnHP4+WyEYImiITKOiFGJCg3mP7kQw1EdKO2K5WHYhqWa2W0Smyvxz8fTL7
F+MydGDjY13L4LGHik+FA38kVBd4pzN/GLJrXQnjQGKyjippkbsREdnWboyTPf0B
RMn8xPjuRprv5dEdTeph2yPjev0yleahO18lVC/NaOGZGXts1PiUkpvRd6B+qS95
ZvTEixr0pH8X6LghYKEqQqV7AQzNQ95NFS5gkcT0ufRDY+A55KTRupbBO6vsInH9
YwpivaZsmTcDH38b/mo/4xvP2WmuVi6pnygkCw4G9m+Qc2r0OGyYl9rI3mz4cS3f
2lswfX7XXE4HQaxa+dv8AYZhwqPes+jgfPM8LjyixppK3wP3w4W/RuCvFT/sj1sG
YfAJp2/cpFWGEo8T+MNlMufYxyJz5PrV4jEZxKehBALCw08UBVqX+vnxK3BnRbuU
b0nVZborWELFa60aZXY89g+miyf15CkVR8fqjcbiCtmdlS4+mzJWC8FBna1tZY77
b0qAvyJ+047XJ8g34ZVzHQlyMCEXKMp/ERHeX3YbBGvzdpnCfF+NAiahhH5cAqG9
Pg/qCxZaI1ivG9h/RiqzrgfJhLjiyLvabVCjKPST8d4KKGhKZLnsso1xn8vW4+wk
llwVtQdW6eNsvM7/md1gMsBD2o7dZDWFzJ0sAfsSbWj3CuMYi+QmH2f7FsGDcFoB
JWIG1/DkhMPho0bD2Vzabb7HskC9//Zp4OqITF3FX/ViJ/f+oxDp1RzGMU9I1wB5
MphsppMYDr1alugxj7F3siWDj6CJgEclhdjwB6xXRUglPdQpWXl288MwXtHC/Nxx
o9YR1vh1buU2BGploHIPf2OS71s1REPd5Jd1xaI85Ya3/Nc94uA9DjI/GK8by+ZQ
ImTqf/KJTwmzsEcwbG/WE5u+wzmtIUb7jtlJ4g1D/McOKt3OWoiKVXPu7he60GqY
u414/ZfYZnyYmMKtuXs8ITBXhqu95pjxI9xlV3og197Vkt7jr41zhDp9J7vVHfGU
e1AgmZJ/sByRi5tTlBwzkX7XKj7Uo2V6WezayVALn5YeSA8hmegPmpswkthjnSiH
PloBE6Yx5nI+t1wXRjKw07j5XTJ6LFwfwwASFB5DUBmUA+qBk3JnYOrF4UaFYN44
kXiiXLeIHQIEOZVZcgUnF9AMBMC0dfxG0bE+6OzIt6ldU8tYRbPbm2MCRQPKlDRQ
lMFEKWXK2DzMt/q61/hQD5NsqX+f4L6JAKupaPNnR0hMYNaxvVFRSAH56yO0lldu
Y2bBbpGIMEHYSMSzjp6e+NozofvDprVMv2/D/llsnV4Hp0KMaGjbmPX9TJrTKVRN
Vnx37Xqdy96h9uuS0tKW4l3WaUhf7uFLpT17ea3CVCKWFpuiayIriucJ44cPiMpU
TZ21XDCDwarn+JJocOkOjkqztO+LbPGh05BKfRB+KHlAMmS8szk1laKqYaD3hCEw
yZHbIeHuMFX5d/mlfI5j3v91lcXIJAnnQvhTpyMx/CwQNNvUvuHsKKnoLqJDMZcr
n3xN3R6RDKkxYjUP5i72dO5g2OCtM2BE9cbyu6OB22k+CXqQ21m4o0FgtebWdYsc
0eTsn9BOMKpsqFsW0Pwsdy3nqjUGgVF0ew3nVelw9WB+WKShAB55TJub0F+Xjteq
UgdGoN0vWkk6CV8kIuycaz5UzAtVArATvY965330ltv5DUYylgPfuWG25jmgJRlM
FiwGf+szC77p6voKmh5GqRYlbzOpkQrwT3XaJGZnAJUZqK9AJmk5d0cSbtFfxFn3
xrnOeehf0g4vuewUJlABBjsObW28PiWJt/wuPr41IB8GLbWpUVvWhdOTp0FJlP8m
jWXjP4v/7nmlQyw2yRMxb5NL1wInx+VIaAg8idSnKjUe9AOGr6VNUus4XsmGMuVr
/c+H+KVxokZH/lx8HFZ0rpYhs8unNZ0K841E5jbY0Cgy+kk8Qw01NLzmb3eCyg3y
uilBfgHHdAOJQFptcJCtfg2+DI1tmvEXAsW4UFYEFonR5DdoD8YAh+14T7F0oCkx
Yf/bdEXGc45QV73fkX4QjmcRflwXaVUrQoar89OTUAe3X8yy+Hjk6FhRCxHiyxC5
J6ecvc6j1uVXXRgJwsH6NFp1rlF/zrzThDUnvBku3MCZpHmau9Cbo8++krh+zj2j
fsKwpEEs3ne4iC1Fl1r66Sk4wcUkWOo+Ag8xMyRueltz04Hit5WMx/cZIoLo9TOz
vpB16j96f186RPc4S/fEBzIH+ENOMHyI2O26s0Do4zfB4QR1egjD9kc43Nmsm7hy
/x4A9YOGvzYTh+xsZvyvO7Mqa0soyHWvkEY2c0OY48vbBlvZvCFixjzUy933mTgm
jXfJVJPV5rKs5zqBtSp9CMbhHsBeikTrB/7UbpdYr9Y+bYERTbiDCBDFgbm9maKs
mQTTwDYdIT/M49uEdLXUZgU6mIQifqVbtuoaEuG434B6Ytr8jN3llWDBlinWzFKR
x1hqb4EY4uzFelUVqwlhqP6BlJ+kqOigdqcHAPkOp+oQlTGX0N7neGCuEfJMr8+Z
ohemMjcqVdyzt0JL6Age9JNR0Z+GsidgjfUd9mhJxHWjSiPQunB1rrFiWIBT5Ddf
ZJUiRKFiE3EgDx+tOIaV/lAlDheqPiB8+sy9auaMN922L3QCVfFqgSaXjWn+YSDP
UuDpqJsMX0YU/hPEr1HS+2K0Xcfd7k1gleZWzQHpGewU7uSN+RT585khugSO8kTh
lTefEF8DuggQ3Na1pvE6ejpTVZRMUb+CDpiqJm4rprTj8D/P/k74yraqvA+s7ZSR
HyOzd+/X/Fb4oMvdkyZmi4Ei3gDP19564NlaGbeUoDrHU2fvIPii5OOQlNj4a0Go
hyJpnRL/osFFBF6acgRkYgJlJl4tOV2r3RRElNI0e6bWzbdpJdW6mL4Jyo2vNttI
RF6mqiEgvyQA78n2BkPAJNWoWVPl4MO/htloKifd0bMK+9T7Je3vi1g5tvsFzULd
rj6tSCdSYXJnqdREhHH8QwIFudfJSasm2KRBdntp/KUkJbK2Fg3fPqiXFKNZjnN4
zhvgbMwVUgo8d6Deyfk2x7nfCfwK+HMxBYIr8dGuYeJQX6NmIjmfuY0GH1CuRc4D
RXvBa/19sltl++h3uCYl7oKUfNF09Fo6tp+u7SLPl26jxy+RnXND37on76UBKr7i
oD/hvuQuee1K5JVCqfeUJHy4yoNM+L/dOoN5hGQkw1PVJD4wMYE+DgtU97B7QS+0
Yi+4aU3rNNX/H03A1M9FtUZpSvnIxAJ7ud3n2x1jimdo5nKtmmshOtFktc7+Ee9h
dtRcvpHzp7+yEPwYNx93PgX/WcCUiXEalKXVSQMTeio7fs5m3FNRN/xWGmuoIMhw
0RQcXp+yYjTnhvoT5eCGN48IdKBHJQojFBfLuKW6HHMdnQtPC8thtL83yE9lnQNd
ziGN6N6n3I6tvZkSmAVxN4rwd3iW5pKcyFJtLkxH7po6IfCBfqHHdRYhS9V9h5Tx
y6iD3RqM/YJ38BbaSnOn7PjzqxWDZZZBcvt4cZj0yIhI/orz/JbdGmbkBXZeTDo+
dhU/OM04jLSDPvlRJzbhJxthMuu+ohypZ4VpknYtsufw40Cb4Sl3tTXIVHgV3YVq
y+9OhsLs05ES4Wgpupux2AKRGHJbKjUKDmTuCvI3WQyauwMN1Tncby9OWqlVnSV7
/3paXTORmmr1vlsflt5u30EX8YlP3JYEgnqePKFsn5ieU58aXnJJmsJRfqCO7ty+
HgEXKvKy7A/Dq9hF9bdRNid+6/CoEfKQFWpVCv54zP9O9BLPZjZwrx5Q1f6Zb9WE
/1xHnTbiiECeOZolLIA274A/olxSF3zx1Rs+MV7rxr7dtrOLVw5mKpFwnFWplRHE
ZNshFsGkbzUAf4jJY5gy3AJzRyOdgpv19sbPQE2ZEZfZcat0CTOORA7XF9/UeuKh
Azt4i8p1zJ//mnFiHamjognO6P3YAhhKida/wA4MKa786kKTVLuqnHtmUorMjStR
OhtjWRAR+OlCFGamTkIyTEsrGQI6RlEvHXasUNSc1d8U4uRzWyzu9fbmGNH8DIsq
uTGipAoYuyMC3FW7FeJxqs0eEZI4jwvPEbfz9vo2nfZj6FiKzLz/lt8EGHbFXx3k
xnWNI2Ql7tKTr8CfvYWFV7T3lgAE9gcGF9Dxm5gySgBWUeLnoRVM+SiOFJLYRrkr
7ySqZ+tG731OyzYORcY+Qe7Sp4VVhoAf0pNj/W1a7ByTqhUpH/YiRNb0tPnidrOu
FhFPuEIOz/d+Q7lgI0N5MMf01i1h5kIYMjbCsD4QW+n05YsS/r6bQc8cuKWqUOzV
RVY2QY31wnx52bPv5GTkEG68eXSEAIeKDNjmOeD0YEMEm+BvRIkmgWxpf/zFR3kN
g0Q6CYZmGf+GY8ngDzKEZ2HxlBvNC4dJQ1gh/rXhWvyfzaYemoCVieMENtR6Q5C9
G1Y1XSJoYsTA0QPgx+EESbH7wBXyjq9O7CHNazo/YWTLC9riiaYsrGxxgfdEBrZl
T20I6m5yXos2U+TSsHia+2W9zz4QinwZCZ6YP3dVrOHdp0+/wk7InZvR9VGyEYiC
tn5aInXLj5bdUtMLa4TLFcmmx2jbu69epDCKrlErJ9yFdTA6zkk1OTfm5b4AhCsj
6MvhnGvLAy7nvbAVi1V97CktrWy9aQZQenBonSNyPFSoUXrLFZ6dL73pZRu43zD2
CMbgAnyTpvskE3DcTOsj/oiIWJOwlvqbGwHXrIY+bpmNXH+n8xdwHKlZ+MJ4qP+1
n91EImpKEdKTgAIUPnpAAE/H/jAObr146X9KejhbNKp3nDY71xOUhOX+w2bRZDkD
zwvzbpJ6v/Y25M3k8yChfuHV/CTXSfhChax5JaqPQSvUrQxCWExD5cqR1W6WCv0+
LXH/1trjMOQmCmO21ValMmswbB92bUZ5i3dTc57xRgL/EWMnQFWaimPILlUp7wsn
eg1mKNvJ+LFTJW6ay2qck5i/KmmvdKHhl/ElSWqrcparNqjTpVDYLDteLiM3Y3Nc
6DactWgUmFlXiShHCQKksrNGquZWzvkXr4Suoc6f667jLAb5QxCjEm+gk3RWHmSf
ZDvsRkaImglUrzdXQY0DhhOudF3NCTwRM04uE40bstRNOMwkpiccBL609f73mKm5
85vyH56wPSMnORUt7NynAT0b4hqIRX++AcHgY6Qtm8/lFJ3w3IuDlOicEks72EVK
DX3UZ6owbPfowzTfV9Ve7XUODnbjhirj4AsbmuuPHAsEEctt+pLEH2LgCKNFR7DL
rJDI42IiNi9T50onf59KQWtKGTE0R0A+Fs0PULPDcuViXjuBbxa4bSKTQluAkf5H
bd5D76d4po6QB7Gw1ZVPqdJgN+ZIavoPk6jNTJ6Z8w5op97rBzuXn4Rr88tm65nt
dkGDi2u/Rso6j5RBpG32nuTsJwgfu7DXE4+SyD4G4lu4rY/vqqSfCWKi/SBgfiq0
6p0wqfUzubTZBGLbnY2GyLIiJzTpy0rDuUDzhWaytAgYXrJmzVXj1x5dLrjRmNPb
kLzN1dEeFxzJJ1a9+fuDGxU2OxqNA80aN6H4338qLTf+v6PXlFIm4d81JnbyE7RW
hEev5gV0CHif3UwMzx9rcrFG2+Bpf/UEm6N/XGqm1T59jGUrGGbR0mxSx1NecNbh
VcklVfiCzcWGpD8sLMiZJnSPF95QyTFDsm1HVU1lOzltojTg1kd9kgTdBzv284IT
vZaCUUeTYrMnEGa19KGiLZoyptYQbkBfH6M74w1nUPF8xBYZh6NaQXlzFHzkHNm7
V+Tkf3Vb7oNNBvXSBynsfXc70Sbtxc6S8MdUq7gHCBtqLyjVvjbxoXU6zN9Ko2z9
eWz8ORj+cB08BRx6IHaTLFKl5RKKgDLfLij0LF5NxLDCIerKXOYCmsS25CHvADSw
WL+YTkX90ZIwERcOqhkvCVaWevx5s/bkUpZK6aCo7hoT6rUBGVOZ6yFvPQVam1P6
9gtKKwUWcxc+AAKy57MrI2EEUkKkJY6F14x9mNk8BkTVi4ecschQ1dhDBDdLd8dP
eNQ9l7uhdIScmWlILV36yRr3w3iUu9qvzpSjRTP5+3ukiXeBNC4/jHoZKlRWcgea
Rp8JZq6KuZ+Htgqba1FCowkhA4JsQbR6fE5vFgEC0hk2o545anT8hKdmzx8cG92d
HX9x8LYqMxP/yQjNWwVrEWTpYKdnYGWQr+L+dfpQHg3guHDS4cBrrSbg5bUmAL7L
7HNA8oEwBO3x85R9rcrgmv0IZp9vhZie+FmTOi9IxEhuXLpKFdGJxxe0xk9pbwPy
5IeSwapjA3fChBYrwYLP3TswaHWL58grH9hIi+485Vvz79bfIU+vpcCRb3P9KTGm
lbOIZEwf+9OWxvLfN3h4TwyhIKkoYajYHt1Fp6nP34sHrIbeDb4qJk9D3pXa1U4W
Mpeav9NxMlCRiliOxkJpWKhghXWFK9vIQ5V9R73KmCR3+85In0NqZfKplXuLNGRU
wzFJMq89ykZTJDGCvz/WvVl2+5GLLsUgVrreONuHpN027tscLH6akf2jIxr3tpGW
mEyOO/BUXAeivxLBlge3j8QhhCB6mgS/eBr0EDa95Vab1IpCSxE0UKJNmGAWc1/K
pAk81b2beEwGYSJllPS6q8BOlUP/DbmpE3hulNK48+5D+LfWA/qswy8F9DzMr0Rn
vXlJgqBK9OnlugMN76/+fHjCyqXnWv22bBJroh++aB6CnMNXvVFfCGDP5Fy2uEb0
HGeoyCaf0L417Svnd3v+SnFTMLnZXqTscGGcM6Gc98InS4Og4Vm+c4SpypD+2aOh
EqFcEuUPRz3FHF8OzBq9yY1vHXhtAZQQovr0BZPP7algyP0lSWu4OIcA+jO6WAQW
k7ObDYtUodo9dsTR10zlmQG8BDXeWvj2OZlLIG/yUh7dYHrsvQdNpgLkGua7XchI
yKwU+SJwXFawmyUKeO6iJQTEUrel3xCBMglbztdUvy9ayIxh6CFpIUY42RamSpST
uzJNE4+AMDeb8vdaYFlRBeZ+fxQHXKCiJCi2B9baZMW+rYwNkPrwD1xEEEHvgAB1
2JhxhTAHWQan/B/nmH3MamPnf5gECzzmBKHnohpBUE6t0mwTe5GHvMcPlulkvvuN
Zdu+5Gis363fKdNrmCwbvwyRIrv0o58gPxqkeP1tzmqPdb+l+rCaA/ukwkmxoWUH
p+EBPCLDjIbCyZL69di5ClP1Vj6gMfFjuhvZG60EA0FfSobcWkR9LtiQXZH4fuJ1
iptfprDYZFJr//8VVB/3W5SVP7w4p1P9h9p6ElqLJkiEa5LbSi2yIsvnhAEYFD4k
G5J4kDr5wIjuabef+sD4OyIrIdhIkLihfnE9WiDg4edsuRyX5JZpQE1PkPmIeCEE
TcKc5kibWbrDSjkiQm/DEzRBUsQ7R7e/Zoi4G9Cmast/MqEFAy0x6veW0AqCF3WA
q4q0tRMzqamxcX27ABuXCH9XoH6vY/lW91hJSj8WdKvtnxmco1KEkudS+P0iHqjC
1YhjkbHvbC2IR6u6/UuUd+P/mvxSK0knFmegSto7t8jFQCSzRrdQQyGl/YIzEF0M
rPJ8BtLopPXsUME7Zi/r8PU5zq2Foc4rukbSV9VpgNTOpa+tTA5h9JdZaZiV3WHP
/6MnvQUcOcFvtE7bZvXNbQQTHpBqqg6ApkqAcmuVwMAUG7ttVjkWwq+ptsdumsiJ
HmhZnW5mO7sWtJH3HPMapeODTidWvbVO4YDeG7ZjB29o5imOj3oXsrRBluaD27lr
MEngjRq1h4OxUlRxOckqoSPG8HDxJrBefHYnEt+RJzQ10KC3HwHbyVSBPxzpLaxf
0kcFOFT4F5OgmRmMO63aC1u73Jxfy9k8kjaxiiNN243+SLQBlCE9kS76/mnmkeJ6
KPHQOAcx0pHCHX8djkPfrb/cUILqaad3/pWUO87YPt97PHS5jOOCRj0V2/ZILkWe
X9cB4arVltvCRWmt2JRF9Gix7YoIZnVJdSTqDgsxTWtkf3jxrqBv1hUNMXboHaaE
l6NHI/ip0P/++iZaRhz0DWx6cYCUslW1iH4zljsh/BPW14Rf5JMb6zLzKY7Rm9hM
axPrsKtI7ABqXMF+/5eWe47oyn2Yvu7bfTlyp4+/TmUWQECjWUM9OnT82Mhad3z4
aqNZGZ8wGsL/tp3Whaj3oQt0gJBc8Ps/FU112JPWBBYGgWcsZuNXf3FpPiEg1fWa
ZSpGqR6V7VkAl0p1CWVglbEFQoO4UsJDmrT3PDg/ZNzTNQl2UEhL9fYLgKlBxZ2d
9Ih7iTjuiywZvNkJZrnuvgXHVpAlesj1g+2fq9ClibVwRJCOU5Mx6BEAP5M1MaaM
5luLotPP0o6coi3ATLZMJNOWjLLsvz+j4DFjohekctqQ1W904FQj+hqL6GzTaqKy
Oh8tN3GPYYYl/l1kUM5M59NVrQlAUX0bNMlUzK0Z6huybxGvDcK3nbVjPdzs3uIi
H010Bxu8573Rojk1bnYJ1oCazGAkFGmggW5DMsDyLKElbYrerDxGf5I15n3OxUzs
QmUgwMMkGqdTmbbSUaPTiATXYh5pxM0hnSFsS2Pdr04pXy+d2yWnLv2ytTWzg4S3
b/8IYuA5Kb6rn/HBEYDTK+fbZD4ud7Z/dmUnOxECdQYvdQAiksDKFeSya6CpNkWg
f/HDs7tGuVTlxIUdSJbumVQauw6anWzbpgc4U80BCHQe23rJ4cYYUn6GojFnWhl6
ndMLmILGxL3dADhPIXXnHTMkPz7rov2UZ+ntCqLwUzzBLPoO2qdDGaxWtbCIybFp
y8A1c65JDHhF8Gth9XWziqa+4MJ+pJapRP8AxAQZ9fuNM2qCVsZM/ptEaN+02T+O
U4+Zm5riqeMYo7SrkN1f3fEVKsI2UAPp1/RkiFpHxcyPpF4MBNwuL7r5bhck99ac
Obhpcfb3CvXiCJzFY0fk6dhjBpcTKFoRuFnzw6RCiIyGUglOeqZ6Lb2sEkoiRZxV
tOCM0N95LgljEtt7FjJJ1rvyXhG2+fA07+Hb1HvEh3xE9WhYEZ2BgLZYcIy6J4/P
mon4iyE5pt/5N2zFw1RbsZ4wqHLFz/aL1aIYkz67Ntr3aE7gxg/WddcJ2eXtNXsZ
UpDDvDf6t8yVtZRg4aDNHw5sF3IC7nxjWud17TYSOVhaCYBJslXGjxTgZAjZzaXn
5FsOOhugYuaP5OkrfNtY4awYui669mkiDIOa/mUazyEcOP+ZWTCHw18Soe3j/WAC
x7NYjifEmT4rUXGW0dPDwpeKSF+kqoA+JWafIhlzXy45bUBJNe28RDrQb4Zms67J
1uO+XquPxcLOpKcbyGgc36DfG2gEpusxZCiphaE0K1krVZB95tqhC56UalGJCCEt
+yLMLbzdgQomJ1YxQJUjDY3K2EhAPk1Mh7EJI3BYRJCcyfX/6W95Hi744+UTtx7l
zX+fkn/q4Zi2y+xSexZuJsTqZZ2+Ti0+z5pAy9BPQg8Ldy1sX/lyt2yCV7UobKYe
3xNweZHJKDEN6vMmyoXn5PeDXEQCHX/b6jry/qutq/lPIsM91Wgbzvb3JLT2xaHI
VH4hIbYcSFxRlmBu3EZ0lP0kq9l1skBMQyem3e0256s11zw/GZpVkGxjFthJMUYr
SRSdJktJqB6bNupcdadAyzdS8zambKLHCyGZskoHjJidHo5SDQGzKVHwiE0PJpw/
pYaSBYPh3FlWGz/WbTkY0IK0aUliWWr75I8ETsBASH3dPC7H2vXdKzsyd937UdGg
fmEypsiwatEgGDNnwrJnvnQXhDx3ioVrDiD5Vb9b1maDJIRcs0FPcoYADwn3+hLp
RpPjhEXoPNtJT/fMqucGABlY0dFYgrxo3QNjOzZIu01SG0Nrbva6QbI0xh65wnWZ
FxqkttZZnre9D1JTtd/vRUx5NFl6uhdIZ0mz7c7eojNb/1M97GRUxiEKc5JJpQ95
vwPkQ3OTJiR0agH+IO/NGXoCem+Z0PPtnEmCOdUaYQnv5ptV9+DJVa7bkRHB4rez
BOLGX4whpS7ofJIE7/O6GfGfljVbI33elxKvfA50Kj93BYEa3E0KanIH4t8qI/ZE
NBSXoi/cJEa/Na0ULMgblnKRNt5tUBmsJd7BT7g3AtlOJ2lzVfMGVrNMc4aUCXVp
/vp5Kw+A6Hj8lVY0JlHwaWRW08irkdDsJwRyye5IIVVrcNspi8i79bybPcNFd6LP
Wnc1YoUp3o2VX3iDFQa3fKeXPVYIJvVIDo6HSpGaz/x2RoipIS9IGxelNqw0TB5b
xTjnC1V+AoWL1WJtQDA3QWNOzy4faTFdKXDak7xSOp+pDDngwYnYLUGnIxH8LYco
19feFJmNO9UvN1EiAG/V9GxQwOYJKnnbm52Ko1uUL/NCzMERJdm3FYP9kBKjhG8i
KeKkWvfHwJT9MUmPt65rOy+P0M4UgRcHxtXsIFLLmzS6I2sYCRIfHLOFYOpi+uQP
pNm5PE7SJGfowwFVWckxQakPZNc2/rB0brorWSumtgccu6bZinNcpamznwmngMSg
UAuiGgQFYF/WAYvst+AA8Q2sI+1IDjcO+sZE+FmxVY2f3iQOpkQRApH/izpzXIk/
dZ1OfW2T4GOmp957DNTEs1M3n7w8pQ1usTvz6aIgoRs/mvDjQPG6tYlTEUiyzrw+
bDAVEYxDZN35KDhUt1tnegpY2Jqu7wcN7cka2NYneFKeO24x5dsVBpP9NC2yXJeq
iC24mDFcdsZijkncwgtuV+ACTU1dGzTXk7ASyh8+BxJzb2Sv+s+hOc27Zz9J2kvv
MdJvQhMv3Cu+/8lLEuELX5QE/rJHoSr+XkAOqBBlBXWdXp4JhNc+b1GNQoH4wVld
/hqOiqusCcaaOWETKUpSXum0RBgl6eg9yi9mTuF24Qls1wetPLUGXbcsbEbZXdIk
o6as9AtgBGIRoDJZ9oPtBFDn0ADRhbkIU73nAoy27PrEt944dHUDiHChmPDRAJst
ecQK2FXsvHt33yBRKRExsXpzStf5Hq1cpCmbKh8PGmh2ClTWZ/fbLbJOx30wo82v
fLcqWo+4OjP36BkaUG8jHqYPyTwaEuKvSsfl4QM95nil3bZ1bFsb/3ID/33bRMaR
+V0poz8mBdzMcRaokjs0P44GmMZEJyt9MbztvbRa0b+FRdEu4zomDMvCbxm9iWcx
6t7gLccQ2mkx9NEKGc2ojP1aFZt9wnlQhQIFWyVuaFlXSGLEWRyEbXei+iSyiMHE
YMVXxsprh1Coh9WSioxGmwP7IgAB0tmIKl7Pq+IqOB1tf6ANgcChCBWZYK/lHPi7
pBd6JCmuQDlej2RyFgFptGAAbGxm03sOHdgPbzCOYRU/vye6x6UVlVinoBBNicKd
eNdKG4zY0rIVmstXbFg9r9sx8FsQ5iqLvv1ZIryXzZC1crd30d01GKK9vk6UZ3vz
bjwFhlkIDy1kK5TemYVctSqTHhpFFRnIAsSpDs9W4GLnGOA4Af2oApU1Sy0lQBfl
n+y4FM3tn53hbY3UIXDZWEtFe425dIaXypSUKffdP5VeV+B1HY57KA0Bv12VsWxj
ZKQjH3IZHIyRZnb9VuYeTxl9uWBQJAaJP4ffY1yylQ+cirarRoqgsFALsHitPcUb
lTmXJwHD/IfpQaGFYhVEKb4SU6WVQf+XDHrlQug7daY9SVrHLgbdzpXjrN/TfwkF
1soFbMWhfPallp/5SrE0SkHTPhwM1IPebZqab+5n3RZ8gBw5IeXp7aG1e4Gi7bi7
LLtaRXlfIe2IgNt2WZzDLgAA98O0cYgcGme8Bewkea1lvIsfLGjQBVnYAdaeilfe
yufzYjessjRlBr3UhSqmtV680bXBgpdw27pOE0Dax/FJ2PNl07iTqhFqaHdz93ma
H/v0tN8W5AKEsiqmIQxtn5qYaC3SekuGYMJH206TXYXXZE01Lln5OmEeuqr94zD/
lrXmIra2wBRmo674yN+aUOTZo81TpjGDR47l8eSvnFjdzyc8vYOGvGrGhsWm+wLY
rGAA4BKdy6EPELh4gjWr+AmP2cJg6GHDoSNJELsLCxrl/UaZwoV26TedNfD/nmzr
D30A/QMDqiSYG5or4/i6m0DdNh3R1Z4LzUaZuIBzgSTr5/cxRr8buiMxRhrNLzsr
ymFPOwWCpXpDg01uWuK2EqoHz2ZGSB0Mk0am4DffoQzZtW5G0toAwiUlxWIYf92h
p1ZddZ5q3sGATQr11IZplqDKjHgMr2H/dTEIJ9kBgnr8z/j5Lpnw/GN9bjYDFzRH
NhyRrpJcr3KSF3k4Lb9I9IKnBz+/QTPPk0oojMp0+rnPMeAMhNtnKQwXsatN6fZm
5ambd07QwNZrkOqcHJl8pNx3uo9VH0gNrH9rWLCvOgigyjlAKcUXgWlU+g9hUQNT
Ebfx82auuhRfi6HGRXsxo3oGqXp5SiawB2ZT0HrVEbldGmvWGgs87btqfhduqlBZ
nIPFL9PQ0AnC0deOGZEZn8m2h4OvhV92rUDoNwqSIQnRsOK+Cg0kIk6egWyXh7Oe
5mIE2d3IAYgWdeUOZ+TjUq0hnawoCYke5kCEFeESBUK/kDktx91V1lkGYu3TjjiA
AJK3iXp7sxNLCN58w59Uxfdowdghj8+AIQdGDcj/KDJLbe505GT+tvSAy1s4/aI9
E1H4NTzzMbOotIyG6qK9U68CDEpyseNVGFCGPcncmdfXM/PpiNYhrhLlUPdiB7Uk
2tlk1+SIs9F+m+1Rp3H+89fYcfU3IkgFditD7eHJ7R5B3QhYNWnm+49uMtTYXv3t
eRv+vKtF2PoszopDPg8Y/CAHvKrz5C5/TyJdP6hAX1DYDTsKNU4z6qh6B1IAXUwZ
jLI10QmV92Og+GUz+fEkMP2zxyzRYJCfzaypnNoFExhngaE1WHBPr2dxFOhCu5h2
o32OmC3eUb47fNzNT6tnc7+Bycnna+CrIarU5KMO7OQzMxOc1G08OolDIDW6HBwE
DIkyO+PvNNe1yqBJ/z8xSd27AXlg06uFouSTuD3doKQ9E8SsAnT5vYcaZM8LXaSp
OAUdDRr8D1OJVltZ4A1JKR9gIrI2Sd+2fY9hCsYH1kjZX5YGjMWYYr69yeMZblvm
bCgMW5w5+o2OEioRFDC7Ra38shAgmWQl2CXiOKq5hU1OP2sgNypiH6qxdJJpPNtH
2V8fnxjkKELfWDKS3IFlYv8heTu5x/0pDnyy2Y8uioE993ALiTLtDsldD3TSfOv8
tvLSfS/Q+hT1QZ8rk2qYq5Cyr6hTQ5Ot+DXAfY2u7ky451H0ihJ/8EdW7RVtYk2D
wivJ1qy35gsHfc8KKnIY18C+UhWXW6sgVg5ioC+nQNl5CPgUbaAeF9zHUGieyv7C
/mysHF37/tPZtFpizm1XOmFupy8HlDQ/OhqYvj2cj8soISejU6CSQ5ZQ3BVRehC7
cAoou4kBWUNCqOwpBOfzYaN2FGs3Ne70BnAvCG0CDb8xCn346WYnv0BLaf+Sjlsx
7GKQB4xCGK1WsNredK1IqsAxe/cx+7soY3KusuJtjRoh26SxuX7QSdPVJ+bknU4r
ANn61bd2/wT6d3cCmD1yJd0q6rQ0g4186LfMGZI0azZGeGvO8ReCmjZ4i79JR+4j
e+z8EVrbBB0FXvZwjroNim+Y7frK+9JepKPAy8d2Wo+rz1YXCImGrxBbq8E0Ujjf
bo8MN2tKgd6ety8j2AFIriSpIZHKuHWW/UVp85nBN2vr2j0T7+Fde+iTh9cquM6A
xhNTWzraZ4NQeaEwoEj3OnZJP97/rIDItGWMkRhnQr2Vljv4cfy3Bd9ktM+vjW0s
FJDdmwrq3hKx2L45U1wZ9XIh2tqQ/cmRseQOlZzfivDhFzTEpEhfRiqCYK1+S87D
7kACVVwwdYYVGJ+/BE79OZ4GQf+YmdpuQUmkLRwrPLTJer2bxPCiJ8JeMtoq87Pp
fLQiGfKO2Ovd8X4VEd3z7tADcxObF+mK0+TLFym2XXF+YS7JtYBih4ROJBl83pi4
387NnxrrDioxZTNuRNmeXKt63NPZEHEumJi4IWCBSf1z1yhk03+HIRrycSX+d68u
40kkQW2pXPrSR+n5P8uaA6F8as+UpLMmjWJuPrn2JthuGpZLKbDaeHV9kCf3qJqt
YnEDAT7clLrB/YL/jUY462thwSB0fjcHZ9KmhwGiEtneQj4B0kGAcRRLsiVYMvnz
1A6kjZwtsaJvF29mRtGcw1guJi+XZYHUmrHNTzGNWcuU3KV4cv77GSmFq9f3fG0V
N7HPdFOMjDH5YtmfXN6uhWjtoHwqRbERUK+RyG3i/mt/LWaemqjWMjejAoZpAjw/
vKEYsmVTv/k26CwmNAoJBJ6kdUdMj76n8C93LuGUk4m2YpAK2ebwVHUVaxZ+yxEn
FWAmhWHrV07KCsteIRuUmrUvyC9b4FTHBRBoiKSMxV4kmvLfppEF+wSSnSYE2uLs
JWuqql5lRl/Jbm105jvPa88RwLs/D6s8Sh0N4AmuzrKNOcHn9BvaHQT00aLC/sM8
O6NWGIi1Y3mtifEtd3E+4lBgskXBfn5Xxb/G4V9s7lus+ntiS8OdffZe6a+v3okK
hvf1Jzii50oW5lghBpmkEgxKd6RC6kjzYJfaeGSgZshA7tJQADJhofVbw9vpmoue
PFyP03PLZdBaB31LfEYEdvg9HuSTaY9UcVK2GfBCfHb11abNRvAuYc1S3MOQWizo
vgQMQyTf7l+mNbXpLXH2gf1sCXSP2K6FsPyMjA3CxLS6bPuYE2a0aMSG3w9WPz0X
l8QNkTWCpLj6XTGKvDRsrtOLzbNiWou3kNlHrt+NmUbZkgFhiUgTYIAKbI5MaU3H
hOvmkhzRyam3345wfiwzYihV8Yu2IOmKPxmTne2T+LPUQCeW89Sx6Eq1AKH2AFfm
hGVNeekDIxpxIy2P5S9fExzXORuJUrNpCL+PzO64LjzuDciHBd/huSjZx9SGmsRT
MwY6mTwKaqgvEFTuOgdYNP42oOxAT/wkbwpc2zHmPuXqQbgylPr45mjYxFcr07L+
JUmLXgT2IjtJWM/TDdZLwyEweHOXTjwgcLslfDlOqUZukKcm08Z3+h3BMNrcsKEY
QSrbWdp8AsSrMjtcnS1j59IeK91+DTimqz56yUQi5B+Oe8FXOe4kXyuybJwtYnEg
5OJFn8MHH+3u2Vc+rDJg5mD4HXYocQDJljdtvOEX3RDVSqTXaIP13tFmOs0JJh6u
34IGzjbeXHZkAxJyJVTAiHrDWiWmGEL+g2ae+aNb7K1hod5M+o3IYzYYvORMBeSd
Z2WGZ3O0xl9o4gcpcP+eqidzefUGTdcdpQkNXHAA4lSb1wdt84swQPfA2v1Ww/p0
CThqp2cSG2gLLFNKlkygT8h/Z8jP8BEAsoVxpU17DVMXkamEx0o8E58o5I7reUrw
s1t38YkUshwte32WmN8lfaldJ+vInc1GDs2XbjPNP3E0tszm1Ychx+mB8tgaaU7X
Wx6L3LcjSPJVcjZTwsn9oIaGGTLdgUHhybfrv3HMbvVStlEQfnxuYPlq38zdvtU9
rJBrv8lznVAqiKp4rovDz1jryENsV4GMHEYZkek5VpvJOqia9ZbYWuXDQ7RAeX3k
zLvKsZoIxu561c4Nhcr3ZACP1QTMqwNXxsTYJGXAOV8CEguNG8As7hKJAifvVWV6
IIwrqC+l4P2v70OOU7hfwPxvBIpVXsJmvdyJOhsRpLZnUhYmWNcVCL8+2aX09mQN
WQ1v4OEYoJnWNFzpkRga2Avl4JEk4oxVc6fd9tiwk8A6OAavtnt/XM25wkS2Zc1f
omLwiPBPJ4d/vnl3SbiU3cB4FS5/zJfPMQSDz0w9mqWVid8UptZivfxSihRJclg6
uJGvSBY1/GwMNEyRD/dyPd+P9PdhAwTvzBTkdxqOqEVKytJfTA5oj0rzjoE+47/P
vWmj9kuzoqps3vvL1vCrmtjcKFFEOpPAg/ER2+x22z6r59Vm0zQSACx0/4Ixheff
HaPPPlpKRUXcbqFTCgm7TVrKyPBJR5sMBGg0Weu7tfjQREV4ET0xeIF/t/OB7KmW
cCGe3G/SfJ2KCtkMGJeVuvrH/AO/aDMz0WMuU/28E4FJBmcy+uSEhWGFlpaR0Ht7
jO5sI0uoRvKNBKe2V0lm2JQNQV94xvlNuojn8Hcz6U1dUCNfXU6FI3uW/TsXq+Q9
hqvW/eBcl2iv/1hKZsW17rE9dE7081BwxEqKeHFPDr7d8On324upnG8NJV0ftxyV
SOhcCyZJ/Q+dtXE7V0Cjl5muk+WRWQwCGAckg63ESS5rPgjjPI94iD9A59XX47Ml
AkPJYLoBETCP4uj9CmwKx8UKJlgdo9jwjVg/4mmGB7Im4iCEp2kg/qjGRfNh9Sjw
CQuasw0xM71M5akTAddEVpYAr+cqTJMVs2C7bXrkOJ5KI6eKglI9xcePLNExWEwl
L84mfD0SnvXT3IYb/6KW4kyCngDr063qi4VY5Wfpfbk6n3RYY6is3ujtz1QEz0Uv
WzAPuipbr88e4HvqknEATwMAu+BQ6+A5m7jLRr9b1P6IMGe2hFSjp4kN8VHXc9Or
ctSOw1Y9sW6nDKziQwRA/f3VNx4mkv+DB5sCG89L+nmUNAp7rAhyzcslRR2Irhaf
D2DWsQ1/wij8Lqv8c1KTl5O5VSF5xwUw0jwmxtUJkkdrKsD6q9sIZ8j4Wvz+CnCd
dNcBDkGk14jTk7jRmRo/PeVsmtDxHHiIOODO+gXz25j1u9WNJqDwC0cGx1mOK7D7
gX7370gz5gT+QYLeThL1bsAGAkMthHNGzi+/cBswje3vo0MO2+hHJSwjGuWHfZCt
bEztdNHicBERFdi434EpdiaGqkuJmuddLSCjqddmoiZCkaVJCZslcBEf3UIHe3i/
dm13wUxC1v8swM7NSJjsqH/mJxhXJXd6vNrvNLil+zMWXo3/X/5jdS77N5H2w9Vs
tdhrq6h5kOLIavo8V77boFxxeIH1O3bBB4Dr1EMVDtXWU7LqrNT6kV++5obyDpn2
S7+A1q+KEPgQUaJRrqcyq9XGyOisn9YdPHkgkaSyGt1Z5otOkUFb0zfX0u8e3d0B
qqMOObE7gROo3QKaulDysrITcMC8W/Dg1utECcBstjUvnH1RPGVvEcOlZY8aMA1b
ufnUd/VYQ+7NyBZfwjcHfh3P+BJKBU1cB75+OkJsse78gYOOoCfmo+NaLvfntQDY
VrL6txs8sl+H1Rz74FmltqgdUdrZiEGD/HQyy3sXgqjf3YT6Ny0gHDnAQxBzjpTS
DMAA2yofa6ozW+AZNTH+KTyjcV45yuBw5gVm36uvzsjqCMnq/r11rhdxIa9B4hr7
Bma/WVZBvXxGnsv5aN1DwvqILqGLhJnQO+C57UiV2nik2DB/E7VM9NRu+Q8nal+K
O2NjLpQQLkDf4iPjfj+h/vopX7mIVGyVjjFGFf8OGq7yUZ+UpbTHt4CWNpdBBxot
vG+MeAk7dWt1ba860TMNV8cDjeIhvYcwY8ffR/EHi1KNujxGLIBYHLSLvrrmUE2u
hUf7mw1O+I7knWuik6m33HrGIc7gTrMPa9ODE5bTEB3mQrqg/Ih30eLN59Tz5xUR
4DgHpNl6lEYXtlIMu/C6m2psEFJtl0t8XJQe/ZxIvsC79tyMctHi7VpcsBgmxg2i
NifcstjNIxILy48T43EM3D6nR9DvO2Xqgt5jQQJwQt4ZwhjsZqOqI5ly6Bu/OrE0
HmZYE0cV8MN8O75fX2IOONOerbcz21h7b6mzfa6t7PPv7ZtOgythsglZs8R/n2Uo
QZslDtpPpZHBXG1DDcIboVtbbWKVUpue7M+juwaIsOFQxTnHgVK51BlC6auE97w8
sjUYrAIvGURWQ2FHSLLPriBTF5mj5KXzP/n+bSCM1J3vsrXRhkt9b2XntNYoMAbi
Sd+ZCY1X0iMlTMhZ6O+vbCUT9vFNjQl7s/HmfbRsps+3BLVxPNwPOB1pA41+x2yl
t7pAql45r8D8s0qb43zLmooMr44EiiwSXthIzyoi9+VXz28NcUCuJdie+gFfqH2t
RDzaOghHTVFePHJ2jYvbmNndZKmYRV7koPlyTRQcglYKX5bjo9jfFIoJ3JmUsTk6
BDvWu0mCZmkIGUjlJRy/v8RXHczazSU1dfAtsR1y2Lu3EnqZwOdAjfy/s44sRuu4
tqoopDEZfVTLxTfBmvTmt741NOQseXSQB7p0GGAJFa8mY0RVfmgi3yjTRc4Kint6
eCvLT31c6MZksVByhkztI7WDp2oixfGyMMSH6MFkPn1mOUQOvjOykKDwR+u/Qipu
swK0qwqsk33rvb3zaCeYE8jvxqd+0XioYnlPs6jvJ8ADewMtJxOGVOK4OzSdVH7s
5EDolL5Qe8RVw9qZndyGhRNs17yuONRwAzMVw2ApL5RufT1yx1VL4gvdYSW0byKU
tbOzUkI/2mq23I2MN50DM1DXtVFTUmj8R9UBzL3Zm6V7JQea5tUKnmu8dNpzKbfo
0umr/mUv92dC6OfxptqJtwIaPOmhPrRWi2xu3Bey5obAcLdKgUNEYb8HEgS8+8aT
FqF2QqfpSLs7QzWWTvsB9E+kC8kCoy+HHQj78gYsdNzaPNZDTxwj48ESQlsCwlEx
x+pc2ShW6LjBsGjjBIGGQvQNWBRabCColYfzo4Smb2kCAhnd6PD+d6iFoVNd/QgA
3PJs7J6+nlixmUuzpaBGAp+uTSt5sSbiqiFOnql6niUvGDkcpeMOESZ50OjV5JjA
h5YCyoiMQmFay3F3m/OzeBS94DDfzMVVsuny9rzlw8HXHElo6XbZ4SDyNgSFfKwc
Z1Fklw88Uvae8ZsZH1oDfidOc9ixXcIkRW/njmCAfocKnh6+C0BKvRE/7kgkp/TG
dCZFgp2XcLDuFKsLgpJg1gCD52iD+MdGadcGAKLupVf1Z/1cHnVhWIhHqd7uvBk5
G7CQ7Y7qOE/04U2nqNfk/ieZufNl7r1BPsaNNgjKH7Z2DUFv5qSe67daNg1gDbih
ZQFrQC9O+RoqLCk4BzXWdjPcHEkNeM480TMIeIltiv/uE7iVYgx7ah3KQB2UuySy
LDQCC2XOFZtadGKAXTEvZd5pNRNJS40mVkdAtOgkz7FxwGeru0MZdD3IBYrt4awL
AXnNdKSgCnaWtUGuLfZe7SqvmoZ1JpcqQe7yRYHpwwasCYK8+sEIOah94rcfPf1j
a6HCreOZzgU5IN8QyTyDJCrh2JMlgKTxfRVGmxSnjkd+k2sVhknAp/2ZFs7ADJtY
xvg9X2Q1b9Se72F/3iy7jdr530dHCrcd0FHZ9jJ9gL4z0Ac/wxMpWQh12Aug6VL8
oErjzITrB7JzTFbG1zUdHa3Z4hEwqtLbU50XSk0NBNIbsLPeb0TA3Qf0aRL+Wmfa
NDLmOoXFWdsHwpVWF/0MjSGlXgM/pZ9v5KU8X7v1ESqpZGRyTtlAPQEOtCgIZoET
MVTW+Edng5ildAHf6NmGOkGB9IT9XDigC2Bsa7vg6u4f42147rGf9rLyfvWZfDkA
kDzpf1p8YhLbzcaFZ2nbcgLoKpel5Fl13Bp7U49gg/s/RgxIwI/F6VkLhraj8VVQ
EOElrxQ/I7ru8O65CKRttum9JaMlLI1gpBHWMYw6FJGSxFzsoH9gx7ZVywIZX0Uy
QE6obhhk1KfxenOlFN8g3XpTknSxmvhjidG0Ex8uNhPXzmo/7qL55c4RFxi5+VsT
AU/8mGl0+U+J6GEq5XnwTVq5qMpRzlsFseJkMgLmi1irmkahsD+kvgvHfj7EddKT
TEiHp+BSV7LOU91KspRivCmWQqmnX3UfL0MMxK3lWWeG56XW9dVCFRTu3EOIlqbu
jIp+ejS2uy/WB6Hss8zFEnUhvVtzmcLTx5+DOE7EUIVLqk290GlzECUlmrBbT12W
7nvAtLyDGNODk8l3R/jrOfFR9Mm18E8dWW2O/yitbasN2wopnWdNjrEDepLKU91+
xeWEyFsZUvvyJhjIYaN+LCB4ktH89yjlt74MlDjgjIFJNNo1HYvrOPtcBx7amj6C
dhISxbdU8LhNjTiljRWHwKvEOgxHp0ljJ2ehzvQlbewercK1DGPq30XaLCD1KYKa
5wasDJceBy/Gp3aFv+AUFwyMrNN/NBYO1A5gJKBRuNqku/8YP1zq8T3D5bTIn8XC
AEgF+IzhGA60HHo5BS3q3zcSt+/xRmjeoRCg7mGx8G5yoIFAxh8ZK4i3cbPV4h+b
VUs5fxirsIIF9jG8zHvLPSwnkS2wH/0JpFuTqJ2fcsUNJRg2l9NmoTWSjfF1GoUw
4q6jEY9TPyvLfIgyL13akumHv750a4o0n0k9tCYXOmgo9GpixDyaVgtSZOsZ7Mgs
XOK5dId1fZHZ1NXf4xLsbvqqvtZIyD+2ZKACemNv5vN4sm9hMGE3UKEHcpmATEPR
21aGlvD11j3Iyeun3PTQIdWpK0D/LNOeuxvOJ52+I4CdN84o7WnLS640fkZyXusW
FakZAt0YYQeUxZ3vverTFaH1X6uspnlfmkxeBsq8ckV54r8LuyUj/fyWccej76Uq
B3crelkRT9zH2pOdDEHA0fJPfpTfZApyKkgIw5JSzXPdZVCPZw2ldjFhC0yYaaIQ
0kQJkcHwhbygG+iODZJ17MMSJ9/l9CJAsqvK4w6BuwAw28grDqWCmycV/+x0v4aS
kEf/ZQLmFHPhSWWynXuLFBX2V9rX4ofCeNVb/QSgUBFZs37RLNdlWN7ZaRMqaDHF
epTvTMUOWifAJAXUHbn0wBcrqBU7IyrzokdsdNJOOgDX81np8Q6jL0kXCbBjLOyW
7ZP6QR+cn9NnI6eB1af9X/dbDVwaM5IFBMUOIDyoOzMCyJH/ZypLVab+ESahB5Up
Xb6rIaMblBpSpOqvhPZ10xltrK4tJxTYt03v2LSqO7809hpy79PnD5LP5XRoAxug
lEd3fkRnVWo0dw694pB1s1U47igp4SXAh2y3Q0UsbL7EGuygYQR1WWdu/gmVUzk8
HmEAYTWrKzPoWYO4CkyX/tj7RQptoiMHhpg5hEyYMgw8w7yZUWDc64KY6M3Af5l1
8jiY88BxwnJ2iGXNcJYNbFpdOhR7zSrf1Wn7gXLGM6L5IeyYL/8ZaAQpR7cecaW+
5FAwwRre2ICgWmpvZZFFBrJvVOZ8quJEFkElv3jQXEXOeO9Pegn3EGAu+HIJQfwX
2fh0Q8nAqKjVco+9v0biAyVGjR0JnhwqF1Hf31HS27DplgCo9AeShLyCRb8qqVCi
PJKEgqfOQ0/0v0nftZ73lE1kVOx7NzWIJflVPXhMyE29w9Emi0ieNru3ANz4mUi9
yBg3ku0FIPkrkTJ9aKom2pzEHcmla3gujWLt0aEkHtG3DgfxKd8z/tSLOTrK2j97
shVcKIIRYbNkqTOAi5m/ZhJNr6xCgvt7RxVicoWf2Jtg2ZdjC/93x5eCxeisLc1+
v+7QKcL82uzg5H7l1PY5iDui0Iqk6pKXMQgiq9DLW4Yw8ZxlDRS8e4gdht9l3nKO
lbdB5UysdUUyl1Ok4jbIXW3GmKBUJRm4iezlnfHGW/gtmm8cX3sTM7HGNArS2Vhp
SUiFtdj99+X19AhiyWqMfpuJDFkXAY9ryBEKV7fhDy/dNvN3ITK1Ww0BBJ4UwZ1t
ra/N7v1/lxjuGqxCZbhxWtPwu6e1Qn6L4UAz3AZ0pryPqtU2AJX1VF8i/FL6lngY
b81vXoV0whBzQoA2QXSqsBZrA09XCK9ew8DcQQl8yZZHT/f7H5rOj3bGUinHuXSN
kWqJO+BgCeI+i+cYWSRbp8FyVR0etLg1u2Azg06D8WooXEx0IAQtpsjRmon0/LqH
J5wEux4+ar/yeO5pUv60cmIbiuoJ6p9iC8xA1bjB+2GPFcLtPTbM7cYfwH5g/zWo
3lMEt6Mr22jRHd+aY9TVkrFwSUTxFSamazQSKbNAuosyAQvg1xobYvGU3slRgztm
OUHQaBgfVOSJzQwte5tbLEVwnhlXCSyAJOcpAddvAS3OmYvH1NUejC1tz94meJlh
LiZ0Dz666O3OY8DUqhmLjB5Q9ZpXWPu5CXkkhCyAvDrdcH5VbBxFYUZ9NYy+ZSCp
TNt1NPjqi5Kss01VOJi1EO3QimpMebNGSsKMH+6RvWHw2JdUtcbImNSq0yu3sOV7
gbc5/tT7ir3AcorzrPk1jjF73OzY5kiP8xjrRQ2Uo3TiqWaWLdS9Nafpvs4tFYGB
ABtmJo06mDZ9hK6eNowFxhn4ND7/nWLU+j4e8U67X9BT0LssLlP+7PxLJujn2+rI
o3052KEIgbkbat9XjF01UQ/s3XmLmqraDQ4QGu0aNHnP3ffdL0OwZl3A9CEUPQKv
GCVdSIUe2cqIJQWS3CLYZjon+hkJxdPCtkblI/WsQyKugfnX43TbS1K7IIfjwjJO
aT99+PcPLo3x2Ft42umoUuxFa/Cpr308RKeYj5NeyRGa9Z9CKBjpir2h3Y921Vqp
Y//Xr1nLrV+JxG69943ijxvVX8yKh68cx4U7KEjIXL6cj9Hky/QzX8CgVHLUXUCz
ZKzAs+hLbAEkMsG/o/ODD1lumKxBGIyI6lUcRZKp+kPLca2qqFBwGmapYrh1sm9W
9UVZq5/M8vLTWE2wm0T1zNWMOSR0zu3keEa7g86LDLM2h0dGDWQsJ0mvc7TinVBe
a1nZxEjkHOscLW9slvZzCK602UTQgW3+WQJy5ocKUrD8vyDZWFDUL4SMYetJN52o
YooUcOhvZzAnJqpDTZEWtFzfhM0qIQj8y8axkDziNDrg4e2URnsBUQQLx0xbi65/
CJfK+xy2few1PJwV61ljH6T+MeB2rfaZxLNFPZJk1RI2xpRzZ+0Q0raUtbVuoQvt
g+oQvkE5tSM09Lmdijhf7EyxkY+W+IgkBw3gHaPpn/F7TwPp2pGzxiVdi6ugB3zn
kug5hXeeUFbTzUhCX04+8ypfctJxzt8/W6X4A/Gp8iJZB11FrrcsrcNHHuherqGw
IRTyDNGLIJRE+4kj5VTWfYwM8m+P51azEMBEpxU9w59QUpZ56QRgQ/6RwSRo1m1Z
KQ+o3HtR2hx7O4+o186bw7hKsOjqnan7Kn+FbXVrnFoiLP5BwEphxPwmfZtxRhqF
8ayT2Ul2pepaaLCUxgQTSc+IVlHr0yOExQqvzNklmuwHSi6/aL/ZBdsOGmsMCUzp
euAFvl12kF/Zeu4mdCtP6OAYhQNymcZgIAmHTa+50yDrzFd7RA8ZptjoydyzSaaE
1B2fI4B+ba9VPPGGJsLWFQ1dQOuv7JLdX1D6CrNudu1XLb7H+htzn4LFebYYhWXs
1t8+Wx7SwzPT7HOodVp8swFw1IKDqTx9fmOW1lOO6pgPrJP56RE1+ZDyBJjljnuX
/FG40wcNj/Az+SMcrm7B1JGPbdzc/pP2etSnOeHRgpcUY29m77VpCnP7lReuva4q
D5eN3jPyjlV9irEOI5dfaz1qUosf1WEVPxHD3Z9+rT4QFaDgOf0ByVzDLM4T3zGo
2up1ongmbAAQ9E5/vkm1Dem4rhlIuv+Tb8y5x7TNPVSjfwyRHXPRIN8fINd2cZUt
KifUCrkahDSUBE6QeI2Q6mDanm26gDNVl2Bybtx2aUVsIJ8IxBoicqPDP2fBgA1r
4oFQVp3XV8IhrMdGJbc+d7Pin8E6Sdxv63+B9vc1gs5IvttBGjALqCLleVkzDCDW
fzUCNGofp8RumHKxVaFyXvJ03orGvODLzS5FiuAkjcLo8vJDlMUfmFbUbKRjRk8y
gZzEpuZu0xEGUs7b1ZCKaN1MhkMQcRjwJy+OMtkUIa1XZllEWAGodb3s8jDuesEb
o7LITPM7oEliHgQ8OwddA6qXj71n9y9aUfTLWgftRyhhsLfU56S/K/dCiRBn2Zua
F4OyUfaBGwETgts4MplJi0wgq65TbLflk8R5SCgUN0NUYNClCBIuxlyjueKTWkUm
HstPbAfxLIn4jFyez+zYgfPRbhJLjP92gYVmHvqAHaIBcQfkMqs4KvuB5B1lxmiz
h/EXzXQ5dyM3dEdaIPq2+dkIrIaNKvkBM5kbOoupqhhaY6DyxkS9ly9ys/PuohQ5
ci0n5YhlLVTj3O/2WGK9jrzVK4oY41t8GffdgscNY9bN04B83mr89XDzteRD7hSj
g028m48wRuHu8GjUhm+a+AyPQqLGCVys1r4dtzuvn3ltxYNXOHzYzNFC9rD74tj/
yx2jknRj15PtLeYDSBtq1gkcND53GQaPyuYLI+oSWstKoOX4K9caqSVHVEBanK8l
hNZLY+atVZAYSVssN5rZ6FLpRlXu/3M5i7lJ16WxJ8fon338QdBz9oLt8rc1GLT5
VVsirTnKrazL5LLOXaTctrJncNOmDVBXFmTDpnHhqjs0IipZP8KMAvAw6+mWujLF
XlNUdDHlwHypmKYeoDydYbwvjuBAxT05QP0Yb6ctDZnwmJiMbZHWY87/XWcwjH3a
WZ2/LVL90uPcGR1ssLNl+UhcTn27+nVDR76i5NzN5aslwsR4zWLAedZqPCNZzdSS
bwtnVdUiOgip5NmjbeRzJN6D6vF3o41YNoSrGotnmYzoxmR4eIWoN6a6wATe+r+E
5cZNVf0FnfG5BIbgHADcGd5mqsyc+OpP5qM4Pklse85Iee9T2sP6FseXzWBCgMZ9
axmV4DGTyTjXjVzbNh7cldaNjAJYxc8SL/ENYgnr7dMcnHyHcS9c/1aDnAS2xqNF
Suul0NslNr7Y73bMwqmKLFYCdqbnmtq0lz+Ob5yCmgK8lGtC7bxXef3Sfp84EvA/
Hk1y2VaNzdbBYvlatl4sf2DKt89vaxlxE0L5wV/ZO2fhwjojaw8qrvpMoRD444NQ
JeSFDpwLZUtEd/dbjlb8banZZ4cCuVE85ufq6kvplx8UJB7JuCHRIAu87JB+utIT
lcduGrTYJSbwVIAVZQSZB6wjWeT5p40WOEkFHVHyJYDpy/JMru/e19bonXHugC4Q
pzBHfGVUA1mpCDW9zfQildHpAC2GdDP96rqPLKt7r9xlbpbDOeqEOiKObtcCeuce
QtXurkMAQyrYUUnWNfelV40gi7yH/9g2/dNWkJfipnDGrlinTWPXKL/zmW93N/+m
8C31WktJQ49F/ss84yq3CMYs/mMR9AdOrZC4kPab4Kc/XrDd24SO+u17AKrX24Ud
KxaAxwWZm60BsJeUmWbo2+TNvHpQPkXdzbzCqQqLV6/8Na0pHrfh9EpSQZ13zOs+
l8bk6KKnSBA24sywpPnlWLM2ob258kuQhcBvaP4dtCWJjMXP0glqkk2FV7bLt78x
scZS8pitqdUWdpfTtnkgv/ueph24lMhnNdASGZxFPFLXMaCF/ykgkSjMHxm2s01J
KubMbOpKZk88TyvjCyxMEjZG/M6Pe0ng7qJebDmNGtD5+/bBJAT6rs4hn8rCUDtz
tARB0l2GILufoXrYaQKJjCUbK1vXeFPYMTbFsDxbhwxDsN3slQwOhPz3jAKPJn5b
hHZ/H/XWLWdQ7FzBFkoDTbF9X1pAG9uy1SQEW9XJazaLRaGw+skXv8X9NpBQdV/P
cRNBZl9KBQfpHGUI2Ec3/ViA3KONPddFEQfYzT9nhwY8uMZPJsczyH01Vonfnbcq
u4FUmDUEXWGbCuyDPZ+uaI4v1GRlBDrPqLRqXUg2/VJgrimnbS5urJEgG2L4j28q
8+2iHpAz5quoOumbUwlArWirxjUCqf7x6rO/4MCejHlz5BPI34KiAKVzNnqVTWN/
/K50hehz/OJnXqy7WGqUpif/R3y2qL9yFz01rYsGhS3SX7rKeRkOeOgbt04Wj3jC
R6Fr6MALeRSuQFauo+GrI50Am7kX0v4yFnDYahvkKa6qt6vmZnIn/vBlFdFkg6sw
XkBDzifkZOKGHKVbafGrs2PBBtTEc1GSxHjud846Zxb30Jf6IxyliqGJgOIJg+6N
I0s0N7QKfW/xfQkcTlyVKgktuoxswPrmrc5B8tgi4nDmBuN0lLr0gFDsE/lwcD+/
ArZlMeqmz5UPLSBlFS3akkiVaWzyP8rdC/v3EmqfirmrnlKpdtQdciqBM9e4MPA/
eqdskpewL7PCkyf2nkRZIcbMBYNpN1aZfIjs3/g52CmrgkfXyOPKuXdxWrWOzgNF
0u87BVVEuCN/DlhgDx3Pm95pQKWKKXOBx0MSusuWvC1NpNIEyGUJTzRq0MNe2Uzs
BBoQG+T4yU61DzIN0cAQ04NS33ztoPFB+ZpoMQ3uTDWF+7oxgY9DIXf6lCuCtBqD
kKcTT1Kb4km2r1UY/d1vbaHYz/lJB2Y82wyKyERcwHYmOII8dsCxOqnZBAJslkIi
CrrWENV3AkZ/7nYfahHuRav4ugafrD1VHStZ4RwidnyvlUbHbpHfzwME5YBIPbsY
rV096l6h12bYBVudMeacbceImMgPutkx5IVCxTCDu0ZZYUhUu8QnQanTXmeWYOMi
q0O9E4QnVsHts4pOT1MG4HOhLdtZoQavZL47fPWd8zxQA+JT1pBn0EVA0g3oF930
z6gR5PGtwY+EWnawH1MBzulVKNcey7alqqt5qm1lBLq4bUkmHA2aSIYDEGwxX3h+
iXzKm7wtoJfMuEAkzFUkXBqE/rNffKZ5Uyxts7coAqNSzwcVwWP/qhnluNKeA8hq
OD4keeZPEb5RboUZJ+jco/Tgahx67tWxlzJjl054gCwVZVTwiBAjC9LCgSHl4d7w
IkTwgm30EXBNLslU7aaS6DHueLSIenMhRtSFej8Wht4WUy5RphNNXQ+y21RSxwRz
3wB6RMhajvexnkY11tLJr9c0xDymiIwDiw1Skb1d7wrO8bVfcKWpZLgZWvSliAzE
f9Fx6N+OXpa5Ep8IgvKTUVEWTuCbt3HMhv7eEcvBkHqDhsy/mhtujxlcaaxCqbbo
VhiYTye4q1zTZtmG1vDCBAiHiUbxmS06MQ06fIG2ZBTDW4H2FkFnhWrpGODWTEel
CKNrM3GnvCYRr4aNQbuN0NTrTS2/vPQbgFQRC49YLkeWyH1L/himnS+ACc6Rtfcj
nTFsjCSnl3zZwf/ujqAjw+QCdi+MaKVaeB0VCaUBCufFngY7F4SxLcQLaa8HRcpt
64HUuYbPWHQ5blUTH9CtiwYCDK3SBi8gNWGGhQCsMEB1Ezd/8b02uXCtpppDWCXb
t6tbwcWYeekmjC+adKeTJGHv8+drYTUlp3amAgrJddeUT7uRipzM0r5qqFiNpGZo
SiVlh1j2a2P7p7To+Bn8oE4NVUPuwkzN1UcMgB/P0BKhuV83GPKBjG23uWTfIO9X
Be822TxHik4KDYwThurZ/iknQ3x8olm4vwAOYKCrgX+Vt2BK+lDzrArN3jKRC5yX
8IPd4YH612T61ZJJZC/uECJEchnMRoZ4WcNdLX1qxpV8Iso7mV286Ymgc4iSbH1k
Mo6pRdBOQYOgAg17T4118Ebupl2yewnls5StplvxMkYiu1PVuhoHtaPTi4AYMNQK
j1FFIh3CERYdtGMlHfBxsc9QVwSYHg4PDv7nnb3UBnK1D6tHeR3IqjEncZtfYERL
mEpQcbySvU2fdTXak7/yZ9zCunPcBXavmknsNjWUXF7lWt2WH4KQfImO/NuKduKQ
y9Db6DaYdqFZR3Oz/7jFFlO5v0JeGO228AJfencIoysPoifV7nxHBDVTt7tbGPte
r5eDhlUkVxjJ2RyI5jnBYDSEWL34yuUqYVtxOC0BX/OUcrRo0FGl7/8R5raezqH8
+PgfKwNxZdfbX7ThS29xo0HV7Z7zlpHEaSSj1ySoOFBqPjsuHC5RguQiQjrX1HEk
9Cfd3SqPtdxhC8br9n589T9Zlrp2lbXr8a9aY5l17vhZKiTAABe30fAuXEViNfg2
j1LSMACIziaKIWtrvGEV883BWMtl+Tk4LO5DnM7jDcB/N60E+YenN/fEedv9fe3B
h5wPwWcrkMjIHrMWcRzvhzrvnDN9dDTgIkxjEWkyq/DkdjgrhcmygqgXiQJDdXZP
lp6ygtz1aCocEVJ1b/9r/kY3uYh86j9bOLrYb7XKqpDu88nkAttXS5lLvyXRxmLI
QRFh2LQtvPhOkR2NLFJvwA2OApS2izkXOVmrmsYbnRLdFcOgj77pU0nHehgyLAwQ
K3HtMiLsnWoCnYVq/+9DFVJvYJHQe/19FkiuweuZs5YnkBLpjORHx2T0Snsi3zab
/ja73ERS1Sn47aHZ0hypfZ6Bj7zp+mqVqO5YBynBh1wnCFu2pp9QixgalrFaTQnT
ZCx4wIViTJEoOpOhw0LF49r7qygxqONLlpbhG8r+lZ9Pt/qmkkXoBR/8OzXrvtEs
EC2ZGhM0dSOkbKN9MRGnqUaeNtj/W4ZLkf+vqBIp3sDnaiLK4/l+izjSVu8Xnw/p
oCG4wtMVy4FLUbKxqoEzIGufiykbqcL/YGBDru91ohmvzlDkH4Nz1RbOCv2Kvu4J
MEUNSChrgr347HtDahWLAgXBOT4yXLhwOeS8EAY0W4tjoabyO5cS9ePquIzpZzcB
mbpsUmJCCMhRxEHcxH6L1Qdab1M+bdgT797aqdigYQox2Z52lO/2oAkMU/CZiD0c
CB1P2gGbg6ws3REN7izlj1kEsxJdn7Nr3mAOnJ/KO6dPkwBRGe/461RNO/McVsC7
VxeH/Xl004Rra3qTObYmomf3G0hF8+mPT7Tenbj1zeT5bTtHosXQ2Z4UuGlFQujG
hkViYGZhaz29JjdDrq1lq9qeKhlygvfn7APD8WzLFCMUF4VPhqayp3hFEp/gl/zh
GK230S2OlThyysDA5AsRf6tb1VUsFXP0UXsdapsELMeuSxkNOUSnW8hqMSmXxrwA
iAOT/RPi+lbTFfQyJKnksbLh5T/x4cgqSE8cMnY3RpDmTfJT6bGFf1ZcuNk0HQjF
nWulPxn9ILEom0eo6zjvDhGJQtgcszK1Jt7+ymIeNmMLT5qk+94JvFNSgVqtsrlW
IN/+HYrv7Gx65OeEU72bO2y0NJpwS9uJ05OzAqb2ntjQaFtap7DzAMAcRPc+KeUW
K9mS80lj+5n270GH6QP2mYDpSukPvHTQhqpWE7u7KmghKm3YGTcLBGKDws3Ylb9C
j04FtmrGTVs+cLL0xhlS3mzVxpTO0aRczLz8yfRvrVN5YisW6HuFqqCJsEWPw+2v
CMsl5havoT6UFT2/br/mrm3aji78jfFZ7DZ6xlpovyPaRk0amps25ua/aVW56U/C
z9GkXIrJ34sY+jLFI3pmED/I0gxAx5TPVZvX1XoA/GLnnY3HPidSlcMStWSD3uig
FxS57jy0xLGl2sWPxIBeOZTb0Z/C+x1IZI7X7tSvFfbdwoQdj3unIH5gqKt33tG8
GrYiW96V+ALAgXxKBcehaZLP7H3A/DQF+09HUdShJLZUVno8pgT7I8+7rmpEuO2j
tUdQncBcxtQgvzNQPr7hIMksdtbzpKtalgPhkUu6hkIOe9CAI5TcXg+FBMWMnwEp
JfmVDiSZ2JbVRgb4kT0PLQ5mbNHnWrJoS6fHsoFu7NQ84jBpjscmIRlGZh3YJ3Va
xHSr2G0nCo/sa5l0rHc8JrzZ1+T3dMD5WbKVYSGLCTpl38AVU5+CK51noKDr5Czc
HomkU+phm0wOQ7ItP9MxaJSe4v1qvu2bMfzmZs3+FXNVSeTg+Ug5tvWcjwBr/J4v
J+6ON6qdd8B/EuhEAkwAGqIc/C6CIv5qH73YUCmwNhsPsmqHo81Ton9eNzgc17iN
M+AwrAHvqQzWifgitNge251tAiLknsBo2lCSwhGGBJX0CBabFdUVUwWaNkmYOyJi
3/SnHyGF3a+r5SJ+IVFa4l7loUZBggI3pLcfnoj7RDt2tGVRn2xCCeRSyCWQUbhV
vDwiU/562ErhRkHPTAt1bH1XlX8vtnKf3D1nz0Wbr5yBSXUtaBzDW5aOJQhYrCaU
AlGDSrtsfG09nVDrf2t5fnw04IELsC+vfpDyvKSg6pRvSvAAfMz2xWe238+yZpCV
aK9rlKtgwn6a9NUQH8Hed0+z6nBjPQyXvNUk0+HOkc4VBtMQMh/XVx89Gpy7oiaN
hB3sNMUQu75toLB1xenMyUa5Yw/ps7Foj+AmjeOnMmYZfZqZT3sT3ChidZPNXisR
uP3Qv7KaEI/ziiHoBOPLqzeaKLEHuWOX138zL0uyg83Jowsbs64cDHqise8vjSlW
M6/XSC9bb6Z2YodijkM/ngLGKAIL5cLe444ynWzSGGMy+ljWm2vVetznNrcB3GFa
zIDCE4OrAdf4SGDYRUTME0j4fY8+TlCuGhDVyJp+xHSt4t4DD6SOyUgaCQsgV6lh
8VpEciwZaqsjNZwr9soo7bY5JrZpFNTEi1spkVS0/GZcvTJwn9r5Ams3XGDuTyI0
kcPmml0Dchu4fUWu5Egl9rYi1+IDq7vf372HXGL88YAfL3uMDwpE3h8B0pjMBIl8
ttJaag48DLwZIgbUOXiB0NVisaHcc21jjODAglyKTjIwrOpbz6mGdVUf/mdyeBNx
JZU7duPHoeL4FYSPP4ocb2gZBwj7M5PZIXEmezoqygw+RGyS5ANFBpHzRejHw+vf
Fiuv0wHA7fl8CutgFC7IIPVBIScrlBzT1VznBmaZXOYLRwZQfQz9eLkpvmE+yNPQ
ncAteJ4FEsa+7bHlJHJBrteeYywh28MuFmIpjrye56cMGIfVal+gURyrhUF0pvDl
/hC+URyg+tg/RyHVlf7Z1cp9O1PLf+tM87KyOPfqAp8swduYzRiv1z/3QfI7hiE1
56m+4/4HQN+0Nhf9eOKoHSCQl3oV1bDDHrs37qkLBDshlGDMTByKgTnx9WcAjJdx
p7ajeLntrJMXh9j9eAN2px0axlFKShTMJXo7TxQAZZWme989KDtmV8w91rK/2rz6
H89EDcLjFW9Wuc1J5FeqTV6Y5q0trt21UqwlUcmaUkTuVNMeWpCap3lddukbtT5C
wYlTjeASRwLMNiUxc493HUQlt65dhirM3RlRBSRgaT15BkxxvXjB0cY7DqIkhDS0
gRtAEq0PqWzVG0yGlrxReLZi6YD+tGDcJ1UmonQIP2pNkIL4t/o8/a0x6yOhh5YW
kVx0R19hTEyXuvpWTD2Jy16e1g1jUUmZ4aS2whOSn73BuVV6BJ681RJk7ybU1nQx
09sMBDJINzAW3648sDydcKyMEoqiT6npaMLEWSPxpt6jFJGFQgumd3AWj8Y20GLF
mzGy9+NNEaFdp3ZzbFRoqjRzQxHlcYrjsvwi3GdMc36RPu9CM/2hJwfFXhovRBBU
eY6iFLyUccpzL2gYS2QuOmZrDV2KiQ7BbQ0WPGuzBf1Cn6LH6pfG3DD1VqfMPquJ
HkqEhP2unHRQ+4X96Zo3C0JkgdtMqCGLwhIxGhg9m0ACxpcNzx4/kpkSNLaEU3oF
I8qnQ2+jMDdVNBJRIn8WL29snAerF/nus9GR59Za20swR+Nq4AkLesUljtsqwTzL
ruk8/17vRDrzdOMB2B/mxAg3VhUZtKZ7YEGa6nq1GgkHI6TIGUklG48u9VVo1g53
OS6kIPLCgU6DvxClkIOU5BsZ7Xe/StmU/9p6mDnuxxU5XH61dqJ5pkWYVtD3/sR6
SPv3jikchDSB8GcO8CgRfMwAccTFUefoq58d1b/eOItzH4EMpwiMsd5bROYHlGvP
PQOIV3Cc1ByooXpGCl6YuCh1aL7C1FOA3iJPdQohk1HnFbmYicW/4gMvAz8lfmpM
vW65WYU/mpkPjWoRRsMvc6N1caZv4ZvY6Rh74vo9FaQ8KtrgaObfaQFmJKi+aMW/
CGLnoHPaV53v+zTlNqOR/s9iAU6jj/tOuq95huOSJGVZQbjUtvpBGoNGyJ8kzsZv
N9CXWRLvuhShKdZLXsA8LGlK0fhdDPggPqB6bwsP3K7qHKGmqWdv5F6E/nya1lmm
/pbwtb0zvgoxAOdRYSJNuql28WzEsfChRemnsRf7OVi70kYdT9yljx1yOVBsMxYd
HRc3holrOqXl8HKB9qCZeuA9zgScCcODkR50kyX/rSB5tTHhyCs4cRcl4OjVtvae
wnWEMmm3qKZDhHQYxMc/ggwGFx2USd9bAVXquWxcOZC2i9iVFSQXeT0uNw2WU5ow
mwXXEOUT9hyu6VExiVPZZx7hBY161H2+6eX3lBzFIzDAwvSoWOlDn5rVM8BtF1f9
FUSH1n3ao/jAL6iqJuLBoKK0D82toSstzI11lKx1RaHVh5U5q4Tgr2vZhPRMEwzw
5HRA/3DG90Wt+yfm74Q3PYj04kGfmJftE4SQIq8RSJ2ATnGNNv6WtQLS8JGyjS0L
MGXUFPD2xK/oxNA0vgjq1lpN38GBcT/ndEkZ//9JyKx3yvf2eGrkavGClq9b7acw
uzs+Tg84MBZVGmz2UmnyxXchdPMF2SQ7W/ffCDAi8EMTf3n6urRXkv9Cw20gtmdd
BOwgIHH8QVy4on+qXLUlnoiRMk22NHqjj79hROexnHPiqr7kDwubjd9EwUpozsjF
ZWcJNPOBYCELbXuSZ2hao+RXUoK4rCS7b7sFtQTi3jHU+HDkkPhu/4znJz9LvNd+
AFDGXSpQp00mcLJYNbn1F7VCvVYe9dKN/POSRBJTFbvk9k2BKH5GPxA8J6JKFmuR
99llPMQMRKvEm51Abig/RIPm/088v39MQZd9fHeth1O/w1fwY1aK6tVyKhi0aZW5
2cZbvLvNbfQ+m3NA2ljk62BXF4AvyE1qzmHRng6BuE0a1FT/4CBnk+ZqNBIM7EE1
Jq5wilWTVyRlscs1vUUz1mlA6onPD8cqIY7vDz8tk7EsTnl6Vo4hU6YEOhyuexlc
HQwImZgg6kH0AKD8UbRrOCGBon4otbvY4KqnEruEG+vLbFQIeSqvo5IkkulHi0d6
kmbqr5dDSXRX07oupX3sGLeIzf1j9bN2LuF2XoqUfXNLd15mgKxbv5jGqKATOn3S
Ww354bbGsK4AZy857TaWys4RviGJ2FX2SGrXA/dGdmsAd8V/VczO7ILm3By9TMEq
7np6mNFNhHoWOq4wBP5UsXQCswTCajoML7SXCu7/aLd0Yyy12tBIQqGkicxPE9s0
56+cOE0+qQNIc4KdC7cn+D8rvu8cndLJzfv1a5O2eb43myp8/JB9HLaLD7pFKMe3
szX1LYa/D27vrM3JR5N56KmOzwe5JeJfaFiUeRDJwLCuGCB6Firsl8lifD8gEWDX
dQnDH8KjoidVpK06bPKgIYd6etSAzg8u9UNkU072ga0SJlBl7ymTUksHbOmNBKTb
yAyxzsNpNGUUrKro4lNbd6J4jrfZ/85ZyA662io8/3q1PAwC9WJpDFtD2BZj9v0r
MIzp9DLg9OYYAvefy/P5Fsq6O/7KH6PcZ9d/NxoKDewNm1Ha65LZ8UPdwEOBDCq5
rpasTd2KqqzQRP79R294hmpAG1HO5QtHVs1ZHdxeKCFje7TlHH79R9I9cA4i3C0H
A7GHAzAINSgcC84tQ8mwpXWKFxmqHpmOuus+Ix9QXEj+02LTDX7ip7O/xERt+7C5
s3sDoE35bOvr1Eau0euE6NdbpjhlZ3IjB89ZbJPZkPFRYNgULAt3kjdCjRbKugjX
U19mR9VrxhfCR9YPSZ1gGTeYhUhOCDEcmP7QtCJgnJZ+cHfrGwI/uR4mk8RfS8xv
zkjgj1RWm7ZS455dsLJQvX9s0l3mRLO2ySyMfvmQuQLZ8qsMcwYGLzvKQd9GAYxB
lLrjARiNdoPK1/nEA2vcJ+c8K/jZ+7tW5ndD7h4A2HGG29tHjtPeoY9rEUjAKBYj
2QOcw1I0w+S7bOth5WhM1cK531ZDBwcJtFgJqrENcktie/D5Iil898oAUiUdHe+J
fUDs53TkjhDEu8fFGeKRPSU8I4i3v5+k4YXCZ9DddnMRdP4Q5S3M4FEMYCVr1nzH
R8DIdT5ZTMpkR58eQ+aCGV3Cpv3VuXzmcHfRpiEIaEpnGqj6Aeltxk07SFLRmFbg
mEzteU3PyMWLdBmeSA2UCzWoWRtr2huZJyGvQG3jktUAQHPwk7Kjnl3oZmrLRGJ+
o8A4vhW/07sxX305F9PSkaebFg8U5+hJAesdrgI7YnXFkiejrhUFYLI/cwwVmuBP
3idhzf9/hymRCAKyzHTrYbMpG8PuKJyqwlkfqIB6BV9axcG1wAsCqEch0HF/q+OE
pobR270VUDAZLP6Czjvq/3E8wuLsel7nPSHnfNfK6QE5at2RiQW41U1ayvyWVZTw
De88L/R1THS/93ca92DpOZtjOL9GsAdxvcC9jXT0V54cz/tDa+lYoD9VqN0Fd88+
WMvMz1sBRlZxWDF4gcKzAv3KwYai4hx97klD+46Ar6WZ9LiP0GoahjVkDZAj6Ssh
Euvxe5K3tq7JhXsHBd0yiQangB9d2lcQDX+im2rm28CLeGg7tn5mzZ2VvRxBY93Q
MDy5Jk/Qc9hLsDUaesBnWV2cnkNjD/WrlqD4QfI6YkcWBgemEmTVWlyRkUf196WO
UFOeqibiHTpSIwjDi35zkaJnVoOdloED3SIulMPV+ggV4CCWeKzyhEG4xqcr3JKA
oGOgpPNTrKJvrUmzMEQ3cLSof4xCbwbhM7GxMzHT7Y1zkrAAVUWxY5orHPv56fjt
MGd8t+iMlxtVLpwuMVwd8EQd518htr/mvwmi/ErlnRVKLjfIHBwQmpzA0n+9fwGX
99Pq2e5FRRM0qAFDsbVztwnvo4hOftZs5Bp1ffJpSi0QjdB/6TB4DdpRXsZMzaZX
QC8HEigmv1xdNlwvQW1kxxET+qOHH8v1qgzYPHOIyY/S4or81f05qrgodXCbyAqv
cael4vjdl7Sv0QqiqvqaHiUAAVGPid0MZtW80ulng7nLLFuqo3DgP+JtbZRQQm/w
vJtTI0ZNhS4iVVoidTupyXkQh8xw9AXw8PAt9UQVIIs021p3sdbd+TBxjdftsrCk
qncvAZSIXb5qL4N/BJgZiv5PwgtuxFGuIV9LX7k0ho9Ni9zdm06aPHw9fr77386g
BIu8796zRpfunMTX+FOcKG40aJX1b2HB0p/Z2G9pZvrpd2W3Uu8OMLqmJzbLcHAd
e0QfnZRPHlEfjqnCtlVGaGhGANWKQhCMtwkn4sfAosaeUVEDLmG+k1Ca4K+dToKf
mZksl2ntVtjWPAOHK1GH/wcKbNWXwyuLaL0KAPtzZ1Q/XA0TSoDFnf0ShUmfZYV0
38lM6Kta0dsEV5A4hisARfyKQUQWSUAaWto24BAr9ri1+JGuvxBBy8ILru6o80x4
MYmPAefUReDgW7x2ol9INOtP4ZAAn0F0l8otbcm0I0hgoaplvP6HPiVJBHkqdPPn
CGbbO+7njxVXfKfKYxNxKali6W40BGi/uD7g860VeU8CW3yCVXtLnVwvtG3vDzat
6R7nfRwq7oAeRYm1XBHSnpO4sLYTCP4U3XaGZwytCnC8S983Hvn+hz0V9MGC6Tn/
9IzVQT6OSxXU/T0adZXBcogxinDYR8XBYI3ggLBZ/JiZWQdSvQVVxskdBtSvsg5J
Fn2CRnQYZuzrhrVsYLiam7HLuEdaYbvU4FXiS8yQ3MjuawP5PIVl1NZXVJf9L8sg
zu+yM2SbN6W218TzkcpVhh5isiErGYpoXmIQSaBMvWtkyzq/gAEhsxzwnGVCIU2w
9jvmZINGK0DRQSBOTp4fcnIm4IbtWLUnvPXjh/ydAtGPWpnXKls6Rjym9/WrrfSb
Pb+QZWLY2QrszQ6B4GK3xgIWuUuIR588eXM+pVirEfp+B1g/qGj+IiD/kPbUwXjh
xxNGX/vhuO1NJpO18BZTY8XNaUEM498OuBhQ9Vd+sfOPiBNHExjyYPVOufR9QJW4
h4zW4DPkXIZBSGEthvP7vKlOIFz8Z9i0/qsnVgyxNBDeyVHDldla9CPLzLSnztuE
8oxU6A02QNEU6KijQuE5UFIDAL3VhFJMxi+OwQopmelMACtTi15aGVY1fSpwM64V
Qg2lDYGEC+VQPHHDX8tWeBmVWUOvr/jBOhp7qTz1L0mmqRbwfhOM+d3/TyZmfX4P
pIey0EzTMbRhtXQs9UtrinJdXzBlReGGpHoe9ycuguWqKPTIhdAGUC/7bPF+Xq4d
iTB1WVLR8WhJHLrCQHSGm2yID7BJkKLD4F7s09gizxJnRuvNyFZ+i/lhMaUixVC1
63kTWmY4bfdLgTAkSeFtyl0E68EmJcgcOAHi4jCZrJD7HACBqbfaETbyQPopWPCB
CS10LogUL/fiibKgzHRi7Rrlor5GNtVMQkds0ge3VHdefn8IcfEUeMAkxU4T32s2
pmU4mwnAJqDmfz3zItnzlJazrF5t30vEA1Wftlhf2CFN0lTVCFIjIoemfhJhVma0
Hlr4W9MiUKdAKE2FQIUORmMYibgT9RwubKLwDtm6NAeZP9Pa6XT1WLlYu8dfwx7m
155jWvy24wrn9JZkmfQnIIRiApor1xkJpxPJRQ1ISucElKmfoKUBBjev+uFMMWKd
WsiofwgeMKEUseIeDjhEGDfHsD14BLq6w4KakxfDa9PK81owsprnUf9AMTItH5Xa
WkGMUe4g6FGe8p9ZFS7RhoSsamPbllYJ7JEjjGw8ISkoc6zyuyd51jprqR+SSJP2
j4+C6kUMCyCz/6oPtHoEjKso3VcjxWXCfiMFOFujcqA4ZOs1Oo2RR/6/LcrezQo0
xS9bwZFV/J4uSLAPdandRC3K2cP8PfvnQ3+eQsxCPYu/qY3pgUkpZJzLbwwbLoRV
qUGktMZH1U3bfUOgmMluiciq0FXs49wLrTbHV4yjPfHYkry7h96aS6mu4vDUMk9s
R7d90XwZgnwoytncwRVLALNUGkHbMEda1ZBFmW9pgk3540NKG2KDcCQCfUjwZQ+2
EbPgzE829tBGhDiaSjSojISNi3s2nSz+nZyfB9a0YKl4cbN9Xb8DIY51rzh6behO
4h9oocMX7v10fONm1U4Z2GISpVHfGOJYKETL6J/sgyA1y2ets66K0EdrXjnF4L08
blAlVOdng5MKWLKx3oobc8CyLzO7BRj8yZJA/mx4QEnNwH+IYe9zR6CdHPG0uwKI
ryY1wwWFnzZGCKa2nJ57EtoU2TU/if74jtgfMY+mJd57xjZ4hLj6ZUkF4HClJE0o
9kbc/g5G6b54fNrVxGeuA78nCN5oD2AFDihaRG0Os3sa6CpAEnMIwCcP8EXXs5GD
VuKHFe1gv7UleuDfekIBWiuwLuGIvlGQKowdB3mCuysrI+7jEvL5vMXkoI4cq4/Y
aU5b5pajhYEoLuLZNM2koEsz1KodiKhjuyn3VzzPxUhlt9Bzv4qdslxbbdeLyjwP
3Q14PNqQwZCHkHZi+DmUXdzy5HR0B1lGZlofCmRtI7TAxTxXKgOmqWCD7J8RsR+H
I+0zhaWoaTBveg3vON9x8WnCl9LgZDpo7h99v+JB6iSI1JVTYemCih3nNWj8X01G
56cphSzRW8svsNOCrt+kdEhdo6/tvGBt9VrQ2/Ji/l28QEUFeiCebBMxgzlbcFoH
U1TnZMl2GIwB/XQO115KXH1zmHGjoWncB/DNK6Hoi/mzq4dwE92p9zjCouJLAkCs
FyCibmZp1FPB1iZJRJ9wpDyvxJs6C74zI/PtQxhTr8M5mkrlqcQvIm9JWiAb3C8T
nFiiM/aVTqPgQ+lMBZPtbXRDRj+aMoj+WvWS0H0VJk34Q7oJIiDhv+SEBtnnYe10
g4zMMuW2YUudeG0EXOu21W6nbunyvHo+IadtO4+nOcRI/ZJIFQymQbwlwCaadhXj
AAr4WJ9nype1B2cbAzaqwPIyE+YKoVa2Zh2/Jr8JKchu4O23TErg0Dv07VTTKc9k
frYJYyYLnHyiQkL10yuorhFDBa2k/DIb3kEr0lPGbIxpLjNayMZ7oiX/rZ+M+Zp5
jqxxRzzTnHIZB0+bUuC4YxogKHC6qrVMdH0y9+SSgA4aZtnnO86mYak6hfyaE0va
9Hj70a/Wpos7HiqAAG44bbqfT9CZlMtGiYYDEb0BQKtVHQLT8MAXTzPybvN6MWvk
U4xtcYsp6KDkY7K2aYxvt45UoDe+8Bht4mZhXM/Xf7r+/QVGzjAOHArlNnbSCGGI
j1XbjnBF2lvtXYFwrrKDW4vxYEB0AmqFrst6fFD3/2G8hVRXQe/CmZVEzCfYmzCu
44uFrtu8hg7gp16zCufLJuUSMiFCM4fX4l13Rnz05QcPVeGHtV73HoXsBG0EYRSm
kx0SNpando/WGlC3tRSh/CpztDjY6cQa6kGYuEE6OV/sQZcR93L0ZDEqI0DdOwuX
vmDfrsCA66ec/VZo0csItiKBVF6Pop3660KlC8BboQJhKaJCCBCCu6Sb4NnMbRut
9h4oV5+jOLN+Uqb1TfrqdM3wTyLgF4qhxfqvoNWvXpdCFglj54b3Gs5UgR51zkY/
3VO63LwYdVQKQYRQJLpUwcR8UnJgxB4dt065BtiEinBTK3vguK8hujyDk3OR7d9B
+s+VsCUa3+BkBql+mdMjHuKo1udl1FgH8mGeqOkJKDUa3j31OoNLLyEXtLCZ/VsC
DV4Nh2tfx+MHOLNv6eN92biMaiyaWomeh8DLywtaveytURChrddoFMQE56VTepeO
PA3eHG+TIYcv15F+mtFzXEj9Upqpp7KSp2g8M/jhVgdRmzVjdAsQLeN97vdKvjDL
7xiDqOVH6ES0l2e9amjSOyebSo9aAqosdz12dNa6QbNlK9ih9Ek2jnWV6kVdo12o
+KNVl8u9MYEZ8X4pg0n343SuiiRelq4ekTJrrPdwYMD4FJbzjU0pFZmI4Zpt6vMm
6DFOBvWaT6IjEHEDVltikK6GJ5WOv1SoSkBWyk5bkL2SpYY4ybiLsroqAda2xgD0
9cnozZ6paLxYZzEGwKNJKOjYtqJcV2Yzx4j/xlz5oSfIOvsEpq/PSF6JLI2KFct9
h1g2B/6irsPxkagOXASFnr5kpb9CE+BZnY4EEU1BrO/pXPskUpSnNknOeo0bXqbB
qcF3UilC2rjZaUsgWTujNydOjaNuFE6tauqiQ9T3PPBDfCJchOy0hibb4AMMWuC1
81443xdfd8SAcb/fPP81yhhoi/9gNUpNXZ5fgCiubOwDtAarwsGQyDeczHHEcSsC
BIzOiEqCKSPKkHaYfBUd8QSkHrJ5wCyj4d2brQgJHM4M+PM+4iC4hAjKkFnPJqRk
1Hsz9UgmQohckfb+4h+Wyry44fIb+qdU65XfcN0xMSAMwjSPBNjrSx2sa5nAxoaP
URbBGwT6OIM8FEr691cSQq4/A7F9u6nSi1SbuwfXK6Wo7+j0k+ONixt0CVKB9NDP
h/wVBm9FE6ti+IZFiRaQ4yx7V1Ep27Hyv8/oNPowX41tdaLvQD4ZrytErDSWJFVA
q+9DH+/XvUNQvDB1bI6OFLYmFvyOO/gEO/is4h4mvSl1gnvTJyES97H7CThdaBpB
sk4Lx0A36uFxM+m1RdBkTVPqXkGo40+2ilXr9/LGmqc9jZrKWUJ/jw7NBqNwfMXx
ZcHTbM0vR/3bJm3WU5fwaxBZt1kI3YEDdif5UAq+ZaJxM1DLL5wsm4BRkrzEwtWZ
hC+XgABRdFk/kUT23frxksrX8Z9Zn+6pIcWMSqHujxM2JYhyBX6z5zpJXl8Pd4uO
Zt+Ab/rXHK8VnpSaZFVau9P2SZbPGmUjChZuoetAQ+bDRNUxksL0n742tLb1IQ/b
N7pkQznFccQB8XMk/r/TP/14ywsie4nEK3i2zXTwnJmdcq3DsHM3v0dVou1BuaA8
Q4rrCOeh1KQhEOCUnu/ZokY09wKnJJgLNSAxxclvGUT5oSWjU6s3zHmsfrc0cITA
ZoN3pQJErE6Venm6P32GCqdGtaU03Z52+XmfUn6kAtsX6bzwKjRGRcFJQysYV3PK
v8hk1P8bHr2Zf7p+klS5oXyqpauzMhNKNMCD7Q1fYlv3NwfL+s1egMlFiDGzEKYR
WdtAbsKNaebNBkWb16SAj1WVC5WBnJUVKbeRjJ97sCyZW/wkWrLo7B9NiVyQN4Ip
eEBqHPWK+64s0tXh5puvGbIMMRRE+PtavtXb+rNFbh04ix8dZ9uc4hxDC1roW9XE
NW+b5TVQzbI0z+pbyjvjtK3jgT9XLoXUD+gAsdxKiUF8PozzrK4GGUZ2SdVP8hq3
RBBLhuh3sMWd3HVvZI/OOX94LwT/ioas/+ofyOIaSew/yaO0/P2876U81pgaPjas
uMDQyZPR3IuftMqQuSWIP68isAPnZH3QXwLFyB0CYkZ6eIGJSwDxyonsayoESVY0
5VzZHDMaGUeLHcOIxgD9tQVGCsu90qHqxeKRo6F2I/SH7EeLiN3jZxi3Gop+Gqrt
xeHtBq8GsWsxL9iULxqyEazphCxryJONXLKM69schIZRrRfiBGOo5kuCx1YdP7uY
6psVodLJzLegnlk2PLNM03ScWXgRTnvTrhBWw/78ujzJqcUJob6SxzhIj30FrrS9
iFWZEYinWjkThV9zMYWNY/86YOLS0u27L7uwMCXfsADZgwy2b6Y31bVMvvZZ4k7/
kbhMNSwOgexRuWtMbec7kYQq+wgS2Ovel/+cGLR/6Qx4tAIsY+l820i+Gvjk7kCr
GKnOVhx1pum97DAtOXmUxcKEPj7bPgRPG5f5D66rgAQpKLFwrlDi220E7GYAZMIO
cHWzu1qC3O+jxXtsaNka3+zN/Ymy5tu2rs4aCNoOBMPwH/mTg0gh1l2w3nMzqsE6
2cMMeCWmjyFn7N3Ys1fF/DIF9zL7ACxMCspofHXuuz8Xy90Hr2TxJV+iLUcp1N5W
AFRZ09gmXuRAh1B21bTWDnswF7VjOwPDsaKTEY3jMcnEP5T5CoRsYlNuEEcvYS4r
1qC4S/BBq7TXmqAn65layFxWVi6ynFj1eH6uPxeoqhMsgq/DJ9nVDr9MUG1XViRD
9vQ9wH9i/fGQLXANbZvEsc5eilAO7RVVcn+p+uLSgThFAlgqnLTWj9nIlUGMmTLX
5qI81y467ukmY7FXVoB9nChNMsAFYEndXZiEcHmjlBR3fYybo5kQZengpHmm3Cg1
iOVkyLE8dzzBj5PfXV5PRH9HVnI2VEZx3xUlpLGAefTjQMHzwYpV/zbyulW2i1X8
9Mq2LwTrOti2+MFT+e4xTXPkVM4k1ce9+EdSC9BZEZZN6CdxcoI+MkTosuC9Exoh
WJIWL6gRP30FN5CFGGzq6V8n5nZHWIt2M+4uPUBTlSnvJCuqdUr7TmhvvlGGFElI
VqOU+hGDQN5rcMBwGwpQ6pDoQpLINpUp8j+pl4S9kHgrMCs8+vp2Nh8cXWH0ZVT+
h2+9TtTT+M4zMqfgLwdLRi8TPx8g6fVc7Y6WE6CHJpWTSuxJvEFu3fog39TAYXav
mnFj7Xpp+ohbJ/3xYQSZyP4pfYLKFEspyTCOgEU2fS6rsYmno2S9LXwAB3snsmPk
URptJDPzb7QZPw3sgrPIfjzUBaZ7Mhc6go8L3//pGMx2VYfxHppEgYArJf46gYXT
Jzpqi4YogYKuTMudXsFpqO+Bo8I9m4vN22l4rG/CIbXrbLdYjbclCR0oVQE9IHrw
W4BOfwr9JUT/LRhGJXiap1XV1YQWI25LRlnY/KHVbvPYMex3FDBLucsoAUX0JyuA
nHpXhp5bTpRgmUJ8i553aU199Miiynqkikf3MMWLuck6usLj44OIzsMVrbLwVRqe
QNpNx/1XfnKaxzhNowR0F1OerX4UEUJitNeflKndSS28KtraSvvCe8foUXLp4dAm
aIhvcPCanVIFh0NBKjf8tEKwNX+THC0U7iRltEFjJ1Ppf/K89b+LY1xXQ/98xyku
XLjzW/gPPJvqCf2CBZ2KzzAXS5vuM5lrY4JCHY2S44wY1rfgcVnlhnEzPZEZ9rCJ
fYrwk/tZwiFLBVkYtHCxdX/W6UxIibAXszolFoIpOJRC/Zi4frZCoE6T5NfvIy3w
mSzefS/QW9ulre0hRRJ65Ya+F+AEGhF6WtcxYjXBwd7UgKDatCLiwL/LCj5cEWBx
8LDlCf2DxdMuXoBh620VAVHsFc4GU5gD4Do7ALOO8XV2dwiMmtD9jShsZxq/x7ME
NbAKPfAsEFC0WMHrhVoHHCiauG1h7fdCvJjALaAnJdYKka+vvpa+qA2LQP3z58rJ
o2Y4Nw6IsyY/i+/J1Lek3syEtQTILXrqyCe9clxGMhaFwQ2q5ItRyfA8xS+1gZ55
/dX+3QxzD3hOZTt4HuRPvy0I8IcYw+cWxxL5GZaMjQtCWnI9j1nw7tLmW7OlluD9
JrOo8D20g2LMsVdSR7OlKa0Jm+14mpvw7I79qcka4vvbIeQ/I0G1u90SyuXfhB+k
rlZe0G8hfYu0fIqz2djlolw5kpDF3j/4rqNk2jXn9Kud+K9lCkgEhRxjpsF8qTTb
G6W4V9Wo+QkxPXwKJ8LegcQI6v2oz1qNCFGKwTVoL7Y1V9J3XIOONqmuyfXaA22y
mEzLUEkFNHEXfWRQyfpgW7qzK5+vcS5RBXfnTuRIWKULbL6G3z5sTcOylpLEVGhl
e61rAAHBsGikbnwpk4yFandXk38Sbo34QfVFNEGW2gcuLi+9TlKoJsFcPdam529b
aeMmKzHqSIHfuF3kNzvbjwEr3FZoPOGVgX5HXNYkFQtXPr6PDTAKsNTGbl9jeC/p
wJ4lOBfaZ4Iwc0SxrTiIu9QVjPbNOKY521a3b9nI9Wqq4eOq2gSFzTWAVNurEnh4
MPk2Frl2bmsbJvZCyzszduJeL8IBjnaXj6Y3ez1ezU5OsCYGF5lT3MNRHzoJpeYf
7Xxw48VrtZVGoRB9sBUDbZxR3lnqWoWozAK78nYVQFbwEjJBBCmVXD5ANe6oFgYM
yF533dSEfiqzUvdpPArCaPkBBOanELP/w5cbKOSoOmrYB/Jz953Slx4ugMp/WfPh
Km6Nf0v08i7giq34V5xAdmNBD7WmMAWHnxlcqtXg8Dw2obhoFrTy12vQC9GJGbyu
TKUNSgmjVTsvLD9Ij8P1HMMeV/LC9PviHiFhZMGcQ2YtWCK1lDYQAH/lKh3X2m7y
7+ECZ3BhgTGSlqLtoYwhdev8SgbEfdHtzMo/cKuIxqZbjchnS+77zIPZyxooUSFY
+9OXiCceznWq5lABpGcvu+8DGXF3s50Y2REewI2RlEWo9BBuxRTNp+WFskXzSbZz
yP/GLP5CRr8H/Tvo3X+HjsgL+dRW7H6DJ6wiPVlixF5W2jY6bqmAxboQoFqfso5i
DmCsJpMLSbnsmrz357Kg1/dzo8D9f/IXmH0b2dRv48v0zW3HAmQQeMeWMIMvDuyj
4DQa82+pg2m0MxLWgcfPyxTwTzc3IAgeR8voSOIppDtsOMEpFm8yFxWce+6+4gne
zzC2xdOjpnrfb4kExULL6/SNny7zK8dse2Ys1b+QjZeqQ/6VZ4HcWS2/g2gr7Gvk
uldhYrRffCW+czyJ4IW1OCuGw7EUe0MU1O9rmgNp8hY+Uu0M0smRZqPuQHxaR4ds
3didF5fOe9WV3+1Z0MMXfCS7IyZ1KoA4tghMTN2S49CERQXkyjCahQ/USmjYqZxv
DZVcr4zowErIwob/JMHVwQ7fNEjJHr0VbLvvknmIYPyxmaz6o74amU1/ezwVmrfH
wUX0UJ7vPTlka+5goHN7JvoKwDbbTMaz4h9gseqe/xrD0ZzxWTQKJ5aIwfLLox8E
hJInq5D0kBJEtO/TBU/u642FkstoWL7hGyxVBp4xTroy+hWRzATIDmqn2D2k1fvo
fPl5faHqQQvkcMCla7gTJo6H81bexNuuUgcY8hFdCqHr8jvQPVjN8X6i7sq/w7AM
VBrKogC2DiYYUXAIL0bNyNYIS5OCYNICIaJvbQxOpShUG9hsEgqL4Vkc43n5GAc2
UE/NZITqIPoeUY9mk0Yi/6Vejgv0C5Cj8xqr7w7Qckj9i284BDUua6qvHaDgxoXx
B9sNio2wOlA+WLPQx4m0MFuMNnxqk4ilqrBfpriCFVMS/+3Potbeorjevee+LY88
hX2X7SlksDSINLyz54i5uWaHN+z11aZZiRMWTiLm2OwPqc9sjguj3w18BY5nLFqs
+Iin3No4BqcXw6C1rMXXl7bMldNkVHDV/kfmDXJUJJYKr1LBhFFAnJsvdCi7MFZu
GPpJXFI9DH7xzLbaQNIsF7yejeJU4KFDVKvsBGLKmItESrAMk6EUmsn/rTgG/ZtP
G3VIypWCz6v6NprCBRZg4RMk/t8A5c4qBt55u1knRQyclX0+sI4VXzRbzSIzMcub
Z4pUarAl/O2OWs1CU8TTuu4Kk9lNwuLWe6dQS0lvoyBxC658fQ7YnAuY74TsWFWB
MKoFQTVHcdletF98gbbQ47F2hZouYArPYHJLZhyLt/v6wjXkVncP7MzSw+ZQQI01
pVW9Nxl4KFgSmyzHACWMrpQnKW8Im+QTikTaZUjn2FkQTohaZelvHD54HWnPvcUZ
9STISXtqsjUW7rfMGtNbk61vF9ItCSGVGGTBTrWyP1VmqhxkuOYL0VDz+oXeB7T7
RCtbLXvBWA/J9yuxeZKvyH8x0Vx1u2LkhzvHruQDnQ9YZ+ZTd6QV54TmlxvLtpOm
0bib80V5DkmklQpTMLZ0LExm0jfLwW59syOHhycNONR2vu+V9v9gDEg2qKhPvy9H
wEGjoUNnlVOoHeKO3CN2ss0pcNevRPt8ergr+mi51CRCsyEmApnVftZrnPm8mxpQ
JFzf2QCLXgDtIFsww6l5s3u4I4D5RJPO0656JZo9a0t5IIe4jdMXAHji1SHwNJi6
m9mGqw+EGV0ITY6bBL8//iJhIdRzUA/Hu4+p3yPssDB4qtkM7ilxeX6TlLQ6NgZF
TtaqW6JuqCOJFG5RztPe250ezTptiTdFBcRtLjra8ebXpDXrddn7SvjGMA4XjpZz
K8vd22A0VUTeWYZtwIyXD+OGmrBfgU9SOv0NNa8PQieMvUTt/fWucD822wWpxFfH
Z90Ge+TyhNd2YxWZW0WpZK7LPfyxVY3RAC6lsgTDA3lxg7GvGTuIFDkI4FLawF+C
29hvQ8s+D3NDE0I7sZ1vuqAEEgoWfQzDikZDWMy1kU1/WZFRYSGWfZUcYLwSfhgs
wNKfXvB4aZr9vj8SZDAt8uzXs67/6l5/cgVtXlmE1s1gJQDpRLQlHCY/bNS7xHNM
yf2upKJtmZU9FVt7613qJ4m20Adk7JbLKbqbzAkpA9B12UwQb5/bbFnalF7QjNgS
vNTVxGBfMFL3nRzmlhHrqbVasoMTpBPya7pU8nCE9FIKLH1UN40Qm4gLoadnJ+5t
ACk8MsdqSRQg8u+dogzvY3oiMsRVnJ+RrBPL24Yz6ViKMZqumMkrPCoH9i31Pkuh
pVb2UxUSJl0UcoASIXXJLUfX1OVuUCGlOlEMatVxlevw9xbiSSyaOJbu/8rEOgbm
Ia/2J7MgSU4GVI7r7VWPR7sz9fU6X9+T8VjrKqHnu2kZwXhKBaMQ24r1y5BUjkay
EHk58e2s3jdaj3m+zGqRUdn5lN/WtQgYOjMj5K0l3wy9RIE5nqX6IYvSUZMvjw3P
Dg7tIqBCzcptuOnLIYc7U7b0hddhSOcd3IrWSsAcZjvknwV2sOVR/q9bAVAC1ySS
JZDRex3Tbo75S7SQivupfTeuShOm5PH3SFQroqipk8zjRmn2RndFWD6pWhjvKV1b
yuCOCSHeaTZ+P6kn2uSLi67ydZ4xl1AnS3L7EmslWwXnsoHX/73RsVxpNrPHyykc
X09Ie2WRGCJHgqKBfANJe85XK5tZb9SXW17dQ4lj+rAkJiw2b4J6Lg11E5/OaU3u
eGpDEd83AxHpb4LmzrDyHhzYD7DKOLlzhtsDIvpetCQkw0VMNQ07bgCZA0rq41oC
SP1z+dVAJVwVmrc4XZMxuYidrpmeiWX1PIYeq0Nv24HbVBw1SMtpi+UT+mXyv73F
VJHw/c1O2etVRFr/tqCZrRGHEEaHGy78JRvDcwPbnW3bDBH0XhQRIdQOpIjLASc+
FjctPRXkIEb2JOqBNMuBJEO03kfHw0AGH+2MimfXpgwsi0lP/8p3AjgXOo9Wutm0
CV3ZFhe8Av2FAJpmg7nUfONDos9h/Z9mc1DY+Dxgq2By0PpuAjxMXw+4s3F0/CSk
1SeH1HEvhGkEI+v2sbKXX8SsFLGu51sjRfSxMmOXKyjfMT5YXdy+/2XEffc1hS5w
UBWEAK/bwqMW2an9EK3CRkNrzlkPwXbACoMrUFyMp51FuKlYlZ4bRY3A1ZR2nhp6
mv8uIPBHGNgHyqUB5Mzcy2ok9b6cZW7S9kxMpGDyk3teLeC2F8fWj9ZNCzxEOcZd
xsj4RUMAy3TT4vCv1i5HUbsnStu7gTrd92wkf+MT03ACTDrqavgk+cUkd2SB8HFF
flayEppgfwVh8EQnC9umwiIVbGr/V6oa9AEA7bI4s26TnC6bbeEP/q751RpwHvMD
MayPjhJLoIORnVdLUfAQyteb42OHZ+MIkW2ojWlRWSc098ECMWiRJ/WP8q7G3gx8
W68rEkY8AB9hxS7kDG6yBpMQ8SwfEY9sWZEzsASzO7+808DoMTHcZfSxEQAxsQ6k
kcA+G9JFVZQUYPBNAVNLs1lynjGQrJEA2ghguma3t7RzKVLCqCns4MxG05vXEHFW
6EvBD2zyuaah0szJwUjz+JDFv1pBTTEsS8ynOH7JJvV/UVVklnDdBdaiakq52ebF
6DZRPW/tvCVEObn5+zMAgawFFtCWjjut932hl4Sfq4TcdcxrYBgNXgPwvKFPH5Uz
L1lwebf865/ecddVE5yT48Yv7mlmDlG6puqt5Xsx3GToWmMazeYh5SQvxk3VAbvI
9DkveVg7QAb9h6P1aK+WArJMVj3f4u3ReavCYkvb/a6cjohIEAf5fK0sD/ZocrZ8
y1Q+LJOt6ZD1cmN8MsjbeyRJxQRTiLO+2F6UISb+F/QcHdT7gJ/KUtOU0Agjr3Nk
3a7UeqXsCqDKHRhGJ0TTEwPJjAXSfKvpjYeYRf05/3ruyqq2NAtqjTn4xbvVPMs/
SOuQCfoUpYgJSyTAX3kfXA5xcxsvnb2SVTmfWweXy7Jwjgum837WTtkjCV9ThrS6
5DMBph+sk/NwpXnbCdCo/MFhe667JE+hRUou/FOPJJoXaZrSabot/wvG6PpzrKTI
ojHQCADLjaJia268Kg/Vc7ebQSAJ6B/5k6gKN5SjrMumzyOPF0phENk4IyAQYGbH
mqG1srvQExHbxnVsjZ+Zf9e6dvmCYE+w0TjgUobRHReTTVJ9j4a19HZ0I59d94eh
d/Sqe9sGQaiGbPQENXXVgk0OBVOiJU7ltLmHQOPcthuSu/ODqmyKX6DbfRB2ZqNz
CGE+SX7Zc5Z7IX1kk1KOLyUH4aXOu1Yn5IyOx1+1W2nvtw95Sdc45Lbao9GNZ/wx
ZQ6waLWq4+1whRnNdIVR5+bMo4vIWzVyV44KNmmn7d8=
`protect END_PROTECTED