-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
u9LcKn3CaN7NN1pap6Vnv37NP+vcIkpxHuzoFvLglc2Ss7m+xugQ1v3oervJDzFNc9JZ0XZhVikx
n/AaKQj5YlV/ccjcCO9Dk9b/GCFaI4k3CLxVRCdS7khZN+FTkmxuS8TKPQNNtHZrCxfACc55EMI+
zPEi7Xf9IlNAQLDOOf3TFEJmyIRDv5qDs29a8n9SgYUQyJS54yqx3PKQ+kV/vwbNtBv22KqqS8iA
56wVRnDMv7Ab6yeniXzAJcKeL3pF9bjaDmmgDSJCwhKJXd3O0s9eb/Am3DWYJWs3zisQfS/toCvH
J7tKrsnYbgGJYiMsRd4Yqeul86FeUv6gAZyoMg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6336)
`protect data_block
4ESqVSJ7g5Ah3sYEA7h5cTMQLNGiL3xWv3mt2qo8SJbLvBNVTAU04K64VxN1CE063PdGOtddrHQq
TbHGAY4Vqc0O0Ugd2KEwCP4UZvHqNv5wRCtu3mnumAsZ8MsDeDDvl5kMZ9m2Bdi7kIeoYMUKhGmx
DLL0YYu1OINxcPhQTKbp2kMmchPVLViXgg7XIxJj8oTbbAOBQZPAJrXSTa9af4ctrjR+Li6nJOIq
+pU4mqzmMTsnqmZ1uf3NcbQNsu9jF8Z2APEwnDCD9SuSSrvkCwVpFOpHZ2mONlAq3ylU1L2+m4Bc
T0yieaxrNPfEVCuZLsUFw3WyI/6LwLPkOi99ZKGaLsDW8vtESD5J80IMrdZODC20o36C7lY+xdzG
l5LAlynMosQ9Wz/nmPCOkfakhsGrGQU/aYoXLxkEt0ZTCy90kqcA4lUBv3gufdM1QfwRF8VigeVy
2ZTpQN3jVoMJJPBc0Vj0eXM0a+GRuSK9PmB6uKBJe0xkgn4+SL8GYhj1Xy7Lk1xbp+Wgs1k5qmnb
ldAYEl7TpHNma2F6Cg5fvIEoUX1YIn5HPcMyIbYQ3BiDEPm4rR5DiXJ/Wo/uN1AsIeoDFgsoVUqe
2Vm198rnnPxBzWalpDJn9UZS1LdJKIlLULsfagX7LZpt/fBHPElw7lwT/OyLfDm3MR3gBERGhBdH
hl4UQr9FkyVtV24W9Eu136Hq68E4NJkwGFwL/QglQgF+tMsbwec7s9LS4BQO1r4BAvSYfPIu4+qM
/STWzTlhTPFEbb6tS6rqEOcrKHa7ETL763/H+XAIYt94ZOTCS17r0TyPn1yosOAi/U/zT4581T3a
yT4dD3wguhiyjyc58r+1m1m/nLfinruQMlTjCuPETvHkiZT4QzL1JuWBFl/XWBZru7/EkBAgXGKV
HHNaH7R/HjvyyRQgnkJuKdcSiAteKdg/bY/UGf3vDADBMYk8eazzql+JboOOzi1+x0LZE3Aex5ln
sICoUunVRFLyO6q6VNKx1GPxyf4pbByRPnsT2PmEqb7cOwTsYaxfenV1TaV/WTFM1jAiaQrEKqoQ
ae1qTLcm6nFvStRp8aFkUCtWRVKg0n6bHl3uhL9Cwhu71D7XQo8JxeGKmdYWibm15LaMjIaWx3JR
opjkulM2zmfhataACWftNlrvMMvhhKzMuWSJ/GpJvrjUPrc7/q3QEkK2K8tuUzJQFc/UoR6XmHRv
kyxrHK+xZoGpi5xtVPxrerT35ONMkbK/DCERHE+D9AvDAFOeRqKWA/isUCDXXufBN/BZXVTBk+oG
YBqwK94dO2heEWPxTw/aRrVUPVKTlekMe4GU8eoL9L6InlH/6sXy0MUkW06QmXXpTDx1ZJiHXTu1
uI0xjmHsdW5mvu8ozfoDqgzPb6qI27EUSVsL3TBqPEZEbIXehqFOZz7YjTjrYAueKCkPJlWb5caC
t8VZOjn8cu46vkHLkGn7ZosdFpxvldJWSZkNxg44bi/4gfoOvHr3k75azOIMTZ847GLW9lBqiz6b
PhSEiIAMpYQFZMgbP2rMeMYTq/hPZ5U1V18lDmnMQdSNSTk4Kd2kmH00kkDSa4zECUJnAZ4QvD9+
a/YCz/UXMH8GkrPwIhVC7P7xq6dgaRwjv32KLuG5dP6EsoJzOO9+zmJyBEKPNCqoCpDm8QnG2cOS
TyQ45FY2bBrDcgEA2GeC52SOdojo2BBLTCMcUs5lQEYIiYY5m4oy0BtgukVjJiEjtE9cVKEWikR+
GoCOJ4BLJTAQ9CpuhpxVGH8+j3XnQBy5s26kDQxtYqGlSeQiM5eie1cG5xd4yf8m3QzyJO9hNq+Q
OLpPOWIf6XCtSbK5VaL78EIGKe8YW7EXGg064ahZXF1+i21FpFvCb9yWeBk8uv/36gxnG+tP5Toa
0MkcECy/Uc/F/39C5ayTkxaiTZFkKtouEN17z0Ssokd+dN4g7mMtZfLfpMfF2Qk3n+OeJT6I4FEg
xYB+NvMgKmE3AIZcDrIYbvF799IIgDlk2SLyFsyX3oiU8g14Fnln1iQoaZcZusG1De1gNM1usKCW
gwj5cEq+yjGycqg1lrKHdakf/mVckrROvFo6huApU/zGj83DU8ozqRetJ98FCAZyZ5e5lesTAIA4
l/ddpIKIKyKpPxzjhJcF9Z/0InHjQvDafxePknCu72qX+zkK/ZG07sAyhvaS/MPrmbctwEYS+lom
kFE7FgaeowaMFaTkSRVh8oDwCNPwPCGGzkGs7/YPVqFGI6aCTh2YZ+Dvq+xNaatBvcdBgvQ7YI+9
lMPfqQMALOfxFztp/XbTHDsu0OgGqHJpfcnxSA8r1Dqh8rjA3WSc1hKu0KVvVxL7P/6hf5bEb0dm
SaXUAa2jwIXRB6X+2Q4jSi3uRiDUhJ5SmnYNiNAAYewBhiAyFXCSLmqkrinRCMOr8u/0v+K6cIIo
0YbmUjkBNltJ7BvgVcOodT3ISVbCcEXOeJZGFvPHUtphnwcinHDkzOoxAVzivF8n7Ry0knm4eEj7
PQc5zvyrzVS1q94AdfMf8UO8JJEu38tw25GmlABUwCUafqel7b/OQ+gr/4tfMdPXukh+F6qygEq8
e6FhoLJFXhHKskpZPROTJnKtziAFCIws2U5b3LstiJMiSV7gWXeE0OxwuKVEzJaUtFaU9snkwqfE
YoBmX37nnrl644tzMVvDRUqSQUfXUoQyxb1fjwAcyQAWDDVpe1+fGqV97up5dLdzSRvEtExf4cnp
5SOWgzeuyH609hZcgKazRgdqMcmzHR+lJ1m1hDCbXUn3N6WceCZb7HYMau4Uf4BdmPw3YIWclJgB
hGTUyyzeKgz1y4DfT5cIzD3i/d1DdphKq7ZsS8VAPNAmthjIJyJEzrUmXUn8bkC+LfhR17igvjzK
oDr2lAFBXJCZ5ywT8XTK8/OXYIILOLFDoUMP5ngelXK0/N/MAJvrp4PbjfCaZu5GzjANm+ocnakv
Fm/ocfS8tZ09rnPRkJ93w8ZtmbJ3x2QHiMwAM0gvFxPokuxav0DFCgWAJqHItsaVvGlXbYurgkSB
xDoEmXOGRjk8ZNfiWrN3aiW+dGTRVK7l1lKnJWdPFFAAJfzbuxe5oaOeG3CimoawgWYyaCVZ9zzl
i3eEesRVf2lMIa2KYJ1KmzNZ26uPF2OJ/YGTco3+1kVl/bwMPgrKaT7pzVGc4T8fow+mo5HKAPF/
pumEElywY3FvOxoE51CANHQvTzhIJgo3SebVKrO/jxF6Xma+lWgKQGEa3qnEZvs5A3xfCJH+fYgM
1piMzM48Nv2Xwq7ZVxHk0q5lcJFDm1Sx6c3u7OrMjABrpPEVVeU/pY4XWlM/PDOWWttGJEEwmObH
3Syy21qOJgkyke+jos+cd4d6UX154cBnlMd52vUzN4YMY+QzxeZa8Nb9de74fSEIiIlJhsI+s627
canB0nw9A3dpIUTFjFsrOtnLjAmwK3zXI0jiWm8iRc8GW4eY8jMPcGb8yCzRrCbgwe5HwA1b/mff
OxOn7UiiQRNmL6jWRzMoRL9DCn9igp6jf9kvZL9mDgCN64K+9tV9+/9cOH8hmIeHCT0W1udeDi21
Hl0M23v9zlcm64eHhCLtxHAFWF8L/UV8QPPxsTphNCenCjNHf5A6rIaii+XNVlyrb2BU+iw+jUr7
F8uKiy7vntM/LsA/w5hYIkDLg0XHUq1axvchXDw7nzA0Os7s4T21l4hjaOrI42LCddIAppWcTqO9
0LyRnS52v8CIU7AkGipLGNdtB2Tc080N+Nb+sFUN1v5WNPvSapcTlwQXnZ3fits7v2tnYR7ZuQWu
c5vOoWn6R29Fxf1vfzXNgJNbPsEvwLQmoucGPG2nZuSPrNVOS/N2MtcjzDeK6NsouYneX1Sf8PSf
V1+4MVbrfJgVLtxdnQ5PptGdWcp5/sPZD4Ow0tr34qH/kbPQao+qGuX+b6k4/pJBpdKyxNCk7vmS
qy9+phmBsHyyuET1uAbm8gulOmA7ej+ZGxlKoOW4kge+xCKFmRr9v2uNbQ5aFBzgYRwS77PrAJJj
sxhpvCCv1e3OoySmAXqL5CPcqhWnOs30F8qSdHSF8SufocEnCO+azHD/kpPxYVh3wzMuLRFo3oLm
W9yX3XB3+UU8rDEItWLHuBDdCVjfpoehOCBAHd0yAlxIU2tdCiG55AmtxHNB4rq2KaJHnj/6vMCu
RN0QH4J4d1yxSkf3QueKB7Otz42fQj9SCZYTfxtX1sjXAAR2LcdT4uxT94vQbiFvQpk/pdomVqYZ
ra9IF6YbRI3wE98DZyRhwv0Qr9Tcj3nKJcO+rHunsyvN1Lt5Ad9heFnKLsURxpZ3/JtmXvXOcX/P
SEy4gM+FpO7o/s9fp/BlV5KwqXP0WL+QKJrBGo8en5QKz47XVIqXc8V4DeJSz6e2dhDnanlDwJ6u
DC3PLsyxHG8V3fYQX2SD9kXE5c/olVVSmaAI4hOd9OTPzyD36wpScNIML+eyWbrANYLir0YmH+dN
95f30tKh3rhIsCsOoVHsfIdMxwRX/JPqyCBXYW50agBmBHgVX9XzJ5lhNsZzX3fi6sbwIXN3W644
c7J6JCWmzl7kLxoBkG+s0p7hZI2knWkm0vmZGMRwoRdtigs1+jaF2DcyJDo/NqF5vaQeI2H7dYVK
Tr5x45q+IofjI7OGaqpIUDRyLJyMtztozx0MSTmw21dr7O5tP8kJxvnrlaCsQfycOrrmuSM2fXJb
k52IXrGc6K8QFvRkjf68+ujFkhXTe45Q1tc0cO/cEERMBJxANdilqBqSODwk0mz+oRzBY7vwMep6
NTpa7IRGvufEGDcuLAnHLaja3P7Mqjs912eQB68j10uwln9WMlnScd0VCfjq+cY3KXL7c1rqOOvR
HeTYK8NrSmZ9IuyIZs1MqxfYjyZTI3f8kian7ZjBf4TPeRzAcJ9XbqUEXjf1aL2yu4o9niKQCKeR
lhK7syuAkTGl0Ta8SW6r40E5AbUdgOe4pQ/2YMTdKENwm5vW/PyH+EBsgnVKlsSkvwB20babh3jC
kr1CPef5Ei7A3Q1lWBLZGdeugWC+9EW01nrHUJIqlNbsLdUyqCXGes82cPI3IeGUYTt0RoGcNDrp
23uXw3NWDn8KsBxJSPbcJwQ/mSpngaHTD6l2ReWxrBGQmS/jCkSP4aiMP8Vsx3f4gY9NBzYWOWMH
1n7ZH7hHvneFAURnpNn3N5KxTMSlO3vVtNO7v53PUhCQLmgH5TcYRS1mlpFmTfjAsp53dUiRWCv+
bBsCP+U9UA8IRrwv4Fch6DCyQ+BeLrKiZ/vRqN/Pt6V/tV8sJ5+jVOBbEabB/mZN7QTuMVGTom0T
By+KKPg8S1JvWZAN5OVG0pCRYSM3OiUJfzRsDM++Z5Jvyc62w/JnFltIgG+1UivB/YpWs2F13JVq
P/YljgU2GFIsuy6rq3OPhue1mU9+tjrWg+SY/bqXg+864xBZjwybVOmW2H7cA9IM1XW8yc4eDi6W
EEH9gRoaJj7jgM3Gfoz4guVCZXyBlAEiOPl96HHT/BTdugqrxJb+DHbICjpD7RiSAttDT+YQ9Z5S
TayGvsee/zms4b0gRPQ1W/8wTkaG2gY0Y0mfHAEi93z+mVsa8CCDBMAJvJCsk7IHuxI+NN2BpfzX
oNkgEkMqcPtStk94nqGbC16M0h3JUYL6lr2VwY1+GMXiyNLNBM3SlVbqx8b+BU66w1KaLTqynKqQ
EYDQmO7ok/SHR/q9OgR7DkzVF8m1z2x5kfkVM8NTEtDFhu9Gsfx0MqdJhNhNfrBUvdAEC8l1N/+U
bop4Z08JdplOk87CvrqyA596/tkJ9sp701PytcQyacINIqAdDxcysS0x5VDnfAj7t3gZSniuEPRZ
9sbQF8v8Ep1MPa1bpRaU+xSblMBP7G5OmVsgOYw2F06fGdn3+0M0A0csBt5IisPFYvapexrdGupT
z9Bd/ugHEbndLvug985qoLDXy1V4wobgYwiJwCOA2dUMIw1TRSQdY9g8BcP1F8S/2bvy0NnQsaSl
v6kSw1kLzYqi+d2TLhwlfmVJzCDUvaFlIDRSpb8Disjw5GRrnoNyj+sAcb7Nb2yFME1mHgoBWs3P
sv0Besy42S57NGCCP5ju81y/aHwCsoVjaRWoWFvtX2rPxvVEmyDFMcOkqkyWF8rt21PIh2zKCcz0
KXPzr8ki0f3M5Fmo2Gkup+M0rqfSEjGwtBx6fWzXzIe76bQCDRuRkRYjl6YTFcKtwCHpglX3uV0G
LwuZU94T0dLDEMIV4kKyoPaFDVlZlJki/A/JEj9p27JeYzFPpISy6vvsxGW2BdGW8vC3rArPoxRn
vy/My7vs0O17/xPDx3w7xKlDwUysHdEirkzMGtMQ0oS7PGc9Z1feU905XZnpPWcV//8a3/aBmjEi
AxAE9jtGJ3/wJruAWAsC+Da/BUF/V3/MkC8DpBtQmvCH2woVBlpMdUxiiipcfNU2FP4xQomiJcFp
fo6V21ScadnI1L7hKDmNW+ZKhbOIl/qk0MJDs3gQUy5xrBBH+GRvGzFCwV/IxMjcBJ8RAZ+eRJCL
JLvgl1+wlYiqxXBF7hBIX3o6BB1NUOS7OJevldxPN4qMXlD1DolzJyKUUod63LSHcY9n2oCS8AcY
BB9QntIclTwp2nW9kRwWFvEYO09g+XqPEAroYuRKWafACyqIoTL64qpu98pQ8mI6GWO5AqHqhRpD
6gD8yLr8gCBdAYLjdc0zi/gj5wbhATiHF1mL+HJ71rKqImYpal3Ao8eTAlWndDzNTmcMgIb65NLn
wL6XoC/aKOwZNhK45UzvkM4ddFSe78HRYbU20xBu0A/l74U33AZ7cZybaD4TUqSHUSrcmfTEJomi
m3ZNywejD83F0xTGO/mLWLyOGgbRctaSoD4U0ifmMJMBk1qxf2nc20cKjjjpJqF1OWHjo1xDONjh
9KgVMNQGBkj/UPTs67IAZaGXCo8f6rjwBVndsgbrvOqnjlc0g5rOdj5eoicj3aehc36pp+Q7x/4m
xYvnx5HQ5WolmJdEIMfzsV2J1B6HSmmEuIC/o0M00hKGMoVKPutgeNrlo5w67vmdHcZI5EVhABZx
/SaG3e9nDqROHKxVyF803lW+x8ct23OtHdQ4W8smACmoyowH/DWyJnuwmyIoFk5wgw05g/UK/qlV
ZWaatk+ckxiuEy3sU7ORGSyllZSZQvYFmuRxpmsJpAWOdSTADd9jlNLs7sWf+yn+Ef3YDE115RRE
1kYFeZ2ogorpBGFWTyTVopF4HnAl6ao+Nf4bUW/4vZUNZiVn/4H/2+Ob8JJh6LugNQlkCpUh/mmZ
RhDHfLZlrjmf3Rl/Yf55UydiksrG/fQJwo1lpNpXR+LzvgwdMWCO3SuXqUgzQxbcumT4lcWGtg3+
HxFiY6Vuh56XwdeHXFULS81+aMQ26oYtkvjKv0yCDLEPYK5c81rlsUHobyj9/uNqoklCfs7lmlCX
ZV94M+AgRAkYHzdnGmYPjhwICXNoV5MFg1g5xABQO8UTUemuNYiQh4at9WSYOXO9hbSFTeoyAfem
nqAYaD1zL0FmjDrQ7eo63PvyKvlxGc60/Vydbeevwf2CB/j+RC1qSFI/YjY7LFFhZBpzh4brt24T
nWLbxQDNvc5wSov3fV06D3jKcwfGpSqqm/D245KioCHegpyCHwB0/FbcS0VKgySnPxVjRZ/v562Z
SVWSstPJNwa6VgPIRV5REKxOICf56UG0Ri4ot/7Ado5WyKaTDUp0eAQx9hXKAUnzGmjiRdzPVG9o
THeyZbQYyjY0j8Y3XODaYmWqYnWb4Ne15SHRdxEfCNvZ6JlA06nn/TtHQpIG53ZU1vny4ZP1T1dZ
XcBwu6MFw1z8xSXw7W/O3pkO+g8u/mc3VLHPDNsTmQVdz3RzHGglCdjVTBaezfvGov4MVaCiJfYQ
mSmXWO/vVyvfz9kOhW6OQAN06Bz3d8RJuzlxVriGgiHPBgurvUlSDHLdMB0EqhSvci86OvrxdXAC
QgjGj0ZG89DPEHiHvAHFXdUW4m/wDvtCe6nT8Jo7AtQ0pKxVZXKFZoXVU2Fi3+ZK6EIYZ91eJJ3b
xdbkO5E8Z7+uKu7U0P9S0wsGHaXPB/fY64niBbH06NLdBFp4ALlQGSLvsHLddZYV39OMAxg62rQ0
oBBDUcHcefmG/3Z8XmCvofYIcx9C5NuCKm8tSBScvsAFkI0+x5RWt0fcw5i4TjiAnFxLNoB1syU/
MpcKKnfjBWVeDtNxSMm5HNAi20s+lrBB5Sbffg+xW+A5/jU5SWGdRf8sKba70kExhrWgAKKXX7TU
YU3C8zqbsQj8aHKMUmChyHsIMcPR+bvYNPIXXU5MsH1jsnkWmSY1eTzmuHpX32vt6jJIh8zOCK2U
Eh+A1RWdD2ta5jrfmtFH45t4tK1OMqrad7hk3jlxIuPKcmXO5G7tSuYUIkLqxpFCoTPnEoHTA9SX
3Iqewu0BwLva
`protect end_protected
