-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
k/OYi5fH/jJ/UIo8bK5dW3pb/Il2SlMjVaG0Ee2GfPcx3i2G2TAL5aGmtWHG8c9J
db1Qt2DMKKZHs30Rri1ElkRpCasDcjOMFE5rypaFi52NGUDeUoww/1nAZgEoNmKv
IV3C9W0WZjpI5lLuW/egu36xLYQDa40jMMiPkHoUlyfgo/c2q8HTVw==
--pragma protect end_key_block
--pragma protect digest_block
cFisLxDKiq7gSJ8ztPUgcM6f3I4=
--pragma protect end_digest_block
--pragma protect data_block
h0CCvc4KyJj1dr/gpT+LPzp+IOICozWWx/vqEYBmsjFFrQpK+LQ3yuoI417C5f9E
zNKm5oUEjr9HV0KOCFqRg7CoVYkvtNP05NiZ0uUvbSMB8dQy4aja7dwLoZVbFyzW
xLk0oEwFMEmKHE4p7PYZbw63tLe194sut8S3uN25OWmzgogT6rR79d9HW79jmoPN
nx6kjf7ry2oQWldReH+h7Ppm0JCProoHEWtp3EXKWASk5h+VI+65XFLYCraucBnP
9OCQ2oB1Zc1CimaKO16gRX94BfmQ35G37glSqCtdKUO5cEBpVkC77nQViCrri5mR
x6Oz6yQABFCBMr5XPZ+3nGGZvVLzTmrnv+eu3BVqh7UUn/BL6qI7n0x6mFWZNd+9
cmFQlOdTP2oJ98sRik1DqOE/rwF186rxTVxL0BSrkMmK5eMGHDkfYisqCzbpmJEv
ukAIgpQbaxwfB0ltIvucDcvU3sBC/he54QYG6w5+ulSVf5T3XlGU3eO/685B/du2
geLYmlO+UclX6nxSaeJKyQFwpbXf1IUc5q3p0zt0Rqn7T1YJEfs+OXXU4eIzuDS1
oYZu/9G82sJ4ed7zDvY/lBprQyyZ1ydzHzoCD0+ggl6lIZbTjNhR6gKgKkFrKDJd
NZhQHyKbap3K7wNnFbPE5n3t9miK+WYf6J7pWvSXa+KzXRIn7UJyAXAZLV+Atloy
31hpuYGy9TU/SNVCdOBuvXKSusYS1CfpiVdDmEeixzvmJXBeOGQn1vHov22sCfeN
buoc2UgFIGu333BLmyksjaZJIZsqs+ZLl/ivlNvXLvBVm4guFiNOXpahMk0pl/WG
B3b6KnAa3iGUsMfEauhTfP9kpilh7YvUDTD82QcotRAOMwaPznR6yWsE7JggzN7e
PYLRRdInLnW948XLSuDHp3yNzSvrAizR+MHFZ9TfmlnAXLhLA9VbXfLuqKLpomPp
E2aN1f+frgxxXBoiDzO0C62whnDHWwf2xL8s0AFURHg9aqEGJz2uTjTzigsEXGdA
h3xbvPMnUdAZZV8TLMaj5n1kPMTsTNYpDuNvkK31YEja+cP25rzDZ0G1nEBPVdGe
ZZyWa0K4sujMnbAy9taP5cBed6YGTxNUWM2MAGDC7AvTuszudHgM3t3U7WNMnv92
t7fgaLoVScg14ZZXPEkZ7ePkWOz/2Er+6WHUbwXYQMnWdQrWTvNPowZIZ91jj8c3
xeDFPg7dZsfsXh6hGg3ImZfrEeM7LLDqSfI+SVgwYnGIXM4U+TGUHFprrlfChxJJ
/rlSSqNnd+pZdr2EL75TmfsHWb9KTzlWnPDWttuWB5KZDyjM7Ae6Do2U8w90cYZs
nTn5fQkswxdGCam2OGTlfaQfatxaalGVVBvtlXf+8zZh4gK+g7SIyA4/0gRfN9xv
7412W2TQdMsWLMmCsaDLGXSuZAMIfyeCuCdpnq3HQUCv/8Uk1oP13JBK3Cavb6tg
PYbVWYpUAspz6NIUQ8xtU3VCU12ux04bvNkm8RLrp1uQTKhjGFTtaW2SYk3NOy+l
2mcG9FGhFyJEVjL7ggvP2TLM+pXunVULDdShQl1jIqw+e9wLitS7m4b+b5KWDwdN
YYbxY97/5GuRvKmEfSXjITsSgVi8T1+CS/Seqrk6nfg0+I38B731k8gKwyVb1NQW
YakfFFanyHlW0g9Q9hnKWE6/n3NRflEYL59ihm9cm6KURsTKlOtyOE8vj0FBvjAV
0uBgUvX9//k7VxJZdDtW6EGXE24mvC74ljlMexYPj1NZ8/Cg3pK/YjeR6d0xYYws
jj03iBRhh1gzafNYeU/R8GU0wmg/Zv2cHyJ44O3dqTFkz7DuOVw8Oisl6rb3ZbO/
Xo7ZgMnC0oRCY7SI9MkakafkHiT4yweqGnB/7tXWR8EnlsK1k23Fg4WXIr2OJSo8
xVZf/9CnbkVuV1nKPldtZ24BkSZahL6mZ4JuEptGO3s+75xYfOcTfM0G1Egoq/44
VPpS1mHpWtTE8msiXx5lC5zg2pd4LEHgXJFvzVyvuxYLOTP1iaaVwSMjM/5qaOcQ
JNIpjNYmQ0IOZc6qz++IMZjE0oOB7nHtfYlh/6myehFjbGFlB0khyTv+Gr2S5+A6
ojcmEIbBh1FmrwBy6RmZxnArASAu25Mf0m93ZNfj9CUMEczLux/8kYgRf8jGyIbC
ToIvUwQSHzG2AB7s+1w/+1VEYX7z7345WdhNB/PUrKnVs8qmnRvXdeO7MbDj8bvX
+Rvjw31t1DDRm6DvA2bRf5YYrPHtQtKtykoVYD2bSuv/VTeGX52iMI1PEsCssEdK
YUAyfgtwOZmKwahoe6GewBPDJLjti82jRE3G09ZTu0D9XnvHXxQqzUpWi/eSe0Er
6STDob0Z87uljO0MYb5TLATCwh7tCP2SlBB94r6q2eX941to3MOLzdk1oklmiLyv
rYzfuHRYcVrxojTbTNvRxMRh7vyXSAUmCuVG473/d9uBerA7EUm1bp1pxWM2LS0P
mmZj++Tqd6almTsZ8MFMrORar0xxkbuLF5GDzHJCG6Lv/NxWOiJdSlusMhPBbkPi
yovKGCZTH00eccmFA6DFOXk8v1K58QLc/6p5N339R9eF4hJFZJQdLQhqBRWCmCa/
bFGlen5zg+zecZsSbUk4r7ll3/iH8RYq4V3u8lkgV8R0Logs4+sbhhbPo2vz5QkF
tPKN/W+2NdZtx1ectbpoSTHqwApIw+eW1Cf64C2XF2e820agN686DdjgkmpSsjio
CSo7mUX2Drnsq3xUZLFHXMwo6Kvrid5JLfuuQWm3SpdGyo9ajJ0o5/eq6NX5UZC8
THV9jAki0lmilIfPFIsn3S0/GSu3NnX/igRkq7y+CwbCeD0oup2Y8ekEksIiSZYr
phbZXzxxl6rKcCtygOD2wGXHw/MhjuAjkU9euNGNgj9n3w969C/KSW6OdCOfCzXA
49aYiTo8kbUxU9FmJg3mNw0GrytpTpC487N93+uDRb9nXXjHyRC3jq2mx+qaVc+6
idXgZhaw2pzcf5NF0rW2D4e+bt7O2mozq/Z4zxq04XSzGaJ/609RkI7Bq4bQHMI7
wriY9/IYRFEl4dpzo2TuOIH6E3lVOAVdqgJv4OqyxyIxda2kRc6Nbnlu5sGddQBJ
j+DabihJbf2y9stC3p8FXfPQQkMShzfXYAFsevy0Cky6ClT+wVlXV0Xi/DZFB/u3
+/X0aUBXmC687YZOlUVmM3nWSneIcwZE0lVVFykHiQJf45O6WT9fX5EgCzSVTSKl
wKP3bdRHbYz0jw0L8ob5+vpFRHTJ9BgEgEfdF8REwx9FaBg89ObBtn2L+YBbELcl
EpVoxVmcexIkSSqtmwbryTCO2gGPLtTn/ptnyVlfZR8mc1u5Rp64ozYWYrqUgOr0
DBsekglII+Q24sgwswTe2Rd9q0StS/3ubshE1TUar/VEP5Fflido/5h8jvK+bMpS
KDWtCLN0DhT2foOz3HqGLknBYlpf+PT1Yr743tnLw65TxQzazZwCBCp5VM7D+GNR
HB3KkNhES0SllLMVMriAjq+Fa2pJTBpeJ2ZlRciFRYsyLNF5OrzMG5X8T4hKMGX9
CAqpyBjHZmsmbJYdZafKC2i9tkVao9+mUGdQMIYlAPr1joGxr/SXjNAw5C8/1CZP
eMHJFksmsbown7nf68Es0nw7sFqDjh3x4fSbxZohowjYPP0ya08LVAeb9Sbd4omX
w6ePRPtRs8LA51nilgs9szTA9c/SxIYjmT1I6TOsijYebBLp1yc1CdAKs67fYfzp
JjeqkHAYJuFcbtlJmU9TV2gZG/+KctOE0QFGXT8xLx+13Ge9qy1lkenyMmIwJ1BX
ta82EHGgudn544LsBMDRxnJJGbU/0ZC1vfldZQnJRIjmNbunHYcRnExG3bN/FLer
KA5+9iaXLNjG2gFsYM0xlBafbc/UNYA+rWugX4zXGR4F7nRckxwVz/Q4G/sp/vcf
FcFDxiDJ7NVInXl+4TzPA6pWcbfwLJ3vYAoKD/LnGXSkNo9j8x1SGtl7+2zZxRe2
u9cGwtx8g2cUVgfcD+ghwT4Kb0wvdDyBAjWuKHdaTommLVtBmoPUvyfVd7dvXPjv
Q+E9eKmfsOwQGveNOFhSkCgXUFwjXntEGn0F/pYrRoabOBGhwZp8LY7uaIspGVHF
yh9PwA3a9epe5YlgNxEHD2y963Td75hr8DNX2QlmR2L+eNgQcdM01QNvvD60fyTJ
LgiLFza6NkP3u0hwrAeoK0LQAet9UA+X6rqi1VWsdN5o0VlA93UAgZIJkwEmnmU+
3S5IQ7BzXzqqK0pnd24QA9zzmbMxCfmfrmAi7V/1OTS9DtvlIVyvVSaFhbmpmxdq
BjO4NFNgv4estNDUxCpZWqWr8tZk2ml1rnrJ8tnbdwIUyZAFPGefRXMgDy40YJ7K
zDaskgQ5OCUi6Y/Qo6tiW28OUP6nMzNatNKiO20TlT9SD8lGgZWlnVfOYAjGQpU3
29sp0VvMDri6IAeDonmaPIhDVxQvkZ4wVnQi9e3unY1oZ3q7iGGX9ZTB378u2jOz
8QTeInA8iLmsl+geiHabcvlzGihOJaKvq/9kG2GMi9+3pXUrmLA6yXRcvF1UMjpw
gVy+tScFRX2KiBRKkRkpua1kcFLPyWWFk2ByNrczVPEAdB6+RzsZSpaXV2JUp9ZO
S9+Z5DoU4zYbNnoCuiYHsitMOuNqWamr53KK71ywOYxmkMyfg6bTMvSijoaoBMnm
IhH9NQvAuWCw0/nF2smzlmFgCUoNchbSOb22wmfRcMB+dZ/2YvEIloD4EnxyL6uO
cqWAlw9vv6rJ1Rs+flm/lYtf5t1Plt9/8tou8B4NedWBw3nTrPzNIjnpBiOOmW6E
c9LbiO0GS3YSjHF0G+1J9TcihkEeQio6E2K7DwwZZLCOoeysKYMkNzOa03h+XHjE
7X3PaPzrxMxR8HteMwYRR/05DQruDiV3PDC24tXhYqWQkNG3tuvmKrGoB5Hr04dQ
blmUWu3u5ovvAc0lDbWpDLskI9saVWZ3XAOIFhFwnDxEIONB5WVq3rkxYJ9ROKxk
LCOuSmLdutGkvRtlqyr6zd+B2BRhKx9LOX+z0075BNVG7Nzu7fQTNDERU2uxRKZb
kwiqfWS7dUgZXmNlkkgXGSHGTVLvfgd0B6tN1pv3CXDMDjZs6aEPy3wIlNK9it5x
umxZhcxZkh+a1yau1X8ULl4MoH/IDcm+P/IRej0rR5xYYycxb1yb/z7fHlxR8rtA
eh7uu2c8UKK3Nk0ShO4LAKDIqzuDtPAH1aUBItgmGLRmXi4KXa/FvyRgmkWtJkyb
i+DZlC7T779hApdqxCFH2pCc60jk9z16DDL0KZW+FlyBJTkRTaImooPp95l+yv4s
t/y0i7zbquykdBY0i0zRMk/W/gIPO9gpG3n985U1/ME/vlTvwmMvSOUn4pOjnUrI
Ephiig76EK1Jv7vSQLPmZIlub4kGzJSSWVkoPc+HE+gCfwjAW/lymcBp98JHdKR2
+Y8S9zN/NHc9jt6Poss8XLTfnFIUgnFPrTksDfQjgG7bZXwzyW8QMv2ntmBpQE9s
5bRB3yBOgXFWs28MG44XT11/B+fQtcXoWN26Ym0WAU71Km5iObwiO7t4TEGN6J6x
GOEbmQqy0+PsoDtNESfOW4LUyKpKO7/grmWKtQ0nPRZZ38IJsTf7FhGWwt7vfdzn
ni1deJLJxVNgBBYCmvCB+um9kcIemNMQo/jBpbgV64QtHAhJAmXbY1H5FwI63fu8
Ervu/6CGdVoay8H0/KxsGVYm2hJahiSHzVG+F6Pfik44zS2BuOsq6RHbrBGKF3rh
kDVUXi4dae7E76SNDwG2GffuJiEnm+JJzp4pJvws66JNrq8KWHvJXf8GrTrkOHvC
eDwmUYO1JYK2RL2YF9LznT9Z+A3bzeB95KWG8VIIsuNBdcVedr0NZB3YmjTwsyZ5
uWWmsY0UkGgDK+AmwsGqc+b6B1dVhndv1ZmBKvigsm4SIpBY8aE8rYjiLWuyBGk+
BUH/2n32FWQHSYI3FC06D6E0Z9/hQKikFbiJ5fJDfJ4XX0f4piL43tV3NglgarRu
08beIF2C7Ejw5PDz3UO89X8O75yupHFK91Pne4VR5fkXSfIYPihPlUd9DiG0sTzk
H/C5AT9IZL1FGP+rsHw5oEvtRRW8BANiJJg1+qab8Wlp+dBfh+DBmWHxkUxcLiKk
MG7C+kdYVPTKKcCgA6PwxvwbILIBYXUmJcgApPcCb7+OaIkRwLaJaG02fHuVH+5T
Bk4frFRI3utJGd8+0L2bsE3Ta5ebrojMSyg06Gj/TauOCABZQq+L7rSTCidtaYby
1DPBg+C/9fnzx6vxcfJ67d/4PwvWdGPdTqr8N1rIZvvV27gjFRJe/HXBf5oeReGR
qmjtIX8AdI0FUi829qBsRIZ/ALTrX3DznNelXAujaC7n51jDPTAkutzft2AsWDmM
t2qBrb0ot+OGOW8+y1dqWNa+n+EiVgbVmb1OZgdQ2ev3t14ccXUJ3LNbtS9ET08L
eGL24YhBgipHsXiXu/xhkNMhWWuO174vUgFnTr/eqpnqTB86IDpxHsML9qh4OwyI
ys2lXCPgXp6hGKJelcBrlIyBM8l5S+jfIIu5XMeNMo2CNic469SErBiFUUrDxcY6
8v3sd0O+B8MuOZxXjyzg+UeAdljN5usDK+Rzi5HtJeoCtdT2c7EmaPaX4G4a1/12
8vviGwlA3yO8IdCx2Iqc0QHU+ntYivPwgPj3tFd/mVK9F7MC+qsw4DdpoiMPvYe1
u5ZjUW8tm8pq0ackOpK7D/SPpB/UbWcrEG+ctuZfT+7Dn3ImIv4wMAAIgjwKpe+u
QIdjBnhNzHnIF8RENKgdnvc8ENYUEl4AUzdkLVC1ru4vmNshIbiaXL3fA/bqS7xW
rVvz4ySNPhsenohihpnHLHKYAgWW5oMGd3uXC/WLNOqPmJI/wOYA4fY4WAPfEWEq
NHSJ9SJsYixmbNyBKGE9dGd5BASgoVKBppnCaBjKslmXwy8yzZCpUB3ioHnbhATI
Tk3WJUtk06HSZyNrD+I7iPo186jqYduV0bP8WK8Dy+laHjhcxlY2QO9rZh8lmLqX
0fFq7WQ9AychzPlfHMdy70iBoJhySOcYVUn45/D2j+a4omz5GES9nfUrzttmdr1O
7Y46VmmkmFFQn3YUrOlBiRMs/fV8sWRWd7CgtPii/CyPo0mnPLsw0ZWInVH/RChd
ZvVDhDW5Gmc9Za+U/oeba6GtAiDPv37yRXOnR1MiuFxgUviMiKtJ8O8SQsw1Or7k
pOObWGwrmvrOg8o3XtjEF2Y7pWgkpXU2fdnTrXta9Uq+a2sxApZDjmoU92Bzk9Hl
tAFHDKJ5LApMfD823n8FlCC3oW+A+B2T9O+58zzQW9VX3jddL7SJDM9DgFNIo7rS
aH+8q/nGVGCHgp3C6Kkucju7Mt2t6eCbYvWjFlMMkigBYUbxmtFLe+S1DAfdc9U7
94dUC3xy6ldFIQjxgxYy7av1/47k9mkn2lbI+4Bbn+02ufgjkVJDY8M1dnkAkaKA
0DTDxDGxQXUHZB8cH+YbfLJFIsddTl8lrrPHG71aKHjQwdPlycuswFwB8ZMD/ZV8
E1KMC1S5EI8TxXum9AXVwGo2VNHtNtwe3KceLag2QOJRKuWwpzexWHxog0UN7mef
9hf2qRaH1eJrgrA4QJrEq+hu/ezVdhMYQvdlmRvTN72H1VJ+PnlpqOFU8+AiwAuC
Hn/waWB/6Rhs7LrKh43WT8C8TO8b5h2214wIxN++tqMukadOACwnj/M3N4+8euDE
RtYys4Z3sYm+n2Q9POBW4CVWCgA2qA5a+eBcfymEgi9MRoNUosU9mvoTjdfMmwxN
g2bNE2aiOf1V++kGcWAwwOT0Rt0vMrr81AuNYjc5B3hXUGdm6XSX9xnZAa2mddx0
iEZOCCIVZQ2hUnI0GfXLmc8pBY7OfmWuKP72GGoDyV/SWvudeYEchFVUyr69sQwF
hApTrMpDAJqvXCqIO4zzidp8919Wih2URHpcojlhiof2twAlmTQUzaXFyh00MQvH
Afe8ahDuNWBJmr8xPErq52GS7BGUwl0LXKTDZ4vsxagssG0SjBWeQKP2w0m3gcjt
lBafdg+UUD/sQjAGqmLjRR2npNy1AsAJmGCii6pUyGz3q97dPTrka9xDT/iLhynu
yt7EAXyXz+Dh/xuwikrXq8vQceh70qfGzSJ+KBmYYG4NFl/f5HBCOosllc8/VzCp
oY4arQQihtUctDA3vz4ImGUdLGbWlxtwE1o0FJKeuWmCJ2ai+ccRSY/IiPq0KSkr
KOPci/ja4hDSpSoBvNLr9marKs6lQori2ZxAGwLqyV0dQqnOwX4J3w+tzdzW0Zmn
KcTG+zX5dNS9LKNdBRspJXrDDlvmQwO0s8ZIsVWt1ZqKzFno3t+Q/PAylIT8XuJR
EvJeP7ncx90xO7UoQfQfPxApDtrHwmOtyeQVGbdtPolX/htin9h+Tf6lu8ve8xVT
AaZpkeHEKxMXwKpYqy5glbyyeTbICVHefSIhy0ooKEkDdzi6xCeByRrC60lBdxO4
iiXaO76/UoU5KKOAHf90zwNvVVTt9S/eIPYNRiYzqkbFe7JriMgXCIe33/jnRi2Y
h+67FVwEcxffXO3bHgJZhTiBjZBQltjiBigH8vW974+HFUhwJVoLMI6H2mQC3Tkz
Y4rXZvwzgdc1khpSswvEo09xTOXjbOINL6aJDmdsGkrMFzr0NHHZ/Cjeb+mtOkuV
mkPHXXOkix6foPoeKCTrUg2MG8mr8Ht2bgwkNwng1U2KvWZV8txV83mujR32mT1v
Rg3icKZdrfniESfceU3n69Tvuf0KmPUn4KYMLbxGwRDmMTVNCyiZxe7Ckf+tiiST
oNpukCPhJ4qg2btZC+NfFGqrL4ir+ZN3UTK9L9EeqhOy/DIUNMl5TDqGsFELyb4u
4Du2tN/KLwPXsH/L2a3Km7bE+ZhQU2eIEySwf9BEnL+xDNQDCX95Pcp2IT56bobo
zk44YWLTepPR6+PXtjG+gFWeQHdEOq15LBIjtm+XuY334F6VKE2F4oKWqWidBHYs
bjNFGRWipqWMie+90M8xchSsb8Vta4WIm1HrOdq4ycQn9PxpDyamUeuv8gFzxviY
JMvT4GDzhANdLWwbGceEycX2/0SqJmyv2XF3hd9HWFxxqcpmYWniBHBV+Y5RvNT2
kJC3KB0I3vQDVucyToZvsqIDWUownk7ac6BCpZLOglViltJGMfbeNSoaBGOJyEmc
gXcmcEmMPXPmeO2CK4p7EwdRyjPKMYTsJLkxqsCii2OtPoMzgX5vCrawmRdeIcOY
8rylCD/yXhHi1Q94jHURLeDHjJQ0QScIbYtrH3gKJWA5+4iQyGk0snChxiUO1073
q7g7+RnHzZDOLqwYBtSWaLOTNNNDsqZ/3gqheJw/w132bMQCWE4XkcI9VfNjoGb0
PZZGgsdk2AysohXEmxJCbHI17h9Wqq34UtGZkJAH/ReEPRONq97f4EpKEmoVVDVB
Fw5u7Ux+6n5mTItn9MgL1rMCcX5yPSh6clcUG0NE72PvVBqn2p2C+cnefHVqJrac
+f9C/bisfl6lUM9A4vyluSyytZWxrfu1R7BiIiWL/1Ld/vu5zbHCzWHJ11WTip4g
RJWbdLd2Q6OtaDBWuZLiGMXgJQgsc8EgjL5Qot6mH34vP7nKM6Gd8AFy6ilDkHuy
SAr96ihDLw748nVO4bSc0aTIxRlkXRCOXeKIN1OwE/RYU3IwR7ARiaWlUXNcvmLw
R7pHckMlX0rSzyU5H3bA8Qet2MxiVPgNdFt6lahw7DD/Mx5s7w4A+fy5AGD/6bQq
NTJA/qD0xds+eToe34L66hzi1fXbrGNwVbk8pzfHSOgDM/TQqyQPltIkZtgFZEPB
go0iddqkoPLJE7DTatZS0lVJhGk1VcCkYUC0MykcHfEFVkmXFua2vhZuRqSNqvb0
3LL2AzN1PBlTkWlzJx9JvDJUpztbP7+Fel8ngPjgjFZYjaPLXbTHNenms5kNqu/B
9snsJsqVT3oxm4uXIn+cHlKF+AKlFuxHgNPs4JQT0f1+RMH9YNFrcDMy1jg2MAO6
jxQTbUCo6oZ382OO+Jyj6LouQlGcLKp3KJopq/H5HpxgW13KZkpdw2w6Bk1ZZi3I
e/jfV1c9DC8yTe4slexBl+VUL0elFahMBRVdV60j74VdAC2jMfutGiimqHFfe+Mn
LW5ozHxjSmyPS1WQXLKTdPK9neGHcsOaGpgdWyJWHztj6OXmwNQBHIBvBgTiGyqZ
D1bEDwfgQCVTVpbBWq/4xxPVOyOJp19s7AE1e2EhsjM4BDImRY/h/6eapmLEUwJv
TFnSBh7VidmNFmOnmFwuA5DbewR6ajeJydO4A/aEw32NbiiJBgKeacyF0W6ZDxmo
6b42hzk9xOm0Bm5pmARtRefgWPIP7W8hoQLi9f5Evk2gtQqkHae3iRekBViJV0k0
BUhVjToeMC5j9KhN1iRHAS3aB6wwDnaRue1zQztsKZWbLDGzF+3xawA5bFsaqne/
jgn8VOcjO4k6Gvob0L+McZd3I8e9lrkpGF85FZJzZm4CKFtce+Qf9cKTkgCmkCNR
Bqp0QX13DAbuVFMrK0rBqFlDoh1PmXBrYnP318urKHBeg4LkOG5JL+TVSubUgePQ
8Gxf7J3/4AQP6aGUIy8IjN+Y2YMi/Lfxe+yWHo1pA/44J+NbeT2mGftCJJ4pXQOr
qxU65pq9ErLEW1gZmGhINhUFuAFWTJNDf7ox4fZWS0o391d+SVkG5wG/6Pxhcv1l
jbtzogGyu4J6r5w8V5/nrWGgX1J/mKeMLnBAxAKsiC413rSvHmtunho05MAvuI2i
mts7jxHnuhM0idObB+rLIQERu0aDGb1T2+MOJyzDOM1Izo8rtsidlD5QfpZrLHDq
eSO2Lk+c81a9O3LXJ/y05BDS5AZwlxjvSOlEAST+ygtQ2qcdp4YMDORChKbEw1Hk
F4JwRNPzzmAAFMNX5Fui1cP6dPFXneOapKEum0ZozbfPpUtyKtO+NbRSwUPfARY/
RJYBv6ObVkfBhYN2PBWQ5qhX8fTbXVtgc4bbJRNE18j/0qF28WZz74dQY5mI2jqg
HQxWl+DTgwtG6OUOgTjHuZ80qJw7gBDWTOqHAExqbdeICRxqtQxKmUaOUEZOiWPc
D0A4+c9Xunmb15fLJZ3dqlAzaC1DKVWuxN7Vn1mMwx87dxb8kqY/2dW6P4oVD/NT
BNE/faa/ApeI1Po0aZGwKf94fIVgzquogiFCCLRe6Zj2tiBu4ORNMMlF8MVSMr8C
N3baVFiSrwdeTr7+uuXczy3lOYyS0xNvGIYS1ml56+0i4yHYK3C5s5hVF26pYCUv
pmMKBGRqeJi3z3PNS7QO4dTpGYWRJeegKudIw6/Tx5kcG7SeCaXFKI17BHHS8lb8
OlC6GEI75RAox/uB90F7vik+ih8hwS+bhxtomoVlAb/gEJeAo3J1rf4o57VuXiPs
N4EIJ21WLHWkzGABUtwBwpok60cHPF7oQSuwxUrLEQYr++HYxeoRTTEDxu/4o1MP
HAVhMk+N2A0eXftNd1a8K5o9p//0QUrZ0E7raqsdvn6N7EvlCgbVrmbGnqYIVBxy
yyha4IQizetZh5UDVKDo6fnkLBPCSWkxy3oPB5ROYS5jxNChgPKMw5Yg212IkIDH
DcvxfsuY/UOh8FoFaaG7LtkOi0J+NaEjrp/cbOM29ofo8CFjqSVUfb/HSqXYZv+w
I4903D81y3NtSda2BvoGleRPXeWXCQ4CD9ZV5V8RFR+0L1ERaNjvjyt4v8Qb5OZT
ZqD3K9a23Elwd+Byb2vMLpIeDWQdWhDyMqUf2pzL5vJ/H9Du1yu6DlhYWav+Q+4f
jNG7uFSHZnmq67kh669C9h+QqneMO9lHB9DORWrzWw5242DQSX1lp7OxE9qSdGZi
4mSWxNO4b+cTMJoTUWQKURbo0XYTqxVMXQwn44o3YA48oAaKxtA5qsTbplnLTAEp
1oGfi9yoyFqX/OHNuWqE3LlpkZTfraBV0JGjabja2b8BIvnEv9eVu9guAX9pq5qQ
TwWrDuX6LA2oNl/eHKtZpvp6fO+e2gE5BQ3Ziws/eswEVkLxgZVPIg4TP/sj7/pd
2Suv4UtWhAnMZ56gXCPfYZsQYy56utY78OGLAVzsaGd5uUy70jimJq/Mt47YnFnF
8dyY58h2FzyF0Wo9iRZqBk82HSBQqObcozOI8ZrwPxwGnzJMtryzx0MYsftb607w
Gwb5LHiYOofLEGX/oXnWwlTuFBHJcz0EfkRGS6tL5disqcnLikNPWdqhTsQdFwgU
2oeTPB3OjuCHriiGZRR6BSaKbw5IXPPRuSjGC7wUXYk3E1YQNrRhhpIosDVV2870
MwaycHKnWRBESpR18kBOlC4oDNfP04Vp5lP54OgyVAzMQxUWsF5AWLVq/xYdfPki
JgaITsoflvlJPh/FwqnhNq+rUHK8M3ogZpfepEKKloH2UQa5JJk1QSg65lQj5S3Z
CqvTTSdPeM+G4Jl+UK1cwAd0iRbLoXJXS59K7jgDZ2jGgdxAnxDY+e4n2Pibq89Q
6AstOWjH/na3vDMS5+lrc1uQTVV1kCG3tcTEfb21a7sjFsaOOK5Ng6kGvsW8C+oB
4jjgM+WgAgGxSkjQg1l8kYFcIr2ThkoAtqGFxbBl8G0dklRkxkNxwmi0YhCSpDc8
WGxyNgNBDgSDAxfp2PTGiCqI5QDxtbMAkhOFBOAYwlX//T17Vz4WUxGNfk3Jt2NJ
5T8bighByhEEvLALwa0aG0zsT6+0abfl91ymDOBG8dRmdlU3bi8uf0RV3TiF/cOe
eCd5H7uTDJH+f80Gb7CQac3aeaUssnQhMggxCAlgkWWIAgqaOMo+Y3X/epKvBBCe
zJP83e/VVJSgt6Lsk2af9lYiQnmEFSzql1Aly8ZzQaoHjqKStngr49BJgAHRs+S1
fw60YzCLt+OyO9AC6G3vUOk/huOMkgdWsaGiR00Rp25gK/3804Bbc8d8SsHRwrKB
KXWLRGKihoLdhpGR72DXbyw2cMmNWCiRRvrrhSP/Nrlj4IVbgneXO5WdPaMC2iqK
cMLXFLiKsQMsckmck3uXOjiWZmZx/0EektnEnTQgSYxcKfA9r4b3HhbSpHr5Q9US
mFdROiqjFhev1oxnccrpfiEne0iUA4ux9k3X6DLi9bXd38Mdgwi+XUvG/ljRiQ1I
t/0rUelwzXQyoV6ATrBcV8FrNPWBUA7b0KVUYTAYBiC+W7sjWrVJ/lTSknDU6RPI
YK4137DWxLqbvhDz09fq4D31IffTAWaAx0iX/zwY8ryPPNfPUNGwsfhf4TVQhCJ/
fRaVDpZdFXlT9+oIvh6CfEVFZF5Vw6eWhomlTYmHZfzc8lU+emjf8AHMtYDuhY7y
kXBqlnIT8zLFkuyUREzwTWWBddlHA63ix1l6L9/Bnck/5lwn7qo4TOIS+rRPLT4z
58/rZrJqoJkAcSm3VjojjgdICagYegEEdsoU0foFm6z7m+/AxaqcbINKgsYWoYdZ
7dXZj2R3PZvPQGWJxKDbhJdjsPe59U6sB9rKfpsjVw85Q6rGTKdHV1F01hmt1U8w
kYmpeGSMzXeceI2EmmIhHHRLU1qJbeLc9eHL3hOUh3qxy2n3o2uH83he/bCVrFtm
Bx/QsRhstZwNuAH33s3YVCaQRFJ7WYqw3U4ijZ92BbJyGkD16/oLdZlvT27P2qj8
jqA0Afwu+IDPvUaqaUGVkyDIVj6YqYFCPY+wCRYv68zTo5P2/eNClGZQYMlbJ5IO
+RiXCULoyS70kZgrQ+ygE+Jv99M4sUkGZFS5FkVNmXInUXXTPRgxXa1eGYGGGxxI
qv4FGHZAYe1enVuiZte/WqmCaMxFcedwHHLvOAJEkqAW2sduxtmNEdKL1OybAju/
bmYGmMY2TVne5WKHSXU4CU5rO7P8GeNCL41gEYo5LGRdhoQxHMqXoHD3NrrqW2Tw
+XkNbxxyyL3tK5+Kh2GoJU1AsDx9SfkPwFer/OW/dhtJiqDWL74r06rz3kZ78BrX
z1pOWUGkA5eBbnFVnXZBG1SUbKNpOgJzq/9HTvvqsbweOGk5XKbzUfigplRauGf3
JjKtomS1K0fV2W37qsZa5FdTvcywtbHP7tSF61IB3oxLCx/NnK8pcMC7OmExiSAm
XT9/wKRsBzH0cnBuqsFXUcVJSbSUfjiCBpKGXm7JGmkytXo8R1FWp6vUsMop56cW
Jp/z3w2nwvfsTS5rB7QdArQqAMplV7H0mdSS9THzPS+v799Y6ue0jOf16MomIq1d
dnfj27Fu11Hkhk9FnXCv+lIDclDJVCxqO5ASfTtfYfx2SZuMmyfOTgVH+uCnLdsx
nU0Vj4DZhg+NGXME3qFEO/Z8NDbFQqtbhCsHW1AUlx8oOxvs4MjNp1V+DDw67xKF
YDaCy/YLKjNzYxmudtz7KF5GDNuOwjMoxOpLXChJNGRU52fx0Om0ddnu5QiReqNs
nrhiMtrG4Z6cd0apjLCv5w+7q0K77AYb0K3j44QGvj93y8Jw091Q9EY4edZJkK5Z
pXXmsu1VsPf9y/HFy8SeOIUFo5bzKRNkeiYsal/tQVdse+lHSu/QQHPD9PQ6YiLM
ETVV9qES9GQqIYdslLEbaC5cV3czppiw1gV0SuRcrAcSsjabGBzUrqhxcY1p8YGz
vjmajIsPJkQPARZs+/LmfiJkwM2MtxqO1RfcCZCNeN9m/pXJZgVuf0FKcj0saDME
GR9EdFfxHr3Lc+LrIPgnPsKdkhE67ceBK3+KZqA7TZVjxqb6daMlRaqE7CoMhM0D
9OqM5dA/jPcjvAzU6PylHvp4WMV+sw4ftunAS9Ixgq0CKHty9/Va5Ke25jm8coPK
UPK26acjsdp6Ph01FXlcrAWrIDQ1H3cEfxtYYNc3T8lkBlCwpfnrpHjxKX86gRHe
GvaTlfrHIYYozACxYQD1mzIlewUN7yYXtofDG+c1IlWTaLSThSdzemKBs75OAAK7
VpvUp/okBCtxSBG6KsSUndxpMPYnhvZL/PPjrTEaS9C1AJrMO+5q5vLgWnisw4fj
l/aYD7uiO7cMBPcg9nrU0XXG06j1AUjbmx8f5EDGVHgbJgsalmr82H1BxcJvpGAX
+oetjbR5M3+MDzRNMBGbiQBOQmLzMJtRNCOtdXiOI5ne3w4u3e8X2eoz4XCfxmBP
80G59xVV8yVMNk9gPASFxmuCirt292NZ/KqbI0KEo5oYraTpDrlBx8VHBVRKk86q
mlAUY3tFqTqAFdf6uXKSIN8MRr/Dj88/0H9oulDJBgVnt/48/F6wwG6B3vP9i0w7
jI3KCvRt3j0Zm7K4dKayAzqZHrFJ8BegfjGLvuklXs/U3gtBCnDqNOk/9JrZfKe6
jlVHpEfoXwjuxw4dcYbyJwb7FoiwyIElCDnvM1ym3J/b3wq9+KIXm1dFgB/dCall
gD5oFot1zkIZAfObLaBfMw983OqErFvN2aXmaCdEMf4va1/Ta+wnMkldtHXhVL5U
SQ6Qi4KYxK2zfe1rSFViLmaFd4yw+nWZkTJA/Jw4g7y0fGSSCse+OWTTN1MczmIh
NPoU0aGpDoN1u2UuMJP6yxEuPuq2KzNvnFdxIWs0s9CdWu06K6Mx/9pyI/rQxiEw
ZGXkpvwyshzvPU4i8y3kXaivJyJBmhE5VZoNkLrVZ4JUe/GaqAqxZfwTZqw5y8pL
kQ0sKaxNK21ZhW3Ipkk2orHyDiYRIyL6+bLmTViuwmkEvXGYPX8ocUi8X3TdQsCS
IqRatsVgw25XG63a6KGO1TNWsZaCDoL/554Cb4zrtdPjyDr2Tm5wSxLynAGHbLn8
vdu2JYvxh9BfNGRbQxBooomD/Viy+T3sHEgc46h0+18Kx2Ou6HH+ime7metOl4AY
7T89PWyWhv9gDg2oSBBCA9SYSg1OphKTiVm/nZusuZBteQM2i+6no/3baD0hDfW4
2bGmruNlZyLvIWZ71j/XCwSbrtCj9d4Da57f8/+D/CpHrUCmIsbtOVaXgqjXE7LY
Yc5fFO7PXj4g0GTe8h0nWGYRq8RTuAOFWROL27SIwDtaI4NAaWF1snrlIN4c2v5v
8Oe/zF5goGd/G+zVjSJ0u87HnbbfPhotRx05GeeCQDqNCThwS7M8mxV939tdOrFO
lyee6Gb1A/NkhErr5Z1FIK0MEoHfCh1DMhoOX5zDo9dnsI/ltTfjs5caC0s95+IM
IHCKwa78piE986S5S1I70GVRYVzVwu3J2Ee75ZSe0PehFXwbqyz6ny1+kKftdeJW
CE5nxnMmyKrVoxz34gwJOguOhV1JR4Jj8e2cLqJK9ihyJRXVkkzR8MymrZA/bEUA
xmXY1jAZ9id42pVdNv+UiWOgM63LHtR8BwnXByPdaX7PPnOVoGMPXcY1ZCPTfJxV
+kgi3A5kvQ9PCwWKcMtPkVyFAlJvDByrJn9AwALognbBUGne5j5iD+mVZG9dj3UQ
3ekjOVEkuVTUR1gl8jGzJDrNk01Gpd/iyrqoC7LExAGCXl0McKPs9+99DHbeFymF
aBCE+j+5ipXPO48R8sVOgnKYXrc5Tjgsdkq1c2Y8rC3yzIcrpC9AGfUBWGmOFkgl
wi1gM/VGocLgwrBvATvUv+W4P330be4T3N0QWzN89f6+byj4jdHiPX5C9n7xFwAt
YCPXx8gKduIDo5pIqhk+ytlKKic4Xo2aeIPnal8Wki4TE7SE6ItS2Xqr6/RdJ8wh
xITMgaLs+wdGygz9EAGIxnEcTdJCt14sfroEsCD/LXxkyNcegDI+78cn4RX+KiTO
Ht8x6NeuGznYnuCuf38GNgRhUA3NodW6M/sCjHLhwL2N38uOkfpo53AqbA3B1psT
KFNrRK+GDd4s24Qym5fJ6C030VB0lz6MeQFqIOVbWU5LjVOHxhNT/LpVkas6+tj8
TRYI4CMbHbJiKMNjCgeCBF4m1D0M1AbJ+DkQAHe4N98SLtslstDG94RJOgqttufp
rqou9KUQbRGdAINfYh6ZvRSNvcVJAmlptzppu9VvF7Aue7Cmn6RFvjuNriiWlyiO
uF7oyRf4BOFDpvCm8h+G9j17t7TKNkLKaoX8E9rvOIOdsEtWgJ+5wl9bKs7qipKQ
TX9kOIz/z40urokpN0j/xPVgGa/XszL0Ttp52oB02pdWG0rJ8gsLMZQM5WHzKwk/
BAQuv7IUaVKliCnUGB8y2UFDKeU1r6GUQNpDijbe+em4K+s9IQqF5dXbOONahOg4
BjkCHkNfnh0vOzYUFKULsWpaoChMncaoVVuPQJN4Jd31i+/+EAyzI5MhhJcSBvNz
+iVauOOUPqYzOFey7xA5X7+YYnBkap8oI1kMpBkYasbATyLmeoCozdwc67kPmbDW
Cbe6EJK/FPDGynXxavN+qdG586kdwIAiuoquv2DPMiBqRaXpuBLI1zxAs+ajugiw
oXJuKCOvdqFwTjdIO1793IUdyUisuxpJLMdgVjWRVU6DpFXejQUD+s/6YEJHl/94
JdakVBPRfhFTZ1BJvrczIQssviBQN2AWXJg8FPyxtiXeprG+cMyF//9ocrd6nloI
eE5IZ4QgFHsjbBNUra7wyxois1wzr+sc/F5U78qTDPeKFk7aVBtJ8j8j1agSgs/j
2iZ4XHfzG1gLlfaM36UOCQvLSuXXTnscJoav0n0iJGyG+wgLsfhobLQKHeHJwOWx
2msEPhC8IVMUkrL4uNZqKE+zZLXMXEa/O+vBGQsgNZVshNEm02xpYroWE6kuUmqF
rJlWtC9PRq0fmaNzpDlZWGEILkE0IZ5Q9rrPN/Hdgo4vLeqPaaftz+FsmlmTETVv
2UTntIkFUZ1tz7oUwcJjHBgm1O8sVqrxtbD5T7QU3O6NR6Qlxv5Ljj25+qR/Ofm1
lNxETz0S6jnUe1CMV2H+6S8H4kuO1WVFMXFlTEHs0u0YDOgLEMK/jzBkMTL7ZoXx
c8KQWUVKQHMFlLebCHuDpd1FUsq7bzvI072kFb/k7rYP10rWZL4/LgFV73CUOAfU
I7cEIs/tMaGmjPV9RNDj3EnFh6Oszp/t3V+j2+HRcbRE7b1kJ8kymWP+smSkrIt3
ENpE8o95Y7XGnPWHUa2MaxR2AoB3EKtEV1mDsVPpD96pdpSnY6Bg2Mu4mjSN2pVs
kGXndPA9plX5wHZXyJHXQiZl/Lr0dMhWduqmNfczThQbkExzJH2hlJ7FOn8THkRw
wwZZ/uCV7VvyYDyvMwIpnqkUy1rxrJcXm3KqvIRkgTBQAlLXJlsisHRUf6b0l+VU
fP6Pr2jKVCNw34QgTuxjZMCwT9mTZvjhupPaXpereui/4852hL7wU6T2ztMVWTy2
07rvTwHo9XC1XN78QjpAD0/6rIwj6p7TpnjM8N3vUyHB88BRZypl0dcUdnuIuj01
+qhA075zZQAYLCwi3ofHlWbZF4YdiAkDSDbDBFdxcQR2M45+hLsl9iUp1H481htu
jWxG2A/85F+5CckYfqupKHxP/as3Z939mzwOLUAg9YN7JUai/RsMFfTS3hXfa1+i
bhG/Fxu1bhjmsBt16vtNnwV9WWEVJobfQj3EwHPWsgpPtgyq4HHw6r72bFhpTZQt
UHkQw9z9Oy6DNJkPD85TgYckT26vP2oBTxIuI/FSNTEHy0HCD/0VR71ltJYsjgfE
mt4MDyMXRXuzG/2pj5HlkmuSf0rkS8asyoYz/ZEElc0JFKSoxQiIonszYrDL/euy
pyBoW++NKiyxbw1GccH3ZwrX9++fVMPwnkFC+GXj1y2mKYqsZ+JkExPDzb7zAORl
aRB3W3vRJxux8Tg82qCvRqyqGt03nm2TIwplLwRQ7+/r2dOtS/nrWljYLkexNQnJ
K28vB4uC5XdWKOnifUvo4ere8Pv1wzoStbeqDUKtzeXyCxqthcmAsJ/3ghWU1dkN
K+Bg8gPh4ZMQprtHci4ioTmKn1oozNnjBjSCSnHkPY1aQ71AJBD67+XYm1KFqe07
u9XlimIjVcKkBtWXZhRqxWSwsa4u4HypSQYdgtHxxpgzUkFLMzjEeiHohqjEgD+w
2QtcZJQOhkSoJcJkw0xbqX/7yEgmITcBpM5sv/WtibXVwxhmNrBnsKrB531CCXlL
lEzgos0W7PeE2By9gbxhj9ikuVVKtOoHZvB4XsyHnmLIm/7IrycPoS0mxWAU56Vd
HUCDEK4FDD9PSaY/Xz2FmXljFfN3ZkKVYxJY8vOU43caIyvOePDm/ggmwqol0ncE
Ls/1gw5Di71urB2NlHGOCCfWG3rUwJ3E3Uu2pz1zk087FrlbR5eTClx6VHKbJTTy
mgR/Z12S0VNEQxkVAR46mdLD2SJQoCl0xP8b0+DNqbRKvxhmLOLCmGmkaxGTZv8k
gwXzU9tjKjMlAhgT8P9KKRVFKdVf1gccLBozWjcQ8HHZjxmX4EkzU0FJqc9QR4yr
xgGk6EOBIadzUozsKfO3Ok9YT1wF3IvypTzkI9uetwwUEJ6iUzV/chePsXwKxDzX
/6Br2CFugBCmjX9Jt3xHBCQgcDpqmSmdwoeoL5ILyb5qhIRsl1lYdIK8ytazCOr3
JtEcyUlz7Rg5LVbXCUEZ+ESyrY5Of5FiiI7Ap5U8iRodwB084JbzfqJez1zqZhjI
UZKKFh0FtOWWZC+2Lyv2r09T4CfHC9rHBzL0eJmyIW7hJGY2E0WZINpJjYrHB09Y
+L53ds3blnh1lBD8kSNYRfLYEXJ18brr7Tu57rnjWttXjBE+vRN19ckK8K+n63Uy
BjW7pi2H/vhHHI9/d81G7yC3ErvMgbdxeQFyPoXUJeK8xUJRHXMnTMQ61rbfZWvh
UNw3oln5F5RKSth3VNt+XcAJvBgV3nkwDFBwvvnsKcmD0uVxb7k5oUQxfTk5QNJu
l4cqYoBDyPt+twy7Ni2j7JD2DIU0ZgxkrxW0Gq1ZFpS9FYTr9Dm+5TR3g3QskdX3
5f6cvTlIegw1vfqUXojKOkOOYQZA0pI9YeoEBSCSUBWvM74A7r9F4lg03ExcULGt
HP4CD+C/8MQ2S/YdaTQMbkY1TEitrYa9iY0QvO88PC+QccvCsGZjPAr4ScOBfu55
CBanaHlCN4fUndT9dO5Py42pkdyry8bPbIjtWKOEudc9tin/RMZLvkOcs1yB6fcy
ANlDlFvYtY9YAp8HB8HQ0j0FljCx7OAo0Jw+PiWu2TCE2jR80FJDb+ePrSnlFy4g
yTB1yLkmf+dTBa7dmsHAx7juVFDiiCiixjGHon3OAj0GR5j3VIQIkHkQezlaoplC
lykjW+1Gwfv37bh3ySjtaXXZkQUDHY0GvO56tOVRdZp8p2BxbCykgH8dAb06vLmz
fFJzCWqn1UybgQkED8z+e22q/5YnZCM1ckXa6ur1rz2T6JK2FYNEyPumtJSiFuU3
jFUuQ5F2XL2FpHOjzcnNcm7JhbuoM7uNVmkl+LTrRR8CQlAnwFePriQgr9lW6/DQ
0g4Hibe/TL7WhRhd85LhigONUszZmuPZlKO0L6gV4U3SObwvP68bRwKQc1ThXDzQ
JczdY4GhCGQMsnoNDzTEzD0A2Gn20lzz3FNngD1L+j1PhYFDo8Cucp4YDCYUsuMQ
sKl5NtCvNY4+0IRf9jYl2MNXcfe8zOglIw1CYQlKKm5ZrK0N6dVYPCM2sWVD42Fv
MHAMxsx8m9+R/yREGHo4k8He/cGfFTxqBxfmKn0CZiQHALnr2qs4yFtRGZNTnNPY
47ZSvVSnKWLu4S5ZN/0kV80wkB9A8UQPKwO6ER0LpvvYQDJaxXpdBBuSKAsz8Ypf
7wxg/5PS0pcqNgl9kTrK6z4oAGCI2fU3/w8SoyKYwtxIt2tCNOTNnq1LvVFpVrhH
lk71shdPZt9J94Q/oG9fnpHDcol25WwXI0voiVjHncXX6oqP64qNFlTkm8KPJNwe
nsgHGTJ1rsd19Tco49QTlcuhHXuENWEV6oFRCOKUWJk/N9rZmngCQm85G1Csuped
jPsejLg6FkM5TzwPqriIZCgu6hkHYi4Jbl7Ar65s14O3pOx4WosVW+MEgkGTTsFQ
6lP6mnXZa/L/B2l2ysW/bJ9cUBzeb8j3STtGlMB0TGs2+Xv/7mnCcvmuiJUs4MVa
VMBrlLALs8DjeM/t74/0rnCxRs6pME2l5fkAJQOwJbNc2YDma8gy7deGwoTaf+0J
EnxbcG8MviNQSqDwRcwjmOfEEFsM/Jf24RdTKoWfQaKIKEahCbBmiSkvvnQQUU5S
4D4LME6Ba7N1p5thKLG+F+A60fp0WeVFRVmIZBZcmdcQkZeMuQltbo0r+rl6yhsp
j9Wv0GowEkisbYwoHBekyIG8jlNfbSekebkiN2XNXHBQsBvgxpjPGMKH9WpC2aS/
bSdAXAXVLPinL2s7uSmDPCEdW641CNmVm6FXetYw+vHF4d5cEEO8sKgSbbsyWBFq
6E8brWjNuPyR2tLbtSrR6GIe2eVNsUc0vAX/tP4rJaSxtfJkJ/b90pIg0n8y8/Ed
j99GOaaQ1kJHwu+hhKXiq85TF968sNHKeAda6JeSqyH1HqNXeZly0F4O1pKav0zP
pyshPYDHtpPqFeqvqsHPkGMFEVG8ZyaUacnW4MRyEFbf/KFMwL14jeC25JlcH5KF
Y/s847ye2MVlfXoo+ZHHf55Pq3w+zXbfrcuH70j8oAYQIRGeB6Wcm3weVYZMslnY
NxD6SKBsKVlnYgIlhjO0zJdE/FzkjDp+O3V2K4ATZfz3Fsph6GyYCT9zDfhByQcC
TUA6uC1wHaR1/H9IMKNF/zmB67iWpsr49oRMvp9J2fpkvPauQBcYR6+qDQXdOnyp
VqexmW1/EZ6GLI1BCd7s6Q3G9ilYiTw5AIiK0APWTPMCk/3kg41MGUqZxIpWFMAF
OmiHhTaNigLmkp5yKtUjSJ+HnfpySsoA6NBQiEwbjRACaLyUpt3jkUoCidDFxoXr
z63UE0/XXi1jVG2nJ91PjegBqN+pxxOXKGBOyZttX4gX5N8PiNjDD1UpnwUgZZgj
Z0knX7f7MZK4I00SSAJ1HtLIaYXUMQPqFtGdq0abHrpTx9D/woxNoR0mXP4IdW2F
3lUeQShVbvS/oaTzz+68Fm4ZO2Qwv/LnlfhyV40dS6AbrnUIF7vow1kVBwOyFDPY
IUrMxVJnnUXMckRrT51k/O2VXdVZ0U1uuJ8poy7OxkrbNg2Qnff17og+6ZKDYRCs
4JGiEyCmPPZL+XtEt49n2QWt/V/12/k3/bXUt+ANe9CouFK7afWDGmzBD8ZvZ2sV
l+9tibUPBTXelz/TRgRgFDJa/Vbf/1i7IqHTHeKu5y+MjLBd5JZf8nwVxK9Qb0Hu
kYlHXAOczKx4w/9L4X2+rkFsO8HaLGQnqDSBoKxGDD35BcZH3ibl2+1GTqcfQvTY
tMh030XWTyASEGPg6YcDpL2VVR+snfo2TnnIl6Ufa/8UKDZkx18DQ3GnQWnRqnPa
Mg5nhY6WIJqj/kFHwf3d7i2Sorbl78pXxWq5GW335xHwa6dzPoYmPJUk6LOh8ORj
0fMj8VmV8i31YiWQl2LFzfL7HWDH2I38hq6Z7Dpm5X4WKqK7wlW8EOjiCnvq9VAT
vx8FzygteQUDzgTuj8Qt6dDw1i5T3hi7z7Hl/ea4qYcnfJnnxR+wU4g2OO5EIW8D
PgFBV3MW1pfi3fR2Kl4ToMgpk2LQB7mMaJ8WwP8U/1zXdLp74DEGkOVOaJMCWtw2
Yyrs37dNLQ+395Sgu2XhxiMQHIrnDAQXzBAQ0AM62VRDwFZ2utGhrolwhKEf+cio
IZZV4Av0MqqTeUfLf8RiZC/dXSg1YB2h4O1URaGI/KO2kX+hkZNDvVn1zfQ2VMlz
nf838dIyRdhVRRltiFiEBiL5LNbMrPZD+kjlkNwN0szXAsAtYUG7mIMGV4iekGK2
cesiZJFs/e+MH7Ag3xnAfOWb8LEFUqW1/UfjCvvSxRB2WBlLB9VeSP3gjCKzu8Kx
VweUic4FGiH8SVi45XDCQj/+/dTFqQgDxAZC9Cs7nSjYhafFo1j8noiqIIGOq5hM
70tUFxaJwZeOXGXXzMWXky3+IOa5MMOHdDwQ2NRohgQPLExQSKqoal7MyOk9ihNb
Y1Su6f0BT7JJBR3G6csfL0u3jDjKvBiPIsOft4gbMqybbursqi2Cb1b9koAsM5s9
oDF2kGGpCW1cMZTRhoEL6L1T7YeNkp0GGKqLhso3B5TUkODsFKGiohZlgLO1/Dhz
SkD/iRiUkUzavBlzTRYyfbjSCz3aUAwR27rf448wlO2udz7r9rFY28QPlwhqICgX
hB+Zi9zRsw8Yhwb2+c7jtjWqVn5YWmHo7f5wFjt3cPMv/4nsXtnoTvJLO0AxJqHl
8cGiQiPDqzUgB0P1hV24lBBgTwp3IYkH7+fdEbqQrsx8TF7C/AnYuaFhBN7n1KIR
YjavjFp+5Hs34yhF2yX+qxOYiCDqNAffNF5vtO6qdlcbN5JoiyG6ialQg08KmR35
iz3kWRs34Oih8s3rRpGrYlzRF9cCKoSH8E49Y9h7f6lgVbn2ojTjasB4MHglD4/J
Y5mrpwLVq+odrgGWx/RYuJj6BPvdqErAh7deThONVNE8ghC2RlgdLHnqB7L2hwwA
QCeM7D2UFms1CwNqRfyEMwhgjbRqx4gDhubYh43zvC+vvk/CrpurrT0eg/HK7ncV
uDimkFAt1JKnqbVQ95KMz9wnNi31tFEV3e0QCE6RrKB5HUcV3LApwrpIoRTEoGqL
UzmI+Qfh1T3cPzvsdViBUkrhmmBKPcmJHvwZZUfwg/xNSerx12laCTXPgcRFTCmL
I/jvH+LkKC7eU+sOp+lLsCWgxPRkxdkQPAfKv/VbM4IsUpzuT2a4gE2oZGp4XpET
iQoZOQlNDHO/92tI/93yPDndnKt6Uk6pHwbh5gdngpQ7WZ9HmO96JcxlOQZwlt2S
+aR9noXgePAB26mAYMW+eYqruwC9qMrefqJ58QcwLgD3diSDziPTxRWl8qe8SFVQ
NI0hJRgXioXeHwR3gKqghO+TSJUwNYyD+jfj85fcnTjAlefb+xlAWLChySUf4jif
nQhAc9baPSSb0YuyYvp/UH+NZ6tutYVorOYCez8eJvk//Io2B8KVPwsdygN4TzaZ
2lpIFbtc3Z4OfwreZveNkoixzJaXr8iyriahpf8ESBUlUrvVnNOkn140d3HEZXWh
3ka/NC41Phv5LFomoHuQO2Pw2kDzx8QTfszAoAPZVLbGA1ol1AfT5ILto1ILfsVG
uOFRkmBlvikv2t+qPJ1DTW7n9WHHbo1ROQpp//W2bdBtw8WNkaJMzsvUHzmtt+xn
GWK1Rt9Oi5a1fvXbrDp7c3k7aVcESUHSdRMAPjLwiEk8KqreApN4RJ5goOzG2D28
I3WdZInArcDti7P0SSje3NDhFGZoBbRwNVnJUOL9UFDEwkiBW3iBIBhQfzfV6f8e
HhepvHhr2iXH8pEVe8enR8xQMwP93aBDvjIbCjfVYTYDoyMyalJ6nCAymMugWTqz
bAWPgSUnpVqntvl12GclHwCqrnYAGfyQFi7mNSRvR7USH7WaaAv6rfU8ZdwKr8eW
YeRzhqS7CiLBCo3vSRkI9/S4fFFaHvAJSnfuFWXWkK6B1ZeTa1JGtW6earmqAf6C
ICt50pzKjIfnfQVbOhJLnWk+u6RljoLGLQrwQRB8kVgYwV0GeuTDuSLVUtOir1QO
PzgezzEba/S09bYaRCqI9gYo55igah9a2pveTvBdzUtj5bYUPoFGkDzyPW5KZdyx
w5DdjHOhhL7yzmiqclSn+2Omo1g9ZdkVmHqscNUCflNehMYFRodlG8aHtQE/mGn4
VzKapXx0LynluvEmeWqorANGSB/1CK8dHv9+ZpahB3PWSHWSDZRf9DKU9xoo91WB
BdBwlok1vzya9VjqA/inhML8gtIifSMcnXkwO7wdMvP38HvlokZXXBOFP5mrSNrZ
natfkb/+xs9bqOGX5Bdt61jHBZEXZuItBi+YODjHL3szaOSnbgsYUwfl2P0DzajJ
w66KNx9Va6KvjYGoyZXrm+fQczxKTQIYPkRNU6nSbmNOgD4X1KYt5uVMDyXNeHDp
Y5Np4n5pGDIBs0ITVYLMMLwDoaYN+WB20IzbFcfS7ADovj+juQvDyo2ziEmzVvgX
Fx//Yr+sgKRDLWR3aq85CdvjVWQmJGcM0h9XZPIwaAnzz6HRNiggWgb4HD49dW46
V0WQ9JLof3BhwO39FaUn3f++WbnCwatPFA8j6nulblNhV8bB6Ok1k2xg3sCnsdpq
aDBp2VaN4r+8rNTlQds3OPsteuh4r841Wl49+k8iJtvJ8NcRmt8A3GvFRXCmTUMB
kbg5vxzpzWQzXF6K5dtvI8AeI001+vcUEb732WoGg+fKPagffBPt8pQSQEWoNqs7
/vMcifiYPee46XziWhH3CuqDVp4aQVXsw8+XGrMSoajYD3Dhux+RkuS7UHGMZL26
7iVaS6Asv1nM2/HKUz1i/AtdzTbhg8OMGECBoXI5I5VFdOHbFE8x3u7s4LdBCW3J
AF8JH8zr8LZiyQ3IhHCyUd7Ko4QjFAKNQod6Fi07C44l7jbz6IgtniLdfgi4et6o
FxAqCnAl09Mz9SFQ2fuGKIstIfzWFycHFKRO7C19C0CfBkAjrJCAYXU7keXa9K06
rHepPwLWbxixbaAfXeWM0Ufdus/2FYfVpzrut54gmHRFy3y8sB+/80fk30NI+t/U
OOhz8ZT1xnhBtjqqZMoLKIaY53jp8qlDbKitKuxPq4dyxuuJMo74zOHylzIQnFcI
WTAic9iF6XFNjL1VU+ly2gESktkGkH/UJct5HCbXdN6DX78aX1KqKpnenS6sghiM
XONK5p/egGtHJDoBbZzF4mJaoVaHiz69OgGAuliof7HNMW8tDZKHGCUSvo0zXdFi
euwHDD6uPvVmzemDkcUpOA8a+gjpXBwz11Zv565h4IFI2IC/k0411chNNa2zH+1n
USX5evo55TjmIZF8wBipjqLJ58SbScKBRj9U44WmWXQZRJkZnTN5Ee2/jr9Wpv5P
C9jo14DcflIwXfnVjhKG981aK9JWrb0i/LwLuZPAsrFNPSH2gDFUJMsY5qvmmfl7
Y6VEfr8K+wY7H1SGpE5dAXKOMcajkV0ti4viIsP7oFLmEyWwUskAVh5SneLwn/WT
sCbR8wkB8bJqhRtEaVVp9RW2yLO057ejCCsskShFN5w7Ge4QH1scT9B/nQrJa4Bj
dLerVXsidX47t1GQSWqtTvKC1C2trrAuc7QaE0iraRSVfAC3Rb5NOdka6UPrzB93
JS4Wa5ZXn3wGIFyzIX/OgD2s2U/oEAZuPvGcoRIeaOJ25a+KCwr0CYqMgUga7TDL
pjjW1GRGzWS3ozs/dhis/7KTA9CvdsbXLE40LleEJtDfUjivc3B14NnEQDktaq4O
IWb0pbBJbtPF/B2CRMuHeWkUHGEBJfFdsEr1eh5X1V2r5Y/HVYtgrhSGnbBicKVJ
FdpyWSs4URQ/iFy/DDGS/hLsRLz2Fj/VXQlv0xF+vRaCu8kUMdnNz/wagjykyZR+
Iv4betyxz3Ad+qVZUZIeFOuB28MNpf6nJ8zdBVwF4duTlWOW+6CexZjVJQrETB6+
vUG5DnZoGxyPQTNfN/vfYSIyh4CC39lSllYaujw6Lk3LZ3ctLIM3BwJnn5rGmo4s
lRS2PsNJFmrDJG8OhEkfwKf4R4XYq5Fxv6e7n47SEu4Cx520O5mnOQV+bEZRzNIW
iSwJoOFbTN1cMvthPEUEhJU7J4MdFmAjXZXsDY11TES7fs8NudQVrYs8aVtNMsW8
w9US8d4Sroa3+UNInLrYmIYn7ox9Nz3DlwmEoLZ/qFlq0Wu2HC49+mlD4jtxoEVh
FTmCa5kv9Y3Hp8pfhrEiba/ZXPbTiKxQPFeJd/HZJZ+bgFJCImwv9spbHGePO87D
e57fNym6b448BBy4ar8Na3necvYnrD3J6kQsL4t1cBTu/Z79OS3jN1QGZLSLcE44
nsylwYnY5GPPbmgNnp64keqm5DB7WzqmdEMyFhFumPDV87ceLrhRp4SoTCkWiv1q
KoyExji858onWGO73t0W/ArlCGIuxtAQpn1kLLsB6bgVnmtJqNAwQEqbxznHIpiV
gQAo6BKwi8mS7gHEzEifTYnI0EUIdqs5p3Nk5VddarBmrvFwOVIbzsYtdKliFeOw
y0OeocLfkNQaRrGI/m1Lt0KpzT11KdFi7WXqTScpVEgx8cq8FKN3G3LlYo8w16wp
XR5a8iUfPOcMWAXqu9I85kq0RHRKMh5WvJNwCm1R/fnQTS3wDl17e+UZv1a38lcW
NXvYuRvfZS4W4e4Ht5Q4SGhoD2MWEuijaUqv1kGAn38gxiUwqzxVLWcAKLp+6+gN
AR4USgkeUke2oVEUW3AmqgWM4hnJTqF9gq8yz0s3/lzsizh/jE3AAIOCwlz/3Cbq
qTdDy5LUzxM/LVICa2al2YQr6a89KqIqRKKQbmLqoy9lkLO7Wn21o7dtkPLcwyW1
5o9SnqPEE0ud9rpOQqNDotgg2TM8bwFzdzNGro7CIl0Rx1ioR0Ffdkx3PfHHx8u6
TxNMBef3fuXyhMocrawaa+mo6xFXNJx9Bp6NoC7BrZwsXvDl0IduGbHsjXkUPTIh
eq5PgepEWpUYO5/srO6rptXabWFlWbHNEAKibWTeXQjoLqvry7LcpgXe25T0rd39
vQGGycfC3lqeuQk49HcteEAZLEa3/TX3w8Ub0JnvH5nWAnu6MIeuAw6eSV/c75cM
1s6bpnE9CZ+rXSGVHXSGhDH1m8h1VBBIbTRW7vLOgro1CTQ5v/tlxT4h0xPKRfEK
z3dyPAiDHpIaqQWLnxBVdRxOBMSuzJw5gMfJCyqzp4BRWIvlk0rw2GhR/8eWOnjk
oIuXoy7YZs1QHMeA8gjAANcdbPJrQQ5+by0wYsCO9uPDkIosBqO5bRDDf2NS4Eze
+sem7eyuTVPagvN+EQRAidB6t5OnvtoiOyGbUpCZNZ8ocx7IkHxBT7+WW8ph+uJe
krduhs/Gy5NUC+Ss8Z/eLnhAWedW89YSdvcP71Jt9+8R8pZsaEW0D7QqEp4GFbMd
2XrWjJD6gkTFIZbxLDp+clZq6Fkr+SGoMHn6f3zQk3kGsteRxHKUqapfW4MIKcnH
e+EBkLlvuqEbIQNE5VBb2qcwnoww6OZqstXLMBvADczE5xu6pqqqGKkFUmoGOrQj
1EX1q1qIGg7xHJMckpLe7fKQnsmYe0nS092DRP+fNYYVrS0gVMK95CgcWB1hNav6
Cuft19doy72/Ni9cQQqTgSdFtEqENPeOlmD32Hx3NexhU20Ia1XTfxw1HIzCHgGB
MsG2dGwkARBbF+0Flae8REo70DQzXRrZNbG1QRu27HrM84Ur9Xfvc0BXF4S0YaTQ
mT4iJgkEU97Z6HJD0yK+1KDjHyq/1XGYeD1OOt+omHESXzReunPRTvILeaMq1LuQ
us6VCoVzn12QgBoaiGdMu0JNlbzRq/FXL4lvKF5vi36UW1nmhFD2VH3xyRrC96pt
yGNL+X2+uPAvprRNteVOvGCBc7Y3ZZvpERuFN8HwQ341d85AXHKmyRPKUsRIAGfl
K1bPUz6ukvC02Ceq4/VALgsKg/STgxlz3a7Oxf4Hn7q/keLqS2Q0X2WeFljCUS/L
00TavaKh3zfKNTeSrwZ2LcyG9YKo+1pJakytOffeVBBlEoLHUb8kwVC4AJB/fHUE
KpYSoHDo+UR1qLr5ljna/2rTo9i9QmeUblHjGZjYM+Yjdn7jw4AeaVv1e+zDOPMl
gsM7buf+UFDf6u7zPip0EdxfocGsccmpPcIK0JOgMh/WkXYuhuhF8z9o8+RLRuPV
1gOQnBHQY441Ywpmp0WsDy5wO8o0OAGsV8WB/+ewu9ohPLq/UgT87olxf9sxFJeA
H4GbQ4rewnqmN3KEqSIWBPRruCvc9q+6+0iUrDkQVBvNJEe053jV41/MXe9WxESF
Dp7TKNwzF4wA/Tx8HhJsp93GFXkbz7DOqV2vUre8eO++gWNPURTxQRZIFJgMSJYn
x6YdYemayTH9kidJFsvaH5aoJtHyZQmWaZUyi2esGbcKiJShnBKWuaOHgzdCcRSu
U3DhTn1KR68WesOAqanwt1aOF0HEICyh7Mxlo8CXYreW2y+ic/8maPLkwjhQTCgB
zvAKKTZYT9CyyxV6+y1IFF735n+nySn0FU03x1SATV8BYnlx3ZNr1NlCMB94u6Wx
kBNdf3/dffKy1aeq6EgcLcN2pJPfXlofZoDKJZIZLb288qTLoekjKlIJMwXLT2hk
YsNf1vsR4ytVwbVgNXAZPYmbTahFV6V5y6WUuFqAaCxCa/p1Y3O7E1mHRhAP+aYc
HmeGi7tYyi1pNl2hVzuUWLA4b1GpmEU5qD/SIY0lXQLlmjBYoA4//RAEZwe7xIv9
pw51BbWOcNubkWVuDmN2aD5cDJkwV3wiImjpX5AIQMmPaBTO8VKUw3NphC5s8/c0
eVIoge2NQ106jPQ18S3ktSZZShTLYuu7R23l456M1u0Km+yOjn3QaVbre11v0v+B
a48xUJBuNws/9xx/eexHiu/BHtS4Y95GIgv8XHJxfZ0m+iwWaOq972qVF94OUd/y
o+DYZPDtZkh7y2Ro8+sr0vz5KUw2pymbjknyGBPy5xINOyVPwdAx1LVcDZm8U6wh
FctKNm6VgvXpM0Ix+WADPmLtjZydGXzrs7u061F3C+rdikLafVm8QqVeEsnPX3HY
G00vyvBgZ3vxrTNxUCd+cDq9GV6MAH7kh74tRdl+MN15jnYYBKVidIC2PzO3j2x1
yaAIDM9Z5tGIBYac5rTknpBBho/MECma7gRPxod/e49nr4GRSx5dLyfx8cLuPOQg
GJMHERh5UErZGJyWIe+4SGEMQWoQfnSqEarU3aXm6O4W7Y6KXuCfEBBNEFPghQoy
BnATH7rJrQmy/vI5YXdaZTcm0hQlWZLQhi2eTBiKAAKIGBcBvrWYxG4Oh//IT5JK
IHSmMlkam6r0dd0cQR1zTh3hKCzMku2dyPZXYuKQB3Zz3BIWnVZo0oWOdq3E9fpH
Ui/m/Qivs8oAnibToEIU5AUb+FHAAHhYTSUdPPV0Cgs/n2UwOixgyMzmuP/iZNFG
jDRrEVsB1D57LNKLlBf8YebQztttsR6xsNDEltryT/ROO2a6TfDfgZPYRe+49Y8o
FDNOcSEeprUGczKLjcD4fHErwFHpXclH/ujioinVmCGlJAUKRqrBCGkUXTvscQW1
nK00MiRcPZQRFQ+TSmWASA1pAFs6ehF1bXgoQS/I9dk5BP7XmEbPNYRpvfsvITmx
XIeCy84epZl3zxtariFOeShts/HizJJNFXAY1LUs2d9D6ZHmneQM/5SAgc3/WNTi
xCDwgbspe5LIBCHI9oEQlFLnWbAe01ofrXrV1we7vVZz+EfE3YH2ke0/skzIvXc8
yB3F1fLxbRYm0htqcJE8A43sqqzdXjHXbenY2FNIGztASApyQabw+nnRiw5r7j6e
WgtGKkxeIs5rArE671n55sDufl4LhEZgmogya5ykKGCYQSjNAHvzMChqHO3xqgT4
80KMwy7ngSFsUhnvCg4ATZV0AoZjuIJ7y0kIB4R8YrIbn/td4fmaLClBq0RHhhoR
8N+yWXDIzRXUr+kYWUBvk719dg5LGp50gNZmxshqYVkJuPaCKwpY73fwKTaZTLLw
Iz42sxc/qdq21pEsLda7DWqW2tOEU9jjxOu4wJQGUEi8e9EYb6u2h1u9bGzjCrCZ
cEeQcLifmH42S1lzcPdG3Z+9ochtLDjC8XxXrgsNchv7lTsY0x7NlzpQeEs0B6Ed
zBeqU6dwguGqaRvWsCyTryBMnNM0Th/SaOD2P135Jbwd5Tm74vXIgCJ3VwWv4+sj
H3MaBR/z75DDl9G+mIoLNAJsKVbRBAQ5Wamgn0TwMUSz9OOEAnqYTxJc6eV1F0V6
AOMN60pRc91/O8gmFv4IgiPDP8zlNsetf6KjJx9uH/tORLu0aQqd/NS7kPps5Wf6
72uCcCe/9kczyObN4Orv85oFzme84G1zl51ZxnbK8mPb9NwnLpctE5O67C+ymD3l
2g3mhkjQ5Oa7CVWfTgSdut+7EJ4b596PpbnMQfop47mwOWn1bGqWQdYk57sU/2Xh
tysXGuvY5YJuSifMY5Il+63Pb02SiG22/fWXjda/yNFtZmDObZKiy8osV9KS4WDd
DkHrx1GhEH5MgHi8VY1+/wDVvwU42WboS0ShBuZzbeEw20BdJjAEtExuzHlcz9Wj
Jh0VP6ESUKiyipYSo5c+p9aVb9Qzjlp6lUI8TAcO6fu8HNh6M55Ty6xljxYPuFXG
HpIoa+ZS7/0HoT20OseQGSlBya/Aq0lb79LEczICvKgLHczvLrg0kZQNAdvrmiD+
U8N8XGI0UDCiY9n0YH6iITxmdNxxMECv2ZXqigYK1VZhOGgWsgN52HTieglixw4d
df/ON+5i9ZEq8q49AjImhwwQzNPbKJDc3IqGJY+V1uxEiMLxTdmtjN9zsqJZjCxN
HueMFFnHQuY7D1WUd3Z9011/nF2SYN5nc5gsWEuM9gLR8wSAppnEBNFlwKv4sQeo
BewxUImIJjAzpS7IgkIPzEwTnVMI7QaV3BoQkvn7AmUuAso695w5YXKu/0OV0aAy
2AC7t64SDW7SARh5uL2K+WSJD8OfxNBdy80LFeJ/7V7/sq+LGVLouS9ARRviyB57
kyEIn2Q8IICXX60/gcCzR1ge67Ed4QqScLRSJgsnntnLBIxjvvFeyNpuPE0kR6TG
MZrVFy+TeWiJU/tWbob0eIJgXWh15oqgw9koVsa0pfJ/0q4wFy9pDilk87aX41KS
0BXzvskELOrCn4JEpzLMEbD3CpoFpYiFXIYYEjn9ns1uq8N0AQMgk5He/Sfxa+M8
0/OnEh6tVAdg1KuC2wLV//ddEZzFbXnGbJAupclUO95tzoh+W1ESckgbB8RAHbIn
sVTiqvjkVgffEe/TiO8SkF2umHwDSE5zQXvS2XjHk1ZLsLo2jlOjSMtpfEv1aMPK
r2kFaAiBv4qB3pp7t3seyFJwKD9WNRndnreF8Y5r/UuZYhmiYnoH5oNAoiCjr7mF
uXeixuMBrt/9iWEoI2hfac1g2NACh48nEufFM0YS7YV+j9/3PDXLlFpVmt5e+guf
3rPtoUORMqdAhviLcscp5jKY5Rc27UObRFSYLau2FI26gaigDrkMHbbQrQ3z/2Lj
Wk+bkd9+4ZdWUtKD3SOk8/8fMOLyFsgA21fXK972R4J+gPpVU7Uhyj4e5u0uEmix
clD+HijO/UQgWR4qLK8KzYeB000QJO7rwgoNym8ccnlv2yZ2P8Dy3Lu4THqSYhIq
w9zV4L8IgHnPzh+DPUwLVvNpEl0HaI/cEZm0lbYuS3LwNqODvvj3sTpiZZ6lQSsG
1nYcHdsCKsAmZGZhQ2MzCBdeDrpeu88ZDxR62I68bhRs99jgklMNg5MeY/CEMUG9
VqtyOWpgHVqPaZNKnwOcgL9bsNe0HrcU+Khbw4yxsDf8eMADDzq2iWwuh2u3Vf+r
/BBLM7XuWlxbzk3Jz47XxXtBXKNQ6tbbkXbStpJNh4ptb6YzzFB3dMoAouusfF3g
dmqRWTztoY1fnLZfaqxAwmfognIKKe526fcQYTpONBArhJY1GqACH9WaCW2UCfkP
qbyYvkR6L7BhdJ+FXVNojqsWPwJZT2E0PPNjNJatPGmOJWL1W+jxgYKOLdQdD71p
0P7FXoo1Ou5UnOJoFEH8nDEU5K00V6HaopAGCdXBWv1IhkXLayZW5xx87leo6zEP
Ag/wqQQ8DAO02ifAkwNYW/38/f26YfifOuU31oK/1ezg3U4gCk27KRCUqgNVlZtV
cm9ForE1d4t5yAapa0Q/QackQVyzj2kELbRFaw7/nCTKtgRviHBpjDzLWmwL8Efj
Fmw0ds785aD6EVItEVcE/edPN9A3ZBAa0/X+5Hpanxb2Wj9Xq5wr0GktDcHstDZS
z5tUfcHKTsVLW7bkOUuKxedZIcIkWIRkBHYFYxixpIbJPh/0DQ2V0JfO19+pwWoV
bBYkxMWTyrHrzTsNKFJEOZqaf2istJt/oe9XGcyaBU77ae0C9t1NglROql+98Gyq
mTPqfoERg8L/x1NuSvpFwLKvKN6rxuuzAp0A17KsgVN8tgjiUqOwkSLUqfkWczoB
4KvOghj5IIHLTVkCgyYq3oC+u3HcW76Oxm1I8YMzGJdmOioGsmL14+OYsfxtYee8
FZ/L6D/gMqy96hctbTi3eP8MBR3088O/nAvMW57xm5/z4F8H3yNTNKHTTyRSlI/M
ozfN5JbqsSYBYX9lhLcRsKhpIUH//+LUiGpNh1igGnOl5iWfE3UlT0dqj1YQTC2G
hURDiKKKnjj6WR8G2EANf3UBIKG3Nb62QLFkFibn+CSdQv2YrqPVCir1daiwwN0r
UKgURUVHfvtLusUl5RLfXuP1IZebFaU9DTMrzTc84+FuGMca2WL9KCp1itmAymHE
9YsiI8oQZOPsHIRO3OF08y1KjUh35n23dw3SV8HNigWbVJro5IM4Jc5GUMLwJxWi
gsjyk7F/pnoEjD5siTVV1TnzfCGBsVlBtorJELy8NoF2ufARR7HW9WVBMKmdfaeB
cglky7ghzI9mgP4esDnp8FxskkjggRSNDo+Wn1Yb/G+s8k5jjdaxuIc43Fe+wlCq
TrzxHJCFCkMpT+2mvWDQA+FZ/ekfZ3mkuAJg708BLxAYu4FKsmCszMLcnKsVLotz
2LaWZZzci1gS4A71UNcsJLHjG1BTa8wlNbUjGXuAXymlJdNR5NR4pemDCxEX/jJx
Wc2DJTdYfKze2ppT3VKc98u1XZ+FP05trfxvX1tpSAYtcX3gOn975g4OT1QwgU7f
EN0hmokhjb6YGGRNBHGPese3pttxw4a4t0oMzoxUzPOBj8yh+5Y/hoBDcno/IOaz
VjWsHwMFkH3QYRMUv1U7UKsxs3XeZlTeRjMDTVqR6ozcoMXGXJsCdZmxAm5yAM2m
YeLNmd99ODXjhxZawObE6tHnRZr09UlFS22tyGqd16UGqn+8CyHctYgaONbKRgDx
uxphzgQYZG1dKl4UZagAS/MfJCMcl1tP1pTa97B3ve+5FwozRQAfrEeKTrCLGc1e
wRWvH1eBEVfYHX7sLimgId2GvVSCxxUcEgqPbw2Za7y1QPtKOkoPnQrxhIVMKdO2
6dDZzwFpFXzqgf7FLg1JeH4lPxEVGTbK40IvtfmI7x7prRZidxI0TvSEH3yTLgvx
zVukgQ0sd6/lh481zDD8wJo1Q9FTWnFX2cQ5mOetgGDdDYGWDW3/vsVdlasNkJ5K
C9j0cqkVqdHdGSnwmiUPq2b3JcCvU3TDYxsboYQX6TXJf4liVKDs14L82g3h59Yo
AyZ+VFA47+Q/7gxN7r1sN5dKP7adygqBCdpFmsccEDG0safvn8UheXv32Osrfauu
QMQ9O/EaB/MQaXuPyl9MmSN2WrBxNECP8PYo+qe3hbpd+u60OBnrU+MNIr2TgMfT
rzhuXryxf3tc+ZmYrsVdQGD0QakfYAZc9bU7363mYLJwAx+3VxySZkbJI3z0wy5S
HJ7385boU3o1IquyT8YHz5Lh9ifx6K3fOoSMBTyHO1DKLKokgbOOI3R/qJkpL7yl
rj5fCCiPm2ZdO2Nsrv5sZl6QCWUkX3Abd185Rj+VKtpT7dAIWGNIThyWxE734Iu9
i08TXj6Xw2SHP140NhkUx1h43hPB5gsg2cKAFsZ5oBGCn2ogjHa1JkdA+CWnBinu
aq89MNB56R5VNWzMqDXt8x5lq2cxmGUAvdSNlBXQ/DUIS/QP5fdF7HtZ5jMYAWq1
oRsGTFIJjLuiqGlMwTFJ8/ZWfqyXem6keq5GJoBQ1NR1FAJY9cErHYM4OL2vUWzg
+/1X7L2fNRcqFctjMmNsenDd8IoZjNo40RAUqeNceHlyXSa10MYURhQ1tyO435Xn
sJhrOAatRvV0Q+doYeNYLLWd3e43L6eYsrho3Cnj9tZepUDaYqYLhJIxHVbTNdDl
H8qNDqT2XtdKQXR62801NLE42E+KfSCZCS6IbHbZc6b2vbFdiXPa2GmgRXGTdxzD
2xLxZL2K2SKwzaFE5xTKQN5ugp8LqsR2ZNR83freOzbolnyvvqg0Ls5wK3RgqN/H
Rg6EKs9b68F06OuQuS7uawAKHjUG+OVh8XFK35uouxS8lQKZMQHTvRj1/OS8E+7d
s5gsY5a0dvSc+Au1e/17pMwiSfoMbRdInk27ezqmFp5Oe8QPBZmCNFOrTpHq/1Wq
4hc4VkSJaZHnCfLXkyP2I2yy9jKpZgGG/iY8ojv09O57u5GSOPaFCEGZy1h90Qth
baiB0UbaVMGiVtvFFbK49Yx8HSwGO455+XcPVrxSleCsaeFsoGVbsJTYE+KNkTCO
4+f/nDC53Lp7OXY7eQ6aROy/BZNO6lV4IcC4vlIPTUdz6isFt5JtZF5X4XlZMkws
oLau4w6Nyzwx/+h+0jX2Q0IB5shO4dSWHKUDLLgqDk4wKABhauFsokoVLvpDJ37t
qTzW0Ce5/jsmUjeN0ra5CvZyyIKw0lu+5mhfWDiwKXH6zCoeCqNO3yAJ0cF/UmEu
8yBOiZo23TPb/f1Zt65y5DrzeLgjyiov820RFuyEYqTeEeOknZrc9NvN/siQJ4Aj
K2f+slZCpksRvOZkyELg9GxIkJS5DBBwcbwInjgDkZ9dMm2jkCerZEAokkuJNIw9
5BxmKgQKf/+OieltUORn+1+ZmXYwUI8AMtik6AYjtPPtIPDHwmkGbhMGa9uNAGPB
3LEl9qLxe25X+ig8qQmRam/6WTXHlNc8NzX9s6sHdEhefzzhsROEVOpMDiUZi9ab
kZg9m6xgwVyoAIAUAZRUZtXlP8FQNr2x0Y/0ks/uz/0XwAuIxwKaN5iSdHD0vkH1
vVFg2KadLt1blV3Pg+mWd0QHXeZDAL7UdG7wDIEimFAlqJLleAwnYRnPNQ0qco5W
3Xu4xF5iMAytg4jxwvaVSnCHPJjOjzfDLFskosrg8kgkzig0POENqOnLRnsfWZz+
xYfCjKT/ZfoKJdKBmQA032o0Z9qdBv5MQInZq3nrNFY8FFpGQi8Ttl1P2muPc2XL
ue4y+w1AxFePIZ92s96EPziN+V3p8vmiSl4Q7VeeEsHraPFuI8rbdziL6i6BJjPI
hOXOaEhfNSO9zplU+sNjoj67UYxAeANa5t/CC/1ENmjJubFTlGbmj+oA9LuWiPp/
36UKwsnYUa3Tc/kpymJ+1U3RUavF5eG86OEma7nOkWNn5DXIZn15utf9YfmYB3CS
pGdP4dkkZg0ne/sw1bI/cWU/QfxSdMdveIAiKkbLGe/sxZaXh9JV3kXiagU3lrUq
O59nU+xuarNZ1Q+HavAFtPSEjohoa+fvdLjXppw8rrTk+d6mtTMcWnXhEXod+N49
GlLwzoBs3oaIPmzBsgOGvtyvQqG5ujq7kaME039xzD3zYb+TIp/LWAyOUDqlX75P
5s4esQYkbnncKRawQ6LoyeiNgdtI5TxWWU7fzP+ti05wtmD+5Rc6q5MOf9g19YI+
UOezUe6Y8W8b4I5+oYAHXKuQIsmaGlDF6gVLjtuEsH/CuPETEOEGqq4S072s/WWi
zbr6m8dWvZd86OrOwRbWnBhOLjC6R+BnGafsJN7iUDANJ18MbeHPC4qIrc09xytm
w43EG3mtfpecpq8McbuJO4Rjn9RdMbuj2juBF7mBmg41RNPq5axpF4RRwCeUYH/9
wicpc+QDOrzOH2JVxr2TsJ2UuO5l5brE6UAgeAxg1EZMJrtQT1dEgyK4dGb8ls0G
14NVy9XtlUoXOgY3DNf2t6/oGZT6GCsDwjhM4cdSrrBMuwhjG9TToiy5Q/H71fcv
w5kYswzAmsO2SwGkn/mFFukvdLTTojllLLfC7oFYuEggXPjjou+LmCirE5zK0Fi4
9YroE3TC4LlpEuQsFKDwU/1ORMYtjyQ4eFQ4cB8JwmuOdFuWBEEN9i4DmJpYGXMG
oXuhHci3NpyVpQdxPhb8ZiKPBAwHlae0X9JkbWuElXoZRjbqtrhjhSGUPPqHJCt5
239+VauLCn9CS9jOF5kC1eNog+8jpAIQpa9XBQI81rVCEFr+zSPRzWxos8L3yev2
TA3AJW3P/jj39E7W2NEWgAMXuPXfcu146DbthAjs3n4XBf+vgRA3veU3ySlFJP4v
cYf8AGRdtuZD+viUQ1rzMHN32K1fZs+Ax4IOUTGWRw6VBnvrZOYpQAtbKwdBoHNq
JSDAFivXaoiFfjQLHP5CZMTrsY19r5QGXzL08qHKk15rUbJUO6lPeOpaZSOUhyHP
dkh5AJBHbSe9rJxi+rh3x75cpuBCRYW/wXcexmZp43lqOaqZHrpDFQ0d3IxqflYb
/amp+RwNYTSPA+U0J/VlWg7emqHY1p23mZguDckYG9TgWfG5errVgYmGolFd2NId
6Y6Sb3Dk8Qh141DiGmxr7nJsVvGMmQM4fJkJp2KeUJjBkbO8y3c5W9OvBjWijT7E
aHbvVnYTMbwq1lRCpPSIQM6UPKFn2dycAIcTf+ew5jL75hyARGZiHom1UX+1LHD0
kclKJqthCL6Ejty08s/JdbbcgmB/ZXQlVpjUX2JCoLo=
--pragma protect end_data_block
--pragma protect digest_block
lqKg2AZ2FnUNI3jwSetW+eygojI=
--pragma protect end_digest_block
--pragma protect end_protected
