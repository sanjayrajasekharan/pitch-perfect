��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki��Ы�T���!Th��y�*��#,��?���Ն.�Fڂ�� %�gd�e�ڤ2��Y��%���>�󉚙wl��b���'���B�����Ө��ԣ���r/�羊`�rc�'�+�/��y�!��Z�Zq�����6�젛�����I�ݖ�6N�k�N�l,2M&fJ��u��)m���4�ѺJۥ9��=I{
v�5pȷ���������v���
1^j�A��z�}��!3�JY�]�l��-��eD�;��T���A��fqV|n_t� 8�L����;�P�a:����������P)��WƯ������m��FQFuo�#?��&��W��'�����7	G��ҀJL��*D��H���o����wz�� ����A��.��|&�Ʋ���|��X1��-�r�_�Gvu��a��p#�y^����ʕ�.�S}K��~���ѹ@Q_0��ht?L�"�9��U��	K�K
�-���.3)�t#�������GM�i�Ϙ�jā�
i�,�����42P�<V�VD�MF�N�j;/�x߄i8�����V�kѲ�ҩ�|��#'W�L����_7�J�Z����Ш��ev�� �+C��������ưqP�֚��6�lG������p=b8�,�q�~⶿B!eԟ�\{����N�M���)@�ʵ�m3�k�J`5�T��5v�~Q��v�qc����������ô[#k��!ʹ��U�k�չ�a"[�6��R��]MSQ��Ëu�f�/�����y�&$A֛wL K���#�f�ܗ@��Λ)�&gٴ���%�-bI�ێ���Q����W� >���	W�?�Puf5�u=�n~���*�R�����w���cF^����æ��4������Q��,� /��)�	e�oR�C���� ��v������.��T+�K��I����X��y�+oW�٫@�ɇ�12�]Ns��?^�$l�6���������h�1��Ꙩ:�Yb�q�P���g���rm8�n����H/y�d�e�!�	�+�Č�T���ʟsy$�hL�u]��S�0���g��W�������o�n(C�9��H��YaڃK�",�r�P��$�P�3��Zp�����-��ܪ�<�9��G��|��>��|V�-����7�;���=�Y��%'w��n#�x�SRJ�~���?�ǳ:�y� �����ڤ�����Tf6I<�/ ���/)�mS��S�C����J�<��5́2�:��q���NezB>�GЄ�xװƂ+�]��m��4烏�Gg��aW��,���-��T.�G�M��#q�qL9��&>d3+'�Sk
Q��C3�D� 3+A��܄�}����1�
_���<P��h�!��2ޢ~��ٟ�a[�,Y���{$����[d�4W5��w[9��M�w͊�����^�����v�t(Ek
��.a#y��JtP%~0G�"����t�V�d��V��HE���b`Μ�oD��)�"`3B�t�¥"9
 ���������3��*�FIW�������b���-�s�m�˃I��[7B���n!U��ӑ��?&�ҥ�k����JpK�l�H���n�Z��n��k\4�0w�X�q��9H��]H��́�]������ݘ9 ��MΔ2����e����5��q�y��$2�q��������{�߽�)oQ<�s���V�#�"��Ai��^�s�[%?_=~���Gz���)�"/�hb��`G$�hJ��ߑv�'-��;Ib���܃<�7��R���L�(1��,�A����*�s�z�K8j�^e�2Υ6��g���"�����23.d߃}sy���S!z>�{CC�{̥Je�\��D��G��jͬ�j)ˍ��q�ܜ��}��?U�o�V�Z �rh�G�����.[�r#X��X�$� �R]�b�.�7�Cw$̶��*W����X%\z�.�3��b���L)2k����bF�3��i�z��G�<�Ւ�zݶE�<��_�ԭ����-j9�t	.��@)��7WE�?��ڶ5�4�$��ϯ���T�������ɥ�3������X��Ѷ')V��nL?9�G�>�� ���8�&��Zc�	���[�˃���C���� ��6P���-�xwW�n�^��J /��Э�ӛC����LNXSG�l(,zI�Sij�}��_����d�����^�������'`J���0�О�i��Ȭ*���!x~�,'��+\>��Ɛ�D�.1V�`����ڵB1ἳʿ�y`��Dn�d���py	���&4�f?>�L�=^ȹh�H��J\8��l���Ѡ�)��H9�-������Z3.H��50[�b|�B݀�
��:'^�I.3��ˡ�-�\_B�(�D�U������xӓ��V�N�pP�7"(�G�8Q9E��u1�v IX[���g��p���3��7�B`$I�)�A�?��o����:ʹ��a��9�Z�>D^���K�J:b�$�B�>E���
����Z)Z���_%� ^S�?L�=mnwdfGQ���7��l�H朠"X��Q!/��\#�4�6�/Zmv�(�(J�h�e��L������_x��/�c|K�G^���ܗ�4�1=����G<�<R�	�i4�)��������D(܋hR�R��z��DKX�&!�͐��Nۍ�	_Yft��%��ݣ��|�G�l��58�*Q^:hV���;��t0K_��pM���aW�lc6���FO!W���mW	�u)�{��c2����T�X��+��MS
�����m��Kp����HE�N��%q�7+ir�>Z�HE�d���� �ޗg���u��`R�%o%���?YzY-� ����Km�dk׎�,��g��C0s�Jf�%u��҉{�_oY\�ǟ���=h��	bh!��d��*��[Z6�A�f=%NǦ��轨ݝ���=�D7C?���Q�g�bsN����$������ȗs�j��i��Y�|�pQs��R�=;顀�ͭf���mnz���֘��~��eR�`�DKRY���&B��G���w-\�BO�3��y��nN��uXqݭ�����3��/�l���K�@=_ƮCA��a�%X�G�Jd�n��D�]�Dmft�Zm�L��b���E�0�˫���_�0��Jo񊳢��"^	�F�h���~"�W��5�B�I��Qr�j��ظ�����·E�[(ɖ������}!��=���d:��N�~�l-�g��*Ds��S>�d�K�/��(]i���¶�����	�9'+�����P@߻�gM�Qv`�� �d\%b0���rm2M4BO`�!:Ỳ-*�����:8'�ΠO]ϭ[��E)�eDy͕Æ�#�Hj}�x������*|�<ێ�5��+���J K+�HV�L�V�ͤ?o�r��I�g�����=��2bjj(S`oG� r�,����E��g�mD�<a�Ƅ�pc�,�ʫ+Ѥ;��U�ߥ0O�l��+����k��@���l8;~�-�<J1��.��\�E-��DwY�?����O8h����=d���B�O!x1ݵ��j�ŵ��v��`"V�#�o�E�:R^.�p{K���|l��t�zJ"�3h)�d��
��-�wR#W��c��^�c�(���;�s �t�T��c�"�yG��p��VhʄG��G��Sʺ0� ׎���^���P1�aP��u��x�d2"nc���Z��E�H��(�����8J�R�I�B�
����Z��u�D�&`�d�hͲ��b�!M�i�72����GE�3d��|�/�3��D�]x���^����/�U���}���d����mCO�ycY2��7>�t������r#�ˮ��-#���)=�/�{��!����^�]4����^��*i&lRt��&�&�B��b����%HἬ��.VlB��u!D���Y��܏�o����H�*�|N?b{����Va�u%�0*�mLuw>�*�0&-Ӭ�P�RTE�H[���^����G�3.#gGl@�7�኷ySŔ��N�%��>4/BVHm����O �4 �ʪNm~ٿ����	@6"����K�q�r�.���!4��cQ�dl��Ƅ��(�<�����6qN��&�;�z�a�[�:8�����;���_l�]��.kk��߬��)���o#�j!*G������#�4��Pw��B�M|�@S�b2H\�Օ�|��$��������g�JβQ���6�;�-���gѧP�U�p����F�M������3��D�Q])��������.��H ���d�غ�k+S..�����jٕ-��^�����uj*:��'H�|�9<fk��s���P������m�]B��+E/��KT���9rR��q�Q�E{��f*C�󢏃���
�4
�X.Q�AiPn�'i�� ���y�8�z#9T��iö
Mr	���c�������6T����#�����Op3�acC�{�@1���O]KW��H�����-fKٷr����
��\q�{���åN��}@���⇎�7;3ƍy奯�?�9���8G�>�	�"9�)W:���#o(�Y�S��ܔ�Xp>"�+Pon��u�O��
��t���ь��N}��uZ7f�-b����z�R��]^�[6�I�a䜌ά���l��aFH;�n�3���ə�y+����݀��i}C��**��G��k�P;W�{��Hsj�l�!�^�N9B8B��b�F��/z'�wx2���{ J�j7ٰ�ɥ��F�u�X�6=S_�&Yn��o5��2E�&Cf���(K
��y��"� ��SƬ�I$�y��i�>k��o�r�3C$豈���ט1cH�:d��Cy�]�Zf �J�¶k��v���;����ḧ́j�b�փ�itM�������ͽ�l�#������qD�nH)��\9�����S�<�Y&���)tȞv.is5����P�M����B!�C.qF2�&�ӱ�3G��L 9��G+j�-@�[b�r�B�E�N��2�d�)���
 ��� 	
�O��Oޑ�O�$��AG.7��-�õ��������)[�JT�|��u����V��t�2���E�|�öB�	��*j�o�q2;�$pe3�j�*��#m	��kT��t�X];��%^���d ����4�����m��_�\OE�Ѷ������Q��j�):��!3�O����ϊ�W+Y��͸�Σ��*ZU.�;Qj�3�����A�Oq,��*d
5i��[^(P������uՖZ�3К����4�ϧ~�Z��b�֖Þ�m%+K�>	���Y�,���x����{{�|!Xe�`�zѲC$�걔�����E��NX���8-�}�MĦi�b�n����rMamw�23���+��y��Ñ@Ha��A	LR��z�М��{�KX��?.źi�~��+��"�D$�I�O�ϫ���ٕ��2�dŪ:N%4�x]3j���4���m��ɐ�G>Èowyt@��Bvx� R������VcC9��@ъ|�/�+��C2FF���`c��.������1�A��rx�g/$�h6Ͷtb��8%��}u"� �:l�-FnJ��R�5��;*t��ӵ�u�Qr�\:�S�̢�6��YT���ީ�#�>��pmǆ��L2�rGŌwK� |��b�u��;T�p�e�fQ:п
9��{Y����ql���znw��AA�q)Dy������gmWaZ��ʺ�c|�,�9���`[��!����0�� �1Q����m��GsJg?09&�q�� z�@���D��uA�U-� �6�Yf���nZ�Ѹ�]��Q�� R=�#J�mD�ꝰ`�C�0�O�{fn�e@I�{f��^���V���X�v�����*����u�zA��ЦF<�8c���Q��m8�d�g|���[kG���M��D�Ģȁ2��Lu��
Q#���8�\d�S �L΃9�g	��dء��Б'%��zљ�x�~F�m�(=B��3���x�E�9�(V���lP@L�A���nh>_�	�����C�@WS�� �8��aU�j�;}�S^+E[@�!\����+��Y_Fh�3�K|���ڡ�JI��)���F~+%���P#-�y�?
ӛK�c��I�F,ѥ��io�XWy���6p����c���/3�QJ'{9�dj��q$�e|����$;�޹{_�C���#G��D�lT� ���L�n{|�k�o�:�&q_��aF&fN4�P�h������b,E�>pi�~ ����1W2!] ��^��%���^��#Y���īU��vD��|��$�d��N��'淿��������e&&�V{Zh��G��տj�(f����\��\�2K�I��*ay�v�Kǒǁ;3ߦ��o����Iꐚ���'��O��\�Y���Rwq�	È���jY4u��i���.y2B�� ����	�`F��s_:l1Ȓ3c��n��6�BS�5��:`UD����ZP��<*�x0���݈:J����"�4�Ɗ�z�51�gF��8h&���gw/�2c��}`����@o�.2;�F0�K��HD�֛��L�+$�D�~���<�3�k>Zˋ���	KG d�+���:���q	{����'h�~�s��fU��,.2w�:����� ���X[��j03
'C�}�W����	w�S�HI]�������s;L1��������V)b쯚i�v(\�Ҷ�&S����8�v0A.䱾LwzYU��@��j���F���}�kpw�������� �*�M�{���a泀���X�OaҜ�(zs����bnڼ����I���گ����������Dwp����V��,(d2w��G�x��gS�NRS�l�c�N�ݰ�w@�h.�v���2�� �o�7u�R,�7AG�rH�O��E-F�&gq(E�1O�$5�R�tFQR����uj��n�	��="�M۱# [�;�BS�A*��"�mc�|6k�����u���_#D�*��6�E��<%�(>�~�da�؅��$��j����,��u�(�7�o�I#.�:�s�KI�靽H��:�6�����H|��q�`�*��\�l+ӷ� �xtkWwq��2����k^�N@1s�/�= 85�H�=���wYv��r���N�\��Oa�av@�S�'0E�D'�F0G��d�A�������Ȃ5�o��Z+��'���w�J��@��t��If,D6	�_��`�He�J��f�~e I2ț���4�Yo�D#(� l���Z�o)a������7�*%��<�D�&Ӕ�Z�^�V��~�������Nh���	���m�z��6M����_�ww��?���"�,�"��
�����f�3��X[3�$]"	~0��@��xf��?p5JxT�?�Q�OW�|�"��K���B�n�����J-�^}�`$b\�`H���]��@��V�OS� $�A�D'{�
�$�7_܁?K�t� gɏ�M:Mm�\D��i����J���͓���$�;�B�$K���\C�*m�QTɰ�z��%=ŉ����&����+����-`���U>`�xL�'a���-�adg��J7_� b��jǆ�:31~�2�F�]�˼�g�/Y���f�f�4�K�,L=�a!s�Ԡmp��3mAu����VS7����)������Iu�9�/lhf<k"-��>gp6�<�G]	�c!-c)�M�qt��Dc�����f(򬈺����jl}|�ux���G"Y-��p�ׄ6;-k�z|a�(��M�ï�$Tœ;�h���	���A�'����hx<;��W��Q�ȅ�˨goXC�X�pw����4��Z�5���q��iDy5Vv���f��CZwv�$o���eS� )OF�c�)]����Ph��ڑ[b%�I S
]�믙���vL9����8w/�{�>��u��� ��Ѣ^�E��/m���}0��G�+#D��Kԉ(�á;�VCZ��[k�D��;�U�.�x�mI�kW�7�F�ʥ���֔gb�*����n��r�O�L����pt�9��1S��+3�UΏ��0ǽ'p�n)4���Z(W��-\�c��uMn~@�����Q4�(��K��7��0��
�l�m'�˿Ψ��{����(ԉ�C�m��a�_&��ԟ	��&0�ɕz�hTaa�ry��jo�~у&F�����,6�݅����_k6������	�iJw[��B,B$Ɏ5�)#U�[��BP9g�x��gR0�K�8?���Y��'�%bL��&Y���{������%��8-/qb�9s�#$E.�_�3�H�Y�}fp@.�����E,�W&��Ep�h�I�SL[3��M(⪑��6-m�_%�$˕���/b�"��������\�.2W��h=ﱍp�f0\}>�͛d:~ÓH��˱�c�!X����> Q�\�'��p|aq�-�$ƲA��4��]Ƿ�Ѧ|f��!K=JLԊ�oO[(�*��E%l���E>�y~��M6���1 �W ����:�&��.�K�P��9q�v'��fZ��b��ퟮ�l��O���g)�Ō�tu�^��Q;�N=��ݜ�Ot�6{�u�%�G�q�K��`�Z���ox�S���(�D����Ю��x�A���E���u�
�r�!�L�=I��
����[���1�V��H��#<�g=3k�)(C�)z1s0"�&�%����Q�{3�Oo�
���� ���D���W5�z�jVq�;�����#����f��b��A�-�}Ɯ��Uq��5s�?l�=3�b���ga��I��ݧ�ٷZ��l��뼖���)��I�XV�`�vsO��������D8���-���z�B�sط�*l�,��]�c�
���8��+���ifXjF/Vޓ*m�*Zr'��I葢��2�<�?P��n<L��WR!�*Fq'�����z<U>���9�0���{����!+��݌��9����LG�2Za�]���4�Z1tr8Y��J�#��0���U~����a0W�#���]���=���i�FӒoC>�؉��|/[}��<�ښ�z"�q��9 �̉�pB)t�bܥ�ḗ`�sVR�,���4�g5M�[��Pl��ҶUtD�7̇yF������E�}����
I}YN�U�D��i��JzMݩ?~��7=�+�T�P��ne��|��?�
gUXB�>�'�N�YØ�2�Pn�Ee�0ѿ��mh��#� t��ޞ�� axQ�R�s�t�j^����<�Y8�}H[2T[�IYF!���1��������}�ƌ����1�[c��M��f"��j#޽amyoo�I�<u����h�d'�˒�;��k��x�����)rZ����U�];���p�� myv�/dլ���J��0&-g�U�J��DR�T\f���Pf�r��sH�ʖ�����ᵈ]�	�1k��dB�8�$-YB (�LnT�����-*�uQ0M����Q:��=�mS��sn����c�b-��9.��ڍ�V<�C�@Q9���F�u���_鯧}ZT���YGW��������.�y�'(	�3~�Ŷ#�By�ED�{"@K�J�^~����/
��T�J�Q��f1!���I��<�Z�T�)���[epȈ_� ��!�2��7�(���O���� ����?�P�b�<������+����[K�6��rǕJf�B�T�en��v[�1�fQ�67��:�?�S���!,��^��<%�Ƀ��@���廇kDUvvz�i6�4Ҹ4w~��X��-��ͯ�	K��t�=���*�C��L�)�Ɵ�ߢM1�Px��퍴ۜMڭ�E���q��]��`T0.��P?�d��ӯ�S�ڤ���:/D�-,�l9J���]I��۹��b��ésʨ�j�!�����2�&I�����H�JS���.��s�,TU��D��|a�	��=� ��JI�������7E$K�)I'e�W�Tҥ�l�M�ۣz�\�iCt �BB�v]=(�Ё9h��$C�K���|���X��x��)�&� V�ci�]�z�V1��ӏ��P���P��ܒ�~��4Y<c�Ł5��̋X��}�䈫զPZ>���Q�$��C����nj��F�5E��=����>N��eT|-=仏�|%��x`�c	�lE��K�!/E��:|(?@���?N��\b�?�K\S~`+�I��ƿ�7I��{F.��{vWH/�ag[{����D>�Y0�_e�ԣ���(e�q�S;וK��X�DCq�0��"o!�5L�J�J��g0m�ّo�Q5�cP�@��šK+�km�G�O�@�����e�|����al�Xy�ξ�cW��<ǧv���XIl1���b�5�u�z{fkQÞ)8�$�զ�u�|n	w�W&J��cjȧ�J�F'���ѩ��?�g"`��R����L�I1c��Ck�:o��'�e(y�E��ԢbT�C��C��ɸ��4*�=m�1�l��� ߜ���M��4H6���l�ǆjh���ow����6�ZP�/�K^~��D��tz��O��\4��L�1�#�s�9I���U5��P�8�ٰ3o*�C�mhԧ*ˍ�����:��3]���h��u���ğ�"`h����	����B1
3��P���P�aWN���C�*mK�]���V��k9�W�R���ۦ�&2���R���,,���hl֮��K�H�ɋ�]<\�h�:��U��ρ�Vr��-�?�O&.�L�� �2鶅�c_��AS�9�^%L<-�j�<6���%�G���ك)b�2d7��>b�l��!LЯ�H��AZ�������){�C���f�*��浦�OQM����s�{��T�S��~['�,�Y������+�)tW�8�:He�d�D8~�������,F�ZX�����B?<�$�P4�wtC
؜�,�dޏ�q���?"Éo(H����N�M;x�ˉ07^򒩡&�.��0�p@�s�D���hj�ԽއT�^��Av�{�(���Z�$��&��8x������d��h��LQ�BڟϷD/�E�=/�b��:��>ө��������S����{OUڤ�'Y�+��c(���!6�����!&:�zj�py�����$������H��k��Y�\{=�_�*���s;���'�م�u/����*����C~G_
��PA��vQzh�)�6xY�_��[EZh.��Y�3����n�k7T���� uo��^��Y.3�ݕ�"���~����˗{��!p({̰ ��s��n0�FJ��LR`�z�Z�v�9b�1��g	A\_�?�4��k�	\Y�ԪR�"���0�@�@u+����ہ�-�pX��49�O��B�	mQ��<ĲC������sDsڠ�wh.���I�C]f�ʳ��_6��fP\ �$1�G�vF��faNHM.:�g5�WQb���4��Z��9Z�Bn>���+����g|�~�B'�j�4�� T���I�����!��s�H��b�O�5������Sh�4���L��zz"394��q+�|����.<��4�6:��"����Z�ZM��y�Sq����V3>62<���0X�k����+������,��*�˹i�z�,D;X��A��^:��������+�0�?����z^ڬ�e$+����`�S��z 3��}����sK1�����Q���_�CѣXޥ��@7�|�+_Ɂ���h���m���'��d<�/����gl����y,W1n�iڞ*��µ���i&:3�� �7Ԧrm���ɤd%�gP�XV�V��ް/�v���$P�K��A�c@k��:���옆��WMnc�v �9\�УE�}��<w�q���Mо8��ETbȎ��7G��T���q&�,�ANߎ���o*jB�V���d��'�'1��{�'��^<U���;$�������6������.��ŝ�a=����rh�s	ڒ����da�?�n6��;�}�	�~�(��:$K��9Ѩ�D��kD"cg�V�e�b�h�Q<��o���%��Wt�n���4�p��ƜC�I��Reه��Ѽ�k���Wx�|�+z#la j֝��x���^�0��VVn�O��ؑ���/�	O�ż_�Ce�τ����rOɔ��-����aO�	6A��0"��7��۟r�6W���MI�]��`{|���� �L����g�y5���h�����z�`�H�m�kv�}#Ἤ��R"�1ƕYw��R��&̕� +�b�fVP�7\��	
�� ��t�40����0�qvz�nE+T�s>������<o����,��vNv�+Cx���azWT@��)�b�W�٪6pR���e8�ܗ����@%���b�N��%��T�{�������d$��ܼ�)��7!��҂ԾMc9�r �3t���>4�S����`��*��7����˯L��z�C�3� ��祵�~�k;)� ��h�/"b�T �|et�v	��c�I�%e�ӻUs:#	>���q�U�}bSL��2|5ݫ��RT�E_�����b!��i�t��7È�����5��,�������J�gO�=t�:��L�nDa��
��ֈ��SAW,Q�;2���"Dg�J�C�5���W8���Ӈf�R�lf:������pR����j���a�T�ɪ\R�X
�멊��#�S��^��4Z�JFE~BD�e/-�gaUe;dff������pShd#����\�#,�2�U%6"ѿ;i�3�=�-c��!�,��tqC+���k�ӠM6ZhC��jU��\�"����$�C�+|�Q�X.d��U���m�ڊ��D�RcG���
c�Ơ����eq�WM�U8(2&���$"�4g�UW���h�%�$*a�� �g��E��iA����6Rp��`�s��wJq�1B��n��ِؐz�\D��G��4`� GY��5� �g�9أ#�c�ѿ�Jz��M�vXX�����_�|���R�'��Z���}�����q��#���^~C����k�F%視���2%I�tܳ�oѤ�bY�UDʾFG�(�%x���������86�÷6��蒐rKpz�e֜�-��]��_�
G� �v-�;�.�.�MUڹ.>µpi����
P�>�ZC�S��x�F�~� SwhV��ȑE}{�����
n^��
-Ιc�+zO\��M�/�m�������� �f���rF�Y)>����0���G�:=`g�&&?^tȍ�Ih�ĆQ�8Y:�	�x1 ���F(��ƭ4�qW���uA�`�����8}�# q��5J���Јh)f��ڍ�V��Љ_����q�Q�0��p���s��v��2�+��졵H_�f9�+�)�R%������v��̂f�]oj �f1Y����nH��u���Pt��K��8����LݦܜS�V:x���P�d,�hs���/T��SgU��_>�5���=��އ?�X�u=��1�����ԟ0]��;f��m�D�^ݍ���:Th&|s�;�A.BU���+�^r>v�.�̧���M\��^�$zH��}�Z��O��Va��k�:+{9�xǭ�3½�I&�|��K�KQPЬ��as�wG�j%��yx��S�i��A|��3�ݯ �=L�=
���VpP#�UzU(]s,M;>�'��t��>�Sc�'`�bA�'��H7���=�\��7Z�y]��#�BN�����u4l1�UPn�8ӛ�H�6gi;���`&I�b���Bv�k4���H3D�9`'���Vwׇ�y>��A��4?��A�c���KHr��1P<BrUQFT�����J�9>�ۊ�g�Z�%�[E���Kb��1C�T�I��)M-�+��=���n+*���k�@Gm��PՇYY�3�Kb�3�>��� ��h��)�N��v�����.���=�����#�D��(��s��F���\�a�G8�[n�U���}��͖�OĠeU$W�������(�Px�k�n�r���`�6�X��-�Z�3��_b�!M�OV, P��+gG���-�����aR�u,�5'J)?�۶,r���Ө��VG�çM�0�vG:��s�5�{�;$�6��1
˲fvP yBUCM#̘�v�庬�L����-ʄ��iP����rŠ,$��V�L�
����MY^�0E�c�m��<;����v�T����)��d#~%��KP�c�@�v.��y���k�moI�Һg�ni��0�����dO7�ėP�&I�>lm�O+�����M�U��a�z�P�s򓨏�L�ih��X��pb'�B>��Tf#ˁ�$�~��$�o�H�2�0���p=eml	�	;��R��}�d�k�[3}��8����!�T�\���jQ��*�]�*���d�x�;�/�L�f5��]<�o	v>ȹ^M��Bg��Y��r��Z��]��Y��h�69f8k�>�΋��n�Z��q1� �lI/ v�����dzt��m��Sh�6�,��,	�L��S}��2��=ò"�%��g�XHt����M/\O�	�*<x�(��(��w��ܑ��2�PcUM�y1l�mܓ�܎�\IMh���1��Z��� ��mR�9�S6dز%��CYۈ��׈*�3ܜ1�B��5�S�
�骦����^	K<�춃h[eK�Ӛ����ރ6��AWfnQ�J�d��A�i���K�J����Y���ʱ2�a�\�
2�[���o�2��;S�H'&9����l�v��o��/q����)��i����ٗha~�+t�D���V�#��W�������S*��G�,ik,������䰙>���V�V ymݻ��˝�lb	�8_��h�+Ӕ��� F�$nȞ��R%��t���>$ЍY@�C"�*�3��-A�cSS()DB���∝�&	�4��KN]��t�q�L��@iǉ�N9��-jn�>*�<�ʨq
��j�x� v���*�T[N�wi�'P1`�rB�`��wX���).���F��ơJu !��#��6����۶#P:��S�3v�
km�� E���7�P�?$�x��֏8����`T�=Gl�I��VC%]9�I�4���sY�k�j�Q'b���o�7t}�5�E���q����P��uL8%Vг#��T�����VF��'Mn�eK5:�K>�j�
���f�����i1�����4
�v�le�u�����D�H9c�����MV��Yq2ì�ĭ�m�_(M��)��H P����8Ǜ!���dX,��7m
��)���D�6{�h��-���^�n�ג%C����0���FMx�B&���'&�ڨ�Җ�"$<@�� tB˸�I�aK��В;&TW�����M8�DԸ�*bH,�c0ݍ ��"Co�ob������U�ݳ C�Xn�<��.o��a��x���є�u]T�I�=%�������[U��'X�E��l=X��k��f����D�?�R9�$ؗ|@$���'�)��@�fbǉ��g{����*h��o}s���^E0��-�;�Tv�ʨ�v`OC|��5�C��(�U����Y��94��7�M�V��v1�\%��{�mx���=�V]��2	��"E4Ԧ��"�*�/���y�O���hfB�g�u�E�ʦ��`��Dn�����k��i@q���0���'��pp�_�牏`/����.Ҹ$�Ef��N����W�)pj�Ŋ��)�x����~uZ��z�2;5�h� 7@�H�[Q�>�V�c6O��v��h�r��8��c���W١j�+Ҕ���h����:�e�Z�W3N��ϙ�i{f��dd��	��-M����a���4��P����X\����O�C���A��
�_;*P�Ŵ�����j���Cn�+hJ�m��-�u��I��eS�Zi:�
�*�����5�}���F�r�!�c����Z�t�=YF=��h�����PG���\�	�g|�������������g ��F�΋���&��䒿?tgU1J�����*��6�=�-]-6��r+�ܣ��7��r8 ��'o�� �-�G"o�$�ܬ�CLl%�)�+�1�k�!���&2��M�ȏS,,"_�,@-��w<+�F����(�EG@[���n��7��5(��/�0u`FrZ����l�b���O����Q�^���=�KU�̎ '�!��$+�W��� ���?�$�����f=F��3Qw��l��4� �"���Ry��%�9�Ɠ������O-_Cк�OR��}�;��[-�eлp'�;�WmH0����?�VYJ�y@*H�o<��NW��6�:wsFE9�n��om8�蕭�b��U��J�����{���C)w�@Z��R0a��߹���=Rրk3d���͎!2��2��
&��A�~��5�C�����k�5"3�8ch/��I~���)&����C��E��f��	�xX��M�+�t7ʐ��p��}���氬�4��}��;8�����Z_�<�t�Z#ᅁU��k�\9��=1Ţ,s������IY���,��ԛS�DyGl@-8B	z	�~[�uJY�ALǆ:���!Q��}cO�o[�g1n�Rb��L���g�5�9�ݣ,��D���E��6�;WL`��C����*݆�9j�{nZ���%��D��z�n�
..��)�	6�$^T����Jq�a5)�z�&��I}0�|�\����~v��tΖ��W��|�Y]`��L�oR���3�ᙸ��{�jy��u��`އ�u{����>�,/8Y�9X�*k����
O�q|t��f�Ǎ�2��^�y*�z��s�DP������Z8&2�z�a�R�����(=�//�5�N���p9ۅs~�}i���]`"]��]J����g�V��W� :��Y��zC�_�O��Ś�D`�~Ҥ�q��u������D��Ũ�e�.�݉]3&�}�9V|J�����hBK�A9����x{o�)��ml�����y��iI��?�ͺ�(#X��s��,%���!��p�T��
�[�:%�+Ӵ��--|�nTښP>��T�(P쵸���O���uN6��p�����c*i��	f����o��q��V.�	�'�}�Q�e	<�J���絿��v��m�{� p�����ׄXRm�t�7A~�玓Q5�#�da.�\l���Ŋ����ck���u
�w���_Y�G����I=��e��MB�
[��[.Y}��%�?�9.q�ג�<zL�x�S���sus&:݉�!�Xk�_'�dBW�\6�Ȗl�,������'�W��	�(�d�b�X⪰����t��:ڽ]��0�)X����fC�f���ଡ଼�ߊ�֮��췍7������~�2�2�-�F������,W;V����/��xs���w�Z^�E�K���Y�����K�u�f�)	}*pX�C�#Q��r�y~�^��> _�`�V/�}^�/M��!5rJP1��j���'�����t*������x�֕<��	�}z�_��jG{�\��������O�pk���$�]ˠ� 7�N�x�c�v;�cP�	T�z%x����i��t`e��>L͌ up?Ԍ�T���KZm�<]ؔջ���`�$�u�s�:�ޮp�L�[V���,���ЅI�A��3�d�7|�j�M���}�7���b>��Z��V��c� ��a�u��] ��������@ �L�!��G0���.,�k�;���H���W<�� �M����`��K>!�Cv�f5<�a�Y��,�O#a�,�)�}��QƆ��J�8�dS�D�8�u�k�mۺ�q���bb��6v��Q�iS�X�m��$o�Xw���$���^�t�GxڮzF/����dڋ�=p�p��,_��-��:���]���eq,[ ���v�R��
GAxLv IhO�(��b}�[LNb,��ۦd����$$Cو0��v��"����ץ:���/��`���yh�[�{�}<��{5 ���U�	�'�Oq�^�/kbh�b�!�}��h3�:	����{�$~ʢ��n���8�����yK��$���mn92�m {��GZ�?k��9�Ōs� ��I|��&��V"-޼m��{�0$tw
�Ëȼt�c����^�ډ��78A���N �Br�^E�d��b��r��$:s�W�ƺ�h���6ª.�qw$	�;;���\����;b�g^Ԅ����j�����>�E�9U�S�(�^^�V�q��ǌ�w��߷p�9�A�#��v���X�E�_�@���c��}� b~D�N* W���3���_���\\���8 ��i�����Z�'����jĦ�(X����<A7�Rl�����?��wW����u�Y�''6�h2�~��8@J��+����'��VԵA�����6�+Ӝ6��r��V��WB8庡�1���3¯@�]�|����=+�|���ۻ5�є�6�>,=�񆛨�p>5�DWJ�O]����%I�c�6lWc�^�S�n����g�k~YX�����F�r���D��K�q��ӣi���?���E(&:>I0���q��' C�?�b�ש�©i������R�}B��I�T�T��<=D�m���p�e�w-�g�Od�L�)���yL�3?�l!���ܾ< �Z6�)�T�{z�{�Lz;50����ڤM�b:3YA������g�	��Uς����m�E�����҂�����i5��k�L������VLg��[�®S.~UH[Ś���'�7G����6�;����*۪g+�sG ���|*m�����C�E(����Ey�����\H\����2��@SӘ"�\��a����;;�Ik��&���<���V����ݶ!m��hE�1)�� �?+�}=�� ���"7�+VYtOQ���JI`����l;U��<6$f��D��0��OK2ʟ�_p�>�lw��E��v�>�>V�B��U�G�KHXA�K�`�`�-v�F'����ڸ�,�n�`�����=�*�CD���+As��[5�$9k4�ݢ�wi���q��y��;k�Wp)c��|�� &g�D�ЇqUP��7|6�=�e	5{O�&�aʲ���V1q����G���"i��% �-Z	J2[
@q�Wɢ'���q�eCف?vF#�b�R�m"���rZ�-��d(@�O�ll�.�F@�	��{�m����`9�y)YQn3��ė�1�d�n��A�)�]�ؾ�5�T"�xj�oYM��L!2b����R��"��M�Z����O|�X��'������H����S���_aY�Xӗ/�;�}mFA��U���{ٺ����	ׁ>��,s�!��_�DB�X*~��_��#����~�Q6��dU&{B�Y��hI1b��H�K���@��q�o�Z5Ύ&;�"����DT�20��:�-cC���-���zP�=�l8��o�@�������)���E�|��J<�(��}�mX�^j����4�ė�AS�Nd��Cʬ8R��e`�"�jL����&;3o
�s�D~��;�`6 Q�:��I�w���@(�j����i����:� �7�=�Z�ʮ+��M ��b��~���?���?P$g3�0�[`<F��!QM�<�l-eYU���0`��bo����he �«��J�KI'0B|� �,g�G���Һ�Ju���;B�y�:�@���t�U��?��8z�_٥�+��1�A��~�:�?&���9 �Yo���29Nӫ�C ;_�_�DWl�� lQ�L^����� ܏�1��=��DX3�c��Z�xC�`"��m4.��`+i�Mi��ѥ¸Bٔ2�{��A�$��^��(fא7J���5���&�� ��gͱC��+m]X��>~|�f�c��}���A��Q8��T���Dj2��̺,�8j+���L�/_4Rv2O�`���U��O��!e[[T��(iS,D"����"��V�$>;��ǣ��Hbϰ��c�|*�L����0� �L�g&���X�q�_E+�^^O���|Vb
���j�:��wi�{밓� �Zw\Ibo�gs����7ےz�I���Æ#aw�����~&�l����-3��'���V���=z��Ĵ�Yj��\*E�Ȯ(�e�6+�+��=���Esź�9'u����H$�d_C3.��;W	R�;�;~�P�t�+h�\e}ǰ��jq��i��PB����t������a��y8����1}����\��N�K�k^��49����#��q��?�����W{օ�b�/i����Em����b���Jƭ$(�9�ă�-�CI���x)$3�C0�lG+���H� %1cLa�o����_��Yh�r>7�	FJ���
x[mn:�ROXx^��@!Y3�9p{g�L�1���wg��d)�������y��1	�Ʋ>�I��`v#��%���:�����#T/� ���V<[��n�����2a=����^�-�)��N��XE!ӗ���*�����_!̕Aa<X�b���a�����������B�]2OL�;�ڧ�u�������6���d�.G-ՕL "�aF��#QtSR��`�4E0�&�,�Fj��^�&��c�����#f� �{m<�ŝ@,�(e85ԩ*�""c�,e෣
���ܱw�6��������M���f\��ۊ��E�4�T{�E��1 �9�V��Q��~�m۵3O�.:',�	₈�*����L�PQ�3�u�w��_K�GM 7�͔Z�Ҩ���������1��T�"Etx��\0f!Ƹl�	�7��/zt+����s O���?J�hfmS��H����o_�%�e	̑����tjCH#{�������|S���Q0�~2O]l�x,BNs���=*��jߔ4�=��A�Pl����>��Ys�f��I`(���,�,�s�\��| �!��o̳�0����1m���ȵ��s�S��_ L�T�G�-���Ѷ�_?.=�9��-t�d 2�1y�~A��u�{1���n�o����hܤ�T��MaT���G�޻�i�2���I�.Ka�ף�������í@'�פ�<ϕ�Q5�� Ϳ6�,$��*����u�7mx�Žo4��(|���i��>��O>�<�#a]�;X`���.����2��Y��`�2��1	+ȃ�Bg�0�齏�t�9l呧�G�+
�4( GPk0@IJ�c�j�x=��謸��#���
P���t��g֓��3+�T�Q!�A��U�H�5��>�d6ݿ�ʕz�L�څ�@�bO&7���������̗��o����jߕڹ}y�'O�.k ]�0���sVf�[�n-B���1�p��c���E&��C7A���P�o�!h4`�ٳ����J�����g8�a�dQ$}�=��<����:��,�� H
�i�ғ����d�㛥)��p2�7��6�O��I�2�o���f��B^J
ܦO�b����Pr�N-i�O�8*�&RZ��+;��[ʢ"!+NZ>���J�=;��S�e�͞'��)�L�����i�& ����N��z"o�	#�%~�"�wC� ��x^�T��"�/�ޞ����*ƥrVd��$�u�fa�W�k�L���b�3xc��^�� z"�@s�J�3%v���_��I]�,Uq�Nc��c�x�4���KP�(�z7���+����xej��6h������.���j{���ޙCW<�jR�����Y�����(���9���A���&��T�n�Qs�B=�����}boTl�"��|,q"%C�{����>���A"���K3�w���:dRR��']���x
z(bA�P�~Z0R�Y^�r��fhW �u���1
j��V����nO�nP�b���p�-PI+1;�U�ƞs7܄9K�H�����?I��8����M���GHk���/��?�:	�]n�F�{
�GNSA�`�u�\�e�(7oq(<�B^�YI�\�ށW����Hv��?|1�Z(�ܴ�Ź6� G�{��
���������	=��n �o~�$��r�Ʒ)S!_���^4�ia�+�����[�'����3��AF\C�P��ni��H3�����z�Ri��~ H������
!�+�7X���V����������|�$jO�� ��\��vx� �3>������ ��L:�����W�6��DR�{�p�${��Vbe�`��G�<���#zy�{�ttԨͩ��,���'lo�j�)W��{���]Aϸb)_���7RL�]���;e�?�����}$C���[�?qY?�{��s�7�.�Mq%�<��*��U�~��J�˘���{v���f<ڳ��CZ�c�L�4���km9�*ŤX�K
�vE�q�l@~h�ཱུ�G
E�.����L�C,4���*&��k�R�q���s�-Sl�ws�53/#~4H%�������CC|�';R�`�d���̈����=��Ņ<d�;]�ɘ���x�HTY�EgT�A9;�q�~��3S���*'����[����_G�J��%'��8ō�7J-&F�/�͙��^�Ű���0y�0%�^��m�5��Ov*���CO%�ɷ������1/���>ڛ�`�O��;�t��7f%�-Ś�{1-�o��y��_���mr}�:�s�u�HR}���.l��N���E�qO��#J�������z��s7��P���4�{�=
�y�����/��O{iq�c����A�|�����=��2�M���Ŗ�C�������dgR%.�/�S[��;��:Fk��Vo��*a�6�0������'�n�
,����-F�<���,�,���gK�Atk��TfM75�c�@�J���-�LS����t�L���Kƙ�3��Q ��vFS��q��#�)2��-]�b�
�>�D��ԡ^���"��Odm�S�=��G���~�k�S��6�I���>j���#>��y-n�u(�l��\�Z*y}/��&	�2��I�T��������H?M%# N�	�8�'��u1���}C��,�n�'BBnO��T�-��IS�*�&qzYVM}�Fò� ���{bc����{��e�F����:��d
�);}���mױ��o��~J����7tS��f���I<�>�ک�Rl���y��j�{�f�B\�~�F�2�]��!��0�+�(:��7t<o��|&����٤r���Z0��װr������~�m��c�=V9τ������-T�`vV��3O�-m�ږ�@�N���ka<4�>����"-��K�S۽.�3z�s�J�#�ȍ����z�!{���z�w�:�%8�k!�S1Eƨ����FאH�x����Q�1��i��k
^]N����mh�ǿ����4�ܬ���ʷű�{�� e�>�C�}$��ȩF���=!ӻwe�^���6�Km3�j������?�2����VJ�ï��b�QڇA6� �z���X�Ikeepʻ�_ڶ�^�x毒��`�'�x��%��D��/(J�����ϱ���Js���fb���,?�XUSܲ���Ӓzn����Y��!q�|u/���A�����.��B��P��^�����^)Z�g�����?�\�B�|#���1&}�c�a�M��o�?�P"?
�4z���mgk'Nt�ZciZ��g���]
�.jΓ��Mh[!B4�Ca�~B[?�@$����wȋp�O��L�怐�t�$5��#$�\7_"D̵�8 �B'OS��-1h�����V �j{b��V	w�\�y�Z4��Hˉ��i�7_��ҳֺ1����f�O"�)���=RMu�������&<���u��'4`8��"���Z�.$��Z`�Y��z��	Ł���u����V��7�2f-6:�U0���ʱ�:4�E�W��'��@<Խ ے&#��P� צM	�����*���6�l�m��������U_O�ᤶu�%��-n��B��s
L0��tF+�t� t�-{��y<��2��.Q�a|J伤$��8�Nj��x��*��i���9-%�a����˜"՚_@eҖB��"�U'�����s\��c�dH�x�$b�М!�@���pgK�%��f%ø=���;i�L�o�V+z��ѯ�s����=o��E�.�w��#�^_�F�5�����X�j6�����	9��q���%GܩlF���o�z���%�٘�o� ?y��
!�� �Vn�TTBs�a��ݧ�~���e,)��dujM�����]�;/�I�Y�K�2jW��OIg�1�eU�|��ʩ$.����~����wl��n�p�*1�T�ˁ,^��w/`�)�*=��I��)�_u�k�(�]4Q(�I�@S9�9	������Q2��Op�L$�6���2ŷ�nn
��q3�U�qE���R��y���{F�����>�w��~牦c`���G�*9�(����ZL�x)v1��J7;���%��c5������>��{�B��A�/�i�+���U�(!��P��Y�}=ՈjL��n�E�Ec���0��r	�s�����.��-�B����@�]U�}��V�Mt:z6����X��J�������?�л<��ś�?nA���qxP/��ϕ���i$1�UF@���6�Z�~b�+bP�ڽ��^ۻק��<�T��ѹq�j���-�!,*-dQ|M�jq
 c^<�������H���rb�L8���ʝ�ϻ?�݆V'���&tp�a�N:�h��=�4j7���̏[ .�÷r�Kt�I����c,Ȍ����0_u�Z�v���/��K#�a�MOB����So�{��Y/�M���3�{K]݆!�K�S��-p�/.$i$���oLH)e1y�nW'3�=m�2-�8΄�k-�E/��*V�(J�t$���啖�5ҝ��+�#T�	+�JߞL��ɲI�HiV8��@,��!���c~�>���ldXʂ�����$����ʴ6�q-��p��V�Z�4�_��O�^�!���Я��T�H:�Wxfx7���%��?8�T)��q��&}ǖ2C`�����cu��]�C'���_��M�..����a %�UV_pZF�j;�HcT�ӓn��>^�f����"Z,���J���n͹���j��9Z���|ź`e�̫I�Y)�vfڀ.2�7��A+D3� hgW8���ٮ��4-,�s�+�5��H����Ý%���?FU��$M5Uii-N�Կ�1�2���c�z0� �j�ށ0C�D��%��@'�vH�'j����u%xK��-�cy����^숑L�;�_#�a.˗�I�1s�YH5�f���݆�d(F]�R~��GYi�N<�VKܓ�&�Aiqwa��a�.%�k�ny�-���2����3n�&%yb���M�R�f�^���o��S0�#��!.������%����d�������{�e0+��3�Gn�a���pOQ��	�"�)���U����a�c�",r03�H%�[����M�c[��&5�)���LX��i�ʪ��JGQ�6��|���~8
F��3�!�������WYo>�kC'��l�K��'��M�nV�7}K�8n��fm�<s�|ؾ�e;�i�h�%;z�X 4�vr�!����WA��� �����#my�E��|3c���r��:��V�ԅ+w�S�������]:-/������ɞЪ�����:��>QԜq��3x5g�"�(�ƨ�ԟp��bz��R8y�����'���EV�~�����@ �м��q��~��+\�OSڳ�H��K���\�pvwғ�nIY�p���^�q¯���r~$C�@J��G��Z�)%H���q�^�l��#���UV�в�-^�<lģ��Z%&u�z��s�_�c�YF�m��JŶ�/��Ґ����uSB�KB�ϛ�=Er��覶����m��h��cyjuz@em������ڸ�,a�tlK�F�q,t�a ӆǪ-?�� �Y�wd�j����lhĖZ�Э�Z��hN�'1�yi�jA�L��PRc�$}�C�z!�����p[y9��|&}y�>!�iA2����*gv�"z#��]?1�C�}���'W�Q-:�+8����}
O��Q��"0$i�/�G��pl�V�H��B%Z��ZDiK?�\���<$�ʐ���5�.�\Q[�.ƛSVa�����Qޖ����C�Ģ��T�ں�J��d#֫/��h�Q�R%����H20�!^