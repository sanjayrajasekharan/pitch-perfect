-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Skf2gZGxqnbKoimz0s5BaFmNsvoMUYjPxxIgYPEhIfEHbnvJDFnaOAfwvtJYpdp5XDMIf3is7eOT
GJTTSfaHaO9KYSO6KK0/ItarW2+iKtL2TH5Oz+/NnL1WNTOAL46FaHEAswEcS/vF+CycRhG6ArkC
omFOyodv8YQczqXZ4QauAGTF2+QnSG2g95hNI74CaUcSq1z+od3eDByfuI/gknTj3c0WC1HvXDNX
q86ghtJ1ZF05TQBcVRcnW2Nxo+e5b8Bwos82bRH4ze49ylv25fvqUjorRwJKEOVxY/Tc27P8gl6E
hFqIMe/n2UiycsSgHSk7oR4ddcvQfmFTvFMETA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 34704)
`protect data_block
iM5Dz4K4xXP2jVtBgF+kGpbWBFgfzIZsnacfhBq7y6sBBxK++rfcYh7qgQc/MFp2t1ESx4iiy628
EshZZ3ee1/a8q7zoTI1yUUG+R0U7j2bg21zL75+6of1nR8NoYGNCCVfCm32b30UWueq58KBYNAR4
rfY16IGeTYfCXMYvXXllNDqfEi5CnYgTUyAqpCGKFrliKqMt5GnLMjvXPkv8oSeUJRwdugUEZ+Fn
FePxsd0kjTHK2hZ7ni9oDzpDKzp7K0BPYtqYjwNa0fr9DtvGUIQZL3xB8tZ32OCOcUx3fe1KtyaG
ML2Uw0nlyf28/Jfpv2a+XnN4vEgu6ko6i/wzeagJt0PNBygyqTlHNWZc3j/3xOqW867Urld5bE3A
CalGvdXjbPNuO+D+kfoKuNYtFyKDkFOX4XLDVEZc5i3dGeieHTxWzIMMXJbcQFJanC91UFLw4bUL
obHG8yDij7LKVdj9N31qB2NGzMpcKDNRza11PfS+gGI9uXbiNUjI8x2Wuw6Mz8uFLDVkn+ibNZKp
Ucp4GzOZLhfbwjcT5vQV9gJcvcdRiYD5LylFJTWeYax0duTVqkts/a+f/UCSj2vxDO3SGtbt5Ivn
qbNB9KtMHFD1ItPlxujp6BII/TenC0fnickJBj8YjSNpbatAvBaj1BcEBPZ6l+52iKuRtvHIdi63
wZmq9a7L650Z2m1ekbFcO2YmCvRbAFhgoiTu98bn88/OZRitTSJsHNWf/wJDB5du1bgjjkxz2Ypo
HxWcQiRCXg5T3ciFJy1/LvVoyAtoEulB+U8EKzMRsK+sE+Br2Sl787FPSPkXKs1FSZGd/gC/ld1a
rNlPK9ALhZ1kF63Wc3H3ubKUaJxLKibh0wa40mazWhzbrcrYC/oLWbgs//EOPZ1hZk/FdSs/43DB
bLz63kv1GJVRMwseZY/I4grHRJOw0is3qOhpxZZwPIoF8YaMUe3eAdbzheCOM17FvLTba+XOAQxP
u/z0QfjJIXELU9CDVLFnRZtgva5/BgTdwu0Bl8jvRehycuNzTAAgnA623kGZa7HZnMH6CJ7wRL0b
caqXGkErF9rQEhUuxVWQjWzKNPPOKhgocsPYNbrmoJe8/AE1B7YXbiExKynia36XSZEJON1154Jb
66+Un1nroyDbQZ7zGZLOiPLhv9V6NN05UTCZl+BcOV4m/lHRNG0EGl9v0ioeO3+1lnR+1x89BrkS
ewTpS3RXl63NngFGL1QNtix/mC5FLBtnuNGFiHEyj2aICnHahIumFiGcd0temaQVixqKYrN13TEN
WUAx+KnVsZ1BvhE40J9kSUf+FP5HCP73Scqxyu2hPeVuyBxj5+uHuejaKB84IE7Jb7pDwX2Zh1UO
1zuD4XKkpdZ9g5N70x1b05Ts2f3iM+uryNyvNvKeDS/11XcIDwIL4w+VYiuyKjnRMUXPXSPIe0GF
wxfdCK+TiJun/cECMysC1BmRGHb+4L41klZ4DkhLRwHkngKLL0SwwZ31NEPwvHonviDJL4HHBdka
FME5fL2zQo9aQKglDrefp3DBrYYBS586YUhrkeFAaWeCAvKFA7sJB+2ZewPAgw9+H8WpGhJtKEXM
N+TSxFu+H8iXX83TruP7iLAKzwEdDCr+iX8dk2ALhEPWFt4fBJPaXPMdcnm2gG1zJHCakexie9HQ
NbXG0Ebe8vpwHdsyWrjHR5RPT8fdJKvheTkBUcmj0g2imWOEWi+vI4fIvXNusu7f00bR49LzOdJa
T+tzJXNZsYaHTtt0f7ZEm9gUcuSuc+ljsktE57Izja0b7XV+KTrxralblCo1znYn2BvYI7Y/j1Zv
8sgq0CNzOzuvRz9gl7ooMhre1t/KLs3BfXzgVMbIujJ7jjp6V3zRe1m8y13VT4tY25ZnQrfxfES4
w7YfqIM9gNE816lS48M/5rGcy4kcXzInu6VPJBeV04ocpza05KkSqc2lNYi/SF0rPeiU3gnAc7LT
DY1xK2WeFyBvE8ERHXQRfMGBOci6uGsE/HfOD28q+VVvAHRMZmKu99pVPdXjmUpjyUuLj9vO6ftX
7UBC/ylciuWkLYcfMmsFzzGvrLlJ5urgQppm/p3652f6CW8cRwKCervw/LEHnWKaQBolii55fv/n
P2vEUnfb/r4MIEHjeM88kfTXTkPwF3T+sP4X4oCdU5HePZsN6Adx6foW4KaauyYwQBsMgGIkcgWC
56TQVQAUKQG1c0Qv9voliV2Dccx3ah4d9nc3w8G59ew9P8YENQGyKFeZce93VaXu6LdaShrBHeN1
q/I+tzgxe4v6UeJaSy0kHDyvatBsNQiUESOqND3+IRyGa/WZBx0Ehzc2KTedp2nmxk0bApDuAASV
E0jiyY/473pEQ3MdMlLUfcRl1FhD97Io0r5Qm1GyBV3cxsQUyWnMLxwz9sctkHAya/hvybrR9vcG
XHtIzvEBBwQ/cpNdObCaxm7P5BC2fyu8oJYxz0mkB1rCxy9uf81soJBvR5M/bPCaqCyLhb/ozdEp
05TKCfUgkZbqo4McQ3jCtu1LTmWg/gQCmagEfMT42orPm/qu7sZaD474dqdoUz4os04FkI4cRwZF
/4fBx5tEx29DiDcowQipd80j3U22ylXYODzC/KohcxYaXXLGCyXUd/gnTuB/BYNRqRpJJVWddtpF
Vr/9lqaP0Rz00tA6hBwm7ThN1CTCtOHQ0D7OiZuaHWLrc1foe2LnkSXgp2QdiZgOM1r8FBEbH/Xj
2IZs4isIMlaM6ORrXnSCdHKNmFKt0Q/Y6f3tjx57AGHOeFLaEQSaq7pQiVXNZanS8HMZmt08NBfO
O8a13FywOdZjZFXlFTrbh0Zs6AuFRZYfO+25qOTTfECG7j0xVo1CdAoWvBJZKfUpkjMP4yVg3sQe
rg2+AJt20uspM0X6Er8My/2Mjac/+cQqags2N45hwwEDKS7bxr824bqxV6b001C1ChtNRl2RzVFB
Z+AGzb6tZlAwNtOujt/GHypfslbBvuR4oNoWJGc4+O53NdFeZ7IXFtU0O7oCco2R7W1xlC3Q+EyV
E+IBA7+sSQCJ8g0uBQEKuO960ASStmdyjp07Ufm7uGViObG71P3k8Ic+bpNjdFjbMyMFmvw6HSQj
Lp8U3YxGkJq9YjbMgKVW/cnWZ46W20xfJjdI/NYTElerAQ3OEvKsdaWuC4yr5LRZumGTFuLsfe5Z
+Ku1TNqVBdZKPuRcyV4kIcKG2/0/o6y+hZg41oMsha+KB5dJtWc/uZz3hrnHNfmAJ4IRvGo8JTnj
eHDTpWw4kSImWXZEj4emxJ0liCXXy4NeH7VJf2ZA8mwRed7jLCF9sudZ+B9gBji2NgsJwuBLwagt
u0xDDSHMheT/2gCFx2iSqT3rcI0Hb+GXY6+tC97N0u6510vG3H9+o0xP3yn+fAdv5b1mIGBZqa++
Bl+5dctzNac/mjoDJqHtL9GgV7pwo2KQ+ZcLHfFdIys/Clk/Hn/xOxdsHDwLZaLad6QojsVQhgAI
GTwVDX3ToE3iVPQBsge6nHuNpFlnwkBuNh/UHOtD0446Nd9qKVw8DnqMzldmIJehZXVt92t+n2lV
UHAOw5yZhqVqeipwMhpSBk37Z0qIdBq/l6mns+SYkgErGUsLrbl9BaZWmrwH32by92sQofzgd40m
ahbDY7on991pHZb2+vJ6HTVX5hcMufzYx5SCZFxKTipfgpkUcV2j5DwADswqtwgC0GpTiXCzG/wg
Y6ULEPWMVvZwlsyJCxzdIyaq0tB69gZlu3YGcBIwTPSXkb7s22Vgsx8dctH37h8qZhrhV4JqsKux
LS4whf+BW1LjBabsCD12XJCoOgVtFSEX87+A8AZ8b+oLag5TwcAVo09ourBj7xxY4tb01zb78/ul
gXjD27StMEwikWCENtUj80isyU8oIn0UY04E8Tc3MyYxLpN6RJ2kQzoMyO63IjuQzpKhiIZmHwTY
CcjGSIlqj8+362fAm47qLnAQ4+p/Hh4SW4GGtQsVXEUWcNcN8NCq8Th8algeWYjN3+nJR5v7RdhO
9MSZ+t33Mt9mXj6WiV5dGIZoWw8gsSbbp/wwTDaeSg496Ls6QXqdOD1ZZ2MIi97aTVUv/v9aiTMP
ss1mql2C2Fi5B2QuN/WxpZd/FQns/mgQpw96DvCFkbCujRba10odls4U5h6Zb5HToSdp+pw7wGJ9
GL/ZW/4jiY13NY0hUN7LYxLUQk/rqBXYgi10mbO8XaapJV3MdzYAce7ZUm6czViQb2JWI22xgHA9
+QNt76DjhILCDw+FWBG4omdtf5EyWyxt3X+onwkKJJkP1sMcb+de4BJH6i/U7+0vby2w8dlQQE22
UZ3e6dEmJHT4VNdEezUUrWUKfMznMshX82gZwu1/TRh874z+tX1JqkQe1Tf/rZ3P/BnPniJJ88rS
ySdnvGKW/2oYECGk1nMG+G9sjpjLG/MPBvyUJ2SWqVYr2L4TphVgYcAWD5kkJI2MTVe+j0QhZvSz
Mmk6z+rqJV3o3Q+tdxXC2WYlAFvDKSNMjgAiYSZrAWzSQdGei60Xqr7pE4KNK0f8IX0bOAYGM95J
X2bEAUOaIPk/1JXX/R6hdoJe+e5d+fw194nzp/2z5MG7Wjh/jF11KIiE2CxcQCl09zy83csQsWVx
Wrn9nfSdm+3v/vmia2U404G6gBMuRzehgBaLACVy0YZtMX+Xk0daeHeCGSaDbmxtDFk0HELqIQGh
yGFIoJc6QJaCHkb0t9jGrxFfqFX+NYrFJ9xHzYMSkmoGGGNfRL2/ETWHaFCXgRXqd1EQODVTC9D2
XTTbmhVOS1rd8tVuAXA8KPQWR3kqPhDqKSmRGvgiteo73M1HkBpLAApUdO6KAX0n+vWfuR0nE4fG
p2B7BvfV2Gqqdj2rIVhoSiasuOQWst0D2QBwLmmgk+LDKODChF6m8T5VeE9bU53TucJTh5UAxirm
vLVu295oT2fxBYYXdkFLtU+hz1meettk8WTkmr2t/T+7EHyNlhSNB83DvUyO45rffkMxel4bdkKF
6bUULX8TMY+lrtzXULC7pE6qi/ppRYDhhwA2cCKXUE6/+8zNgExjygZWWloIZHv6r4Ei0a9Zc9Vq
7xklbXQTfA+A2LtO7jquljNZcqmcu1e5aYbQwhEAI7YJDa34od/cbTeLobsfx0xRC2KI1DnWGG05
YCO3J8nNkmRFRspWZ8QVFNHp1wwpZJ01UK648TM4U6kynFfYhiYJxpE5uiJqZLYnXrGINLL0fIws
4swsl31tmaTlSkzCz+6kqpPQc6pWXCzJCl3ibLvD3dqdqo8hQqNOHo2IdOLbkwH2QhPnMeRJj5aW
1WXuBueM1V/qk7DlJTFGT7QcDsgFZXpViY3M6BcJjzkfK/HwT1pbgGJai9adDNrWcVVqp+QlrgWm
fL1UjtY2jsRL3UtRvk/orxveU4VggLKNp/91vzRrLxTJNvZihQ7E+sYh0rfX1gFY7TIU8eyvytU6
HpwSodOzVM4BaOllxjh5Pw0XM5WtQXtjuKb8hqZA/srwNYaC47cCeKHsQLSVuTOc/TbtJzd7SMQQ
wJ5zqcRAsFInE0U+qBV9flhwOkBt7Q4DzIzpZlN4TWX4+XetCusiT1YL4+KW+G9DQZuVzWIyd6pJ
SsgxWsSKQEa4CZopFuI3SjJfNu2GgWo9FK0FYyI4j02bEunxgvMnFUzX0CIPLtvkhbR7af2zlU2p
GWWptpUyFTYW7RX29AkGGicsIcK1rozO4O1TW5gz/0ertBSfMljDRS9SY/8auxKEBQ0+7XCSFDt2
5xv5KT3kkTSnlrbtIxb/LGyxOANvO2bcdtdfAKqIrujfxvwHYxPEm6dI4C9fYAsKV/qqOsZWPZv0
de2WXF4rKhC4S+n+BB3qQDRfD9BZiByY8rNMYTHkECwSDKOaQZ1XMXkzbaX6b/p7mFvf9peduok2
lenbFoQhUSH2x1ApeZvJF9c/YoitXX6PwTt/BkpBad+zH51XEsA7V9xrMbSmYW3LxFARjcAdDNhM
OD6B3bMw3gxdggLPRfdp89PSgQdQKHYpvsAkkgVKfhmRRRdcqOLQJdtZeT0NbtOtQczvYMjRz1Ub
8tNgjJ9yP9kOu0xoAnhFSweoWMUgEO6Zinxe3iZW/gJ661bVYXxOZ7CaAEs/frjm0TxbFKGP8AqH
SHutHieWyw/hwcVrw/f0ExnXQK8fj5zvmvDGUybG3n42QXlqOOXX3Nksr88mTklTRFt2lVwOIf9A
bZLXBfGRhljdEfWn/BdTphoLzIOO5x97sN6+h9ttxPyqGXatMUZeOp0kTunDnC6tjdm3AS2ca4D9
5Nb2J1myhiyYH8/t9513iWquPVhdETSPWLBi06UGtTOvYPkkICpptbDxR10W0hxuBqoUVKn9CuHt
zvjSGUYt0DB/Kf47hAdowxGBf6dBiODWiebaMwGkxKf+IE6GpG67vWj6xcNzJWMsDZqBe/hP7F7m
qDmSKXzjHmW6vtQOxGO6Vja31xcZD/7Mj5GIQjHiU35+Ry9kyZKihaCc7qQpPdLFv3QhWRQKsGFS
VjtZKl2qOE7uweGAB8yn12TKX5f0PtvcI5kag9E7LjYGi7CJzeXWs9GTwOaJc+kNreQtSFkuqbef
PuDycZ9Jw03HUIxRW2iD+5tD42CG+ap6+jT6hxg9PuoJT6NweqDffkdiY8qgQGQLVu9FB9U6jCrv
IR0UUIIrU8bYRrj6TSPZiV/zNqbf1Xnpmm8sLqFH6RlWYSctpg3S8suvlthwZOsHc0E7MHXuR6GT
T9J95Gs020q2qR9gxsQW+wPrSZVOLMvIKFY5+ZaX+5oUoeaYqHe3hHRO1GVlq1bxx37bcQnBBZPB
MSWYZINFEsr8dW1pYfmnVABtiVeJIWdGsB5Br8uNe3CGnbIXlEAqyUAfe5jYhmDhQqkhtKn3uT6k
gC7ympxKu9QS2rWf/2X5OwRoGQrAfo5tXMS3vqcYD3choEuWHmHrow+iWxpG7b7P4NvC7rY3Fj1m
g8X/MEGu8H0M4DHCsWSOUS/6m+gpTI49Gwht6AlgmoohTedl5yzq1qYcteg8Pw0mBA8zW+3EIFtF
HqfxcGfduti3oLnwuuerYjaYqMCX7mwnxc0rdzmi0Hgado94V3EE9XBspTToykBfVHAYro13tjJ9
NhrywUlcquXTLzcml07ro7if2ZyBdDtZ0SPJURzsYuZM+wU/bIOoq9pwbZmCItmsAo2mcRefdqoZ
k23XGOk6zev/qWN3VeN0KNUIVY+SEHlMqmIoGaSqRpujrflET51XorbevuZ/8Zj/E+rtysw/gMZO
SHYePwM8x+Occgn3ajM+L7SZ/vkfdheSHxJSJamvGXsNV/+oGwdWjGcsvJ+7US7NQA5A93kPnRqj
C1HdfgXpg1xEzexfsGaTpF6E2p9KSS/pKOAflTOZ3OGWLm/ikmhGbv9cki+4WC+BBw7EBOa6nPSG
Sm21xk0jcZHdcDI9UYNSFEReElpCwhuHJgo+gQ9EarNYZI50NBmtGCwgE7bsiZAlsphEPJv/oS3L
qGuvZDMAJBuek6DIPs6iiBgjAtffupxswaQdXfHjHghLIusHI5a1T8HToHuVg5H+t07lvAIRWEdG
cMEe/kblhWiFjUGvglsNAhm5BkMrKNDN8DqUmgkirQmByzMynPuNuX29pYtKPeZMEjVzglOWXt8R
Gww+3EHmygCy//6fdBpWEPQ1T5waEQEWMHVJ8eAyUlJY3bXSIr/q6ARRuD/eRQ3I7+B3c8ai6nMN
s1pyqbiKrcVS+crKLDbLL+qZ3XG3yIMGvyL/kNMUkS+zaTi6yEH2jeXlRVWPS5ErpM/s/u2LCgnG
TpwGYMnL2wqby2GIQImcgZ0/2ldhs1YxjDQa1vu/8Nl2K9y7FvkllsABDJct16gZeY/0KPyXV+/6
MJPjlVKdQbL3dwQRoRHhcWZhQl78X9ig5c9mfNVQG+VafaKn4InMez4Zn5clxl7fHe4/FdsspVlK
EkQSJs3LwRUkS1ZrXs41f0B/rvF1tycg76bWTzOXcpSxcbQQE4cx97qF7fhD+QE5g+lQS6dg9Wd3
L5d0TlXz94hIXL8RbiSQQz5pLFgq2O2/pVasRGrtRrY28IYWPRQzH7mqMUt74AQenHlLrSYI/cc5
FxYLcNYhEB6wfQeZnWm3P8wqjCBv9E+1HzO5VXhYi2PuYAk9Dd49MefXN/nR4F5Z8MMDWTFzh57+
yf+XCFFlfpAvVnG/XE9fmUk5q5SMTktXm9Ya3M0//qp/so3CIxgAy7NKdpXxjPaVnHYRo4LY91Ze
Sy/KTe7jHCXtBBf9ZmkedMiuXAHdKSUSEsanrZWlFB0uf0sP198sYp+zLKiHLqosrvianSNRfe0C
16oIhonxc0bNyRm6CaRjps2qxWvvoVkbQLhNU84gw8LflTCJ/AY+f8kdnPpveuswj3Z0RVQybvzH
e2lTZVKiMpfrVc0qpGkC68/aAZA7GOEhAGvjE8sFPNzl8gQlRVaKMfhZYd8wChDwnikO0UDCW2tO
me0o+4a9li9h3bIR7YaVcfzAtQQbb60FuApNnZrXka9SttSwx/3XSfFODwwl70jh99ABj42yS9rV
VVR1Tj1jvjD09AJmPiHqC8R78xoL20di90FaZqGlx8ejxHwe6UBUMXHcSL4n3S5iqQcPU+8CAgZ0
LFSYuIfn6BlBjkkzQtdJMj9n7adQVhIL5lI9YgH9j5EXjCZn/mtq77ER2tRsM1XJwejfq/iYJemu
3lLup3Y18R72NI/6/TbzRHM+8JgQxhjKcXjbLDlyxLuKV9bigPidTrwquMKlHCgwjrj5w+lybY6I
8bmsQkKwRbfVNj2f/ipjQLQQDHpVXwnBTAsApNj0zu6R9GyaGmMT0W/HAc6JhxFYati7pUZoLeYN
yYrQZZeIRD7eOQZOJs+PqrYpddH/Abx5EzhZBdCKn9g4ueTFqQlGZQsSLePhCYHWrdPOK9hQAY4O
SUjeJ1ECMKCeGy5IfRLkqUP2YnB0AbqdI0iVRGKoeUq1UaLX/R0vcYtGdxdTJ1BuwyoKU3OL2v+k
6oF8ovxnJfwoYp+wrDLKC8M1L17XlZJlViuK7GBh13igWmd/tSrQEz2/KiSDdLI/OksdnHVPL/uE
fnfK14aODxSeA+ir3OCyhPG/fGQSd+kDZPtfF0s+sRg1QwbWVUURiF2XcZbaFZ2SRaX+oNDuKpxG
bz380GTuAN1VKZQTNOAisw29PqO9ybBv6nPti7jumvhM7HjyvFpVFObOG6mni7rHKJtfu9ElTPo3
56c5sX8Ol+HuqiVsB8zYQJpCnDF95rwlua9PnBx49UugTy0xiiHiOSY8dOS5w6Zox4xYofZtkrHO
bbi/oEg8GnTIAsScpRUhhn7D2ch4uYE5eJupsRXL38oZNh+XncTnKjx9zYnOJCKFnHBCp67JRbZd
EhMbfCuO4pFaShFYkjAnOq0xlA1KmufD5zs+dXM9ZbzujJ0Lt7MGJQMVzglXul3xMMv/1rNDn24p
UQV3UOJ3pDzmI6VcwR8XKGAzoOs4SaxD/oYDy06PTwSJCpXr5gyycSORQ6nO0n+eugupGgR4F+Jx
Mw1vzzQ6iaI2FXsGSmrj8IugBad2t0xTgbrDqapyXVMsIPUhFQTS+C+Ham2PqbsE9AUTaR4MOCBm
EUD1Rj/2MzXIjJiXqiw+UiHtHkPU/PR8rht7aC1199VY2lAiZO4X5FfAcAWJCIEx5H9udmRYTQM3
PHy8ZA80iPH7/x4bhRKASoHTdI5PadPim6IPuqYZTwPJqrQkFD8Pq4tpysebPeNJxnb4KMtswhad
1K5BoIYZFAFilJ06HFc1Y+QPSwsjfqty2czEePNeg/DNQYzvwYBvTaX71wySXER7DLGH1rjgOG4C
psk7ZXN0MoNtOAttWBopj/hXWTinqVDUDu0ZaG7XgFBAjLk8c4tCBV6XHOQ4DlszEaUGpf6621di
imieBlQK4u48yBWYl2i4T1IIWSrA5zxJoci6dXE5WFhT6JYVaIqva9p2YkuRbFsNGoTQADOeEmIA
WI6ApcQ03c8s3KV48Zq3TNn3soQw3j+8QFHs4ghXj//nJBGav0w+mo0JpI/cEYL4i/qstR81TiGE
3HD9sjVP9kW7MIVIKephEGSmcZopT64Hdya4xWfZ/C4LsGs3pI1/pFeytwoZ0DqlwXTvSSuKTS96
d0UkzCDWbbPkZ+9bVdHkXA7z+6ZHhgmW1evL+qmXIkCcVBv/aLugJbJomFExy5e20usE5Iu659fh
UK06g6tDJ4USi0p0+xout0N+gbcHX/UmKNZ925Jjc7WwNBd3wRq9XqdwFhu5XGxuGrdWUXbI5Ipi
tl2GOriSJsM0g/csI9/l16YdnbvtVzVqZNooZjHpIQiSnw+TQRLDX2hw/M3ZknJGxjMWZabWp+Kw
ccnv7hPCH8YvSllSwDa9QLNwvy2FnU+0/sq/wQP40M/uhagBAE+NW83UucpCOZ/Q4Nbh/vOh8f9F
5/J17UXgJnxIsf/maf+XUd70J8lWgf6nzE+YSZDAOHpT7I1KCVh/x1qErIt5FbW3YymJDdON64ll
r/kh+yyK88Z7Te376CVMO/NaJ8eU51bxaDx1NN7D8W5cHhmGpYW78eS7zZaWmGyytaVj6nYIPv5n
t5f1VWafWQ/6/1hZfJy6DyvlpiT8ullSoP0/kRe16hN3P88fIDPtk1Zp9osz0MJRwuSzwHRvGarn
E/Xh28Gypr1gt+UD0JpJSmIS6kntBsE6i8yPO7kz7v7gM6XauU8MUNPJMWXTRKd6HMsjAaiwGHHj
CzT5ymTmwq5y8Jgb3oS/VEI7cA1cDpQrlxFyW730NVzOZa4YYXzOUJFI1lXG1FJgyumyI2tIroYX
MW096n868flHzsryQ6ln2BAndkgtzcg5hEvU/h4qbcFWB9HeIrGwA2gIxg+vR6CiS5LZfHYP9zgs
EwwUYUAA9eUoldkb2rU10cfHW3QPgfyZzXi7QOD2u20ypSwaStcEPj4aJAoZCt6YoD0qOK+CQKcB
l/aZ3f0BQGtTb/exc/Kyj/U4JPR83gtcHimC9XzI63tqiwYnW/iW4Wcgq1NuB41+DW7Zn3dsI5C9
wO4l20U5shmlzDipqy4Xd6VYTYxa1xWhitNn+czCV+F/2mk67dJmBVLWi8KQWciKTTJCtucHpV7y
p2NQr0dpUiFjjCbUQhOGHYCPt6pmmRR+gMwYZ/bbiLVzjovIzFBPaD5i1bc1TNaMEUNbzrrlcnXy
nLkQ2a0pyI002wSQ1+dXnsRhdCUGePocvtqmAtQXOXu/KFN5Ei7J2TAGFBG4WAAV1xn0TKacc+Um
cfaoQVxap0s6PZA9GNVcZSIsHp5PMzuDWufJiYmmndfrF+HiHxAHRQ2wfzmHyaPFtjP86LUzbg7i
sAMIn4NUuWkB2Hqm+K0E0VrXWaBM3bD3ykzUqkqKPdoIZbHV1V1JKWmknvwabJkwHuJaGSqfpsAR
e+VbxY+s2Vzh6da2jfWiSoaqZPB2QVD+kgMXuFEJVCF4YkzSYvgVPy/6wdfsO9Q/zNMOVNU6eBNG
NQVjjaW3U8QRddw7MfpKQoOV3mtsQtZbCKbRpVH9AToCjoB32RMV48Jk0xBw+dpbblE1SZbLczGx
L9El9u7ZAJd2P/avpT4YCdHKdgAW16YfgSD3KnOWqHGHIaHTyJp/jCXUuLdZn+9mYbD5Oh7fHwBH
jsDIkQAShaf6mtEVwyXL/6RSmfC413EvIKnnyOs/ULLaFgFgv0nfNFsFhebA7UwgF468hx5MVuea
roI/QZtQaXFVAQ2u9favcqPCBrqaJRlmxmSs7chBT0FgYzNZzx3yjZhmqmXQOhnE8TWRrk63SiJ/
OumRu2Nn4tyRg6SQeBrlufocDV62RWgOcuPwXV/n817NUQSjrJR7ngSTnBAss7QK3SWj0Xc053wq
HTK+I1Ttah9X4UOSO0YEcsTs62V0rtz2bc2S/zJKV6N8ZGFUFi6qphPeD+OPonQjrtavPWsiAJpP
fl+qIHzLP5f3Bn5GZqLjnJNZrIXXEq2qfAq2p/JVRa4bS+FRVnKFr0zFQkol3Oap5CP1D68GYw8y
yQzhlTTRNN3aj9JMGnPBwJiop2pO6z+BXJj8lvnG2OF7+LqHltTfe2e/7jLKuNfzstBDlBX3N2MH
WS1Ed7kjmi5qVVJrhEydkRJ/E60cQZA3mN7xsIBP9hOqmWRuC9DTWzrQQVmovLay9XT8bhOt8y8j
V9MpfmPSoc211qWtbZaR9exLBRytT8Y4qlftzquEoxe0+t5N6YV1yec3HMAn4pJ1J4zQFcGI1LqD
AEwJZy9jO+tBbRoVkRRB7d9KNsVd8qkI58t77aGs4gXVJSBMcDdLOZ5n6TEBeKyLNOUdK/seHSKf
YQxWZGJ46UgA+EKuieE5v6YFdhfAuIG9jjEja+un9RAV6t5EVFfg0lCW3heR7lGFici+NM5CWNUA
QfWEjxPEJekuMCIx1vQsL/cwLYid/bq2ukX0NRVa4b72uV9O20BYnK4Li/AMwvVv7IGUoj6pAiZo
s6KjBqQwDuvBWjS8XGW3DOnhg2MEEbNyvk1lq3PmIRrvBmtgd5ZlZqW9UW2ZuE26T1fq3TStV0eu
LAFa+kEkTvaYS/gy5E2Ag1eP2KbJ1tTndVsceJDRz6FxWWR3tq3B/2LDWZDd+bjIP5ciQRNDe/rE
8y/kzP7B1Wsxg6YDIGcqqM6RU6ooyMScQ4lg3Vpdqa8I5tCX4AKQkQS8UMBtmy2pM6xWz2cfpcRp
rl/28mol81Q0paeOV0Hp+l68HzUhLczB1zQfnXOwyU06nDFLiGkywJpFxUwD5Aj61SkVYRlznQaP
K0bPiin694b/ZubwAgZ9BZlDVbYnkJKHOsFoFUu0wwWRr/e7hJ+R0PRMcQe/E46T/BFkQ1WrBgA4
WsRA9wfXqV1HYcUeToEXJBrRaVzT5nERfmvloPa+5z9eFqH/ierAhI00tib5bGr2n/K5+D9f0/DG
Fid2pOPWbZqirpuL5Bgdnjm1BL6vqktJPtRLpXIVS0Z0PjZD2Mdbcqb2lkYCAUj5eoH1fEKv87Aq
FAUBm+du8aFcArQaEVmJ3bJ0+gY9QF8r2I4FC1uVLSepcfuvSOIo6G2BPhlrP68VT5AwLhQBxSv6
zi4NfqjHfnckkf9vJEFhtVxGm0sMCjuZGtBufm1d1WlWKR8idxuOYbZfjDjp/YVV+jtkraQ3wB5q
mmKTYNW1AIL/VMD3fSWtfDMYYJiCA8lqdBQwnfoEESNr7afLM9uFHs1KnGH6AskgdDleV1N5tT8e
IapPY5o+xx/pu90os8AGje6MWL9JWtZq1MZ1ufhvM56rW+5ojHQZLUcjmOVrmRIH/m4UiYOcHOs9
KwIMo2JZ9b4GuEDYYIud/sQyYwJkRc/l03xw6puhSVA61ES1rVCMJEH3Kl8/okADnBklhbNP75U2
ER1L2JY9kMrZciDKOy/aUuN5rube4ifxpOT9yWJVjRhCuq8T7Bes1GsNR53srgnZryRsoF9AudzM
HSt7SWY2+NA2l4n0fzzcTStiprWZSwe9UREa9BfuaSn4P2XY2nyHEQWLK+TnwlPLSz+YRI9cz+n0
SRL/w9sD365nVQrT8kBSpOsOSve3Wym23AjEkRIhmOaoX21ulDOa7QfkoU4ZXNJTr35oXAwok/w0
vutQ4Q80DM2LMMJ7BixUp8IN85KxS95igPotqFBXKFg6KN63RHnXvwJzxfKZ2jCrjc7xto1cf8i3
r+Azw8dbJR7TZvkaPaQhegkI7yKTFF1fXcjaqdPDbCQ6BmPTuoL6kOJmJsQfXIyb3zBGnpuEvEfI
WlXXZmGVbzEm/HknjZGA9YobQTnn0hbfBI7IqSQOfzpen+qCGOOQZ8RrWGuEpE4Odm5RuflZPDkL
iOMrbzjqXYVr3nT6V4NQ3uLcZIbTVgpezfZ+17P/f6j8YnHv2T1+h9vtgKrijEQDduLS2a34ta+W
QJB4OCmudzBsypN1EkgT3Jfie4UhPBzY/NzU8X2q4pKDsu5Am2afXuts8vxZ1IuzuTXIrn5eicwq
zGt8oBw2RALMSHmOot/M3RoHObi/AODdFlqwJ3EnM7j6a5deuK2SU8c60N3uJ5i4uRisab1Lklgu
wjZ/YimKzhHSjsL1X8h9YTaIDvCFU6F4VGzYdIAZ4J/MzfDE5PyVw4QS4pCac8b4O+ViM1pi7WLk
gd/P08a79TIXXTyMYcYnGNx7jQPzi7I/Wy4n9NQ7ko3DLxHevMqE3y44zg+f3amfuStrve9ZWbn8
6L4LtuFm1YRWQ4h92Xb+MZbMUbH0hfcUCBxLGdRtdTBCC8lxEqBlGaYpcEPdcBu2d09+9icx0d1p
jr29u4iJuJQZco4uQUbhJEUpDwbh5sWy1C1pDf4xwBVn7srT3CBuU2nZacZHFeTjwv4AF+LWbK7g
A8ZqpY+VxWuk2HfvItpqBLPkVVC21Qw8DJsN4XZajbOzlWhnJrKCZROfYokjW2r9r+sRQA9gvd56
bwM7JIClIiZhabC5Z9MCtpC9KyzFRR7EixXL4MayTt0Cz46UZYSszPArazAMpYYhuhEgGw0OBfiE
U+IYR/nNH0qFbaDvIpB6Zmg6bNHLP2YDWCGjNYor1xjbwrpBVhsLlZOCEvOqDKDGszDotbqUbDSm
pNEw5GuAgWBN01ZRnX6TXVDbn08YotlJ1V0ab0VVXmsvz+8CAbP7YJXhYw5ZnZp0vor4uT1ITz10
g6EkV0WmOG2D8DFdTG2frzs/htJFRrQ2WESGPcNyYtQIqOTG9gvG0BnvK8BN36pRFSQ4UV9YYA90
sZRG2PKx5XjJ6nMH5MiZCixbHjbbFcVVxjo9g2/gTYjVB++gEjK30O6Upj0f1LkTl4K+BOPaG2m6
c8ArdC9FY2GoDWMUkFE9q4I+sDGFLGbPp8IxclUWUCqjFnYwMTCyLpxDhgtHpA4797IsxicmjtU2
QTfoChE09Cp7TGruwuYOQwzmnZx+M34LNIQNzTw/6454HeB2NIQ1imqpM905GoyF8WjUjeS0gdzX
k69aKtlTXqOXV4cK1fUObMPGPRHDwrZ/41CgR5NOoRXcrerRVHg+J//DnoXavSV+YPGmSSKe57fR
1bcT/4pWd73kfQI38uNbJfIGxM8y8Jmdt+cTEzqZrUAaPZs3esVKZPyRAdA9e01IM1cPYBdHK3f1
7w0fITlOx0oWRmDTZ13YCeCD6l7qXL5hTSOPdnN+220CH+4sTCdYQryDnqK819GhnMWRFJHQmpW7
pDJ672caoZ2ALWaNsgbpCJl5daHZ6pjnsGp0R/xPvHBRye08XQwtvD7FsUKNRtZkr1ZRK+Munhxs
BOeGDCmdd7UJF93cpUDUlt93yUkYJ7ukh80VZy+pH+1VQrkgxP7E09n3nIzMREggLdOwLawpgt3g
SruwZoER1pURnLhS3jlcv11g2kmlxbnKgXa1CVwvuR6/yK6R0TnWVljGnw6JzKJx6842pGsLgFyD
hAs+GjZ/B59QJF7UrHi7gMmQXFhsGIVfCcGfkUzbJIXcK9rkXhrlsHARVl04SjAPJTPYSnv5NN++
MZ66VUCPA60kmvMspjjLtzktSark+QDpkK5tBacx2zSXgadFf596ZRMd1TRZLQ0or1DqrOR4Rmeb
73lg2QwXRQ278hb8JyQcQGdqGvuCGg+6MgFrHGDneuicb6dtrHhOxCH7QmF9ZeEfm8dAc6n8/Vup
AMSEMcUxTf1ES9SCK2JbJG9kMs3zRt9zC/kNoq8uta+gDf23COWt2sdxgo3XFknXIUXiwAMBpE2H
wm3o2OzrXsdgM8ka1qsDrNprcdCNXhLV1STvhfLqvY+RuUztRnZU37K5lDU78IjrprCiM3G/EC0H
KVmISL9ntARvCjs+t+1uFakf78ma0kMSaw9EVN+kGZ8zLwYNqAjMCXP4k68+Ug6NplbOhSdLXu4z
YzyofRE96C9c3CiLXSbV+Fe55Y21VjbPDtWXq5vgYnr41sXbkOSv/8HMFhY5hD6OW4S18cbG0WYg
3VKwp4KyV8wkBJ6jw/njX8+admwoErsTfd4r58B95aFUC2QF4ScLgt7FGCbDaT/x8YulzKQcdT/X
GfwL6g/Jwv9BWZ+27Y4kvasd53k1bANNNs3DdXF00thifuMLp9ro43girKYxAX6VyuCVeAomtRjB
AGxAlvL8iN5mBDI8AGNrTffEXRUKvN5ogqqsqgOA0iM5V3kbKKkQtKRpTfunLXCnvRGK9kU4Nj2o
BovLRhNm6Y0Rlj+ybKKBP7PrIhULcTEStZ3/Raju7njJQGxFrlIJ2K1DqEglthwwpXzBKK2Vx5bx
OhxxR8MQOjoQRTTEbL3zIbDGtOWlOEcMBBxKJeDmLoXv3pACIpPmsNkU04FQpLFGy5EY7k9EPM3W
fjoNqNm5TDHN1PWTDNV1GJfOsPEDAiXQSAT4A0LTLdDJveo77S74a6U0MtZtlaptLKAyWUp7/CI1
cYXICBS69PFsFAzhV0AgxfHn/4hvS17Uc4dIg1kBFBRQDl7Gk2PZYhjb48BG+C5VRKVPKuW77bM+
2xtJxbumIHkP09j1T3ZtZz4nnIY3dlXJQJWA5vGhf/vzCt8suuba9zM8xNih/EP3bae6NYUPf9PO
CJRk+5M8Ux1aNvHv5j8mATy3dYXuUzLz316v+Qrh8FL7eaOigejITA0tAiBfgOZz1Vb3ilyPrGDI
he/XhJbCk17vGJws+M+cYW1DIKrn3/bJPf9OZCXQ2PogKQEjXTOcwD9wimzo+jH/3yc3Xjmms5Pw
LQiZZL60gJHfbU8MoUZ3P4anp0wpa2UiTptOP3of2DoBE/cihcktSxc7r8wD+9QmiIqNwfQVwa/d
E5vzu7/xX/GVRBT2O1zRb6zJEj3+uz3yFrtgbMcf5Hc1bO5e7+bu5e8yqtPxGGkgSTlhD62V21zl
X9hXialy7PbDoMX2hpFSZEjP4OI+RhjVx+pCUqLV3lMNnyaEoUPB5jHOopa5zzSCtajEMFUj2/2g
Z2VhKvA5f0z9XSx+Z0c/MUMj+8NKBlPkVcWswdQwKSV8dnBlHRx69oa5VCyI3VgL0fgXw+PM1kIN
vjG0o/OImBPRwS7gwDWC+Jx0m9vQta2mIelQFKexHcKvQenA6VI+z2DNCoBCUMO13c5TBIQFLFyl
eCIFwfIzCYfRY6ZiYlFgwszZbYl+q5cgmBL2AK4pOAaNnFlbX+YqQA3HLQ/NC2LjbYJB/r+t4cNH
ztyqINQLelZHFqbmdkuXpE8xrD8FP7emcSGC0OMf5VpIYNif9ag2D28sTwVVWxppRFXOzAuaJlFb
aqURpssT8ZU4s8xfe31tg5XSTO48OWM6VHvYMVarsyXoRg87aO72non1C/JulCzTwWxZYJZ0GK1h
Sjfl0W1q0JJlMAhLMJIt3v65F95EZO5yF5YsPP/uhO8Wh6GNF+uiEloWg/dMIn4KcW5PWjU3eS6P
1m0iom1gXKtz7TH85A3efBcMY47Ln+AHZvFE+WbdqSvTleNJsh+4AYr5D13h+yHVlSgvAAAiuQ/W
rrabtqVyG22TXdvFX+SEuPfSLiLOobUJJInJIThBjC9u6JoBGafDxxf3YtfH3GNX5vdL9n1vXDmU
9dVMa/oGlGwrmKYs9iRFHlJ5a9VIyd644qUAWXtgMTWvRmyqzWEQFyJ3icy52/pG8gpL329zOEww
h1VhblGNcK0PqrUd1ubT0SmN736VNUWU4Q8dV7RwiNW6KffVgIjLzN9+st9Yzye+RDpxUyxxREA6
BuXCFUqoyzr8Zy/GYZ9KQcGCPHRQ5lQEUbIGlFZ2pJzV62hSNRHmqrTTKNQDOq6gY4ssuqWx5UC7
wIODRcIDjHXk/ym7R5Ckvjv/WCcTutF1h9988vzphpfbJa2iqPuOQ7QNNdaKQC8e3SVAJsqVIACu
ov+EgHIv9kLNVLjzVcPEkeRvjxTxycCkq8XXYjXzrGybb4frGuDJb3v8uHG+v4QYPl81pHzQ4bB/
mJV53fGtt0tEb4JMwcVdIAUBICJ77F6wZecuGRL/QZoSpTBkGGMlp1dNSgFcDF2jKmCV9F1s0moD
57ocC5RZb/Qylm6WCYEtsDxDMyAX4VyAOxbwb59SFw65GBtBZyQszjAbyCrjYL2qtQMIMeqSOEXv
tXFBgvLevxCjSIWT2ggzdP+wD/kokZHZsTf8iyHP3vAGv+KK5Hak38GACgJsM/87peJMF3XOEakS
tJ5c9xccGqZe9bWPjb0GkqaeQ/nHvRtwxElo3yLA4iL6hefKmd8BGIFyIWyF81IQL8zJAed9fu8W
hzabcshJTH3w91mqSEfBCoZTNe0mQjN9KbEcbelrysfXFiHox4+9ZnonHhHr8GL0eMJqmfVkvHCW
Pt5kRwytbslAO6vlNhRTISKmDaggUHkBxCDaJ4o/1HiMvMPorj5vu3cVJeKEE7Li1vG629Bzn4ss
mxyPYZlV15s23CvKMftbJlfxOyiwpip7ZxxBw51oFMcUWoBD4f031gKuTScDAHQo6rCz9Zv8IUBp
XiEp5xVfyi1YmLO84ubBZrxLqLjwMjdv5cS27zeFyk38IyUXpnsy72ha5CIdTFVqMPyFO/RKtyrb
Sm8xORzllrtoGukvyxxc4MGX5/X6o1JdwFFIoFcvlMIPvl6MLSL3paCgEnhR3+DqCLKUgGMWdoWJ
8HpkuqWdZHCBOcoe3rf+kLGTt6ROXdWzOF/5HNbrbyfnWURXc6zTzkUFPg5bTlTWGYLr4lf13svr
69vTYbKjGqGrzlt+IAN1gxqqvAIaRyjkZ1K22Rmugfgt4AlC9KhS2qt+OsykqsWOgpiw8xN9vUEz
O4WPXWwMVdoFcW0EyVlZWeniXv5aPJ8UNJSBap1hc3C6ExCneurMW3niUga/dM4YazsfLF9mXEIR
R2fyIYOWsqPkoD3wfSiUqz/dJOLiewW4P0KZ2r2y0um8Bj+4SigYvD8xNSr3Lu0mVCJTWoYb7PUh
XnKsqzBP8zk8uKPt+gx9/qjEXPVl8IkVm5bLje/9Lkal5xWk1UXKGpVd4k1K4rMMv3noWSt0xGaE
Cp2+IHV4odN5bl33ocknvudua2wiktoHp24Yl3jzbXyYUL/w+d5uCjMjIoCA23RGo8X6Vaqb20Ja
1O4nL18PTRwY6kx6M/kHbrPYe2/9jGvqXhMqPnDPAwzucI5VXI059JybzfFiJBL7plotNTtmnPAc
jonGBML4VRU2AwGiinVnFvgUYpmdrDKGKrNC35911jgnB4ZxbJ5Kpw9t7uduujihllcuwB7Zg0QN
z5GUeqRvRLsTCeiCLNfKAFbnRpe9WNDTEIQcMyCxrTBnP2oxm6Vcv2rMWQYiNxVh61MnxR/IccI5
gj3RxsJJBhCtTqRTPmc49QPxyhAQgjXPdPHyoLHiRAdLXkSrwkxIGYbT7H0lwJ6v8+h9XvX8de7r
mkE7ujbVy7r2p0rOrCFPoDmuAFpUhTci1l7qOEPqzaOzE5pgaPes4pPVzwWL18YDSXxJSwk9Z/e2
goZjY5F/+5bl8FoDDFYIo3gROVDWb/XC/KWjya62I2B+EP5Mc4vrpI2b78FwmEKjGfGp+mujFwWd
czk97DQnqVHHN3IzOrnzJY4D1hgjJenPHHHzpCD4FhRLIhTka2/OS3vVrTF/a0oOZWxMBqO1t8N6
g5VydruXOAnUBTOzHdzJlbJERAS+T8N3JGS/zoy6pfgTN20nRmiIe/iaAG4gEcW4IJlSzmFAe9QE
KU/U0m3LUc+XK0/AxcLdcRLhyj7H6wo8qwwTDeLTbcKCqS4y9LibuQhRJ/v6J4+4mCDuz32yWd8K
04LJD2ZAf2PSBwN/XXFKdGsPAQZG60LTWWC/aa8kNvC8bZNtB1bUnGSiuDH5iZ6hO+GR8hr9zIwW
uFYE0Zw5ZE4C80ME0d3znLc5mVyYNvPX6DArW6RKZnHkAxoGp047jEzUtxd1ZJ9VeMOd7SB+q0PQ
eE7KJLxrikmBY/exjvmYfiVX8inHKQ2j9JrQa082gF5yBB1VBRtbfDwk0Pfk7qCq0yhx+LOyh4f4
NnbN/wBbsxOVgM2Q8ZQiEGCrjjLBIBpo1qeRLzOP/ExYyLBRKyqji/iOdzzbTgWE94DcuztJdGe1
Gnu3Uxz8Otgx8zYzJlW1ThJIVP3KQXQXbSSRVrDx9Qq4luqD1lNxLlkSVSVsdXq19R5c5tA6AbHa
WT0HuJHxUgWi1CtMgupirFqkaGU07FIjxr32g8wUDlLBHU2FSSXTCmP4ZKQVNk/1fFxpWz2A9qLC
7mXfcmoh/QaCqdr+zTpMfaE7J6Ukocb5cnALdHZ3t8nNtxkoytgLXJp9Jn1i9+2bhW66Ot+Kys+p
2npTqK1tF03gkZEosczRkP8pRRy/xHpTh6+TteFfhe4VdTPnSHZQtAtn7Oa6G01zuB7Es7VQ6q1j
+18aHwpckYhwpaWSZvc3aS/NzgQzMFy9eUc75IqZ4JipIdD+w13CaAem56XOhnycaGsiUC+ud7JC
kgKFnGg093Uuhmj+117iCFqhIZp7pDDhR4LWxVRM2Ktar95hytwo+ddAWeO4jv5L+38Wx5F9RSzQ
1pTLdf1/pqzyMCsJ+OJ/Xk0JIxQL0xDxt3Pr9OeA0Qy0cM9BYkZug8bJeDBzuixtWl/YxogfANMe
DlscjK6LimttMec83arAlcvnxNedxbWL3SaY8HnDUIJt9YnM/BJiibVvXQLcgAC4SeDjhDWoXZgF
ABNM/p26x9sX/eD53pXoX0cj0cTCXb5F8MP7JX0ZytGh572KA93vgGFZvrnbEGOw6gZsRAqfetDe
po23KyV4TOG5nSoaaoyuitGndIFy7py4Rfk0qlFaGqzsM1yFqMKq3tNc1n6URa7Mh1+2eTk9fUpq
cOd3oIRcbhbx7Tt0rnDDfNzDT32bwIdXf6UA/u6qYJF7dYhDI7AbrKV8uS/HImp12JQhvNjpx+xW
gZEgVjW7oY2pXsx594dmAptJAeiJzQPl5R3tpD3MbPx6OicWZzmLFPQUm06nTEOb/QSwCRKA+gFE
nMIv10MMe5GEtwCb7h5mrQZ1M/zS2rxS4lXLaoirYpXYFZ0XyWxk2STYHcwKrT/32d27uHGbyRpV
GmM4jhLPakCGxAeTiTtdkVTLQhRPMObHV6c8QgQ2NUALc8p7Vx9MGc/x0lAwIZt1kciays/hpIuo
pekJ9SAMNhJeMnqLkrYIl/5xIqb2mjyU14pvpBIPJw/SQJVRWdUZjw7e5AdPNujfIQN3juulfuaF
a+rGeSnkAQy28oJOCWPXzCchzpCwpC0RhxsCdOHB2XQ+1J47Vjle7ZvaXv5ZjCZWtPoOE6ZV9VT8
u9g+358D7hnpqOVFWOIG8J8iREHqHHoOMxnYU9nrhFavkTSm5wU8s6KSyedvPFiSil/Vv2RiKOQM
E2Ggd6YkCUwRUvoYIY1Qz6xdJdiUZx5h4c2S3WkZlCxBNaVmdQTB5YwBblr2L7uO5IWrRRq8/YIh
xrs6qURHsoXU3plENHRC1ak/qiRabRnJuk4ToVCqZ7Fs4Jr1VoTA//+pNTC78gufTD9ZtTE8XpCW
dCloQW7NB27aF6ycC4B4a74ygsCeO3ZrPQN+TVP/kHi5x0RcP9dmNo/fhcweEA69NWZLgAwAh9Dr
15gYPRdyUgP2mbSXM1P0pteYMRBSQ+wmPWvuwIloy7qPcjfWn4/PJOOMRApp0eoL+E7YbUg2aLdF
55n0tWswl9kHyRWqUurGzrOTGTPhHGXnAlj0wXm0fza7eqNcnBXubOz+VyMXUGTPHQUOE7I7Kx6X
ZRsdJ/0XuKY9cYfaYt0J5wvtg4v2nxL0T3bMnGXH4RImqL8cFPKcb0066O5Jdo1ssr4LXYwVOSxy
LyMvVJG+8XdcXpdqHkzlxEHcGqK71tldwU6AoFOzxwgKkFjwr+aM7UGgRIW3kdZ+q6w3H4C60/EX
zmQ7NPCGqHfCzLlnDezZREcLp+GQOBvQ/iP0F9llzowC3iE9opraU3/zqdLWomRKxyQGyX6gmpLW
z/mx/cxEexFJ6d0LQlY2miAQ9aUR8xjhmaCtgpwsxuQVwvI91X9zcRyO5XnKVZ6erA4V3uHg5608
qa9NSnNaZ0pJn2U+v5RFbN6K9EMJWS74/eds/+Zs/rdczY2RKgyIfEv+VnBV4Wr/iH2ZjrBpyoWV
2PXMj1S0qlO2aBpZE6UFz7dBc57hxO1zVFQJY4ci+MbaXjYIAvvA55XcZXuPHZaEO2OzYmoRIMC3
4TEYOhuL49on9+JOCFNqQa4bmvE8v4qMxqa9I2vMOCGIlLCKfHncgc3JyhxTqGLoYQEXkfTmDfzD
CoRjTvSkUUARscmLY7TZycNiQER4NgqoitFBWMiiISsZJibWoSMbZnDE9n6t84ROY3VypzhvIBjI
CJcMpyMOoagr9qI8CKMKdz+iGiCLwq8m+fWJru8pJ2yGngogtcKfa8RtapidE0Wuap+jffBoeq9P
/tT/s5FPaQfM9VOL49y/TAJ3hAeGkdhCUVcS9SfyEU8QjU8XhjnAPTLg8iVeKs8DgzQ1huv54DKN
wBZSb2yMWJHlVH3Rexj64LKyCbZpc2itvIkxEi9T0+/CAzHXlLtkVemijLwg6BiZXfj13jVPa1Er
e8TdFMbjJcICBsJwoyE+dWEIg1MkQ4uqk84GvIOErnWrTXKx3TUoXqWcQoD/Lk9Pvj3jxuiuvvCK
YAITG9EhWyXhkkSMxN9atIKoLwOxzAuOJdHEIBQHIYgl0nH4zrxImMb+XWIT2NNB02Yt9zQMo9eN
jVo1w1uVJT++EgU8NPfpoXttWhqKpPWSDR/I/b5yvazqdytAbp244rAFA0qo5f8/Ov27rRoqxdzS
w/3DxXv8Brj6kEnReTp+7FYSGGgCKXRt8MMWRMtiTbFQ0xG0T1yDapTK3MkUzvaWRSR0M5GHLb45
G5hocTDdKWszrK17cNfEgHTIr815OU5OakbOQboJeTxiu4Tg1Zfo1vPFjj/mj/DaVYWoyzxi//eG
c5dvmX2zWQK1v4GhSXh6v6avrhOmyHkkTtGdFbGc2D8dwsx1BBGfIRIcrY8UI66Ns1lm7km52XQt
0nv1etF73MsUoK2BPvaF5X+wIcndXsRxUJqoYKBSwql29B5JgtDoF65ia2nc+bOeSYtChZ4k9Vwb
pHTs0GFSaVwffLO3oam6Ase8VqI0byU03VZv01b+n/VUbepUUW2M5X/YRGIGOyv7Fws4wNEXjXjV
BLUtTNvBHsQZBRXz8tlvMRLxiNTH3kYYtBF6+tTLkmhm3Qdb2PUBPX6mUii5cHsqsXp81VuSt4/m
TdhDrq9yqgKa+6HHx7OJX/MEP2B8+EW41J/65msb98srksxqRdU5/ShsCO+45yKcyqsSTKBz2m5B
L4lp9Vru7bqUx4QVr33PQwUBYlfqxFLQMBhQzcBbqDD/zMNhkUfmfIV7dOmXyfWmM+K9Z8o37Pse
cGOdyysX9qB4tNmyDXheeocqfFfUuQU0moM3fNd2pP0Sd/uRnW+nQ7kb102F0t9alr0LUplBXGXK
7KBkYkBrALVQwI7IKpfCXORlxC11dEV1A5lDZntaXTA09DYIXoOltqwn87UHkBpiBGt45Z5Ky3+d
Uwz3xX7B+GOFNxIgXMWuB/+CcsP8jtfBbzywNK7veCwTb9nYn1psUYrp6N3pyz+nOUVqcMEmCOSv
Nhk4f9gECDvpD+9IzRTBH64FHIy7gQ2FsQKkXgU7gTJaSfiCw5wZzCjdGGNvvAkSoYJf54aeYjLw
I1ed8+RsDlpRbVsyi5eRYQSJOt/TPvMFmvs9HsXbibixaLqgJL6X0FlB4eWC1ZtR6KUlZQqo7GZM
7i2/CFiFP09Pz2BjRXGxvhCQhEtljGOeZQ6lLiz9bUV6qz10OnXs2hdZVKT1KjXQP2MB2XfJ+5Pc
/1Q5n5w2eZwE3UOKadu9XVTwHnTv+tY0VOm6M/FHdCORUxCVcy8+FqJGXJga3DpXgEsUSL3NqM5v
Ry+RgXlVLW3WjsaWB5+e4n5YhOdz5ByT2BuUs0T0OoyEXEFrsvNY1vT6BoBkz2/TYocoqWYfJjTu
R+3BWagaK756QF+sYgiILHJ42NiulUJMzXTtxymfFl/65P84qDNQXZOMPcAEdX4uxInCxTKQ1dkl
Shhju7T8W4AFfSVfMHHkaFv54TVH2LI6ehcFg1gX4nkxLKk5j1wU5RyKBeUeGCGazZ7rvlR1z5kE
jgMYEv8cv+kIfkp3GE+Lt0E158gDleuAUK9mczoKt+hXdT3HUgv+9wXTdYNVt7kwvSx257Z90jwz
U1MYZWh4qco9RmM8hN7+mdBvAoY0DGKSi0YopyhDTpNqLEX1aElobfn11FDlc3coVD1pdKcadU1R
mtliuBwz+zov0+Kc6luEghifMFpu7bJWvy/kUzKd7hsBALSJqNkx/Fix303W22DiM72oyGOUpZQ7
rYbJBLLwAZQRVWKTGjH8vyc8k2SB8N40qbxEJbuoo36tfRnWdDuJPws76HT7c4XcA6/FdHH/DQqn
T5SDRXFfqrHPtiKAz54g2jqpBG+NEUr6mjDMT3KXeK6ShQgvulGUSoDhhD8/UW+8vqRUmKf43NeM
eDfHnl7gRkQY5dc/5WTTmF40OYDOpKNQonVlevsOO8ggwlEakHpCqEoXJQvKNzei9F09LhvSnWic
QMjof5bTmdNYra75Sfy0pPS6eaU6Aeq4ekV0H7Wta3tKVLNbvP2rmtDgReZHzkcrr7uRPRKnGDr9
DZSWtUdik59+Ve7aEDAdFpLa6DmYgmIST/lVWc2yE3MKrJuMm8hs97zfgq6dKfYvZoNTSbBZYOSk
qDjoNTkkUV0ygwemVU7A3Uy386bJH+rbfnnk0y/P9XA8o1XKpGRp4GE+0gcN2kALTvCzBw//DNjp
XlR0ZqEcypy2z/fIMEsG8CjPVqM9k9eHCsPnF1YriVU7wXkB0Azhs0F2YkyIs1aatZdPMDO9dxwB
fihYt5oiEf7E6r3MkVLtAYPrEuz4P3nwjUeBi3wNGoiasbX91UL2tvyzSYLPj8WLJVKP70oQIji/
x0JIKW8R+5OHHx1r5mmzYM5HaO8KYNXiPAann+fNuAu152EwAdPFn8lTQk+Zl6wZW/6UAHf/rHK6
fs4lWuV3WUYmgR5ULfvnsq8arvT0a9ea2LEVpBdkqwT6jB92s+j6Xi++WO9tMNdlW1HOFXprS6Fh
5BIddVUkr3L3Zbq2YNTJ/+NlGNJoH/YTjinnB89NcigjfZ0rdBZFyj0z9Mqc20e99QK1h8MSwLaH
kNDc3mZySMmYcJnTztemhyEN2x5xmon7uKU2zG7twjcQ2QkRmFHRSZxCzZI8jWTcTDHKyLdlXfsU
pFDtyu2BXe440iZLf4dw4wU9JqamodssJw5BxLvvaQ5vmHu2fObSZfvTTpaH0hFtv9otO+67stvp
55INGBlCZzDHtj8ta8qaPSxtuzMKcPCiuyQCaOCWI7JwNRaRJ/HgYLS83anlev1OAdqXwUa9nGb6
3oE2XVLP6XrlJg04Dngog5CDeIRxXdLz8bwUp4hqoi2mpu+1HzEvI3JpxwtuSdgUquKKJv8fXBge
Ef1OEwV8Kpf+vJqfkz0oPmqaMY7L72iiXgjfjzgTb/R0SjuLIsunQILszzxf2H6NnXApQfZNXVJR
iLSz20w7Tsn7cBuD75vLozYw92YRPaxq0UpKx1OcwuZgyREHddoIIRJ885M6UeHQDduwnSInXvTo
NPT8T11gOrvR3NXsu+bAdxraAiILXVxmCVhwnF3wnySD7OGArnxNsqA2dmVvY7qbMcx+D39i/Kqm
14gApznuc3L8v7NSMtFsOtTC/876u9L3sc1bYy1tb8KR0lVaI5tZv/r28UzHRVw9u5+i70Bn+vj6
WYV7cntCcM1MVO1MSHZsc1xXoYqkAo/625fB2b8S8YS0P8SoTGS3js306rk8ianOA+u7dUw9pGnZ
nHcD9sthooWAy2xd+Q6gUBdWe+coiKwD5Sk9yucx+o7Cvf9p86/ibpf62kamw3Wph6UGFZgdQgdx
fhVuNWH6LHSa5sx+37lmzK8MUqOvSNsOg7bwwq1UF/BIMQH6OhCkV1N0uA4qBlYwrJB6P6EFBJOJ
PrlX3xcdXvUNSn0OFrH73fcI4yUAr5p5xLsP5i0VrEUaRUxS/rF7kpBIzXkPGuJH/X9fmm97X7U5
Ws1Q0UwGADzHu4MfaK/hEoX8mJGetWRorqzzPsOvZG+Y97cZ1jBWe9nOvk+mjScZy7SNkDLpnurs
zafhAqZyoNFEX0Pilx1qlkFmKhjB7zmdcJueuqipY0jiWpyJaryesnPb3TUZF6b/xnvxekN+qqnn
n0tGY8hFubGvZo+Gc1PWb0aWYm18gSID73Ft8fy5RmxAvxBaBf0vDX1/KRDe2RrKphFplEf9J/y2
smpGTeNN7p6srwVZE9eZNkOj9n4swdb2ZRJuhNtqb9V3Pqczgm7XnAcMiC5piNgBIrHppaE69Xic
cfhiOmoZ3Ulg840taMKE4Tw0L9z4GAFUlsMSo1FL6FqvETiX683mRB9sVSDpO/vTSNRotpqAPqAy
VGgP/4HOWBC2mt3KDiQ1KvC/G39P/+Hfahg7PI4rYxXSfH5eS+Zp85yFHPaLeIqDIVIxSoKwOQNy
rXLAEFtOELuo3ucGml1TQiDbJJZlgZ0/sMOfSyhPYGBVYEMOoEJvivsLY6Slrk4Y1PTsqQqSA+gU
pwsi3YMHf5ysgt1mmMt6btqxx8CTWSgKrwRpjs3hYzanCROCd46wECo5zktf9/CKHlj4IACqZZw7
H/ny9MhKknlJgabZXFErvuSH3dVH975MlkJP6JqztCNFH9n9Nk9DG/Ial/0KBt3znr4bG//cjdAm
tLfjr5FJ3dLHz/GMi//zd7TEY0/hvUqs0zUDPGyVkAGzzgMBqnhvLJyYc/ag40hxeaxNDa8JXo7m
oKi+DmF3bbLlI6jgjdkpGh/N1yDPfZMn3sHA9z6aOO2yDfirrANke6vLASpW2xU6oBvgo3c7Dfbe
9CMhq4K2QqiFul6UHiFJa1RbW9MR5sgIcpzEQBLKdAFH3sE3LuUnZqSvcxvJJxUZUO9zyTLVVrl2
YAIuZMm2qoGnGipNtiYSFNjxlPvzfwrHPinxbQ1J0dljtPNlVCJwZouO4IQhdcoJxjx0MblVGIu6
gLrfSdtIKiYyUZUE7LVcHdZSy/lO6CGSE2jp6Od78Yjyu9WcsZBSuYbX9fVqCxab/SfWhidBFCbt
49BTJ4N0pT/8HSG5pfXUwC2yWlXcIpb7qs8c6OgF8SL9rxI+19ydrifyXhYl8ZtVj4o/acej6WZY
IxTO55pRFqGPp5DUBPzv2eZKqkcMhhflIK6Si5aaTWGk5Z5FHVN4W22JXFhMWLpBVoSy0GsoTi5o
B0nzLgfj0vntwRZaPF1O1h0ZCoaLuvvBqq8YBcxupKjOlfNsBNx4h/sxcImTTKf+6hdsQyRapNNq
KNm/X6SLPiz0opG11GrPyzJU/3JBA3SZ8YOZoAhXK/ZbIjZDHAN3hZAg89WVjBZ8Ig2+MLBV/I28
kcw2wsuTGwZCtx7Xli7Tw1kKsyv0mh7uCmsjg3jLoYOu+GEA05AvbY/UvzxqrVA6pXUiWRbc86EI
3F2YgWehzlUkW+7A7NcCbYh7FiViY0+i9Y2tkWSDOKoXkq0KIOcXxZmFmEVRPiAYWN/y4eDgU7Fk
lF4ebhJXlWWnx0RqC5P9FiffT49SpIbtCzKGWas+1UNeFdKYcD3c7EnPenfo7oAZsIU0VGhAFw9k
p4/dpU4ugKnyIVGpevMdZo72v42EycUh3yVxsczWiJbxyLjSdosyLLrC/5lBb6oTHceHDuICOz0J
AI3VBfTQzWuvWWlNcaKFZnGfJN49KvaiRMDBG6/mCLFmh07SXbyXbeKmJzkgfMbiCi6Xif9yGkAb
H4YiNtb75JXuz1b5z0TQ4b62mammQyMLsJq0fSPELAH1u/CFMfkZ5hOoshYQUQb24NvQJfBQjVsr
y7klGWMKVDrNNhpTzfHyzBlLE83EWmGIXgt/WdkYVfrRiwATPnAUuqm0lwlJKsqa/unXlsi6eZyq
guYMXS5ZeGsjS8YfKao1MzQpJLUzTaXghZQMCVLbWOoZxsUac1C7apAoR//clZlsb0a1mgIWjIp/
xAfk46pTZ4VE+hncWXYjZAxBPnwgnCnA3x3S60aeEOL1R7A9+eEU3dwDFZVnIt/BwDHpowRs0kSY
Kx/QhgPxx5ypH96AR3B1TZ0a1nwK1VwOuKS+vcgik08/FJz5iDruORBZfr+qoAnqT6cIJtJ6qIX8
v06UpKKj68QtnX15tMG/scLgDqU0tpmSd/6OankScRDFDWLxXzDjZerjfNF6kXJVQFGcIUeCkQUz
4PQSWs0fOTRWsJZN3qd+MUwrDLyiSuCMsRmHQ2SmMb6qfncHMnsjlySeJE6H4QWOe+TnqckuoYdI
5Jvil+Czmstyq7E6PAO+4KwMlsDTtyslN88/NeRVY6euLS8aJ+VXO5eIMh0AsVxGRW1nwzJ7Gn+5
zLdO9pGHn9h0AeedVJvvHmePHR4QsuWPy01UqHXN3l2rfMUIEtvfOz8pKznG3gCogRguuTbKjgQT
XK6lGPVJzn5H8Ll7itlJlzWWm2yVuRs0fkiGs/+vV77HfSApdxYlhKuxK/ziAM56qMzG/l+bw0ii
Dx+rGxSxEIhjHB1BhGrA0qEmbGiMYvCvc/74fv1zuUJszFyMJF4M8E2wHsgngqOCCD+si47wX2NG
0SyEHsXU4Chz1MKCPdRSqvmBw9rezAdz1ryymkn0eMZLnSsFO6nmOuFMZg6+MKOUSd5dPWlihrVh
Xd7r4XIVbzE3mKAuZFp+UcWvOWkCOc358glW5rMQ2G5zs8GskUn44ktKYthXoMyR6zGGaTUn1g1W
N/CQIjbF8u+8aW+mI12984it5wCm5rnqVOnukrJb7DHxYQy1aZCmvvL80LdJMqzy+RzC+zr2h3nQ
QtDqxQv3jP1WjsmSuTt0/+y90qe9Zygjfpyzh1vOL/cvr44u+6ae1MdkeO83pWSG3X/CfG4yq0Im
B/4OERvGw6yh0bhP1oyVUoTk63wI8u5c/H5loEskfmNA9SOXrTGCAuTz8UvOIxYLHYuhkcWnOQTC
K3oJtVV9rzlD3aYkKHFBoh/KLN2Y4sbePH73t2cOg0Q/fjSZ84q//E2eg0nk0eyjuOpSO2oP2cKd
zozjB1EC75PbTlkWXz4VgzBW+4zC+jH7SRR6iaPom/be5t797QJLAH/+uZewMIJf6OiNvmV1uYsN
U7kdhslKf4zTK4DhBOjIf7rzepGNOfS6DEjDFzORO1grALLJUspUcs4G7gZnSGj3mhe1TpPckBpq
B3uK3w3Wu6EviQaMalCUPm1kdOSfGSlVC6FsNC8jnyYYu6Z/mqt5AP+IpP4Z9wCPmMHVZBDhknC8
DTRXE2nSM6U4BcWMgLa7qhdFFgcyfgs+tejUin7C99BrirdsUuQDW/c519QlIHErTLN8bu9pKhWC
VFpsKg6JWmINmxkAPtQMSaB+5fhKNmYqSYE3BA291BnhGsq8EZFBBoHpeGTGoA+KTdAh1NZkwkgE
Lr/0kLCGi2Ek3t+JH0KD1OVzFBG8qzJZpBsCvqXIvc6c+TTn+C5E3H0fuyKdZMvYIpMgF+MBUgMq
F8CtvaKxTlSMYnGiyFcFCFtxWM7GjQB9o2YbXjomUBEhcKvdZajTCKt7TQhEClM33xamk62uP3IT
fd7jtIcqGiND+azv6K2gLMGhtO11GvRX/x6J6fbDYj9P/6XeZfjeUxwfnsT6Gd7GrVMS2ZpzEEsw
iqoyi7ExAq6WG6PwMxQSLza9sKwvE/3tONgkQVDx7GNprYVENlqSMpi5LyMOHB0BfFmgwLC2pt98
c4uv6o+hKIg5znWaMhClcUGRJvMAvzRlG57XXhrqNQ13iqyxvg8V3wsYysmrzBRLP2jAJSP+gCY5
4vvUFbhPgmIUW7pIHfpoECl5KmfkbQoPBy7S7nvWNt3pR9EeyP2l7v8ost/8NSgnhL7aogqy4JyP
25Lt+hszrDQCAfxYutSPTxTcDXA0Zz9kiI3SfByaM8H2GXFF2COO/PheitMkKGsf/uT6NiifoefI
ogHq/7WBtNBhzRXZT0Vj+uBUb9Ehf3ICpUWqN5Ew2JrRTspEOLIugz2kVfoOcdhfFn5jbNVo2oU7
XcOknMpCaGtZ/w2wzP+dc1HKxc0xXpATvwwDCbYfJYasl+X6mNtLK8HHXH3X/nZhi2ksD/llG0aF
iDQFYlJpQVcpC19Dqp3uBSa86moJbGIHJzD08KTPtsquInxblofwnG0v5bjnKVZDSLgbmVBOzzZN
AwPjYHJR1WTllsPbSIq2M523vtcyyNWxJabNzn7BlnkiIyimzshrQ75h18C+ZteTslTHP3tFZQ+O
gVa9McuCb0ClZ/XsX6P0wf/u2d0PVkA5hL2119QHbzDWjIf3ENxcnt/uffpS/jdJ2N7Eq2y5ElP/
EKyD/uHT4N501PsKQokJVk0pb70cUh16AkNRJcAiyC5OM49TqVBTICt9JJSEztB+m3ibygEW8P9A
QJ82zvTlpdRlofBtpXX71HIYLALNy6+vy5faUidVmSLp8vxldrVifgwNpQRIZ+H/TRkTBC8cXAsS
cF2zst0A/Cl1IiXHQwksV2qS5a9BB2R+uJPK/aT2t3ixt+e3JfjVptVbB8B56heSDTvlxx6gez/6
ZrN2K469OOw1jg8DaIrti4wY3BEDtnvkNDaoXnJ5w08c6HDbeBRAYLDni4eLTZqkMxItFwyttpiw
nqISu1LB1YF+C7n8Sg0XLYtMtYSPfJfjpaJVIYfUFw3mJqJro9nwXiDGyGgsce1aLWzdcY4i7ofc
Nvcq4rGy2cRM0VSZ/7nNNR7FlcvqKU/seYROOx5urSLHLaFYpT6VSVwF/KXoy2Esbhcz2kx4VUlW
ve8AAjc5VkuYCNclXNLEYZumHdVUcFQWkYb6o4po3uRRur++Bg6gAwC+OgMnGA19jL47uuMcwOjc
kJVa81g+3w8+dGm6Yz9SdQxtzuTCqINU5fde8PxiK34tp6+9pA5avaeYn6+t9MhUTnHf4+OgpL+2
gFqnuN+Ess8FERHjR4OVEHTxeLK9TBc87BwTzFn2lwX1+db4Stm23FTSyqmxAmuYWO+2rP9oPV9N
O+1qTM2cJJl2XZmtDNfXWQqGZN0pvvUegdB9mVAdWfiOE3AB9fLPJhUUyf4FdNA0xN2zDJ4Glzd3
5em0M2jrgjQgDowqzAbGdCv5vx7t2MXQ9ETjWO9z7bHhct0gbU85iaB0JQTRTL3WCiZiQ/wA0lEc
5C7oWtVYlUkNoHlN3VMOsvXkFE6RHHilDCnMBeOGpOvtpbHKccIxv3oMl4oTkL6lQLUNOPk1DWgm
s4/hptjrvMeJ5f+zpgH03x+BdyK9pKhGsXNoFmw8D3ErXdvYI3w9o+WJgl5Z7fQMsWv5fFBu20zV
GwYM/TeEaAC4to2PPGOOS3M4rzTZM49NHfY4eYBYuaNRVrreNA0lOOB4vkdFDk55yy9QpoY3mkhP
9oPfQd7VnRJbAgZNB4VQP5DBxOKEW0cretSWIE4VUVUCE8F/j76+45ySmvDqquFaBpa9FNqjTKfR
s1Yh/yVB7fDcP6tA0812TQ+Oh2oGBMq/hZ04kG3ESm1P8jDRTfM2QGYI+rZsehPMBqMa4/K6O/fE
ORWRbcd6m+M2P4AlZHVY7F1Z8su4upCJ3GauxEFi2EXI9M2wLklo4FBhkj+DwnEEAPSYerIGaiys
p6N4A1o0ppoo8xEtZu1wSdWAtPhZYIYVvMljl8q6rYjf0zxewQQC+S6sRuhykHEsdspcRjr2Dreq
k1lwxxn381aK4Wf2tFojvBeLlNSsGYbSy+WoYK7yWNmX0xSPfYbHA7xxCCn9rDuygeg2lyp9pUC0
4GqIb7Sckkz0TENJY6SQSXgGYmsw3dRpiDYe3VQN/zogoUZwJ347BKKOd6Lq9QtqIZLTJ6nZKjk2
0zkAGdDrexV5p0xwQbOzkUdSk4lnGs2pPZYqwkDqcplGdf9IgAREhmtMqlQjmRTwABoLrcCGXyPw
zPpbZ+8AYb9/eQWjDoVzMnBvikPhEnY7IMxqL/Y1FslOW/hUaq4N2dUO9M7Izwd1xco4WR5EnDmb
sXM8+3syGx5ybn/lNCP/NjyhOmgiOFou7x56b2Az0pNHHYNxJrWefaiYeN0OpmYivUVRkLR+UtUW
dhEVBKF+LPq3jzddq8VcSwg08DNxgIm/WlcWeFwCdSfEKww2wKIWw3vRg8/VbsByXUac3naQrMLM
n9vUZMg5OUr5i69KGF7Rn6y7k+zgfnM1GgnDZ4rM1kuzSmpd3uIMhoXTznPfPYGeXryKxOEPTGNb
tpZGqu7QVwWJo2QDEGvzSe9qRTiYtE4m4r5F2FQBumtOagn5oziOp00Xp+z/H68oIsESKp7hk/Vy
tbiEZau7PSZKjKHpuXYg5sFbYY5Sc+BZSz5G19Edy058o5nJDMdJuhdZZN6NSJbQxOoSwgPZz5vm
BBUJr6JcBwUMfLd9KCs8e9NBTOJcZaduUVrLAoGkjAc4xdhMe6FKVa1MDeoeNvdoAMJVIBI98vx4
XMkrjtmRJOcz4j8fw+CISuPk1bxjhgVEFM8PTh5L6Cybg3kqUvjyD9NX68tSfhjZ5RKm4XfC4jVt
lXQRBCoAB/8X7HyHPVjZiHlphMlCvkHTm9nMPA1f3AKks0XV3tsQGddqUJe+iYOT3sa82JiKbfvI
5tScSGrUDb4gybQrPHLK7cr6Kyr4QlSZAwOCAExlo4EnNqhJBZq9N1mO77ZHeGlmA9gw2h2v8sep
4nWiuL1sF0PuWYDhs4ZHtm7bVxXbfo27na0Hi5n/9p6YqeW6BwC1pXw1IHXXNKRhRlGdz994VdGU
ccLDEBUbrAffxi/v07ZlWRxv4/8paSrdrXAxszau8NgGG2T1y5bVUzkGeRWwir1iDNc3aPcB2kAk
tHT7mBKSt82VWqzA0p+6iEhalmZW/EgnC0hgzwegIAi39wdVw4kgFoy0KZARq9HJF+hAmLlH2fAX
+E2T46PjVgigyIslK8UcXy7BfvH1QidHD/FeP5ybfHZLCbdGhw5JNBaj4DeG+b6RukMahYd0tA+4
aMwIOgKaRmjNIBWxbEn4xjXBvZlTj8VcbLHw3Q6aEJInjIKji67F4uVADOIUgMbmc4uuc0egZBfL
P/1ZM14StZHxaydaLGFNPzBdQ5OGG9Ouo7IuU0LT9gZWeGX7QcBwPI7XpJ8FYg1sI2+LmoQQWQsi
OTYHSzLp0XCnRXWwBxJ1x4xNBZGkOuxVpSZPot9SaquDNI7lT6ZfWteZYvwWcOSBQTS5eKm9WiaQ
NeSqeCz4Eh9URwMxdZ5H3z5smQtq7wDyn9x8OfDqWadJat39x5On59DArv5hXccvmtgCcC0R2kIc
qDCexA4dbpaq8QxToS2TZzm/4i2OExv257uvRMGIizgkzC6MagCP/SsE4g6uatWdV11aD9ulOumT
2+BtA+D5UsEd6h4/1Ovlp/P6beQYel5DUAfpz8GJhsAUIYwkHmGvJWr84CVPjznCCkDpUfYtsN+V
ERuwZkCchbYIrlBBGzP/vBpTbaaM0ycfNsqI3Q7eIgNlg9nLhhztkReFkiVmCwLWh4a9dxBLXO+A
/F+4742kVcQeY6N8k3n1HL53xB6Z05Cg3RH3orX8tkBaGYcE78OUYR/TL1CUO56H+WQy0hz6pzhf
S0iA7GEVzjiKKgTSdvoKBJTrfl7QrsEKArw7RpuxcBwThRJCgvtOyaHjCaoYB67yw1HoDRJ1LCVo
zeNAIAkJ6WyjjDJBLQzcWvimTTh3ZrmFcNgevmFP6SeWd9I4vWSP8dAPw6ixs1/uJUEpKmLCOZOe
34sWgTrO+KuwbM8YLnl8oy1E8heVi1ol/9tNBuQmD8Yf0IyFWV8KrlwamOArEZW4XUFSnSDCIb7H
bsuVWzhzV1SAUy4wiDxJzIWy7ixcpt2qJOynKITjRY6Y/7UzwDp3HjFm67dNPAyfb5dbWeKX6YFV
2AAUmpcIMtyAbfuXA8szRe6S9070x2ViqRfuXZHM7vUFZsr96e1405bwN+XoTDs4PvurtToKDQvK
H0U9R3fkF3l5b7pdxYi8OX4t2fSaFlKkCUsDoUwVkOLyM2tXWtJQKAuduufcjw1y5jGfPw1JuEUd
p3KAAON4mTOo2S0u2Z2xH5/WiWgMhhjRGPRRpJcBln8LuniCUyyZ7m2b8A3XvBXUDj636npwxaY+
DsVT0YXuRc1JDfgD+XWf/MrPQPLmfMSA48BMms4qXZbNnjlo2YGJvamxplHaK0W4DpDYssnT5K0a
8ejjRl6y5TtVbzSRaGDcjg2XXRXwJxkJKXqV5ivwZtovnR2sJscNr8h2Klxk2vCs6jzDVGdEtOvV
qAssmSu9EDEi+gBNqHGLGz1p8p8M6OOyvgRlcX3oQLYe6CFIg6wvvVBb2cNa4JLpH9+5vNvG/uGd
ptQEthrNPNGpEeNqb5mQId7thWVk7xvN0hSHf/d3XeTFnyxDed/xPBJ6JMcCZM7oQZ/1GXyRDNUX
3zMDaC4k9w6i4cE8dGSeA7DVNW4FCsAdqIhMC3oLWb6jjIDRoQ/lF6XnmWEPahA0+5oT9763/QFl
cDzzmakIyay9xYYsTWPBmbKjHg56NNc0OxtIIJELi71jDD0o1BzTlRlvbp9ycdTew30Q4MnJ/KyE
FljqPFp6YxY+Lt0ui5K4Tr3bXWiYBu5r4eg4lqt4XrkAcj2aMDwzMgBWjqC3O4PfD9sU4utSFqkJ
PjPWutsLMlhErSWtlRx33sSAl/xYly1iceTRJn2wVXOSSfxnw2ePMFf1jj3Kn+xQ3NfTXaFR4n+7
71YcwwpCMp19NrGRXu09iFue4V9jMa4ERsQQw/cfKWQeKkIdFUtcWxz2J0j9GUCB6SuzgrLLLuZr
NRqLH2Mh/Aw5/vzh/PO83QIZ6zFd+S6Q0bY+kOd3Voc+h3oO2tx8rZAiz5zJ7p9oBJJ2LTZnmZVp
nHESEMsigFC4N5d1go6ah3EH7wFZmh2j8L+9LH4a56a3QCZ3oNoSsluzmIeifOohmL86HIfeeeZZ
rsHj+0welWVjg3gJhYqAPRjzxK3Mfn/dO/qkgThZk/aQwkjQeONbl0ISTEnxeTiVwTAgv3rgAVYd
YtPFYBZsIDxFigrvPMmM7AiDAyxVUzAt8VRbY/VnoNo8qFnk49tAgNqqO+IFbYuljF+/k64ixNzz
SQ4Dko9NQuGIPdIccAovIQ3iZPK40jgWYtOKfJRVPhlpkJsIvEzLsfjW9S0QIoWlqzhwpmHyRB1z
1vksQ5tHrVs2u1L0vFjLvkpVmT16W2wcMHQfHE7beCLI536FNYjJW13By2zSntEPvRSPcot7gxFg
1Jz7/ZuHXDVLEu5orGcld5+NYEunkNCPVQgkEusYl68O5ywxqLejTU3OPsl1ZdnW2CaieWm4CdyT
qUwqEpSa3FmkgawTLvD3vWsHFIIJTq/sAQ68bq51k/tgZ6/Rs59OBog3sq7wI3jjPBv7PwAFqRn0
0V1dKWx4QS7qucP5w7Br0/WDFtB07UZWpjYwl9Q7Pg4M+WJGWVOXaQwZDXGt1ELYOlUhPiD+X2m9
pLcWqdXHvaP8uCxC423Z8YtINdC35dnG67Vw9IV0c3NDL482M7vXKMPlNHFUjsGTYsRQf854d3Qv
MGcmy+As/0uY+WyAhEMETg+dslQHhgHI8tbJcsS1kZBGQAQl9fEmTooLuedbn/INGczjO6+TC5nL
WpeIBEwOxUQ6fwaPllfaFr1fnMF+x5N1APrxZq+3k+WCHl68zjtdv0MInZaY0mMq+Z8JBL0+h9II
zbzjnf2O2AqXkk867MeLyuP8DI4fIBQQ2oawBzU6xk1sm9l1CqB4Kf0l517vk5TRYqSOxnic7taj
9MH3BNKD6qz/tINiNJr/cNzvLyim1STgAp3usgfjX2j/PwU3uEfabRiLmE1F0RckRT3GPkC9G5UJ
DZMadConPXf3fUbO7AvHUieJngom1uB4KlBNYfGXF2moF6gHvxn+7WZA++8hYncxRin5bzISk8E7
tC/AebqmurygamoJTpny9UOmQqby18U8KgS7UVD0TkA8tSOxwmP3YV/pAqENAcnimUf7PifjQD8b
bgaqoIBQ7vD0I2xydZ5x5AD5VitCUrk5BssNdJCiSO6S0hM5O/n2l6AU0PQGxK9lPEjKEFFnRuZg
qG6PiU2+cmViu0zXmWzjCD9/X8bAvBWN/CGiwNf0+4gRFF/be4ajPwKUbGdtw0Ca9ccUcNqbSS40
qBHeEz5m74XjEWP61ivjvO6xozOa0MgQ5/XTdrs/0CZMDyQjDp4t2vKTkVBiBhtwSmeJoi2dRX1z
54L/i5hK8/VnnAuKbVbOLNMrvYgT+3NVEI4xisR2ity1ijwGobtO96n20IdxdPKFXUqMq1t3OPL5
WbV5e/+W6O6c8cI61XFobcwBJMaiYHCv7fxQvqr9drx2fTAz2cPVMS9RS2hm+rAV0zmiH3m7a//x
22qln8XREhJCAG3KamQX3PXm4+hr/no4UU96/zWsZQQuUPESrkpmCWScRbYu6QV78ut6ckdEiSoo
E2yKzc7+Mz3WtsLWboT2IGn64a9iHqP2DaMGFEbMfnMBIS5Z82/o1U8JTtpKoy8pJKDxVhbYRHEr
1P4VHN5p2MnZQAPjP6wgAsBWiYWE19+Rdelt2IffAHKoSjSHauFcQZW235KoARfacSEyzRDQdNCS
2pXAk1jIBSxCjN/fLV5irEusUkAcs87B/H+qEpZWqjbexgcYON3n4wwVd+5pr4Jt8BtYgpuNBHKP
2E6tVGkNyX/31P6WLuaSzwZk5hbs1pVf6ryjFCGVf+xZkAcoybUae0S9PXw0a8qwZO5PbggQt4b6
oVoJuJgqGx3M8s77zzw94GC6sJMUWll6h8uBkH2+PuZislHZzTeLUh3fwpocB3MWBr9WbmJdXrHg
DMQP0HyV0VbsIM95lwsba0YJglJSV9BfZV0YPJC5/nyahlUAtbsnpeeGCGBXj0R0tlTQi4V+Odc2
Lthem3AseiXQp+BR4KvTw+glq+GHlH1hTZxyk00buYWtArQy7Csxc3iNzBX3hUggcu6N4qSZuDQT
mBSPX/MEZO4d1pwRccYiScs3OicnVvnl1AdQX/tcJMLTelT0StRv/8JEcX/w6EvEfCBidoTyeVnJ
bkJPr3ieQ3xsKE6XpICEQI9LwU4z6eVOi1cgMXmBAR3xuHsuOy6FEL0Uu4mSjtuoJ2m8+J0eJQgi
HQFMaEjHah2pbIfwO25DtTewkDtJda5ZtLNFmYBvy8zwjvFouG70qDx/Pdoha2tEcem1ndce4yTj
n+a9wR2DjVfmk6N/U0pTSsfdh89MAIFG8qI9K64mzDWMsGlL3PaQbFUF1TVDqzfY+bCGE2bYEGnO
Gojj1P68n9DpEPaYHkkYFd9g7gMG0m4Z9e+gEdfWbPxK/wPjg54DCxHtMQYq7DNxPNKEC9NmTyoY
S/dP9LAGeyPxcFosWbQnuFvcTW2HkRd+opYzY5rhMaFq/HjDTzNxgpkH4h+blhQd4UswPRPbeBTv
AnTQJhFwEm7RHVsh/6Nmp/I43mOWKB6ZV9hSVsJrHQYNBAXNxJbYMInJ38cYBsGx2tpZLQHvnAuB
DXFMN56+cZ+uPlXXrGmofxXHVK0JpxXBBtkGDKIcSHSlVJG/atopRpD5rxSmQzlyF0ezFnfYvq3C
/7wnAAyDjXKwPwJpzwq1DZ3nBGH9UH04FrckEPBawXbGVREdKiEspRi0mavSP42ctoEdN3u/jpXq
PbR5n7X0i5o1HxApKau3th3Tv3r3Co6OoRjDW0L39IRpjfrZpH46LgaEQdVj8PKVacHRkzrGZ/xd
ud6EIwBuWn9mWuZoWbFFx2OcFoXxOF79VEBmqZzU43B7rMuDrhGg6wxFvSZAu0Lktei6xqk7USJ0
V7hOr+HefiSUgSrbdVwz6EddEEjHupHFdFCOHcrHHGAV7R87TvPvdo35CqwBx8KMd2c47Qy0Xj5N
7m+Zic5v3k8jM4sS5kLedzm7cd22eKgV8gGlDV7UiGdsPS7ryrTRzp2k2t2Vz859xbZqM4u9wZoF
JGSUFPp/SkUDqFz7esWNAt/zTK5bL/GTBaIh/M6bsXWKaUWj/4dyxLijTB9/6TrPsU+krnanqltk
PVhfBJJc1osWWx3f1wsd21u0c07yyWje3K1btGSD6gWCMwUrkRBfd0rHgJEdmcigywwIIHCOJQwM
VjTvAGXP7SdUNDNwL2slJY+E2z4WQK7QV9YbDkUporDagPwlZYCVnKBsX8SXu1kTVOnEmJHD5m2j
M8JQnUnnvjHscMyjMu8J0k0+fK5Dx+DX1Tf+ROnCMa11TxQiZUounLOk1jrit4Z0NIs3RcNSA1n3
u10B4lmASxyv3/Oz/OXwVvyfcpTLA8IlNArC2egsvwAE5mvJ+eqErGVfToDk95DBC+BKupMg4uJ2
z0qDa07cDKq780J8zubBUxKlLTYUBtD6YSiKhLdGKrxcouAVx6ZlpvtfEsSKqWz6mIp2AzOkgBvk
nGOtdj05yTTu582cjEw4ypH2kTzoiPHMYk0kmE/V+P/4f9EZfPpxDiVt5S3c5qzj9Q/Rr7cAUxAx
Tfw+VRdRfT5rIHm1Uvq2ngGRIYdZoHhZvJ48NJ16E8Gz88ZqWGhjNp8LnAK/jywVbZ6dYAAxVH5+
37G57z5fZPNa1UsLaMoiQOibd9DuQnXAoKkzxXTIWkewcbTbIvgvDECMIUsu3alpMiOTdQgiGRtn
g8b3JVUaOjT/nmFuHx5e0m1OUIEyA4U2VGFJy3X6Ow4IEsERi93oZZ6hkqgTKVhg2HfyXL4B80WR
/rvKYM4ElOc/3h5j0IPViJn+AZxTtGCSotiVDutq2zTTMM6NNqvxNXU966P7MSUVsRvcRhJzNww6
xh35zSq9xZXKW6LDvqAK/xZE7nz2ZUvuLdAlKzn0M2hAjoOfeAtjwY297QF+qOBkXwEvrqxcuS/s
758i3aEvwu5u9/vCyDw0PV16HKUCqlvP9EuxS756sQmzVtj/xqAy9aIxHQ9x32jAhIhCtVsOSRDH
ybUZkU3BFVBK6vNS/kq6adfVXHGJuZ89iXHdLqRaIbqMcjbFdGSLdJhsBmx8uAN3orqfcF2roR3M
L6r99xwNAObKbdsHEVNSKvUod58VU42cjuuRrxBR3cQdVfN80b3VhdxMWvHYswkw7w+EvF8HEAa0
92GPlQZHF7rVyez+1iqmbFGMEwxiV3KUOc99O+6au6OgmuIeWy1FkZK8Gc7PckUbB9lTOVm3KeaY
tDHJHvz5PsLSGClOUyqOOBqrB3Ym6XccLUfW5xFLgJD/3uux3uptqgHaVNewvdqEDkPGakJkqSjM
q2C1Q3xus9TW0wLBx2hCtnATIbG8uwKFzAa4zWe1Gky/HQUFL/fypC5Tj+aGropKtK4pUTzEuIn5
vJc8PnPOlam8Zng9BE6s6IMej0iywPDV2/VADkw5PJ5FdcfoMMu+yRCv4Wm+9N3TkSfxWbdK2AD5
VvTe90mXuq5SihWRZYsNwiF5/mUuFp3mFq9qi7sN/doGIKGhkySWbVLaiJB2aDVwC7pLpvKPYhFv
pXvZeFBwdCctaUSENBa7JcBOrBaAlisp8mPHPYD7CjXjT62I9MqTkkz3kQO10bQZEVBPtxYJu5IB
N33XmZe76jmz5walWfmK/3i3GCbVMptT2arZuG3HjR5inKLFtzyoRfaYV3IeUN1kJX6iqWrcYCCs
fudCptqF25Po70rjxjA/quN2A6K1+h4202IX2/quOiJNo0BbzqFZkORcodkfuTKD5icZDnhR55/P
gHP/dpKPalb/7x9DN+g8HjGSETARTs1qXJuaIJhaMkNza1ZL+qbuOT23ZWuXr2Yjsau1Rk1hdy6X
srpyKjSBq7ThJHpJntqzm/slAOsyoG6GfFgggWH4bPYKWKJ1UJdME/vq3utuNLnTEdHWCzsSmqcl
75rCi/ZACmwTMVoOa+SjGweuQK4S9cfkbg1k6PmS2FztJp0CtTow2Kib92+x/Fn9Elr6q41KJ80s
VVj/jzjkJ23fL5I6LUdBTKW6d1XMKW9riJTBMhNze6valTZubFEqoZ0CvMOQuCRMDz4xEKqZ3/uR
5LVqBy0popuB3Ft9kbNEzScm5Aed3sGyMwkt6Kki5ou5PyBVOndCt7BrPetP49hywZtkUKgUnw2G
oap3nXVXb0C3vqn8c80uowaZy6rHJDTystNtn4PkYMj+9r0EWHDy4cDIGzS6Ldd1qCbJW1KL3V9L
BuuUeNKn1bKQwilhhEdGPcMHy0VQy77aQf2xN0pFGvizgHnlCxe9znbgYIZsygo8C6761jssr7yD
5kI9kp9XCAdoxoIDNRSL8KHBt62USXWb0BBt6aYm+3AMAsXMb8qEJa+Nci4ytpugN4XNgWmFDGB+
C3PAmDrbW0ev44Ov6P9csTjZD3tC0l+FJt+GbXdEWaUgfy2Dd0aOr07a4bhPFuFEMv2k7tmOarDT
bcRvtlZDVyX90IPI7qSGjNSbDveC2sxe5y3lxSAbOGTy6izftCAnDA7bZWXoPS8gkTbZhuonSfNw
pS5m7keIKNJW2cwSclfzkgOiGp6/X3N9kKVGPKDJXE0VCReAtGHdqa65QpoxjYolIuoZ8VrwQCMb
pIDN6CUn4W4VzW7dtgwBC8wg1+TT4UM3PGLPMks0K/MAGbfL+tprbLrXkabHup6Dre7ie4BvUFeL
3QJfQH2tN/8Gkx2gvZeHlgVhvudPIFXrdRxwrqUOZFFMdp0T7aLRnmBwnAGpIW8wHBzt+M1UFt+Z
MkUezkxyIXNM97J2LS0Px5xFZA9DbS82naUxEitFbxPzu9roh0GTgijJ/5V2P+gtnwgihX7FFgc+
30/DYqCdryv8sdg3aFfaTsyw9l/lWDdbjJjHBMPWjN7CN5EF2IhXaKMSk7GtaXcxRYsCoKcS6NkX
scIJ64pEQHZtZjSfVyKMvW8qgpfRkIyAUbM/Ji2H4KIPf9TA6XvIzzyKEh3MGPsv4ygqbTPR6fZc
FRl0xks+B2RruAgcBYIaqF10Xjxzkg/UGOfAQ+gjDXcXjlJxzCa+5Pd0GOIOfTTuc98hqfcn3ZtP
ehX6d3doM6xr4/Tg0l8fLlAzUg6Qaz/4geT+FptcrHrCLxaqQoilBArtzZRQyeBYprxS9yZVkshk
By/1VTMYAfiFjbcQ6S19t/QnN+yf5HCQi4/ubGsIpxkp1PEq5Xjn1XsAPw9VGs7nPLz8SIqQP1CP
NJ6cS9PXi4ueVqovN9ejvza9zOLwbTaMaHbvujOeZ6mwvjPiIuBK3jjZ1vHL9E0ICBtW0k6p+e/8
dtQJZl4AKKpFK/ldhkDwtVk82OnK3zMZTeQwjDOJk2w7nY+BPRNXIT3/JFOpuhKErcoCOYXwhnWL
NljdHfjk4rDftpi8qm+nV1LLTJBGNFIHXy0pCazndyOtrBpMYpREgIQ4WieZKtKfWRjpi1DmyRZu
TDMqxTUNCrIIMzNrJ51EjO3jQQETLfEqCA3IMTwFYgwsaYhqmsCaSShXNQHWh+66PR2bmBqfvYVu
wQdPzq5uSZ8ilzImOburd1VpNRwikq8dJZUAKeCShYhOlL7Rt/6G2jXyNQdIcs63GRtH7JB8nfX7
9lYlm66nA3OtyyuAH58DKtApiK/B4QogOHrk/r0zUtfaXpGITqQZdllSCIUbj8BjW/fRWQjq8AzG
7ibO5E7+DOUSOVOSQ0bTl9YaZgpt/VSY4VMOOzNxkI0B+uyO7ZM/5XkTJoWTzIKgrrptAKmW5V3k
zKaOiQeNVFLdiSQAbAmrqSDUEKQmzDO6xNuwbwt74A094pCTREKGzU/a/TSOXz/nRD8w1QXo8FLk
rE06d1O2Tm4LvWrt4gMDdHCOrhUQYZchIaWinGKZPiUXhQ944/1SwIVe8NuvC+xBPy6b+9nTDJSc
DsHdhU68N4//7xZ15zcOnoTf/+DpLFGpYO2Fv9tdQAuwzs4WCd2yWrwd3MgJU5zRHxuuYGHQUMog
JmVXTzZZ9pxNJ6Y1+9GJlmqMR/2m2sikkP12v3LURzdbJYZPC5WwljNbSX6Z+TrQj7DpALj3MRmD
2OjwCCSwHvbthBaysSysys9so5ecEj6J2Ld3cIT6TvcVegx+ay7tc6yzhlE85SI6GsxsqqRmqDV+
5r1kSr39P+pz2qM4GdjBkpMF9N3fihZe1HnXTl3Njbt0yM4B8uLjxi15oVdl/U5KthMgOFo9LTHc
r1IxDRYfeiYrrZJtUIOwcDkF2RbVqHy17RED2qZys2KlWW4jXQhkQQTvejZJlXaD3aSHkJ+5A2v4
UPdfbSPNb0meO7EsdjJ0J8SROVwvqL8KN9m5Opgjr1Ij9kOc9DmR++VDtlYuzPYGECFg7rXbu9qs
L5pgaLOU2pWg/SO3h6cs9uHpaBKUDgwrMrBnHLsZje+VJgs5hMyJfJhj3mQ4uS1LwtUN1Zo2u5L0
apQ1ej+VhiiWZKJiomauqpI3imtLOaGMZNWoHkUEynBgsS/7YTOxLWQ+x4u3yytXCVvWkWUynwdB
3dt65A+JCrrnNKcrMPPVNSNyA/keioyXGJBTeAjBJbjhAkku96t/raS88o1nBpG/ZciJqpZx3xwr
86v4c6hJG3KUkbR8DHZeSXh5Ec+4YO83paA6DKGpeM8W4aTjIVMaD6CjUsKydc4H8RCFJw+8cY8n
lAoPb2R6MduHS5U9Wt1vhIF9PBe4yrZZLfQUlBwaogc1xkvQvR3lm76Cs3xMZbCYfuIvXIqLGp0i
JWFXlLUagLnam4yTpR0dhOoBtLByFhQGFCBcterUy8Qw5TBXvuhjtDvbq57tZVeGgZ3T7OHa8k3V
w+CtYEBqNvsA2WdckAHdSy550FvJC6sPyXy7NGv6y9SuZoIpnpp7vlboIOErLqQ3eI8xQCKP9XRo
YycXPoMfdq03ZR3iymFW8WL1JeLo6PuOon56IAKH6yovf2Yt5M27Mm9l8Fyw6ysJAZGTtxKdT648
5fesXp/5SUd4ZLxlkcjkzIs0O8vLJbb7F5ZknxSUWo3WuK99RtDlT4pKTqZrCEeFKgKY1b7d7JXz
YTCKn8DZLuaGGnvQBLPsz0HF522IU8Sy5An9SO8TfEpYkzdfze+yPxigmdAwo1MpaQ6BaahqqKXV
V4tbAMyBT0YknryE408ZE1haaIFpNm4XAXD/7LuTPrcDgBvC+At1wqDOcxVQmLZOOK8nNyhG4GRO
GTLdnt2n0Zr9XEYPCAbkgwtKvEOZDESbDzUBaLnTrjPOuFWbe8pX7q40nNsIwEEAyYkWBOGPe7j4
HM1rycWKPneMUdpcKWar/AhMwd2TgEHCwJnMkqVszeDn/eFoPJOFQIT5CzO8gaGp57XK0Qdl7GXG
hHLZ23Fv3uo+fYxJaquZB26bbH8Yh7uziLzGEL+LFUkEwceIlX7H4F8uqB0tAEsY9n1AhOKr3tiB
YsbbNiNuVkHnmwiWaTysxww2HKZWlodeF6nOjmjc51nk/S2nUtpymr8KREfZ8ZuDe1bwcEv44/do
5ZLZePEN7gOxkKLQhWQfQKH0gfNFFwQHJzenXRU+VsCLi1g+Om19Ynit6EIJyCZvX2+Xllz28Zh2
YOsoBqEsJeTNXPmJ+LAgZijfDqgeHrpbip/vHoQW3G49x+c0u8RVVgzMjNThVhjDr0xkU6ELBTUc
KB6YNkGBBuxaGAWyEt8TX/hWFK1c2xQvI8KfcNYy5LBmOmaTq+Cy2a/h37DhbfE2ahxyfEO0+v4l
ghPrYFkg6jFuLlGCRqbxLZHRjf6H7zhrYorxjHN8YWgDdSXhbjA5M7bZ/1K91wlcGHxfk8ZlVqtL
NULLVohlnCIKkqhHY6sUu3zZ5WfvYt3DBAgpY4r7NIJFJuysvgg57gg3U/jUyBhuk3MRTkKGEn6j
lORkqSdw9wLidRggsPIxtoEUg7Zns7Xe4UYVcGfXt0kw+V5mPC7GlesYzBvitNZX1JdNpymXyrIj
/YjHN3/hTaP9m3zpL3dlVIH4J0DkXOVll7gRtOnuXJeSw/NcUnQhKoVeykqhfvlREmxProfqryT3
lftwmvCTTGCpNjK1DdsY11gl5ows/wG4CjoDWmm6mSgBp3MEgSXGlQXYyenrn8BIO2fyKj1uQgO3
lkuJxoWYDy8bLaTJcf9l2OEkschXOl3vuEhKQinwgMHmd3xE5EOsm/v7P+WUqem+SBJQGhaM/ViP
B3ZYpFjGojxwnG9R7KhqGvffB1Y974c++W/kQgbSsuKQc7GrBbSj2aq+6izA7gGH21i+WvLx8DmU
JJQIG6p8V0iUzTuGDJi3cu6+dxmiSKJ/IvGxZRr0TCoDYglBuIzNQR582mMZcQmPQ4A4bgxXIAuZ
St5xDWGPX7wUtzzo+dCoZYt5ogU8duqhggDrxsu9YA6Gh88BZi1bWyZvZc2MaI7LB4AhKvWPW+U7
fSuZM7sEuzOUXxDkZCbcLkGaXClP45UUVMhpIXMmggqAPIIIlE37RRMLg54yZavPO0svCXfTF+UH
zqAhIJmo/cLK/oM/GP1uUf/cBTB9divQE0HcIQA1iR0YvzfNHhkg0t881wiGCee/h/35Gxd/4qPP
NuixwhKdQXwM4dPauD6NEdozek0Y98xqgnSfk2NuNB8dlG5Jh99stoRY56125uZZbG5Ug2F3bP17
QXPg7dxuLyVCPjlHgsDX1S6qbSfaCBGvzHx9c9DL/CWznbQNPyWcxH7gxZeNYgLOm0kkcPs8plh2
vFLGjOLQzw8FQ2Jrd80Rbh2dR4SFe8CoLfLpyND3juyDoFgiN72IeStwcJT4zdtFIVcrZyXZRoA+
JhasZxp/ohv9NaYdoSoQSLvj1swSKmO/y+OptIVudSIPLzFPpGSeuCaOnz0Oy9o/sHmGzloeFgtS
D0XszeVmFURM/WLIJb4APOfAwqAbIVuFkVsmHityp67BYxCjk3FDOZvQ+SA9rxig8P8nWeHXNmwk
evs+Hx/53Nk6BS1bTpdG3JECZxqNbJ0j8gng80kUhUQN7RB2ny7/9xE2bgSXYVoGGiEeqmUThFaq
kNXp8Nb9oRYAgymCo7eWft06eO8T8v3ZzVb6J0vUOK5ansC5z5o+m+A9yRLF+h/ETUBmwp2fO2GP
w5/RqixhVVC/dtwEJkIgPExg9NQJqxcTT85miKGUk5diVEI/8WzBH/RAThKFhKfN6XwmxCVE7Csl
vPhyoKOIbFBBJRtDEe9z8su/g3auAYLbtz49ktshrWKxkwwrUz9GsbbSLdBwL/VPmI8KRtmxeLBM
UFWX7dgB9ma7r2sUG4Se6hNyvZuNlKDFVUtHI6XE8ZSQKIorNF+m+y8m+7FPrTNdG62HWQAhmlOh
rhTLJ3XuT+1/TJs1/Q1BGT2D4Jn+bHR+qQwmUwUM9/usdowEi8O25ZCv3y0BbPQ3qBsnFIuZVsvf
y5ENaZjmojOqFvOhmNyeNR4Hup+hon85Z3szDMbxHvHe7z9qbAkleN54RE4MalwtxdzHh0QfFBm3
U+emivWOzNJ9XEjFF2zfYUhrKIMqG/7+4y2XzptVUPcbe0dA7ElFym2YwP6LNoinMi9H61QOeE3E
nH47DqkCJwh12Omlgy0KBe6RrslRRZkcBjUaHftEqYan1PIO8TZEVcp2F3G+llFJvb5QxkZzviOy
QzK0EniwkdqKbOq7mRcEBkDhcxSJV9TSp0kBdHzCorMx0NNw5f9BPfv7sLmduwrqFnLgGH52sY7L
5Oz/y4BiQ9a0eYDSfci2r8fm8ESYAiuue2awsiiYLSM8A18Ig+KJ/oaNAvnukBggI7hiOBCWP+yv
vrRg6sYt7Eruokfcj9F0hWdBHP1LRx8K2fzB9tVOd1g6ycaI758rnlHLGDo1hfpDcp7xzG/h+vUl
/+m7tIJGmuepViD/ZxPKMZLKQMEQLQ6VIWhRAChZAbEiWzxvI9auWWOJ5PBumXBTXK68Kp5Ctzq5
f4Omz/0qD5shYWDMFln+0rVjcltBxBxYjHPZmPWfkYT1dKijB1DyXNtFO1/6HiP36qNiTICShtPS
w6xzQgRC/KAKOjvd/cSRF1XimjTmTmjiIkrgt1AcIaaybu6PGcW/rZOq4soYcdeK
`protect end_protected
