��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�KiM{͗k穩)j�k���G^j�^lb��0���q�ޚ��	��0�
Yzb�
=+7���^�Ƃa�?��:Y���G5w�њ\3��-�
S��Uw6x��k���K�Xck�\뒨g��Z�!8�/39V_����w^�L΢���f�ƾҜJHv��c���H.��P�_�W&��G	Bq�Z�?��
2�xL�L�x����셄ZA5�K�j˻ m%hh��ǌ!����r�;Ou�L��Ƌ���sn��8����n�#�J(�B�V��´B���������������%�gn"E1tf/�s��BGM�"ט�40�7:�J.�>�F����S?_P���.����{�-�W#-뱙%�����~2t�Es:ɞ�*N�]q0�3y�d|�
�E�� ��}�芻�$P�������.iԾ���#C�HS��y7t�8P��Ҏ`R�D���ާ�f���-��M"���aK`��\H�Y� ˥.���ƗYC����$|��H��%�3T;�����*E$~�L�d�b�g�e����ɾ�C�'b��_;_�$�f6���A��L�P(td�p=e���(b�?ǖ�y���f��Ȯς�X؏4.U��� g�`q��'���!�Mr!a0j��0E|�POr�rҘ�	'���kǒ9��2K�qf!��A���cկx�'ǳ���9T�L��kv&m`9����n$�f^��qs�;6�|>
%N�L���	�ͮ*�])��@�\h�����p�C�7�p�n\��
��6ڱWQ�}�s�pU��ф��H���J�9�����@Ѫ�g2��ݻު/�
NA{����(h�6���w�v���Խ�$In���A�S�Hx�@ ���K�Ȟ�D2��	�����f:�_���8��4Yo�z4_���$�_t&;@x0<�<F0��ʁ&��qma�\2ɽ�4�����I����m9Bu18��K�k<oT��k5��T�lc��p�ר�X�p� '�]!�\+�>�J��������[��DF�%	������[t�R�{)�Z�UB���}R<D)��ROX���M�:��ִԜF~S�:�+�����{�euw�8_�<�����_�2Q��q|�u�=5�Ԗ6���Z֩��O��i�@��Q~�@����������ā�F�iTWC��lf�?����AR9�~/3�&�LqAȚ��/��p�M�E�R�k�����w 
��>�=4"�h0󑍔\���kn�4h;`��*<a�m�V���4��HO/O�r�$"y--��ׄw�(E�B�W7u�/���NL��_u�Cbv���۫Q���|I��P/b`���3�wU�d0�f���S5G�,[�ֻ���[�|h!A�wޫ��U�ܐ ��ԗh�v �T�öo#K]y�D�z ����W�!�i�a�M�t�x�c� G)2$�$A̕�G���5)��olz`J��%�
�*���j�]���I�4�ܤN"ɂ<�~�����ޟfh�i���R����Qh���2���A6ם�o�5�x&�r9G�y�\�DBuv�X��UMH�M�?�����?FZt��+RR%PEl3��WJ����æ���iq��s!-�0Ƥ˗����z0Q[r�E��޻�0�Q|�ա+�u���z����A=����29��xqj
yW�m�c�OY�f�o�Y� �^�9Dϥ�J��O�Ҍ�D��v�}'&@�*k^�U�������.Od*� k�J{���^��f@n4�m�����:W�'��j�%�+�� ��@T���d� ^���$c����6u�62�� ��G�f��ѧ�l�2Jek"p~��o��gi2�EK�D|�kNq�4F�_�(F=�L���*���,f�Q2��؈U��B-tZB?�_j4P����nڝ�ڂP#�i��% ��M�p���ĝr��u�4)�H�SBw.?jZV���˚6������um�$��AS��=Ìؾ�5BO�Cm�Q��q����,���k��4M/�f����	}�2�8�])%���[չ����q&#�[Q��t�O�w>�P�c/%I�õ*�rp���".&��h#^P����˫��9�p��d��L<��TK�D�����LF�R3���s�шn�taH@Y�ـϟn	���_{�KsqA�
�sT�ʳ�@Zf�O��(���3��o�PKxlYK8м�x�\��T�A|1Y�!`��^HC�������%�={����i��k!�z�>[��}��}��R��9�%��ؤ��S�h�\�T��9rI���"��ް_��"�&��F��^5ː�4�SxO��S(5
��i�ª�s$_�[�"���5��ԙ�A�]r\G���Vہ�VX�O"[�e&]�`ݕt�"�2C��k�e⨹���S!�o��)�-�<�r7�����	�_��u�$�E�K�}T;�{��CbaJ���`�������ϗ�,}���]���|���c�V4��� Ү N��Fjj���r����K}6��| �*���r]+֯A��D{*�Ap:;h�'/�l�v�Hp�9�,��뒜�.�h��H�q�2�*��C��Y"���r���v��a1�QSq�T�=�l��dy�� ��܎�Q�m�j�.}R���Q���	:Xkr��u*�ѫ�:m��,븇f6rhf.̺�ܴ&j��P�L$*D���,����j�}��3�u�� TĤ;ir7֭�{�YCO���Er$l�Ν>=����L��>�͌Q״#ӐL�'^���`�?Ƈg1"v��O�[�n���>�W��w��JaZ���G�W���k�\+~�!�Y�����W��z���B�ǘ��0\�x�}Q�:)Y�fP1x�!�v(�f���{����j��*a�p_���`[��0��(��ף��	n�ͻ[��|1��VD�Pdѐ�u9"���O��ߦ��Ƨǩ~Y�_���P(�#����9�v�EC�D� ��O��l�bk�Ǥ�<��xp�+��>���	�!�A�R�t������]���'R'�W��ڡT�f�6q"I��W\����|%�Fa>8P�`�v��I��H����/�m�gj~�.W'�X�|�e"q�F����s$U�L^�Xn��Yu0ǒ��?PYfu_#~��P�)l0	(���.�O�?�]ƫ��c�����e�s�2�o�#p�?�,&�Hb�Ϊ���O^̪���^��+��'�*����j,�2��/ex�� ��*�ë�`q�4<k�1" �`6�����2�-uBּo���S�K���4^l4�[`��`�� �n9�5K/t>8����u�9�>�}�=h>�ٚf(��GCDFGd��H!8u���-HK���q�I�{�'�Ȍx�m1]��^3cֲTځ��������$SZѡulBdѧ����ޓ�Ŕ�_����Q��m�+i_-W�s���|"�U�F�}F�����.��&$�73��?�=�:�������ಷ�i����,%�.���xZ�
E����\�,[OX��1�s��o3�l���  __�o�ri�a���H��k�=��Nb��,d�@�1(Hϭ�A����G������0�[����~�f����I�� 