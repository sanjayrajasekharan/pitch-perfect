-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
P1HciH5OyPVc4JQeyHQW9I/hQXuIn2rEdPLQ84mk69+aeV8kvXaH05NH067ToZC8ejbCnmcQhxv+
1ESAGWk93dYpAp6MGBynypfrnkIUEN86ssiti77JRtm2jEScsYN46s+DZysxHmgtwVK0gL4WO5+7
91ZOIxyFJ3bx9VUWX0ZcgMlm0eSt0B5DkhkE+8tRZmytxAcgULMIx9x2u9fNitrL2bXeDVP9fhXX
uH0bum7TnGurWijK29aZZmSzUvYs0Vw84DRUQgErkzuI2CIVByGrB5OJiZyP8gEDTqhgXnYPD1bI
DtiWtwai0t95zVJDpLICqM29Pp9s6HmpjKLitQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5584)
`protect data_block
HKpx7xBR5Ts9+gc/pw3a5iePGFqEE2H00arJl+DTXF+Z2ZdhGzEakfbMoZ01vpolvjFr5oYjid1Z
DOgAfUDmDB6nbS2Hq5ujaPD0XPjqd4MJoZC40hyFvQuBih/8I2Ze1W4kk4BcKT4s6ZmPrg62jnB6
x5mKEm7jhiW/HCAbMRv3TM31fPFoMZ6JYuSZSAr2ATgfoVgMJo7o+6pIOHW0y7AmvcsXaMdWur5l
cGFdIycIJVIRCKpeI3Dpg5iYMGddRcLVsYSupRXLZ2Q6YH1lQKekFuSLINgRZ+lkk6+CqT6/4T5J
OXNdV4xxmeTL8TgTIc6yiiVYyfzQqNpNHgE5qK8kkrR2kdt/5UWKBisPdO8R/tZkXfIeJrp9vdmG
KlATC9s9/MBtxQoxD6HZBcyYQAggxyhrRzT5oVKvRZcumLl7wsGft/EYxMGhPsb8eMEfawSVPDTo
5xuuF2XsYgdj308aCAETxuNqtRX423dFoDR8XXRnLK7MsftnlPNps/ydpxJGvEmQGFlZdg8X6cA0
smztnZXhRcnGnzJOlmlSNCdEaREeI4lyhucCkoMSCIyEsyne0lsKYE7fuajw5bHZL2PpxDRXeGmi
7x/55a67k/w1GlWSvrshQzbTYJ4raN40i2aSV6AMLsQ+yQ2NCkSt7DmEW6kFFQXMtUnlC/3LH9eH
2s59SvBqi6TN0UpFll9QPk7XZsBDkIiw1oaVqdkITnSQFQn4wCDBl6Yz6Kwcb0PcyoVnb0cJp0bs
8zLsMvVzY3g9OeNlJNHBy/7DOy8OsZ6v8Jn89gZxr3A48FM4QMLPse7wFVjgnsw+Xy8EAOHauFAb
UMEm+kVLm4IaeS8SCEYtnXG5A3ZQ3DEKWRtJFheESii/4baAJMACP/QvBoKkWeCBsifDREvLRdty
0sjWZMRDHo0/RnnBcjLizrzkoTjn3pjJ9pcLYBVqhU7fwm/QKS+bEyCSPpKJUdTIe27bl7RffTcL
/50HuSkmLGRnl+yj7qBRQy1vDqCLhv4k/9Pc33wPZuUZV6fujNn07poNg3ngMOHMxOZGNeLdflXJ
qBmLRRgHwo23gcPmiy/6WTboi6yob1dH5lUNg8DIj0JKTswVQiHhInE9SK1D30LAVfSyWq3shgrG
FmLbU0UNOnuFmj3fwbRtvqjiWrPfIduSC0aMa5oaWDsBd5Vyuh2xcqreTs8OcWKEb2B2+6rZ7E0t
xL9x3VRjvpRXcSW+365VCNc2LNvJgDkK9T16pf4vC3GiaokccWd8ESoWiZR+QSGpmYKTF06kre/m
Qb2ZSwDCOBYysejAd58xx0nuvxeq21M3q8U/FSBUjNLVIeLq6g9zzU3wayr1TQ0Vvl6Dq/IiN3q0
M8OF2qtxW442peaIy5rqpDCZBMcMTaODncnVvaknQtZ9HG0MnLOfKHl02U2rHGR91TQEVb07PVQY
AnB3ZIQBq46Y1qskdxAEdAsNqIMXeVUZ2AnYwdT8piPZfTl2JGvi1NAuUJV+MfjqXLN2MJIPu9ny
+/9n/B+3BY6+gGCHfM/zKZ5mw4N3eMpGl3PkfUmlGjv7sv0MRdAuXQcOXvGmJ3Onq9HBGc4Z8whl
vMhUFJsl+x7W3mB08Os52BhQdReL+0LlfiymuBceCBMpnQitB2XFZ+yo05y9fA6Tpy6TNQCsaUBE
HBfRmsAqvAnF0SdaSIx3VmtsX4OUbPe1tNGEOyQ0C85gsl01xtg3Jay/msYs6Ph1rd7sYMFhclD5
Sr/fvwNT06gFbJ3nRRprcsYMurz0sgryyC/JiA9gMv7+4m8+tHUjH89dS+gYBou/yHxgG1MMwf+w
YllO8p+nhRuRKaK1k9/4EJ7BZvD39P8zWOH8zIwwn37TuBI0HnqzueArvKlVJbPElmZ9EQnLbhzF
AB7KT+j8JkgmhdWSHIgqYjO7RXwsway7zYSLjNBSryBKZNfVuXbbBUNvDwNqFFACd+v7f2vygfK+
8mINq3EggXV5KjsbNwzoB9p0qoe/mnOEcPBgAbWVfOpawSeroNlgUiGuaHr4bNTEygm6VSrywdR9
hWFGhQToIoln+Cu/L4bz1KerasqN6wuP98nugieKXcVcF4U2R6435Nj4Ncfs/LOfC7Iu/x+xu1TV
IZTLlgo1FE2pwQQ1dvnXdhd0a9oCLRWaX0tMx4Jx/LT1j/aBlpybPHUhagZyUUqZjIq3cjOTf1W2
BsmTY4qNUVfqtQ9GYhheoym4be//OvXAuWxmHxa30C0MFoCatbQFpiwC53lcs5w/UHWtqRCQqOJ4
tjeW+dPRGUozHxWPUcswcZiK4dEKH88YP3ROwm0xoLjBlYunSwFu7AR0UPytDbyFtivXpRd9V96p
V7konJwS9bshEYGQ+LLcylxa6TlYAcLQtRmPfCefYVIGXGuK9M8UOG6X5ETug+QfuAUoRAdFga8D
7f53lPgh0K3WLHWN1uPvxmhHS2sQ+JTnZWHhrBEAoUxlv3UDc7WjGHe5hUBtqJnb+9kBuJVm3qkB
vuHxK1pFrsoz30Y0+A+TydwWQkmSWOAPHTu+u2NoHZviW95e5Awsph1SGp6JlRRB0nk7X2TG3NvX
xmp0hJ4pNWizf/NFs+qqJiTFgxFLOZ1QuviHfGV4b7nvSYleSHaj9mggDRJ594IAIIc9Vpr+VPjR
BRmAi0ZF3FjEEheHCkY78oyqN9xUZJ2NMUoi0yGsBfFJYecg/72YukpxYtKKtl7fX0L1tAlQjmUV
3lbN1pbXh+BsLWC7sZ+CHsaaD6gmeVPW/t0y6nM2KwbnNWm5KUwmBnWhVZwFU5Gh71rSZurjbiwP
UeXDumPv1OvwDulpMfuwwCU+k7njyxuM7wV2cKeLRH9f2cNc0JO6Im1BK9vZvROg+qPWuuWVwySw
kFoLYL2pN/wyXTZ0UkvATIZcn+2v0XIMf45SNVpoIvUAmghFn0w5urbV30r537OmDlECJoiaJbr6
cnCpwVFpcHXMTeGJ1pPotCKsdbXgLyW1D/lfU8fi3eV0WLcRRnx/B4j/eGt7x1NOdOA+xVbh9VKH
5Gl5RtNwvVXwb7TmXWvyqjbXZXlzYYe235+yxUSfTrOE0+06tcUW9p2vpWOPy6TERv31fqZhFy6L
oSMOZKRyyeFeuBX5J5F8tvrHCgIFGPJ7dxfx7rtQLVP0yII4r7pNeHnFIafQbeNmrJY2ym/m5a3n
nUWEgje7WU87YftWxL3NCF+jwd0zQ0IqkrnN29UeGklqk4bpgJw0C8TbUrIzaFLFTRkAKf1OCls4
Qd2RMOaMYc66H57eJd+MqORJyK2MJgIHvi5tQVIeeJojVYpQXVSsQojDc3Qz1KvOz14mzPM0Xd+6
6SuCu4Uk9e7ry47utkLS5ifqAnyjn2jVUSRtb/AFo0tyVQlBjxuLR/Gsi8RCnG6wWN4Cbmak/574
bC5nd3py8JOkQdhL4dV9D1lpLegoXm4r6S/F5RFBODjOubUZ6WkShOdYd4ko8j+8Qq7oAF7g1C51
3yY7NK8h4hm08YOUTLfMvV7Npj+ZNsWFd4BbIKV3ola8MU1NQnoOwmpGE/SKTIXEPgcMR2oC+RaL
+O3iPG5dChH7BoEX3pennkoW+njKVfHXn0s4WA4lP1xCS+EgvJhCX9q04cLiYki1+K4CM/7F7TZ+
kc5ozuvSiQiZ7SuS0waE9wJvWplqfpueCgJwKX+MLHaIaON1hmX8ZnYo65JPNXY5v7KuAiREC/O2
s1JQFfGiUX2c807eUi/h2tZ5dnylQQqWr0BYv8WNE+JF91q2CzZFJzw6/ELIoOPcD/NwoaNmEDB9
vZqw/SjqngNxIPS0r+aSKWYrE3IQ9MKQWr46SIRgGssLhM8T2ET8FPkImLREnRRg2xfBIEdzK6Yo
d5VdNnmYIc0xfpVrQa5Ji9MGz0rLPPY5LpZd7Ibr9L+mLJDiyLwkoeR3zklZdm0+jUqp5mi64buf
5W7hipupxri/y5VZtRrW8PUUifEoYwcwyHUX/IUkC/TO/GMAi4ZpXxW7Amt/Vfvdo2yqF3EJ7kX/
HAeLVvK0HG4i8HI6Y1ltu4/7pZzgmqKXQnADAqick9QbxjC0oCv/BJtEYwll4CaD4waaI/HpnSd2
cpOtiOe7XTuYvS+fM2LHOE0Em1vITDiZuRGRFIXtSoFfPx7EzhXE9hCGfutzhEVoTaaExxLvP22u
QYnvTyoQNrt8AI2UcPsvbobpPFb+8On7AwHcWzxFl8898meubINh+nTAZO/oQrl7T9Yc9YYwrMKR
nnpSM1A4b82xudT0+I0Ryy6MyYzYap4rlKFqSY+SvK/Z63jeo8n47IHn8+IL6CR47gprj7qBsUTn
EkCzVB9/v+llpURRhZMg8lRNoluB52ymPQeP3ZpnHT8Jz9cNBlZqG6FdG01xGrWhAtkOmDxx2u8G
Sfq6DfXK1/QPgY5CsjqYRt9eKxNmFjbrZvrwKSRZfKe9QHUhzEXZKLrEbQQeWKlkXXZXtUW3BUA5
kcR94Fl7LXZUDdlo1YlQvJlGZWokT2eV82a5z5sOgNtUJQlfGSIn0I+je1YmXXdbiVAZ3nqjCfWb
HgRropN0WbFLzClT8vC1ZzFcspx6378+FnVgIpxImgmgXU6Qc2jO0pZ0T6Y2qw6jfOZOn6+bf7ma
SMacM9d/2lrY8Jlw7ke47Pv+qP9/jcY6PgZinkEvknhjK8rqjXOKlfvNgZbR0YTmAcadc570ZS5e
DrJSD+Ih4/HOsUINUNGjOjLU6Y+lfRWdkacjQ0rlQ6ci78wWsDdtR/f1oSywf2so4Q+dFDq4+RAe
fq+lZKoYhyUwREyULtYbe6g5/vt6WeLvKjXKQFBEvK9OdURvy3NOwuJ2qZKAhWQ1sxC1HfWV2BtM
4XdNGIp9YRqFgnzlO5Tkh60HUUkY/FaKP0mRt9IDfwWQD42wCXGw8rJ7XGAZ3Yi524YfJrjhJDGc
hDXn8yLL5MYYLrRImT53aK4MpohbmZdo8igTLSIvi03l28lH5JbJpDFiBESI17sHvoD1tlGmmK0i
zeGdH50fL/jGOiwB1aEULA4rucx5SMlz+51eA/kHPZzn7TMxqkj56J5gBeF2WAvEf7ivAvwdSfUx
sZ3VMupKX4IKy80Gh9QcQGww71MItKxHxZ51fx60MnMglEgodD9k3/QohkqycEhjQNvmhOdJWs6s
L282lzq+TBF+3RgCUFH1KBS6Mxxm6EJCotMfX1ZYUCJJr+7fMzytucI4ODZGiQCz6ZUMXEZKFyUR
bLDhpGFuVXkTrQ+EGfDAxm/466shuKy/ROwpuPm/C75wUVSbjoqSQaKpLiCi7K8WShBaFT+fKgLW
bgWqM/PvNJJ0X8f3NOqOmc/BZb+bNFtcgrgia6QzE61lPYyGqcftcS00KNkgynixbFHD6e8C24Fj
r9a69yBlbkboOhh8Z+mYodoKawU9YAGkmSjb/E9SnAkVC/xYNIfDhMNRSn++TzsPXm7Kqo6V33pK
6JIwR7h/nh8qjidh9hop/YUgKirOJV3yWiPugKkxEj7OhDfQNLCbYlxne4BXsP3/wKdlawvMPBkQ
j0T9MonFSpj6UQ4MAvEEhEA37pGxV7jFKAonjvux90A/RI4Ho7ggRXMtl2RHvDdNFOVJdxeisgPz
1uotbKooHAVvrL2nQf1ui3JZpadFir8SlbnOIBL4Mf1elTqNFcr4PHcGkfUHqyy/DkUxT9PKRHJK
dqvPqRDrVwhCmOB2YJkT/TJqjfFTjmZHA4uR0n1aW0V7sdCC/QIP2EXuAGykBJRMc7SRfdKrBEbx
/T17rAMl9FVIK4oPCi3DqwN9U5+o9QI5zqU5AdCoTPQO//eTsBzhJmlW7eUmUTmVc1zPZZvPmudA
ogc2GgUBeKSMBh2yLNpnShIfoEYUSiduT3HYqwP8eKKOmXTZJHUMoVXFJYCPRbYuzuuelkClhYEX
Ib0VIRhLBO8IRIvqh8NoQBOvEK5eupqxE7OKaTUSnLO17ABEKsAaLce5M6X+Ftg9ZOWBMvAX5vM4
n8f0NmWzq3NsmUB3Bqyxhsptc61BHk/iUbkcJKc1fqPay7hR+ri5NraA05+cLFSI+aO6hrKARp5z
rSlsftAL7R0ChjP8exS3j1GolbhpfvnBwyJEEQ7FF63oPxPRSPCym5oq4cleGIdUhrjOyk/sUxIl
TbVTEfBO+e7dEuRGsfmR4EozWhaqghKKNs9ha7vvbv6QTfDK5gD6bDa0xshVPoRsc2wgR4vvDws4
lYuMn/GbYxgOnEzQ/Vzrzyv4Hj6ivu8esCQXP4XcXq7qnY5WL5OxnApK32sMMAetaUaDYDFUHZSi
ovUMJm1O7J8fc6CgGhBQAdSDlKZGTnGTgojEtGw2g+RhyWdbt7PhMCCJGN/Bah4RsLLZ8qi3D0bM
ucE/qXgDjYSUmw2aJjpwm0qdYWqs+1gIkLkafqGPFeanDcUyua1IsGvjtbwlwg66hEtJwQVqAv0M
x/y6gDCF7F4j7q5oMVp0sQ6fb9S2mZ8T41sdSwCztdZSMr3FFsN32lKSsySl4n2dnXFTjrQJX2gO
I2WRS7bGDkthic3+WWO4rdzmEY4BOmfdLbkOpt/ZuNg5nCJRpq8eUH2PGGzmLLrYTK6OdYpf7ith
Um8+j+Z5Y+CR8KyTOya6rUA5+GlUeXER+JacFChrUJz3uZmen+aLnGOcreuX1rOkyOFK9V6nzYB2
gxSGeKi8NPQOWrlriG3HZsAGvhai1BBmCHdhBcy9nqZKJIlFJ8t3Ju/TevX6mqGqbGuysj0BcH1E
Gsz6iX4kqqFAnfWATIlPaMzOcVAa6jfnjyNdJwtKFEHNccdzaOnGhhRFJOIBv5ZyVuhHH0+bGz74
XyJTkCUnXiXy9hvrx/MC9TTklG86t0vMwndDkZWrExdRBfNe44nkvlXCr1olxbTz3vJh3jmcw22h
vPStZxNzFRb7rog2MJg3G6QM2M5/SjT5+0rmiiajKWSqOp4ajry3y+0AtlEkhqHE+Y9lbY2da7ZZ
n20ehjwKMRFHZ8/DRxzzyZGLkFKNtoM4u/d8tE9DKniOPGVlV6jKrE+gD++ZmtyCdL8ZWtB9/ujG
kOBf0+9luavcfi2MPcLmT/7WZyJEel5AhEeTtrGg1UOU7cUgEd99uRo5oNJGLSGqfbvaiZ6UezuJ
3Avz4SqqJIOzTZBW/LCX1jNT1F9FUn2XOAS+0ZDddP4ODt+sG4eprWSYnA2FMxTAxDtj5gtlJTGG
amIHhbbENiuVxoIpX+C5OsbbaFht8HTs5YhVh9pcTtVwgSXo8foeY0mp8kpaKqnSaOJyR64Wbb+b
AoAx/BocJEOurTTva806T8FpFPUxJPsy5WpEh/fwXOiSMi/MfGl7+Sv41ZdpZku/VwYtA0mywFlR
HiamFHNZ0N+OiWRL/rgBxtvQ3iDp5hr8gYB9nVT+ZKXfl2k5MWtJyXCcgBTOYJCvg3M57OaNOA==
`protect end_protected
