-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
X9XIeBJKYfrkFnOIhmAsi+0T8b3sKLjtQICtFIbmoB7v0gjSICj52K0rNTts6TO7
TFqd7eT1c0yNtRGq6VRDzq8mcvWqeNl8D+v4n176gK7Fj/q4XHZgMsBHpPZYIW72
HfcfONVHCS6C0zk3rMNcqJnIssa9YxKrdIjUKYeVdDov1mW2CS+9YQ==
--pragma protect end_key_block
--pragma protect digest_block
2VF3PjOmF3fkRweQxFXHhI2eRaY=
--pragma protect end_digest_block
--pragma protect data_block
nMkgz5xfPugCuceDVm2Obz/gOkyIHRlSJlEqWSsElXc67F66Pmns6nDePtG9U1BH
oD073kCCOuYAaew3MS56Zj6smtdSHdM6BhH5pkyaBqEXJcAbnNo0oZUlINrkWPJr
/SHxXCI+OTKi3Zdtsqa8m2T4hmUkLYISph2Jqer0uFjQ9sP8DSCSEaQjCR0Lau1S
tiHOVxjIs+okkW2TUMkfOxXk3ndyd1eki1RkmGiayeF8HjUae2BNSqRu/YJRZfw3
lMKTBGpwP+qMbaHdwP6K9bklyVfWwHryFf4AcIwXxt0kB71FXm78fOYD8w2ruusl
Mem5MQ3p+A8+6Osfokm0/JHk433hjPBLq/0q+38h2NpdZFa7odDfRGxIYX2OsL60
cExpqaULa84sjkgDK3aPHNoKl7Y3PP9e06HmrUWU3t82xIxrM/ky+jcFXe5FDTQ7
5HYWw0uTeDjYlb81Uhs73UmzyiN+69mBu2z9pEpu36pJYT7G6e39ylofVX2686Ev
aLOaj3gP6NWIcEGVOOOVIg6VRaR3jnvJjhz28Q0ZLn+wGQc0K3S1ig+aQzNHq1RG
5mD/qNUEoqftbv8SHJ8iDRtdAzR4OhpN/fzDuj0uE1GzZNmz7crFsPUJj0VLF4qi
Xj3aujIFUVhZjDw0voK65vmDdg2bf8CZMxZw/mwxl3nv4pE22oYUMEESwQqjImbd
KjR/uNjMxcAS8QeHOlAmL7/dHRVLCcMCAwQVvtxkkciPAH6FmaFO/k0gL2Zs8vuq
9rgHTdJj5+V940pxV1DMNdwNC7JcIn4tjuPHuopkAHieJeZxVAgTmK9sxR203t9l
IvWf+vp5kIAWvOm4rz7a58s7tN4K2EUDeiTqYiwP67AaGlBy+h0IfL+WHEnWrGHT
5iY7PnacCffHR8wyNsVHA35bfDlMopxERiLX/ZkRjzeC8PYpLkFRNkwXUDfdeOHU
LY11CUyUfx1mxxElqG0LPVcbrfuJpgdwNMcBvWFIoTw30Vh1lbrL+eMUJ/BIJ2r+
X1/HgCyoIFgCQcudL4FfX/PQpOOB77EBFs3BtEGM0kD9Vye3pBb294OT6/tLGloD
nTVBViGhpdP8jOapF56BhqnoWSaCM0g49NmiouXd3m9cYoEEpUWN64KO9e0NsrUG
Mu0Xsqv9Lt2XXRn8KpekCKflxb3O50QutoexnQjOevuD/spPcQFNXjBM7QlhJi2d
VM5JAJlBh6tyrOJC68sK/u0cLDZZkTrqxGhPMgjQ995U7mI9SauEulSaI9TsaDIc
s0/v6LCgEuS0veXYLQ/NP7dE3vkyW8RNDHTWEkuaJS2uHL0fCVhc6vtcTlKiC8h0
vDHnvwyFjrPb9O8mZPb9rLBq6mrtdgb3bHjls7eE2jFUigszhYrHS7Uj4t5JcXiy
XNme9oTNBx7JHGjebSSfFm8aWnfaBINCGGqdguVSMFo/Emy+HLUEmvp1b829i3NP
BAiHJNKVW3w3L99kBgc9NMIRZfntRUGzmuiltBHzAED/YsHuhcHLm+Zxg4tKRrOd
nQOVb8B5rWN24wZJOAM8CCZmh5DYFz1ALABApeZqn00fF4IcHj3jZZPUHcjz3Mnf
0Xf27SyUAJS+IpgjiekUDMwk0ky8VFEuUWktdYclpYr25mfpZs3dprmX2uUitaNF
81oV9OesxJzLhw3lRKAZMbYZPd4Wt4icJz/3HbFmTIjXG1TYKUqbg5IgE62Zv4Uy
aqmeA9QIRtbhsoMeQSFCm0AhLlv8hVRlRfCmSoovm8ZL0bjFmgRPXUkgGMo0h6rU
yQElKbjZPw3W3knINJXgu7sDh8xZ47tJA9nb0bEFDjYngAFJ5I2Yw18K6Wh3UeUV
crOlAtStQXtTgZAD6t6IucYVwwwaxRdghbKXQfW70GkqCRrlubljnSUVhmmCR7TS
IEeKkmA98wHtZ3gZ5pRK3apIuoinAX/dhyq5666ETaeetn2PuaG0M45BYkloPGpC
I+k29v8dsdHCaxNeD3Vl8fcU76mPMAuuZxkeVnhzQgYXWikqo+/g5rCLwoSeoPCf
MKh6Ou7hb8ynR5Hefa3d2yYOr+yW4+ylAa/1tsvrc7V6YHhvDQNGhjiLuPgwbPe3
zJKA3wCXKo032FxBB4z/LKjpKWu0ufoK9Y5KZwssb8Z0othu+hUmjD2HMLejkump
QFgUSQQ9ZGwbdG/MqXrB3n9JQF+no5ibUf0ayQ1dM+LzCAtd5vtlktvuV4vWLBip
XOxKjWoeaJMD4k+rTOXakiL6UjYA7/mnRvS7LI0qkHv9aaBU5ZBar446vWZ4ojHu
RErc2N3B/LdcMyO0Xg9s9C1qWe0pAqmeecQtybeyW6ThFLaVsE7wHXLV9UVoeAGG
2QhTb5prNDsDnBL99w+kNEyahjrXhFm0ZCquCe8PyN1ZiVvhBpi/9ITYBuMtx5CX
LFNtpCOndg6JGI7cLgt4v4iDwcx5Xy5FMJG21CGXkbB4T92ZbzvAPVWYZQz2yQZD
9rhLDk7YgrB5IgSeYfmhk2YYOGZENZIngs5ZsmcV4kf2VrDF/eLzbbE3pojtcOhf
G9QK6U1LZEHAV93aK/MuG0UAQmZAm5o9VW088f2nNJE5yjRjdceKJIP293Y9DSJJ
qBxeW1hP5wsPgBa3lDajGyqysu/FA0m/CFnf+5qUWhxVDHXnnXPNsZod7Yq5ngYD
SIw6jwW7pJqFHI8ImePfNS5Ro1Tes896l+nIvoraDmS9HSs8DYb+QRaW28GfQ5e1
ZBMaFmSHSSIDInu6nlXV6+U8ofF1bLAjcu3arj0vtK05pfalxsldgVfEJTRJXLDc
hOJv1z2pMiy727C1c6VNfezyFXMDyV85SIzf2yrkY4/sWg/VqVart7LSJdNai6E7
quzEr2w9hnXHoW1Wpcf4sU7pk2T7ghbH+6T25dv70jGLGQYluyb+nz9SOuZXgwAf
bR4X2rfjO76PnLraEqpbrvhBgfe0yiDivrZkjzD2x6kCdM+W3RhzOouNMQL7UY8P
/d+8ga/NabmPRPBtSiDIci03Cb4i3SbiS/2huBFclEQFyeRTmazN0wZxuqe3b0lP
zHhfjsYD5BZqxGC6sKUO0uCBVscSQ3b2M70z3m6F6/WEJj27pQ1jWRRjdpeIVmqH
PTLtbhCncFdk/uBJN5+aV20UhReKnHrLKMxEgYxHazTdq0xhBsY/5MUczKf2bvaO
HVjr+E9rvE8lmr/EhbWib3LKcgunFy+1Yi/zEEQKtiQYfCTZndLbpQ8UZclTfYvK
CMqdmcOPKtbYpsE5VMeTjK3oZAGgYJuki/xmvnyaxdL87oNX+cUvoNfoVnd/8rNZ
qHEQ8e5pF90ZunMhWNefwmaFSGdDYB71Dg58G4/oM76mV/Mkpt2QpcuQqZ3WF64M
k+cptTDHwQGaHgzVlBpPh5UOIEq84rnmSyvkjbPaUa27AknmOhQMDwQnHhRiSDkk
YIOkHMPGHzLR5XwL9U51Y+HnaiEuFqf02AjfzBsXjjbwxcCTgKS9gAcvn/CW1GZn
Uu5TzOxVGCA6VW4OPI6r+gCt6sKi4bCtDLfDYUmMATLR5kYN4jfhtcA6MLrzEWUO
ONveSPLKDZUP4ELAP4zP4NsB9zU2WlzqkYh9C2AX+uvu7Z59Rr5urvVIBS2nIAov
uSE7Qgbfn+JjIsxPKo8avFLz0022t2xOfzen4IhovyePzosg6AS+XH/HhJlPZzPR
HcjHY/4+1EuKSVMT5Dbtzry+LwsK1oO3aRk8rG8ED+IFAiWjvLRiiCnzzONXWGBA
kOVx+UCspzjMypvUXChzigNgigPrLOouyJxzqGZoL4ShjeHvlnsIcvAwBlZXmJ4w
ISWLxL3QL8Qs8A4CM95sMe9ML/SfJNXT9nZoNMU13g/jjB1kysFjb3vo2EZjrGGm
/xcCH96AqqAvzR82oOsQDRmzHosWTI+APdCSP/eBMxyWKj60wMnYG6IkRyrzq4xJ
oi9xctvvPu+BC1+1F1us22iUS0kKagIsUf/8V+NjJp/WvAROcPZzU+0ah+p0S+YW
ep91qiLp6kPYsxHuT/IXmbYeeS25OYm4wi7yXOT4wUXBF5WblmhAtg4Z042puIy6
PRQl5T+yCzyivwjzr+zMY6TXm/mxN9gl6PAYStg3Fy9GY0RXOtEvFgNTW1Scu8xJ
Sl5xqoeEBBNzmELsPUWcpx7cCGlzq0f6xNpv3S1aDOr3ucnVBeMFtIiAZEdJg/1y
G1ZhJQ6KibRrKoxMnPVJme6t7leatIThY/xKbITQFUDwP1D3cnkZfBKwfkFlYiJK
699NV6zCwRnH4M8I4WCdAI4zWA5/Ph7Gjf9b+Gr6KzdLPUguQm8FuyQYQNvb6a9t
XL4BX59Yug0JRDMHLojMINCPD9L6/LVmeIu4osZTzVqBWo9l0V42+IuTM1yMb8ta
WQPXRKiCUVbaSwHdnXoq1fpL2uxvpcMJqF3Bvk+zA+ZHqk5mD0CbCtGGv9IPAuZU
XeLzUh3Z4nc2Pj8Y2rj2VMD49EVu2dgqjO/1Cl6EcDdhVfRlwKTy18HgOkvyimjS
F6sz7f768/WbsUnOPZlML/UgSzNdsQbnROJFypuTorEkO6H+cGbIA/RsdD/fuVLU
p4RTPmnMjIKp1R01mQf5CHADhK8UoD7hH/cYRHfsT+GhOJZcBHReH8U9aFLu3tw6
faM3bvYf+W2seWa1apars9OiLA2Wtb43ZLQ64JocK9tDNznC2RvMYycUWCNk9wl0
2JsQUUCXFPQVJdofyLAmMlD7Ya/o672etbJAlDIvLsIoOADcKrCUGukoaqvWA3FK
U4dOgTSdRsqOpS11D6Gk9zHb/C+ZKgkKki2L598Rw5+41Zz336t7Xh6VoQaHQw+j
bfZTLP5eO0ENtDjN5y/JIpDBbYXzYM69mjddSpxPF5lhsiTPV/L8K+qpam+ffXaq
nJIpT9uLJw5AWh9++5y5y3CSJ0hGkv2nma74SCh4nmSi2dCxcteMVKNp0KQL9BGY
0VZSfFJoUiZEn2WoVh29VZGSJhqME14tZZ2uTzsCXaKZo022Hau1iMNlfxcY3Sv9
V8Dp500vKHoC3veBgnF5a0j0nOAg68ev1rf7bmDZZnLf4YC19BhieAXbetbvOEq4
m8tDKRKJp+KZaznyGVJz6uN6TrQMAYuBykpbAAWQ0rSp7gg91DD/Lv/z1ecA9w4O
9kvajVQQYBRHs5zASfZiA/iKRxqyjN/S/U7MBRN047CqIMq0qFWTNcUMS9MYhrPX
29qgy3SgLp/Og3gl1g8GjDqypfA7ESP25WR4MlRKNkaBR7SFVNod4BB9U9noZJyz
IYPJW6BHcE2XzaVB2BZCVssvZ4YtBn6E/a4LLBmzSH6uMZNj2tUFWaUkMbTXxCaM
ujp15m5/zD4/s7Twlw6SaQsMEOsFiUCNjaW3qCHkNcBmqBsq2RDXFAtnzgMVEtoO
KTzfNAzh+rZqAh8Bu8w32bbidNAySd1DN16qbXMvrZVwBN28hZ7GnxhtcPWVJPn4
CoT8ivJTKDHQ3jQmpJ1L9sUuT0lY3XMJb3pRH4M9fKMKl1c3hWZJqhfBw3rInmEH
xihtIMtn1NOUiJXBMzbAcgDEJdFr7WdF2f3hTFfOJqBp24KgLejvJhmgLByZPFmm
5YHMhx2yJxqLumPfEIoCexcVqvqh/GnNJPW+4kKzfd+F042WuB/zAV0puKBeflQe
jP4Yq/wDEd+d6ZMFE213qri6oJN68QC2yXQcx+51ecucFJ6oEv+VIf8iD46+iNfm
t5j4ON1x1GTcx75hIZTnxyY3KgVFeY3KpH9JgVqwtvcUFferhWAOmMr6/2yqFvte
PDndgq4WdLoU/TmFcz6JaaZ5l7A4wizR0EzxJVzy7c5AAFJXAyYBPiE21O8JF8zN
u/picndWOGJ8dk6BE6l309Y3FWBJFtxm68yeu4EU6h48R4RkYUQgXYQTQTten4xR
fqbj4LrK+Q8b4pswGmIWgwF/3A7hTwQib89AMoNV9PsbeYMwuxu5COQQBM/d9hDt
d6wyIpvn8Erm9EJMG1d1z42Nm/PXOz21D+FFd1E8G2HXLXzEkWWQcnwpS8hXIAge
xpulyoKClB//nGMRkigZFTUMz/rN2nHls+KEegmfsiNUzDvkF7KPdd46vIIDta4f
VyWogHcgKJlj5jhVk2bFppeezGvTXeP5iX3UnyhwBXohAbhXy8UIkfUp2rqf5d+Z
YVUvGgk3a9z/HidEZkaiKbfZuHXiU5sVEpVmuR5a0ulV6uL5k3j8CRPWgSd+g7Qd
n0iskotDevt8adsRsnjU37I3NaZcPuHpnMeOfdji+ZtoWO/LehwMgMg6JaZPpy5U
XjXQ0OSjCh9VwZXiDrqldyZoSaluup6B2mWiYzgfvQnwnmoo+AE7/ef+UMdqlcnZ
yJIytud+3HfkDlNarXRTDh9+j9MnB8X2+mUx2UQGEf4NnmpfaZNTV9KaB0WmzkOC
2hvnRkHw+EhOD3VaU0virsv2pj5nanfAL6zuDAcmVYFHOASE6oHRM39uYGZqR9Us
igNXcXnyTQ/iPbF6t47ZUm505ikGbpq463GUsO+fQgPSo2cCmoW2jLGvhxGro8ON
d0uY+rm0ToGRSXs/Y5Qd7oUsBvDKRWJmi+IsAYbTxSzBtAE0dnqDgaG3Rov8w9YT
i2kSRx3ROXoTSdOlff7tvp68FKkVvu58IDCB0MXyxLVxV1dmK3mK/Ti/g08cLVCQ
FHR+a0adCT9zrROTrxZr8heLWMTWUXyraih41SnHqYpk4JhkRlAKFY8jsLhOrW8K
HKE0SqJYbhbs3C/LqGTUuZCf41Yk1Hvn9k9mCpTY66haFG+JF8aJUzzEkkWKjKqh
XX5KKmdw2WyhC/+Scj+RPVndfr0Kw2muMmmh+GVcRAQ79IKdZcZnsC8AU4FiArvf
3tL+CbHIM4TErkWS6ABS8CaQLKfibmt2yfGU+khPyroJlEqJu8sljQEPRN1LzcEO
NHaAdIN/cs1/pCQykmIltyF0fZGodXXKMjPFaUrZ6/4dm2ugwqv8oN3R/b9RetQ2
FNvmzeoB1ItraIFjsEcAbVnNEZXJmENOu2t4Hi+xiqtySR4anv6e7Bo/uFtDHizH
m+3J7sZ0uk2CVEhsKxdR3RWi2nftwu0KPggmo1mWH8p6rtnlPyn/f/TfJNg4eWSz
NgYu5QHu+EL9bD5kzNiKt4/TRDpXRDbMMF3pSBKJs6NlH0/I9vf/h9vGpBI6CpEX
AB/MUuAJmTt8jM1nuUqfBdGBz73G2yM6SmNAVQxFDUyOHu4zmAAgjInV8L70jIpM
B3IhaGafqcS0DSdix1KDpCp9yJZsdhFQIjC2XJN6JqLLWOmKa01JmK5GfLQFJaC8
yNcdTPtVC/rhZRNoT6ash5VkMQ948oXXHG8qtNXRayRMoO+mH80WxG+lbZycYMnq
hOCTd/30WSDcdF69klTcSb1z5XopFprV13fYZXWxX93H3w2LMroeBEl/m4fLkizh
LIqxmLfStTAGhRVa30Tiiz/XRgz9uqEac2w61rovkYarhPc5ni/h7pOBja/SwBcA
wvIqB3/iMe5AFrLUsX0jGW/zt3/wfxoaHSYxSXPrzd5uQXbLzH3JPpoyajR/vq0a
s+rtro5+tLf0v+GcgTweUs80TC1t55hbPphfUGoYhdhmtZsz71zs1Nj8JjwqFd1z
PxlD52YWm0zAxX097LoktIyp99jxikaVJQzYkRNmHZn8Fc0x+kWNJ6Q0Csvjl066
o0B5QCySFFpYj7XEIEQS2o3t7WJsi/JK3vgwQ/8bD8JHH9nKA7BQtU8ADZHHAYoG
pyb/MTF9vqQcmJc1b5z+BEtyAzO0AdXAXX/Pyy5CUbkvTlK8ieH0yupoQNvZ3pOG
Uzibkc8d2Qt30Y7jCBTyIvGboNUt16gQMY7h2m6FqGcYbGZlaBnXBJK0t+nrgMtd
ngygEuzGxlHs5D90NUeFoY9qZpgXzM9QgtZEZt0qw5JcxjWFEFdQmhiOQrOEccZI
HgBYlVBQ/nQx9q1lGTLxJhjndXLsXhemLNERCoB6F9ahrn6ZCVJKr9hN5sL0ybqs
cbTyOnM096w71y+cRzHYcILNlhG6ZUq9wgsaPfzUQmGkC6eoC4zKtxiUSnKtr5S8
Sgx/56R3zEViYvNv5zS7lULd8APr/e/vKdBjM/IGpCnya1WoOaxKTjI9QpoSP5Ut
WsVbd0Vk4aVZRrBbb2GOJdmm8raKxNMutDatFvbtiF+fChCcUVqo53iu0hJxwj/0
xNS0qS/5Me6k/2jdjnbfgWVpJM5eRutrnXQLv3/vWbTpZgF3xSVfK/KOuuttd2KL
sxo8SCi+F7p0dDuzaCsQNeljlK/WOfGeye7w8GGTvL5uJH9u21/0lfa+DKDAnmEt
/kxquxeIYU2YcsZLj2qbsAY9kGDiu5XYnIs1SC9A8i+PnLA5K3DZpNP8vrw1ZbJS
wPmJTmkVlRUL38OElmkCw+DbXXjz4Hnb4xygLJUCXBWNTOTKcRJrE6CVsRLveij7
VBCKrbAfYSd9IKufc+a292yfz6ndIxXhgcFihjigNraadAkKbBznYOEUFEACjfM6
hpCQBr7pO4ZuIzM1Paro5rIKsupLu+AiCLg0cn5f094Rw1Yu9ZxxUteK/7uCOWYO
FE37HroCfiyR3aoRELhV60l2pnQU2C0oLk8pH4o85sRALTO9q2USML9N/IX2WCMO
0J1QrALYJv/OCAyxQMuunrYM7THQUfiimCGStP5UuAOdaIbuxAtKB/gj99POGxV0
Wt57PEG459wrdhrunDpsNbw5WLvNelVMQoF+XqjDH8q6mkF25GlBezIGBd8trNaQ
q+hR5hT3BSWGgsKySot9NERh5s5HHmu327fAv8bTQtkFtkWcJvNx2YLJdtGgn958
RwtlLtt0tDqIpF3U6gApbOue8zOjlo4Pzz8nkxUIL4AWzxP+ozMPLVgI2b9vmqjv
K7RXbcO1LeNfFnxIZ6xKKS4IpraDQfjCKqAMgUxMif/jhc0CtPZpX8p19ozCv4o5
uKRKNKT5XT7jGi8mblARRQStmcYG5YMzRoqhweUbVk8ZhrLWHyMvenbAoWHa8YGR
RZ5KSokY4XekT8PGAxrGQIq9E2eV0MNDihBiiyq7vWwMekKalRhPdQ0skeQOqKIr
4vgLFkMkoFuxxPiOVNaFD5VnybEdEmAVk+32nUaZk181+wYt1mMGyzi01r3D0CFC
boYb3/iP2qCNAoA28EyKJeKODPNBv734bTx1U2EJURfyJ17qbWfKPstfm3lWo9j5
UmE5PhLphUcpIHiZDC5OCZDyfAJYnRjyPL0l/AyRZnN9SXL1r8otTBU/gLxQWBwE
8OskXPyeLr1NwnVwuwxvp+oWO/iQfniy6i99NgfYMlBUzYWWHKbgvTUB+9/6AAr1
fH/jvmJQHuPUHtSuSgfvXyCyYPLVqKjd30hQYTIIdH4Jvh7CFIyeHfSkqKnRrP3/
5swb0EIcqfcFM3qvGY3k5MEB8pszosZHmXKSuUUSqJXKlxCcEcsg+snepT1v5816
9mS5jTN0gI2rHMzHa81jmjYBuKpJosMsFgMtDBkJw5p4QbLGWClQg6EKnZ+IRjnl
gGwZagUs8F5rS9IBXGMCxteK4IUenGDfSYh4XOhRxO0Q+imAlZU+0AgdEfvNJMaF
CLIIDkxqOGr4sg2d5l+r2RmmsyzBiZQyjW9r5DOWOigqB7Xy6PHl2SaF64Fmqmbk
iTGQKNbQtjKX0PNsP8N2qFskzurx2v4vnPoXo6gQ4LISmnRxaqpmunTka8TlMg4F
lZCO0jqU1dQz1wXmiUgEtPsOToeE9ZrrQXzOC7NfgKx97nD1cjRxXPA/ZWyNMkVA
RQV0X8L0KhyyQpiw0OuIceASkiva2QXU0rMEWYcfDlycsLomkRfWJqIZ61IKj0Hh
DyhaEhnzBkIEasSABjw4KHiNGR5A6Aw9KE/o8IyOiLlOR1q6UNPLk2mPP71T3j0p
aiVg/CE70dDQbXBBYXtma9Tb+W4JU6OuIRWlYIhrsPiRGqY5ZON0n+TwGoeNT2RG
DT34HAIVw3MN4OfGb76V9YPJQeJjKfYGs9pt72BDFR3YMA53ArPSO2xSR6MsrD26
OY/Yxt9QKb+dtjIh6kTqXaLLCJy/+Ob9VztQ69TxP4NIFOLFLpXzzaSyv237zv6T
XfdYymJCUnIrLWs2+nmGDlBo2EMXf/aIXuz3PMRUTMmwuFcZ1mT4atHBCCwXrYD7
g1SET5UOChbkk1rWGkkj+aPZcgmDyTVqPOF1FOWmagrEa88qhMRWofZpgP7OTzxT
o7fz/BJAoEKvMuRbnX6FuhaXe4X4evwCJJi5FfHDahWDPfS/IyJkpm54shJHzsfq
0n19KXwM5T8rqQYNdDXvPTHlJ/qgv1gVxps85kxnlwheqbWY2uA+V1yoz8dABzPb
tS5V0Ij9nYdLSID1tr1tDFVcv63o96Gm/p3iqdFYlO88d/758NtnMby6QEWy5UEz
TPFRcdRuEcyDi9PGNn1YSfHg3hWlMb6v5+LQIfe+YnpBr3rNz7vGtRzpQbfTdxxY
2gyQzH4fVFJyGi6zy3S6I0O0L/8YySB1xk4kjMzOVOcWxqhHPgLRQ2jAEQTsSwKq
rl8i/Pzu2cIXaWr5r9hTBkpA1MHbm/SMR1O+MzOTIEDoNoHoYW7EFP9yaUS473Or
LgY0fejgWPmnRNP9bh5RZhej0cag/AXLm+6Kvb9v19p0bxIfFrMB0kB4Fz4NDnTL
Jjkxrlf1/q2onUJjmYEcEkeztxug0XTPGmv2E17mny4SA5I1GCqR3Eqd1JpfPp48
4k6T+1B/m1GmDNkrnLO8wTOTl0G36lezGYEegnhPdcLdE3K2t8bRjQ3v0LAnQdjL
mujpYwSq35MbHB/L8qAE6zYER1L334SZla4bl9LpcEXFhL38DNy6K4Rrz/SG4qMw
jlVzhzsScO+JS62mynlkP/9n3EtXTSPe8LcpYR1dcle1lctKwXJTBjQt5FtV/KHT
0QhEgBGHkDdZW3RGalxJnJxFmXbhjr/z72mxmnhUy2mh0I65nY9j+6rlrBMUwNN4
6vWbuSHIAz7yrp8QatROQpNFH1iTlc4fLHcbN+6oZ1SFkxpQmfGyfMnkn2+jXZIj
qPJRaGcl9jgOxPnm3zGFEUyOUp3JwmykGhIAgLmvg0tbhEiwkVS9om1/atLd46tw
LuNktY9HsRjB7LS1XM4vgFhvlafrZWjFYz0KYTnKtgPeuSvdC/dgmGILJvY+WUM0
1aUv8DbZD23cdwpO9LwadoIjQg+z1dgBmMuV/121f35ucxG/vvtw9EalzTLNVRGY
Ncjp8Q1V6g2q4fUUj2n+sLiqlgx0Jdule9r4wgjsacx6whuTbVOLI0+1yTA6K/iU
4cYtbgczble7ryxijypC8MCICCx2jWZIeXzPWTNqjpQP/vmhW+mnQkZ4zCK9Rqv5
SxI7AOkNAAqn8p3q/o9vD4sCPq7fwaEn215IjwSQ4idrHP4cQPAsTl2tEscu+c/9
clE7YM06d4lLEpMRE2HKc/Q3PunGQL7P/F2oTew3jkE8PV4XhzL/IE+IorHHGMQY
qX+rmWIXY7yrpTmCBx64h3eKz6erdlhJpH8bVsKyW9yAx+6KAy6HJp3gE9cz/lbx
Jy0/i5eeYZWyHP9q126QsUV6KiJwcOVtSQxQ6o6yu8J4Ww898utJrtHgrAj/Nel5
bbIkBAn8dfUqeowdkUHSMC3E8IlOVB3hgWjAm6ajyvf2/dSZWr0f6uDFWA+EWdRL
MPQ/+i4wZ5GDZf/SbVpLUy1e47hMmeFjJznA/OlXujv0Lmoh0HkD7Pq2ZQIZUw4y
FbEF0E96jGJ9ChLmxkMi/YxvGmpJ0TPdIBIuuul5XJx8Posf9BTKPYUr1nB5zqML
NVSa3K0gMxi/GNJAka5/rqOGcPbNoGwzTB4BNJwBSVHPvYpZvkP744QXErzuZf+a
jJuU15EVqMVqjA1mliwmYr1QGy3NDLHMJn6nFPUh09tAxe7DeyIJqhbA3fsC50pO
1quwHHhvq2I2haW/0tgCg8JN56BCuJlHvuZ7Ry8IsaHtMvKIr3XdUVMdabyn+5y2
OQwTZAIZBGsI/VM0OB93TLNsVc9E3q2teMSlRV0BK5QUsHqnhEIsDbaBkobDkpwS
jkutPRqPQsAiKPI0WGWhAnc1ox3FBFqNbpuYQwCQGMM3kyOQC1o3NT6SteBA0SUT
JAJ75qB149zeGGVsrj3kefiY4R0M3k4wK10kE7rjpnbrcMEsHc6RtxfAaxWPEJWL
ydEEc7bhPXDqWxHyCnNfufk1KDOqqBE9p5b9OqoJMe5WLRjrd5CO7aY7L9hhMK6+
KfQy1+7MLk1WlRKI4/mTdrSW7BPhHv1MDK9tVzuEiPtFe3iRqsM+ePY4ge5gV4dr
zGIlJgd4TMpVDctBtWbQx9nRR1TGOAf6x/dUnhzgdjbMzVX8c54pmfAOzs9XpKaM
snbVwgbn2QZrntmIWqHvPN/1fVNDdDmuNA6gBVWl56bxZis0Ui5Owpt8tsE90mQY
f8STeZYRC7K+K2eXjlzx/Tqi6/ATcd8N/QOrHJ3z2+p81x5vkYe62FJTWBj5HabJ
gL3E4CQ7nWb7SmbmAqTSUsjeNQpnBjm7WvStiyEaJSUotRsLmJ3EaE8VUNvZBlZ1
hBG0q7Ku3h9M93nC8vDM6FcadYmenAEfHaJG+BebV6yT/3KCbSruNZVyFIXGTP2H
DDVmHPFPtf9eR32Ms5wWNRo+U+DoFHsJ3w4+nn9jav+r5HU3QrjuwWhGiEQqMfU6
+txnlZKUpXzxslldfslyJG2Da6MRz/dXbix79cq0SxrPUL2QYzKTvisbEhWxF5kR
8JVM3FqanNOJDjWvXh6E/fKei6MxyUDv1z4FFBWE0LUWzWn8PjxK2Z6RO07SJBZV
ib/mNmXAHAfNePpJ0ePZynb5eqylm1VUElXFWJsDryKTmKmKkYb0KTa750Rj8oMq
tQOXA4RxzwBisyoGcyYxXmvOggeWEFBvA5nOTZU13a5UGrsOgoSwKNBSg60O6wIa
k3QyE4TTvkG/Sr6L7S7NS8C0cX81hK2m2V3ESMQbCNnHeUM2OjPonwN5pH5cv2Ix
uA/jHQFXlkOThs/5lFN32zUQfoHKVp1ExfvczwrixoxwEPHPQLkt4GWdlOU8VgwP
8dxhIhgOPkTyVOzuMeNYFSlNhU/pTeqwtmaBHE89cjs4ZnMFDJRh/UQFuZXGUBbU
OmUSO2eI5BhzXbDK5IHc7Ob5FbKqOZDfWjhjKZAJ5qRXbEwT6XkqccLDz7W/N4nC
i37MDSYRp4TywstpzYRPLvAbxCt7OPOKPul5t7G122LQZ5Y2qiQNwF2fA3u1LPvt
R+Xpn1+bf5R3oV0TLMhVIJtyj8oWci2thOx8E75ORZNBttdo/0mkUrD5m4MwJILm
mZKUe8UTJlUsgCvPalGwcT1lwkVv/Q5eArf7oRRL6il10fyFCoezdmM20UrkaKqQ
MHdzWCIcp0BQRt8RneLUA22BC3UGFvIaM/HrJgfYOmInqPl0HPPQrho/QMCuqAUM
QXvepBY1dlsaHlpOGQ1rMeGXNIb5xM/ZLq5IIFrj04IcLz153gbKmtPcEJtVL5Ns
BZ1IELFnjnzubUL+AzOFegx7qgEYWBxj+JkWujcSav/9T1Lmy4KOBoYFGBrBKe8W

--pragma protect end_data_block
--pragma protect digest_block
OBt6KHsFurqdw/59qalM5+A1GBM=
--pragma protect end_digest_block
--pragma protect end_protected
