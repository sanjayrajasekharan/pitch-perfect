-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QWWClsYzybTqJ/asG1Tki9VOXJCclpS7auc2H7+tN2ghUBqUxQdZ3aBBr2f0mevr5/Gw8j3NiW/u
1MSxzWZlRg7J1Qk9TtrD1FwLhOLcKi9Xtzp2NuOVP4diq4V5Xzry2DeADuZVB4CSFdX93uYAfNBH
6c2IOyvPxb/fUuEhVtwAJHOyXTpucofw62jpOYUxbsp7vK8jnH1wD0GGUvGmk1ZzatCAe3KBSyn8
sBjTA17Mn16+QFAOnHjIpgwQTC2GZqY84w/FRBz4kUOHOnUEWweqnrKKGRmp+YT0bQ0OM+j4hLdm
3UGXD8oGkxojS21onPfUbj0U2Dnl/q4Zr4hRSA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 22640)
`protect data_block
nRoHaFqUXKG8AD2G98PeNDso4pZk+I75pjuvapEGAwSfUb+w7MGjz08HukPwYf3irJLoA62k+gmt
LlQ+8FlBDyEDYnST6Kb+QuRlHqLqQSYTI+Vpj7x8h4nAG4RFesIiraTMQlBk6Pp2g9cDydZeytNO
PJm+BwpeUY6krKOQgZDWf0k78xSVLa0AIUOxtyoNMXpsgqHKpLm3oo8N5LkAOPQkmPBN1nqjnmew
SFl7ILpSHCgpSDvWTCkiZCAo0DAXCK8vS1hFIaX1YS1cttZ/G+amyItURPTkNbY02f0MsQXAUzdn
4OzGC0Tztl/JZA+xnujvfzp+e+OqBx+0NWmldbYvJ4PPsA+XINh2kwT4mmG6CshV6eZlHfFste2h
+0H8q3caKOqMOf8ZKJptkLepFCI7QOjDqFkZ4AuALMmMHbfx6P2TRG7cEz/STy7Wd4SlLvtRlLDv
hoN9b3ljfOZcb2vKnrl6/wf5NGpc6LsAqe7/6NsjgubCARDXgkQHCok14SDaTWwhNChpO/E5B4tg
k0juIVjvTGYWaPSWNi1M2zf0vqfjYPHietxmd+Zdwf4eRloe6VMbvkuJcMxBm/VyT9co2BsZEGG9
BJh4qJqeNlCZdOH25Pd4gghqhPzFhKRqjX/iXM4Amwuk6fxIXVvU2tnoP4Rjz8EorS14+zgj3qgU
8eXhsAQs/hbRC18Zcqz8CsE+ffVbE9JPP/8pKVWYDpdEmeYGNIRBIincyW/KFv8mtHkbkwEkUEBi
dbpRgApL0k1D/z5q0N94jyHm4YUs9kqALJzVe5jfrsX7AlcTkC7TwC5IzgMP+mMYLTiFtIOWv6eL
4TB8/qBNGZZFfqv7V1BqyHevqhLUm6PFU+7rsveuRZvTUMfk1NVa/SBNBcms3UYulpxaW081YV3o
u2etmL609ZpdarLnXjvjmj1WvmzJJDNmT2bN4HuohxpPXD8l/NPvu5I/lH075o6bkvNCwAeAMdok
tadgCW2tfZzp+d8r+RLGYUnO5Hd5ij67cakU92xxQRTdoztKqct7P+ChfM/ZLh+8i7Mz64C7Lp8B
FcnpSgOfoDP4g6nHnphnZWAXqU8MRCJSzNA3ryU9yAl46ZeNUyeRmvhZbVEWHicY1dIysE/q59lU
L2OaR86cyZDTk2FUG78uvczh4AOHRggZaXcE+CxDWVgv0TGGVKGUpBpkvfOVoBBw1p3sGG6/4X8Z
gw195g6GYMzx+QZ700/q/tdZIg6Q6k/EP0E6LgqfGhnkRfkb+9x4IJh0hOlynBp9xcYQFTMXzwBp
KaCcJLJMOwp1PsVl6dj4tA/4YFsBq8zg10Dw9ERLRPdpHMgkX4srHDFlNFI3vQUq/hSsGHph4q+/
O6vNMQljLQcoYKcN93Pxz7/qvv6azBnprkKPgYbb9TtPmcvqwNqjxSWMwlScVhGD/p+uUH8gx6Ow
178J3xzVHd2G8xNOw3AbilnKw7XBUrUhxnjSFKldaoDu53svKJOZVCSc8jGX0bMjmo3H3H9IIf5X
k+N3qUkvuXmi5QOOnv3GhzBKGbnTHUTN7iRW5LN/yV6T1e3jI9FDu981yw+4B1UPoWdvHubxQU0b
4zZkDFs+JTpycZaTcnmMbXjXW9/icZ2IZrselZuRC2+nX3QkjCayI5jqF+tO1cm2kRbMn4SarY0w
vE/qcl152BKTK9N1hkQdrwYlQX8mE4NtUHDQpQ76CsxjSNVBDNJ/phmmUF/7LrAF9ExIMzsbMpv0
nx+gE3lIdMFWDRZGSqM/8LdJzYCUvWZYt9V/nef06WZJLA65CbpCuRd6iUM6CikjgJy5BaxQ9ifc
L6AB1AZ2wjxxdDRTVbYFCTGkp7kPTV6X+9la+pYaLmg9343M68FR7RljyjlYDPPtZZfk0BhWkRHD
y4SPjBHlIDsE/Bds1Ez6juDTArki8mL+ue9BFWsZygci0Fic1NM/JS5yRwl0svI0j5adR1tubLIf
+JVCCxrXT7gGQtyefujCuv1Lrj9EoghNzZ6FM3i1lPr4YFpRrLW4D8azeO+dUPBH/TP2H2Dls904
qCp8reuAlGIbbp0BRlChND+Z89/4hKEhkm8J8t1r23trXMpL5men6CixsnfLB63n+GkxyZRJYLcl
zx7QtoOvFwAnJ+lJAQnTtAb7/s57XEx6eN7AgNfEqWOThc+9wy9HqcVrprxbmiYMJkA/QJ6mvn+F
+XxnKLExnpaqeMvyXxs2r8bW0cR5Nrq4geV4DiphWQ/LcL+WzQohw9y1/hzY1Ym9FSJ/0h7AGura
XtePIqZvX/Fdd7HwlqRCeydTfkZwwFnWuN39hVC5c08fO7K5aJE2NyZd1WuWHPaJc9fSZVs5lbvW
Fu/tMFa4KD38EsH8JINxgHCtEPGLkj+5OCR/oKHWl5yFPlJvOU1Gv0he747U8F6lnZMHzdIbe0nv
S9mQdyWo++nfFp9SnFrjHYKQZpUQXLISQjeica1U87UXw4ZtFQQIloVMegA8fhhj3SWuNEtUGehO
5FtMJ7MoihVHBkttwbj8Dtfpo6CovTVb1lGkoZQ/wC2CADJOK3hlBnhbuvkFX3jvNNax2R4Af4/3
XbnrGSFxJqFD14Rct3LoDSQMPUKENQDMXoXyxLGvZtdz8Impw+AtSXWw4FZ7LXnqB64ZfpfG9ww9
VkEtqbEKsVyO8hKniztgG0s2VAa3NA3W+YdgH3WgvuSstbWR9LRbIbg4vdWV2WuwP4gD3M2fD2NY
QBRCiMlUzMnDFS8iMZLbhEjrOGuDapI+3+fKV638gIerP8QOIz0TPNLaqYvyTekPhzBmr0MRangL
jcJioJSs3+Ip0oiYZfBB5a7apIiX93fUzikYbC54BjmDO1kkgBtiFbGh1h3ZIk341EldUrk1anBJ
JQ5SokxLwfrZCXP5ay6hidwgEUVV1YWhaIF+me8Fi1/Z8ypti9Tm1mAIBigDrlOxpG3v9M/M4HCs
yyz3ijjGJmJc3bPfviYuGc6w2Ww0PlLFkZcX2YhvQlisSefvfv17G8GbePvR+lsNexxkgwtRAMqP
826tEDl1vG+GvkLDWzhY3VLHb5PR5/6xJX7dHKZ0JdQSVOZzFIANFViae+xo6Mng4i1GwA0wlxEc
GGViVToo0QIqw0l+InW3AJxE7+6hih35mmuihRkCc9JGa7ma6WTowmNOLzbVH1beIJzgatxCDxQk
2oXsBfBZHmLWRRpz75oOm/27pfnSXlVK+kS/Sb5f6+jIaY/+5X52GD5TqXcOIcYuVLkD5ke+ByeD
/OZTPH60R9S0tFm2+cMaE2FS/aPgV/3FhY3Wg3dzAKUIWiUJHD3ioaHSlFDjjFayw97eJbL+Gru5
3plC0gPc0KHA/B0FqwkpWO73aUBuKOTqmgVoEUdbcn8VqMizRnyrh1kcNOwWhfLChIAVHb5MafGv
ZxSXmzkKDRIuH1FdWtOVllBYP8hnFLFedTnbj8jIt8qOyPVqTaFWVQtpacAoCJmKWzh2paHOOdF0
/e9130QSt4UdNCf47r8vIgW5DSOF785osu8bafc9JYdakloZ3n9rki8eD5NUR/lE/5on2nqXPAHP
75JlIbVC2bw17tqDfKFgFFd88Q8hn6ylIz5xFUL7ZeHE/mvUl+bQGJQZklZv5NPP5MWqHgMrDLqV
y8BW9AWhTBrklv5VdU1JfMdM1QF0riozPLd8O+Yq5wEmKmpTKPUan2GbONtaGOcikdxQ0tfW25Rs
jubamz6X5dRfXxRozmqo4RSM1zmRwYmNQrNSnEWxUFWEpEbXyBh4P7nVLaPafSVArXYOA+fYDbaO
SyZ5muPsDGhsKI/v8DGrMANkcUWqk26dInuGmnDtU1bPVwCdfSdWiCCOsdvoMxWk1FaeO3UEgIOi
7Kpk92s8zC958R5AhaVnfooSulZvFjcKo+UplObHpNtm21yZNhh93XdConKbfy8DG8sCgYhTfCiG
+uFA+/lvgoGhAfU2q8N6TYdJfYJIE9XapBDhUgVPtFAfqXaKczO9Myy+enUdBH/wbA2oVvbzf2FL
+sOp7E32GEBUdKrILY4c3m0r5EIQr2yfaw6VkyQ6kj1Q8KAnrVgyrQsrJ6pqRPVS1IczhCcKixJM
dojomh7q/MBb238BEwISvL45uzFUAJ8qxnVd6qwHWz9jmnrvFoB2kQwohuNIEOVaWQG70zKMnHF0
Y5KoMsCTO3edMS8x50SWyKeksPWC0kdBnG3O9y+5ARnYjyddnuMDLC8quuUAFjLrqqc4zmJg3W58
HBhQV8YznIf68tnjLx/aUO8rl6h7WIsHTBLueRZDLo46qlZHjqF3SsNGsqx4vZ+XjE41cZQdEo+l
Cr9vuaIZYqsstPW4pTXYSOGcdcLUdiuH/q1vr9y0qkolH3Uz6dXPZuUe9fby7VmidtubWgABqCE2
MrX5XWNIAB1lqG6/b63gTDuK4rIYDK3Gh2wXb3bRHx0ADtUcRC6zsU+vM4xGfbh8UMTM/dNVCgMs
RYcZ+RioVsUnkLnf1td11ggaVQK84mRNCe7jfEhloB4aZP3tt1OnMxot/uFd6mLug01E4IzZa0bj
yqBfYKHwkUtcJof5NqtActlrha4OSSXY2yxQq325TQmlOvrHsXTSyJX7c/ZVX3h7ogj1eCqu7Axq
zQVdEQmNFLo1B+x3W952xjjX4giLKOVWGwTrA7ns1z6nIqUOis1cQX3eIQ10v1NxPjcp9152tfuH
ozAQmsBokX48Lu3SwF6uX9nQHjm0MxUHLATAeRD+uk86UuuCO9ETWm3LMHiQdwkpvNsQkgwJJ6q4
+1OvGwuvvThfydEaN8rwURPc4Y+Mocz7SfCawhWtmZDf9vClLtjRkqtHTdsc2Jfsx2qmT/OShp6i
E/8GeS0f+gGervk25vVfFlxmhGfJk8qZ+9Va+A9WwdakNBntdYBM04RmevGa63D1/+5+r0QHgU4a
8klPeGpk9suYYB+B7leIoOwOEVBW04J8XjHPOeC53QpbjlYRQgi1FgajEl8jfhtMNfa9KpjSGGIf
JCdZ+KHCxIH1z1fIGSnrNfXAPqNlTgbiofiAtnH3wDNZxSLrgrOI/ow8TARKQ/EN6PV128xraZlX
bZz4O2Q5DajofUUCKniPQ37SjlRhWT/k9Izw79pe39lpsuXMAg8eGcs48ENlqa74hzj6J2zIBpie
9F9EMiqrh5KLa87/LY7S/FTGoR62KSgH/tLLXgFFKrOMGJHOqI6fg4HBwUshCVCe6sGBWg/XPJ9x
W/XcG4KFw2ZOM/iaug7GRb0s3ymAZbyzgg1sgQUFKr+Zhftf/IChWBs9Tz60i6jQII7h14pmgZIL
mIu5WHc7npSofAD1mnn/Oeba16E4LHrMYtrxl8kc1haKSTuLU5thi3bROpdkBXaQ/LJ4tGE7XqLt
FuVqA3LBLb400JC0UJIuecozphOJwUCuDQD/WCzjSbZkrBXnj2C2FRtmRSHPfpXfY1PVeKmCWKvo
TgxqtDnN2iiRrmLFfsXxQ5K2/RryFNXOd/vnhllfCYab/fOHsq1aoZO9A5R6YYI3TBz21ptnceoe
dijoM8qWAWjaReWV0E8PArzwvSj+3t2Y/Z9GaAuRrglO5HP66k/2Ue6pg7DI86Z/d6rpN4/2efX7
KISlZJHy/GyQHfMUUqhxkTVZka5N/25qfATlcIu7yjPeI0ko4InhVWpV5GaGpM/jcv4fmKTWkca3
D1vJxqBdATkpGnetSZuTcwZYOj7Yz8XnOAfm76mVdCoRs6Jopl+9XcG8w3zledyL5EwpDSK6dx8P
kI0xfVcz1JdvV+tYfasGk7yf0PKB99vH4kJAAykTfmPFOageBrOlmlJctylbGT3wyvdh9a86MrUz
Wq8p9pn02iqmDbI3vDNwHKojGMd4YwE0gmOQeSMbgSFMB4G1OVbFy9MfEn0AMDtnngt2bb+G6WFH
JrQy1X6HjNiLidPW4eEtwKiKGyIxeVKeo7l702Qu3/H9nsIX4PuXt7oSxSoTQ1xd7w3neTWrh4Np
yf99snkrfW3ZGm/ZqEr3Oj7PAwaba4v4vJLOr2JbqvZbrPOTpfi7ZTIqHmNGVbD+rLy6x8kPJKnt
k++zI+xB64BKae0q8isj1fN2ToVmXHoo5dEsPBYdmH9fSZq2is4FSJZP4PPYyiqNaSgkTT3mdlLt
Arl79sJ3ctMr1Y48xnKwKLCuW/s7eUJ68IWvID1dsKsUMkYyD/46egGHVyfVmRWDBVph/L2ObzAi
UGENdJ58IHXnwhUJzdoFIkkUYbPDJ+7V7K0JkpvgYU5jxyMgjEpYhvjgNaoGKMv8HErbu8bZkKfv
JZlSTqIrr496FQcucmz/GJ8CMwTSB6tKcunumB18b48VurquDhzkE6U7OHU7+v0/gjUqFinA95c9
BgJXjzgw/mtsafTp88+qPIYUizIpYLUtBxadvUqlXDOdM4YtSFJIdRDvWWgASIjVsdGOQtHqu/zR
94eJRjLxSCEwuVzO8umP1W8xkVLvwsVCzlT+h31/phXDTuYWD45a8ip1iAmVUjJkVZTY4JWrqu8C
J565LdQTuVBb0N09cHVtuAcazdi4Pn/ec0Y4BFu65A3nrplRyE2NW2KR858BrY8Z6l706SkYRh96
50kPv943tWwK2vfk2+VqFyeO6I34vrn6Z0ABJ9B7bcmBf7lrumoCjfXhy5quJNh3TS3h5MXqsSHq
rnqO6G8535WdqbJoIiJYzSPLdxNhNyDxDHOeKby1sDrQkq2178M1b1FcFaNBBzuZMmkmAKsMfkHu
Wdxp9AdnWB7ncqobxK9nVfFAMaiB/9ElF3LhiLq9fElkVrt5IIfc8+B/SYhbJpazDkYOX5i+p3vk
xquMXKYFkfM3dGdh4GzjCb8iMZkeLFbnjG8FXiIiVABVH9gYTTPhUMA1sL6kZIRBR9O7R8NfwZkL
yiUa405T21JxuzOcu+4ehLRLVnM8HZKdxF6mm+Q10UnT2U3rg7gG8S8YKMTADFe+EuJjzFkLltL1
BDCDJmEJRSYzLIpbC7c6hsshOGfYPM5vMKiyh2iNDUh02IzTM+mRAyIPk5IGcHjsUFe2A1lmwQ2h
SDrZT9EYi5FPiiujsZlmcGrikuf+BCBMi+qx4NjXxq/SUOssrEoe3FTw/LUPMuZtKyRw1IOt4GwS
CcobvXpPs4L2789PqJYhGJfo6Kf83uyO6j3nm6VFXJVKkfWF+S2bM7anM521aNujF4iwZizCi8lt
gMixN1izC4izURLt5Telgvz72qdR8KNZ8RABMiIdb7uhIeYRn2/Tt713obRjrH+5GMFYGEw29QC4
8Y4YE+EvYHrvHT3nDfi1r3wDcRGfZ8mlBz+uQmrqJPecjLoKPjT6DW9Evu0bbjDNZBxit/y2UjT5
h8pZRa+0qIsVQiDql/h+GqkTgl5lAoe5j49Z+QSb7b8R4/rX3EJdXaDC/UTWO9FOOyVUJEUUi39m
9Ii6LzRuioL4wCaNR5BylxITQjzzGYHxs8x08P2RjxTIVWH4Cc4riR5jS/cSc4A8gPKpGfkAKh/d
i9/092wHBWysXKo2GielKJmQ7YngW0O8KODRibzcK+i3WDrPfMf+tsAsOeSoTVpQJuAdW4Iu+ASr
ASyIAIS/XeEMrrVljjz4IQxzwPqGCR9LZYLrwFLDJ/+zNijH5oe8U8NVMfyvRru2rWuqaAvy84Kt
NrG+7gMmy87ebL5cFN0lkdsN4WadEhRBolwg+cuT90Ms7oJypwcMBsfajEMh5uv1mzkzWtyQgZp9
zUjdZ951tk2Hp4mpyy8dQVc0lqla1zFhzouYtz9M8AynCM+KkCeOhoNHQxqWH7CI4OhwvjY95GS/
BWT5rBTiHXdF69cSG5kQAheZivY2L1iOrCscLx9dlb424ocRtzBbuvVRTr5qIhdlDYHbzCQN4aVE
8yUx4Yyj7AvkktTmBdA2UFW/GYgpWIj3W5ZvZsAHmAbC6vFEIGstVyu5Q0Sx6zuFZCg6b583tv6O
jzkA/tfh1ZUTP0hbs8DnPHcS8TbJryJZe3oTkSOOjeq41OXRZWWdqXv3J3CDtAbMZZsOIKSI5ERa
bVgn2fvOMIlgKV1S5V2aAsuBoECHEd6HezYX/Xi7sh1gz2DWUc2XsNrJU+Xt6nuXerjUuzym2n4f
MFYo7Lm+mTqU0f/TBYZLXoGo5Ml6PxXyKg87SRr3z6MSJjFybh+ZqMPaQIAX1zsCUrqPFnyDZM+n
0+pX8s48c5K/01BKnZsnGLtZowgwSWMDT2J0Wm5YlKcYx1cacB1WEklLlRMKavhgeP+nxBZ+DcUv
nMrSM1hwVCNZthWda9o1eefkbFXh/toYjwV2NVqoAV0lNuZl+jRTiJ5jRxc0ZIaD2atpeoBEPN6g
muBvthPCsC68R5aP3IhApXGdO860Op/FzkuDQ07b1+q61mCZxQ0DdwTDu3PHyjz0HHb1MakulioY
ELiGfb0EepvwL8qAi+HxtgmP+/I8bcQDngPEyCXZiClLvBiZMwmJubOZiHryxN+YXzJ2MshJ2EQi
XnzzHmTLNThgNj9pD0C2uXiWBDcb8RgT/iwhBy87MRqvzlczgncVIAmvPfiTUFD6Z7bteA/0AcDG
foWbDr9Z9x9eckVWfJIXL4H3MwV9tmQEfGsQo05IZv4ghc8Tit4TA+Wmm6ZN2lS3x5fUNIIPWQ4U
gN4yoVBPjDbrfvSYVF4PwmysJ77KeOlFgPirZ8pbvCx5eLhK8G4qGteFZMwP0zF5dlVFsYN5i+tc
Gn4u8peGX7A9MrBTEP7TVrajng8m/8kryzMUmb1J9OEHFvj6oDvWgHUwYl4V18nugv9RSanoSphu
oM6srNKtE5MmeWXsl87/vAL5d2FJYxY9qGqvpOzvq96xa/yUZMI4klw1VSQCgMlM+rXarLiJivLS
1Z3Xe3WK0SLMDUx+l4Uso5bLXL2v6SphlSD1sF24F3M1rW7f+8225MQ/HLM1QbmWQQE3m0kSLCec
YEr49MRWjgYUdPK3jyvO37PrYMK4ypSs1grVexFdsE+dTEVeNlD6+rwr2dLgJNfBfdIi4NEVa5sG
nnjjF0zD207QakC+Ast76TdrbsLtTuMoJsgB2T/my/jyc+x1IIglnNYng6DATixcDDeOJ4ZeVEnl
I8Q1QjfU2RARB8hfw8iXQ50LfqH84HwC6jF+p9cc07kItiz31+RfLVxOwSICuF3P9aagHXG7x0Id
j3pdPzE8AwqinPSoGe//hVHEAikeHGqVU/A+QaOVVL3ZLYJ0k8MmEDygTkHgJpb+958Qk7zc45MX
oxExy9iuBeKF0sg5oA6w67P9vjl0+Q3cry5oz4BDHIH0WtF6NSyg+lGBrBgplFNJVrO7h3+MNdoF
2lrXF8eCzmE1vb+mWHj2FoT4xyLjRdkMPgFWxFZm5+oWyjeIwmv+hOfdvBpUy0fbT5UolfOeMyW+
D7YWoYqeaP8POL65DYIXgRXX9s8fHKKGr24twEMS/05w4QMhbncqxfoNckPqeuwc7bDdCVvNaN8n
cLV1O31i0vWCvmOR10USTWfzYBp6EGsLAn18yrSJFThlMcp3y3ZbxNTCtH24jKfY8a5393R0zvmx
dVh49S8w/nG2xJG0rbVGofT56OTB8LB9NHq3cUWaApUF08XfTaU1HGB1BAT0Ur2tOUhHm7kKggkq
V5+w1q1LrpXU+WUFyGnzcumM38jCIFEF1dCWaCl1ws9vrbWjm7uxVkjvjzX1siwGZcOX5uNPtPGl
bz3ytaQl7Q8iwxe762sHnMFXEpf5lDPMwlg75WPb3JPc8lPrytDXJaCZsx7oUzZQQvOiincLI1sy
BA1jUabrcgNrVBZx30gFrwrmDvI6ILd5zTEllEofLf38ai+q2uKo2k/aIlLjLNlZRHkq7kS6iRu4
TWQQW/huDgDm20znbpCzLPn30tSpqMUrfLfiUiaIrzQRbsnRXg+aIA9qr250Ebsr3rPDGg9ZmPsu
QyyFeez6Sz/ggdFPBgHhaEVdcHEUP8NwMpIrf8+Xi/hE5r/5Z9YblfOn7iJpe8TDTBdPXL82IA0H
oshBmSknVt/4VoaOgw66ZdMOQs7IT2iheLdwen7C8I3krV3WaEi27S6e3gjnSlwMK4TDHQkOsYe3
IdYg1a3ROhnQc17mVe8dITAopkDClw6v7nvotQuXacmWmiaFe1gaBk0jXwGJSvgYdGJxWi3Cpr5V
4uWDGdK888TSe5D9KWqLNsDXq3MSAu4BPpjVPCpJEBQ+MKcLsBh0YJOBBMpnWVJ6wqxrCopPnrzj
qKqAtY33b8DC3vo39JD1PMPHWAQmd39dO8UfYHehgjSOTnOzX+zDRcvSw6mm5XmdOOVfY9UKDPxp
/Hly5HKQLSwuYV6iTYzq6arMWr7hjwHxsuD6fAWShiz6rRWO36t2lmyxJBEFMQ7n+/Z5prIAAOuI
Wp2psxx1nVM5QI/tvH+kEtMWyEWJBTUXAWzEhiut8rQcrYssGJx9XD9rCDqYAwXMfgJFT/SjsgtT
xYkqBCsGiM0W3JeYMvX90qzyKu5D+8jJOhrEdRnrumJtpfhqU308JcHyzh8cd7bV0u2ff65PIn9q
c7KA2dR2ISzvmeiwNnmOUI5tz6rTdF4tCP/bgx0B1wyxbCVbbroyYNw69Fqrsstk96/6a3PVR6pX
f++Ntnse2xwR7YHOT1BBuftN2/MLAwMd3nCoTlyA1Od1F5utHB0XxSf0UstdVCR6Yfjx4Y3cm1Om
G2I//Xf/T3d78MDV74WWLvDewQM0ko3FsxYAmTXyhOSOAScfWsdq3ZqnbMFibbtBciE95Jy4mPDd
cwNwu6loQWBz3KDxxarmEJBsm1+8p3RlcsuTQ55quLdS4UYWKyQkN3X0VAx+rbAhmBtdDmoIU78e
bdpfM8bMobMwXDkKRxbSum8nVv6QNwPixl99qhKy0hDlWVNIruczxlKzCzu2BNk9mdvdEUQjGnT+
mTZJMKvSDwkx1NkPVHIgPP/akLlTDOOuTyRDOUt1jD1O7frfiT7qj5Kab8Lm8OtZ32KpZYSCnXyo
+t00yrI4m+o10NiPvkfaQ8YNcM5brWJPP1n90X3ym71/BWCIrzs4f2rNDKzbqBYoFSbdW8w943i4
bOrXUmKt1sjKzvBSfWGtkriJUL/EZ1qH/VgK8UOyjATLdPPn7WF+LVIHNqfTFkroU/qyp23ODcTr
AgsMXTl9ua6GVHaC8n+2+C5V5c/WEbZswTkcXUxiFnFHmoyTyusHM0Bp5VK3Gio+ZtKfjje7qW9U
XocuZMf+DPUrbcornjbMsP8UD1P8NKIgmApd4S+Ml0SaLiy7i0QDzptEOtbSS7Cqixp5ZlZgvpg9
OZrcSqAEjnWr2wn8VDQiI5SeDWWN0Etp2PfsVRfDoOHyTjhBvFf8V7zVx5z+hXZwjbgsebGyKvXU
0KYtwV14OJMekVHeOgsG5LFfo6Dz7tUfLMMDDmSiUYnWmEetPYp2ugEj88fqbjRK/g3sueou6Ie7
Zndx6FhA0Q2kkD19zJ3+WYYnrQ5KeJA4jJSziUp5jQZNklFm6Bb15Li8aD0Ks5Zv8x9dQ1TIVq7S
LiNGgExE6yAnhw7P/sjRTmkwxTyQRHqkLuruY6L03janSnMUjAyYZnZY6rClTPzDRIgpypey13IZ
HdeUkcuO+a40usFgh/5pJPWOLXgaekaEli8V0VQvYYxutGB/8cWunp+68xUeeULJ9AJ4uzqnGs1Y
7jc1Wscm8y1Ht0/5iweErckxQopXC1f4clffMEDFV8sXFFVYjmOFuxu9sXIGH0V0Kj+zKgjlX1FN
YS//3PIJ16POKKhe5vFGkiKPOp1WYworl5srRSMuJ38gmULRC/UaxAA4aHwoMESP0oNz9Zqdf47J
xk9VwPhErepEOiYqgvHks8abq+gFEK9Sd4AdO9VyEjDGD249IzE+yqxrSnIjvSuwJt8hqEbNA6fU
hBIV+rhsnCMpZVozXr3lQVEeenudfax/ds2vU40SQTsdoa5w5101jEk9Bo4MSHNpe/uhs7DLJV8r
l58JdzQNnABUGM0KDaA85rY9B8K9rIcvhIc/klVlB1DdidAkHdbxpq3LEF5URgnQAjs+2/yqe8Ry
CLEPmR10vMK7kRDCiZ/+qFEshCKzcwbe/FzV6SvbHclGFKAaiNQMBohORjgkiMQDNzq6csgIh9u4
2/c43hDF0Jih8UtwUEtRqFB+/nq3hcfh6TFR2hy5+tsHW/Ep2j1p88aiIS/XKqR8O3iQvVeZUy/x
PfdRYa3fWBUg0SMWiqKtqa/GU3F+54Awv1cxbs8mZNGzeMc6DZuPa+FPe9b/rDblDQdUCaJvudxI
ZeWeITnwPNORPOIM1tMySyJ9l6X06+IuMXyKp3AOtST2IbkDo5eXLPnbPeNMJwwOTlnSTNJWMmMf
dFSV06LczxnnjjaaaMFlloJ/5HUBR4ZgHaiXcHBmgMSlOW/IUDY2HVeW/N4MdbF0ynth9RBy9Maq
OXEphwSkUc2cj0apItgMiVhubpOj38R3gg9hWzJh6cuAL5pMgRm+XY0c6uoBgJSFuhgu3wcQLf4i
f86j2fyljjY2QEjcbaGsPPh9ZO3jaOMpc/ympWMJocEkH6dRD9YQYX91VH9tyDTCwUH4ZB1KIE33
T+pxI3iWpBLAAu/S39JBA9pfWzcd9/zuqy3iV6+XOTYrFX9dQuCAjhyyq5qvRN8pRYnL58cKr0FZ
735miWhrP6va3tLYoogMbjQM3A3ZGD9T9RGkSZiwxKUrCxKSQvqNxzYJ9GKZkpG1Kne/1tAb4O36
pdAgfTz0srnGLshtNFUaBGL4cVzEv3OK4N7h0/VN1Y6g5V8+OoEacfqXqA5fXcIG9WpVNYVAlKOM
TmgZfzgs5pMH+vngiovs1fXeY5REytl3uqhxPOSmm4FcWQB6eYpKg68P7eJyM5qY3Y2lXoeENoBe
jmVaUNgaArzhXLK90TGs4ZsZlDfTtUeO9ekyDTjdvVNhRZ7o3PnRWJehXWp/npbcci9x1SMvc9U6
iqHdcTjVut63UiYfZ7uQX1BvGa7Im/eXvkyZ9Gcq2ZF3fyVBt4mvPDZnpJGRpyqiEdm0QxM65CvT
bPGmL5uZuSxelCJPVTVo+j/T/MM+nSsswxdPruA7vAvfZOhGZ5rcsMepsKJpvchpaxWmCm+6rtuk
aatjyiOGB1orqebBS9sARZAynxWJGArheKlbYZa3YMfDrs+DDDbQ3MC0rECpX/3fM594lUYD5CUU
pW3IUU+HAonyEOct0G+8citlrnXXQWLjvoZamW+LSKWwekISFiGFkSWF864jjgfvFOSsSysEoemb
NCgYFeTsUsHsU6OQkuv/1LUh40UmRFXWUNN4er9GUGzHHQ3qrN7oCm5vlASXRgFDUqsWVxIUdTam
619SiYy4xTwAtpDNeYJ6eCxLmDX9Idj0uLV4JpcJnsDolubK5bHTvKx8mnHJAluZ3qkMjc58NU8L
ynjjOquRpN9VsNrQv2A9c4bdUP41qkeTzk3FYLwYM2rVB/HliwtuyJOR3RCxcfEd93SV7wIkmV+Q
K+kU8FA4HbuKZIpNmIdW8L2mWLLSbWcHeB3fyi1g+kdpea3g8B9Lwql94ZGtYvlbqI0ETlOwrREj
9Sa20yMRdjvAf11rwZc96QeEgW/s9HXWpVZRqXjXr6t/Z7UXbtBEghJ1hw2TJ3eK6OnmIxC2pVq1
2NzfQDqhrRg/+PBE9Q/o/JPyCdu72LdnpvxMcMSOB6H2Kzz8CDKk/8o7gmxN9+izwK4ZyShkwbVD
4s25JEP/bkWqBSWz36Skqwp9lu4KRFtjLuXcHE9SI0RjOqAsYsDtzAI81FM717xFTCaQYKaSjPwI
z0B/mf8kEgLymdxNAZckOij4sGN2u10E2Sk13kjO2k4XO74+l8TV+hwt2HngDaFZVO0k9rh0KQKH
eqOYUMvJQRCK/BkmhQGC9NlnFmMA4TBLJeQpjir06YmicA/EIJLbu4WlyprEr9VDEO6sZyQM40UZ
3MP0qgrKjFBNUEq9neGWYQGANHxrZiGIfelbvMum9bwP0kCdTvE0IC2HWV04vDocoOViBT8EcIxV
J1LwjIMWZS1z4BRR+8YVjnqQTG+l420ZETb3LmppfFRc3fMp82BNULgkctcct0QVDxyoVf+gv5JK
5XQfpbYx4oe8Xgjt0GFNTi7XEvrL5P+chLzv4Cp4dcPf97Mkw/tLO95YiZOQiKa1Voiwgg376bUp
NL311T7ip23N2foVyOy8ZS9QNOTiwymYXqBLo7KDjHhSsv9btL/mWQ+f6bTWA022NjKwu1vKrjOI
3ptE9NyvcBpRj4cvlQmh73do1tY2XbdwuULp3Rig3/SvUuv73qZmt/eXgf6rC7ZlZYMeZFFuvpKE
P/8S+qsWeMrcHBfU072vhTXAHOzIvtFo0Gc1iGZ9IORYmuCav8rUWYA3WlCrPGMc+fAkL/63l0v8
2epsnNZMAlVV6Vyj9HDP8CnKvVyq7NLM0WvNvDyWt2FBcx2i/V9+XwWXba7sEoFvcDTyirsdIBVk
3/sPaYEYw44IQP1SEnDbfKKDMJNwBh4dTKZk8y0Vr7Sp/pMcnStsy09LVeLdcUKe9GXsk+lfptnd
QE7A1MqnI/V5MrwcNM6mT9nocSsitzJdvE0i24YA7WC2uFb027BlVwZixjta049Vq8Q5EUAaQuJ6
35fVbxWymQ4xMg929cPKHn2qU1m4rx7xiPdSONxXg6wkixAFq1tZTH8XnEkit6yM5CgeOlUBjfPv
2WN1cjlvFyuXSMxu0DwdSnoWaco7rhDh9ouLLxUNQ7YeZUlC78Eyb28VRMEPVdVC4phx3LL2SwwO
MLq4uT0uuoqsiE7yhn0wqoSFVbF8GiMe2kmFhEOjBO7C3gP9BNN23UmgTZeZ/CMJIlsSn9mgmECJ
vN6G/6aOV/q3Y1+3HpLjCxo6ECmJTozhO8YVniOimr3ZaqFo0sQ2qiFihE8J4/L4Gruwq/XKhQ7Z
fha+TiCUSZJLOHu1kPADHT6Z7G0yB7awlcA4/0EhyLD2QV1Nt1OGjqwyRCby4bgbT33HRG/rf6ia
AE0iTMOv5sHCRnoSb74IAPlBPtS86E6sxrOFH8G0oLutDcWk0g3uc/NDgGj1P1w4JDH4Fo0lKEeT
Dg2JCmhJ9ImkGMMauAZLPvAxomwAXPcEQ1HZTbiP09ZJuHKx+rjru1xgXZc3hEq47E+MMbbzbHzf
bjxzCdGa5JpIpoP/ETcynMX6rIpByRkVhThMG6Bc7iFEaRJboYfR+HFcWhzZKCGZMSNOZPrHlSJT
R2oRospGlNpulfIm9HuOS3S354siS06NyO/g0ZJmcn8k/YrsmO54ofiT/isK4yDY3h00QRtkAspZ
Xkv/Dy3hN+QVzPbxiJpj7FrRa4P3bBnp2shN1/JKwGbAp7mg0oNhvQRdHqxv5sONrz2kYCcvEFF2
D6Yf4bnFXF8q9uB63VnZRWtuQPWNeZ4IPFmsdN5tmvsZzaAaPW/18/qtA8q3X0KtIG+Y8cLHt1fU
Wm7Dd+I+xdUh68AHhmQdCRl5fxAfJ4IIRKy68fknry90I65N1ZOA1sxcyF17ZIyxPARc/3HFXQQv
zeh5k45Q6W6CHnLJYUWCLfmvyJodtz8Wr8U1kMn7d/6nA9LWtiVo5UqPz1CM5eJJ+Ik+7UONEran
AKQCS2jM4FWi8/hlhdMflJe0pw5eBhResuau1hzgZi/Akkst7dyb4lq499RWam61mb3+3I5bEYUw
NzMCSmWESvEbsruMWnhu5ZH8uhEpBwHtojTyhvjPT4mEDbacnRyG9tiwjbhtWaCotle6UL80RJr4
OkW5j4v5ipFjShNtDv6mpOzq/aHs5F2q8MdHpymZ/LAnFULfur/Unvkk7bN7nDimU0UcGNsErK8C
fmg2mCY2jjxNUAXcKPGbOhJHKbqqu5/20UXy+/+x4af/UNITXVnoBjc2Qtrgb/GVU6lw4XeYePyg
b7s3RrUfd3XUuUVL3vJtuG11EWKYtv8dBgOt9u7y5AS5qgJuRf3/LuqGFaOTbKDSAlmuFL8ToKKy
vLrGwPFHgalL3t81p/JWPnF0J+N+sbyIJTn3GNY5DCDbHZexa0kO1FDjnnFSarCiALojuMNp6iYr
RrBOkRcV7oKxu+2w6HrcylQuEbXFja3uAKn9AFCAoOMkYsovEimt3apDkdNG9UJDv+Bes0rv5rcF
WVCZeLzkfmyu1gAK5dCIrjfz7c/lBZP9jy6WzrLpBsO00d8Pqc6L76bKFZ3eVukeC7oOHbupDJ85
wxEJ2WfACPXZAcLn9Bz5onr+sLgGlrhivHI2R/W6tKxUC5Avm3qqYEtbvStvre0pU8Cb/vXvKwL6
1JsBzMM1CdyVVq6RJp/rzpVXQyZtSTjWKCDVhW8eQjPJcHUQtfIWidNGv6pXlb52YGjfOx6F0miM
2CVfd4sDhJahUt/rI49gfMhyUHDrVCeWlKJ42nDtzi8xcVb+kvqUv4vemYL94NSWsetYp+y0/hrL
rSb8ZhRwevKYWqFa6/6v5n6SpCB6gIGR9W6m332+QjZ5SJv4r4Ll/DiFkQ5ysu8b9PVMTZBhsT0Z
3EBrgk5LvFHrCNtI0DFqgqcLCgFwrXys5tZkLLFKn9alskNPH3YPN+eEkB+6kLPmeyRBpM1+DlWW
ywMZLl6haV+K2fPbUvMqRPHsgtZrCRJ7VP4my/pAwZADVUFU0fNMQuOu0YxVaPWHEAvEnzu7JCxI
QhUhUC6AfuoHBBsf9iE4jcJWnKz3JSAhQgFXzwpMsU6G0q+JHw/bjmwkaCVPnDpWtkU9k22g/xCs
NczEj6F8VITPgv08dVCoSN8ySEdAO15jUtg1ycRUrn/Jj17fXsW3WF+rQSdtH4LwSjdNOlwKK4Ei
x68GkLttJgcIO7bkUcxZe9bzRlXqLJTpHa8lMVVHQGbke2diEhRgFqrTKf9eNn89B3hAktKs7Vlh
KHck8AHOJ61murpgIXrbB9kKO0THfAujwACHw6Aaip3hOrotLDSDWkFVZPg88YDlHGRolmVd7/Y2
6dhadcjjyxrcPiQPDIWIApDrOke8wNOEjyqPKhzx3nQWDmwFJQVqzdMN146cvqxgyNLPx2yALY7I
r0ly4gUyBqbxMzQ1+FUUue0r6QkI2JRME0wP8bYHk9E2xL/xWeGo3AECyizIAu5Mr+RBO7457aw8
2VB0C2ryfLXxI0tq7+o/jRoUM+viP02HfeiIFxYrskqBQMLZu0gROYKlWnN8EcHl9CmiSx4kEAI7
+BWjX4HuqWfodduvWpvKhd+m/1YWEDjHn4c+9wzUEGYGp+xekAHOEUFu2kaF1EpglV4JzXo16Prz
H4e6OBeMIEZt9rKceB6I+kGW/6FtYO+G6Odlxb7e35R6wgBOmmJZRzVbV0Qn/HHEnFvN/4GV6rvh
hsOgPicuH/G7PA5a3GG+4+XZ2TezLwN/Zf5W7BSN4qHvxGVCLflf4LXqvwSlaQJmJof5VJ7jUonY
tiYs2C8dRosrdL4k1SEeH4lrneq4EesQ5OsDl5MuUPhOnPPTIuTh1s+5YbE4+ff80QefbmnKLnuo
Kp66xxIWU+2Z0NRMmhjsZExZpeZGiawtwqwgjEeK8ZkSCpYNkGerDFvWLOi1tu52W2e8lFLLAhfk
tcewv8/C3MFdRtq6Jd6p/WDq+A0RUS8CGJeDmgGDgKpj1tES1WeR1VzhNL3+6JlEbssZKxQHaL9C
u/73oIvxIubb6umSmcMp2TF3TkDIS56w8gEoqWUFPk9peL8yKXZtcZ85C6afMo9m5EExGDNi5V8y
7VaNTXQNnGuZAK/cEcn2O/OoFD1cXo+v7ib31tgujolCz0enQCmzXylfdfkM0cNcHtG6sLMRJ85b
my5yCC4a3HwTkEIjhBg9Vmgqo/wHB4C8DR37+iMS7Qy26ZFdetJ8E5LwQLEGs2850ryAYlF7jilY
srcdT/UoByceisJgbemgNftwhyDgO610dtEC+aMUKbRy5wtEWU0sXr+myHe1mvbOkn8vSrg78qoN
KIJXkfKwyordFUlCtZUCl3wZfBNyXypCFMSJyNXO+k3g1A2U8QckCT9G3V3XXAw9UfM+xaqm/k9t
+SqpxwasWWfTv7Bl/G7hGHQ0mq0FhBmBQUp9c4XbsxA9mX+EEzHy/zFWdc2AIVkRkipQ2FC/1Ev9
lLJeK+Yc0QkGA38BtusuDJH3um6ZEit+qgmbL6KHYtgyUigkM8e8uTuGwjym/5LevlGLcEZyTCmK
kAe7vX2Jwo2odw6UWVPz4VsUL6hCZNwU896xIb7Elxm6nXyuGR9y80Qqh1xgOGw5usX3zAYxP9et
N0bHuL4HM0rr//M7dHRP9l5PEQ8N0KSnPw9KwDAFmU1FiZIoUZxHgyJf917BIpnXWQ6waHdE/qap
gX48fR+meRnxLjt7/e6biOD5IshZZBildGGe6CNSlN7RS98eELQxybbdLq0eo/EiPFOxCLma8tTM
PLK4MyZNjyUy8kKBdyjpx4GJ2KEpO6OR5VbC78mJ+IALjaYAlBS5K0PuzNPiE6w2vqvn+K9snnzF
XmrBaUIWlSnl7N1T2xjPmMeCNRal4GakhDJg5ZFismkpcA9BYYQJoPSPGJ1vmkP0RDdgqALHS3ws
rs953MYvgnQMWK0saeFbD4O0+Iy41sxFYQN05853RXpjO3iM7VE46dlX0Bl8lUArNgT45AbO4VW1
y5rzxSFXOHjQupbzJqO/AhUAjEwZW5/xJlAr38SkavA51jFHiraNYzTGFz4Wkn+wVfv5LQOSr1xj
MaCIMzM21JUca/FrQrq5Ruo1cWubhr/5Q4rqCdQGho8QcMTE4Y7nQryK8l+6UVjoPYFjTkNg68ax
hYbLx6azhekwslgRD0FIO7g5QzYbQzbTQJv5/zvQ89QAgqML4Jdmf6ImnEpYTvrFAtsn43CYw3RR
fitskJNtCYZGz1spmjPTuRprxOuEm7L0JemtzaUJRctfhtX4dVcqNnn3TcXEn84Rgm1iEpdSeM2q
NOVjm2jE4M5PhCN9vw5CG7iFZP7LIXdNy7SGel9unviB/N2qDeGe/YzEJ7Te4SfKygquJ+oZNkoM
mL0sg/d6OwqQQyOJGsTaOzmZiuQC5nZ1veZY/76k/JZI1fd6DGOJz6wffnaVTWRan66T6eVcnbhG
zGolCKEtAALtiuPcI8xL9M/kgUro6/Ovvo/0gz1B1CisBk5XmHNeurqM3o0Jq8sj+nFWl4OcGOPz
buDJ5fZpw02dN9u4HlBZfbkJtMiGCxwVBp+lyQYB2KYPE9KjDBaVqKa7yE4jgrh5cOl/GfkJ4HgR
OogSA9lnQfdUyIsINdEMrz70coJaf8UuDlIkSYPrjV14xh453vTF4t9UQxnY+ZOjCNitwxXbE2Wq
q3ZjjTPWwBdgaud+ICvwI+JQ7emipgwRxbb2c03+kWo1ZpkYsh25siyt/1RZQB60h5ckgZoQJHi6
r7YgeKiDpSO/FIgDf4/7Ic9ruUVz3I8YGf4Lk501RrDHAwnbXPgtAEP1+AyKz7mHzvP+1CnVccT5
PfDOOHeUk8p7EO2HTdECguby3SvsNlvVfMtcMCa+tRCBuLFxBv/im2pQ8lmXI4yjBNKigAU880Gf
N305v1TrVDSIlsTQwnbpD+viFJ3PvZ5WXlap3e5blK1Ngc5+jzrg6e8oFSFGehrEB+5O4VUFIMPY
aGewBuyu9ndTd2b/NJsZd2En+V3RIICNP64e3787D1ZHBYTjSDzVXWT6lNWL6NUWD9QVaHwrc09S
f5tDiQ/w8wsAfPV5PZcR4Doy80gA6Gsg28h+/DZkG+WRrK5VYa2IlDHs2TJsjA2ZU53eAHU9hhlP
JDdaC/ChSf/IV887s2638mewg5AK+SnCQhQ7V7Px6vTwmjTQ96P547uoNmf7/81oA20a52DmHk0U
twfuhES6nCC9gEnp+fZ8FkJJhVF0wseEO+J1AVTT6RJNo1Zd/THcOla+FeNosj0rZMZGnmdplJA2
kpc+p3OIrSK9ShXAvR+g629rCOtFzCwhnA3heRqA8UETEv3Jn94xA3+5Ndoz4gV4/y+Elx5sXfPl
6xX8cdF+3AsC+KpRDvCsaH/4ntH6rdkWLDut+G5dzUD8Q+85PyV/aWZGgJc9uLeUTIJK9JfRVXJD
qN3cy8EzKKF42aqRgRJGpNmoOeRtlOyrAmcn1FJsbJJOGt2B2mKC61qQBGzj5uPSNZF5Qab+G7Ww
Eoed3pZIAGdkAuiLTkbj0zD3HG26Y+fi5itIZa31nuztgH3/CFSaq8pDiPRseSjcNzVel14Dekfu
oFqgM5dK/TORBSr9VqoCTdhC6Y5MBHiU67c5XzyiuEIP3DxPPBCAsNyk9I9WbjH/SfQk2JnogyVM
OnHwCZ5WjS2MgnMPEcoy83caTXSiqhlPaExl9YDuOjcE84gL9VXSOZSfDUNZlH8bum6PpKr2Tzpq
gUkPG7mrCZbkou1UpQPidyB+o5s7/9vdYEr6FZzLxN0Ksv6DViX3RuCfsVZfqsMoS0sV+nAv4KM4
XFblWRZD/E/pd4rra4QO2sQxU/DhzBhW01ZSERGkYS6ci3xl9xz0iqNl873bX0BrYA2Ma9VpnG8q
A67sUBmB35+TsTMeje32wOq2NsoGSEWahlZm86Fu2VQFYUMfdDPZJAx/x/bue2mWZpE1scLfnueE
ksXrxgpBb+vU9+GHT01qZphlWwDV2qYM4EEq5yidPsN9OnORIX0/BrR0fKHLmjYR1eQSh3JFb6rC
RJBzBspwrgbJs+fEUEWY7/5WOdvjQpQQd/e1GMm0bHCuwHccMiB7V0VB9DkD+AL8j4L2icvvKgx7
xSg2VVm/graoMZgeEx4vccCBAjbhp11PWsC8A/KyyxZR7PVFB8i4xYtdPOTrHwNy0JI5u6VTgirT
da81YJNfoj742H7vBXjHgtoZwJjYV7Y2ti7wTlzYEuYQLTs0X9euBUH/sYH+znZgA7sIIPq+e9jv
NeGm7PqaJKh3sBJffs+CmGvR/RWHogCT8FmHWMa2UHnbyYPoBgJKTwoQNsfaZAr4mMA0H+b85Q8H
OxyXwm3Xdor+jtDlvusJyocuQTWPXNqssyPfhELQK0dyC+/6/BIkCdWJnFP7LkxQiCEpCP/c7o5g
YFApk+X6BB9XODBkgnuVeoH56zlRhskcJt5J8nc6Wm2EZXV1Cn5x9icnR5IxYVaWF3v9LjFcdnaf
dtxntgQQTg+VN/S1zVEeqizoo7WXyr+P65mq/U6DoYjmi1OmCvpk+srI4cTZoBi1N7ym/va/AthC
zVIojQrfynNIixyaB4fV7dB6u1pWNO3IAUXrJJteJThytDeR8m4IJQVUwZMKu6LX4AKaTO3i8Hc5
8ZUIQQKynt+B5HwONQQUNgwDpbQ5W6J2SaNTzuL1nWdOK0JTHy6EZ8u7qQE+16L4Aw6adyYeLMSL
OmUS6YnfOTiEBb2tEz6Mh9w9kMpxNa7kzeaUZJwmfqNyo5nrWrJnt7lx9+MIgN3TESo4WGF8gLWG
VqQyELr8nutqqWXGBUPoFeYKSLY3lIuymfsgfdXbErfGUYOe89wMSBQ58+JHbTpaQV8Y45koeyaT
oJ2sYB7mgOu2879ofONVZWfsLvIlycT4jSFz4EohZiFmlSODlQ1/6bn/Z9S7WtaJRKN4NzZiCZtg
b5XQ+h4u7TOJchlbGLnmF5TuGlQJWff1gyLCWeHEcOP6l+A57RwZI0Cj38C9I+5X1qUa5bSHmtvm
rLwavLT6LvPQtfFRIfFTRZsgSeF+kzEoLgCK4G254ZIaiUotCpKa59NFD0+OT3ZujGbRrsSHYGzj
4ZIP6pdstRB/m1Ms8Rh1E0nv2TQgKrsq1OQ8bpzHEjdwuSJe7aQz2qVxYKR+1M6glVFmzB1w7Qan
WRxWtHKQ+xGBOp+4ctryGtSM/fDz15tqq++zwPCqmPVfB+iPM98szTyuTaz+GN7S5cpzSyU2PCan
JkaPW9vm5sv4Y5ajSQ4HoAC/SDOrYxvVCcFtcrvAV9H6RGOnPMQfS/bzVNCy+czE17ewyJILVOD+
o9y8qNVP6pypficsgwU830ppITqL7gtb88cNgd9+jPpHqnYbkcDZRivLnWtyP4bMWvbKWWhEKLNC
KgK/RZXxrxg+uFH7nNmNFqndgtkj7b/K43GVr+J47P2AVf5y9hhK4lF1GCnjI6bGbT98CYqqTI4l
RyJ8n4v/6Jm6EXL6RbtQQGdcJOlZeC+rkHouiZqr2tMLvBkVVCHsqnplqG2u6MJ7iLxgfVi+ZGmz
S/n2n8X0jfuaU5s3eMsGApXP0+ZEcsOBcyhqa6UDh35HXhrz2ImDU/r1xylmIsYZ7/wLWZhlrHcH
ADwXAT6/PU0gjtQQwnu84Rxap0+1hKs5frw4RKh5bGmfiuf6m3RzggN5uEtTV4gg2jCfcVDuLLkO
aX+gar/wkeQIg1VRbqGewi83JgjdPo3mjO/HzMAuJuW2Y7BBrB4/OtNgFjaN2r4LYlx3Dp3AA2Ri
doKc+nZz8EB67h9f1xRYNhh6cykroUJzJ5qfAPQBVddd3AhqaAoUunjnrVO/wGzR93UIsXj0F9l+
NxuI0FvRrKR/Z8qG4sX6tI5KTanbnyoQwvoOYBX+8YjdgQaNkcg2uRlLlLQBuX1mIyy2f1itaoyQ
q/Yir1+Ifb2vlFauvyGJvKzzKiOncqIClt4dejhK3gxGCVvROGMYBifGzr9HDfJLXsCFumSy6H0+
DIIAPbbHMejNcHir/aRvQnGbrPCg0MbqtCJJi37VzWfLgjgLljfGeX8EYKfvNNYGn3KOh8RqbRA8
ht2vLiB6+f8ddj0SvXtqQc93aYpET+AYdUizWxWSl8o+z5H7l5TXgDRYGi258fbXPPU7ErzlDu7e
FiMi1v7WWSJfcorSxqoFUOrvCWxQ2Rbr6Kd3lfQ24KfdoHyHDNI2AyjGdBjI1LqWUi/1aDfk720B
nWWo8GvHLNPyASLAcZhPymmmq7HZ8YhANU6baj0ZfPw98KEiNstcRZEOqE5WszXOg9r+00I3jfCz
FnVMIaCdmcZITUQeHyJM920S6NaF5+FGlgepUndhBcDOQG5FTXo8ixvgvfztli/wtzZi4SPWZVRx
9F78CSo5CqUnikdZOFvR60P2gZKk/kwzSyrWF9kWT9FSvEyACoNNhlCNXDS7VhcavF9xdPFmsZ7z
fr2bvEZv2Yusvu6f3NYXTmbKCOx6Bo+1GBVCjIY24ZA/zz9P35Zkw90AOdHI+iDI9gDYYTmcSv+1
YZXQk3n3gk1S23E93TbuXWL3XntmywKSiq3ZBGyfz2r2POVCptzAnjjEd06Jsr8ShVLGy5Di3flj
00gHMazoGUESonaI9XLDAa1bdrB2GyRdN7L9vmmUD4uzKQ/mQJxYMeVquAyEvkTqIDOG0HtbwkIr
iN4ny7sHFKSLcXNzJZoowvzKqYj7IDayVsCo/XQUy/Bia2tW+8ibAl7X5g9KF0yUDS42QfN5NNn3
S76cpSnF8kIEfhsCDNrqO4I3kkJFUBtl1s6EgPtCYMsAAK4KKW5FpuR8RDJ9S0BMVgMRmB6ewsHx
sUUG/h/+NyWI5LR3v0ouUMK4Szq6QUimu6B0o9byHR5bv4O6DkJ830HQ6eeCxpVJTOxCwJ7M6zig
nOnWWlViuPQWM2DFo0lk6tYVFed6Qn8gYzDtIdf6huDxT8otoVM9jyU5IXGY4hUWRJQ+4WpGZKsX
9FoXiNbwjHWtiFjpSgRbt+5MRwCkMHW8+ARU800lV4Mp8cqLjuWgvgP06sAepNHnXa4p7bEmRYh7
At3vjjAakno9Xw79a55f0CFs1ogd2AyjkJW2dDn1/n8qwmlbMyEm/zcWUgO84SVSF8GgPgLSXUXl
Q9Yiqbu74L/NMfeLqqbeud3qv6HelXTQ2wVPvAptIlLb9tVpuMHPsnezj0AjwjBQGteM/TjCVkCp
iv0O+69gJhigJjbHN4ChqWVu1eiuZuzQFRWFSiV5VnLhU4cyMKt4GzfuJg5uoNUBynd/xhfcFq2P
AjP4MH7MdVxbpRSFaPENt6Me/3v7s5Eqy0vWXNi7uLBSI0QxYB0PW8U9z49hWsrFFKTRIW86kgAa
CyyrO34Qx3cVglAvf9LdrN8L4rBjeiC+bdrJd441rEyUVuHUfF/MX+C5Zq3RqVI3wpi9FNOv1tpP
d8Hi5tQrTXyZf3YuMXldvjAl0RCIX2P1MrRGlD/awEG+a8+3UJxscEf6oU/CYn6zx9JBhWhU6l+G
3XZmRQsybAhgjvv6m7/nzRQ0t6mxVptTjpe607XX9v55J4b6CybER17jGQtWz+YLCn5Ds/39fJsv
ZpW5LkuOZH+rIVUtEqBFL2Ty9w8fn2upV2hDHVif/8VcWDPBWSrYyJXbN0AZA9cdgfKplrjsoSIr
zRfgC+VY9gCZlDGHvLYg7Qm2lYw+KIPKbZPRxJJcowpHM1Hhs9nDe6WZ8vvS4EZ9CvwVZSNDWS6b
saHuhe0d3sAWo+8RFLI54hSnN1JFNHZc2TY2+qY93hLfn3q4+5Cn/NxTMVr4KrW1mP/JTC3kJe08
ErIZOQXlXHO0sVqEZyqu8Srn+t+21IuPwyCH03qhmmRhrNvuUlJScePBiTa1jjLP1P6hgj4/h4Er
RTiMfg4Knh7K00B8B/1V/7NarzzdFKqX3/IVL3BRPo5dL2Tb4lT3+/W1xpyIdETpvVgGYTEoXq71
FVhoJD2GIES2qSHnXrZZwdd2ThY9h0kUDnezuMs7ufgY1QnxWhB2EphZEQvO0YMceGz8dd+/0CQQ
9LnrrMpPJv3DFNp5iVpYCQ3tm8cocNfI1qQCnladioPs4lusuTa+WffliUlz3bgdDA5wP0QA9S5r
ZJUW3Qygicf9EancnHVY6Lzau8EG3I58w6r7709owRnvckAsZ6DsaTIsA9ENgCH3APXUumbam93d
Ut0nt02l++Px2/gwAVLE6kvx6jr3hu/5iaj/ybqcGNcxvkbLgzkKehtYBjrsvQBW6tnFDfnIOjRG
Io2pDOfDAwUzJ/XDqlmTfeTEAcGGSkivDt2txRBg93bh3+aWb/B7Uz1whXGtdIGEcu5t1b+8yd2d
drKfHPgN41CKM3X6AignZwLZAR/mfei2NW2Etvv91kAScC2Dcx7ua7ermkQGb4n9jsoh+7I4fj50
tqGy7m3p6uEPyUfDMRmWWTt+jkcVAx6JNg7kdltEmTifpKJlTI4/kkr4Or9RX5PdLQg+SBe9pNyK
JkpZqJUC2S2J2D+fuow/lAZJ9mw9N6BzHFSWsiAn4YYAtppWoERXZTUfXdGOHuxoQpKZGeIWhg5v
DjonDNpglPInBPbGmei/rAFjpAVz+gdy1Mi6eZ+vIksm433Eno3eUIJ4CzG6DXsNcnNbk94HafIL
nL0Cr2DPnJFS2ZYCumsuq2waydlATPHLC7GPQHNNDU1yniXHSKgLmyqqYuYmcJqtO3Hcv14DgzFQ
vyPscfd8t7hGpXbMtN4NkhABShsXkpDOdQQ0nZrTrF3m5z0/i8ytas9br4Ce79dW2d7+PWGpyu6g
Nam55bmmUIwqm2u4vNosItHBSlmfxVMXb6n6W1QAp9zK8nYljoqlL8OgHbraQ50gC6YCSoDjSDbh
GQu2autvf0bVZlT56R0QWwtnkiHRhVVtSNji2j799KDGaHjIn1QEU7oxrb3gOed2C5kodKFy59yk
T2YGKPiSUakAroQutf2vHf47u2GaxiBpukvcbinriNHkaDnnoIMgdtbMsWlf65NSDsRoJpwj1f+Y
SenR8lc3Ur4huk1tM8pz9aLanDKYSzpsj4tPMTeavPrDoD78gz+whQqGUk+RdVBVqVbRFn8urVR9
fSvz/m9DRfq5zZgPGK8E1Ac7OGSpVZeUNwzfiD46g1BlWSmdB7dLQsHG+0NdEW/SDTntOQ+x+qKe
A6KPBn+7qQ432YH/fUhDdA6nDANuEcfU5aw8NAn/MwKMhTeF3dB3Eyvg6iz/2MvY8GEMDp/yzE2r
s/E0Es8u+I+kcd/H9Osfc6nmURXhB2puiGrgpZdRYAIYOQhcSYOwyQ6tERjjFEwWwT0qbwH5aohz
yKHPcMz4If6ipj2XlBOgFzTQ1wcOw91HFQMhcaKcXBDS4FLrCdlyLuZVVKQ9Gy2eEpC6+3rPaktv
lQZJkH0dt/JYwCs1jAHcllDEXgUFN/IoD0svpCO6NQckZctecwznvjApCc7uv5pQBDUoptkNvMex
RExJztVWLRZqN68WX6web4KRXYnqiAsuM5D5heWU3P1/gRsnB8yZN6HwvWNCm2X2mvfnKgGWqqen
2mXcRxK6YXnjSSbSGai/RlXy8zZr9eREjj7YaPVise6wHpHUDSxgcZ5A4Ba3UOsiWlrW8o194qYH
mvwEZ7HQ8IIIw7NBgsqXZIIDs6+uNhw+LFPZPNJaucyt/uqnUnboDTFuECYAHiffGPo0N7IFmLyd
EuWMyAuql7KtgEMqTsAJ/RzNSsQI2+dOu4bNqhilDrBULTLVoBFW56uqlo+luVH5mpH502oz2iEH
G4haGcnSkIedazEUqaXyjwVkuHcJRZqfe/CCDGZkRRZIeGnDJdRZ745trw9SG0TcGCAMwtO5n+Nf
kjD8XoonHtJXQlzZlivroHPAQWfXwvJgS6HZS/gZOtHIQDCcPz7fYPvJGFrKxa6iz/RY102Y1mje
9zQSjIURwj+5fmVKqKcncWPzEO5DkSaf+CA2Wy0iMYB6BxEZgPld9xOI18j+S+x6LnO0QEtA8uXF
PFq2UM3I7UTmDV20OnAxpFydgQCfcvauVbeO4qFQuUeHvqK0zLjs7J5yiMnnnSuRJHhJLU1EgqlG
maqoEJUJjFvDy6iNcjh5FymkSjggnMmP4vWc/chKKaUhlBTiDvq1BO6J2Fr4dbk+BzjCY6rc3EAD
71vTMLnaONw1S+eLoEn0upoYoo2cBM7Yh4lGtexQCYcu+JFVgZdwlRAcQQ82KfkBLD3WroE+d8wA
w/NUMful2KEreO/UdRQfhnu+lgFfcgAlk/Aa6dsqqO56HyZApaZITB/NkWRTqubSs+g6c9QTftmW
fpixB0AKK1GHtUEDXYkAxwO+SNR7Lr0orGP5NLSpFcUPpLPFDsq5ENsStC2NfmLNxfSqOqXNWNhi
rxOB3l4wVF2Vg/WMDXU0HFRQqIQWuiKMSL5FJqm4Uv7l5O8Zrj71ShHmWOkz/Ydor5TgJpuVIFsq
r9bRWftHnO4dSQqsQxG1FGjdEzu5rUrYBObk7IN64T1nmpxCYHw+05c6w3nX/1/m0lhw5p387dEW
ljAVatBcOndJru8KrCxfY7vU5h5dagbUB/BaorZicFjYocqy/zPIkLLjoFRSTESg/5TK2hakIl5E
TFnaDWPySovlRV7OqShtRQelGVjN9LGFjguhuun/iHPTJubVP1nadG3gDBhi2LqFWm0rM5af4Eo6
EsYhgga7bNMZoAGFRfVNjiTKMybX9bAKGzT9sYPQQf1sIwMDOZZHU2eXsAaRA0mNE+JnvD/xQDmE
uZ5QiTqdFUVX+1doM/q43GLhdswzx5tlowjcvDNHBRGTvozSda5XTXPE5Qy3qDq+zFXMcaJ60tH1
YfWIDAhgCiJI1TOgyZFIoB43Z1rSMYbeI1zuh4/IhsGVFLBLPwkcF13jLPDJCftLr0n9tdJ987ma
1mV8TJJhYUrid1PkcNvTzZrZDbC1T6x1hULpO6G9NwqSxKLtYNZ3XhsBWwAoMtr9imygPsS11mDd
Eoey3eDvt32Vdsy5fStzq7Q5qMHCB0wHJtCsZkxthnWbPZs+692W9kTBmeRBIYNeIpzeWkbC8NwF
RT/t3jd4IKcKyKyCwZ+flH65aJ6dtsdfVFu7K1f5oVPDBfAj8QqHsJ0Z83JXTnFP3PI69xyCriXh
JWU22Eu1ihJ2ay4ndcMeOPo/29FXMNN9PqlEvRNuwVPBnQEHwb5VoHjEWU2Acad2ZCqDvuBppV3V
f/FnoGOa3B00An7KRVc+9sOFfaSZEjuL2YpWFiP6KU6QsKFM7Kl3KYnZp87+p6jsk0NUOhdb5C7d
y0LIZ6jb+331mqgGGVP6vHNMskD4dkFfd6q8K1wRDorPOXOTxukIMJKgR5dDRtKqQjeuvi4t4QO3
r4vPP6QRF3WrWbJEtHXOEoyFnkMaCyZzxA1/JN44XrX9uCxWoTKbqzYILYkh8DtIdd+/dquWzLdr
ZsQPHUBNGTeYJ2kA/WNf4rcVkq8qUFXkFehxvCfOXTb8nBmblJt8HBJfyK+UJnIxd7BeU0EJcqgc
HRrPNj/DYApifUjXjBUSXwpKRK6foYSoVCKRJK/83/VImII9qLYPgM/omhfwEbCnY+p2JOKAeUOv
J2pAromUkSJ8zHmpQiKPpHxGYhIAv4NhFk7KEcLauUvsZENsUPdBXnQSbaF9HzX231ElZdflNiNT
4jfQeN6BwiCHywSG+drE0MKS1C+sTnGvHxzMQ6MNNiyhO4w3XEerdweIQeeJAQAO3dl4YFMfN9tN
9SVHXMZ6ggPsxoV4jdYqNnFoa1aSkKiNufZSC0iHp04CspH8axmRnLmFFWxxMxaLBpx2SrXMUGFc
xU6fL77O4l0NBbqV40FkARuxkPc+v1ApIrrkr7wWnJB8rPSybHHsb+Qxoulob+Jcrjs85NmPhjNR
hCyKvJ2m84/sF2Vmdjilfrmx34Jfj53g26f9ggxw0CwM1qHLbWpuWTgcYEmJiEoZ4gW2mEqsqASV
WUYGSf/afW04S9TdT4wrnO6NWVzpsgZprzDn0n6BoodXlFZMYrVWT+stExAYxm+bltuf6f7/Grax
OfC9V8uwVEWvrLQRSCWaXElWJAW7d6odxNpRQrvM8CFbQGO00bGGUxF0GJ9OdECOkR1pD+gNpNms
xtMxf8JyLoEEBgIOiFr0UW3QkA7MkG5Wd6B5tHA/FM4Ey4r2/nXpDrDIOsFA7+blYMZHWxcgWyQ2
k0pH2TyXqW0SD76/o/p+59GvoiDw6z4YHt1FFUVoWMi26ETXW79S/eviCYaCoMXZeEY4lvWAVZKV
AIJZbPT4QFJhzGCQ/qTGDQWjq4K7z36J5GDKuP962jVdyhkshInYRRauHwPDxr6BZ0nc2JkfZBro
PE4ZlzI/cGt8BjNAoN1a+FaxTCBjcVWAx+kudNKzsSAI/bTMeEl+gJIKCyUOCjaRUQv1SpReg/ze
S9ucgCKkyn5sSkYIlH+fNzOKqU76dNDbHkJFqBMq5W3YbnuXLAr9f50f8K2ePMQ8fqpGYJMWQsQX
CM2+MaVtI8b2XfzCM9FYkT3EmaTUyz/wjDtviHbBw5qC4VdQYDY9kWenhJNkuIIimp/ygqI1kVRE
jnBJBzrJO943hQgxUf21KRLt/SRBEEEAaA3u5comb8639rxY3Fx2ymgJLBItDmCO5CDSGzLJNp4W
WTKL3e0t6DzL315vAifPV+iAEdrH1ahZa3EUHr7OJrMpVuN9Qw1svepiXJl+tJmrJKraquYWqSpa
c0RMr0vogJpVd5ZvmQIDMoKPy2q6wsqp7JYpq0HN1JZQ5fT6ZjV90kQM9wV4Kkxzd/bfpQv0aZc4
dnYwl6mJFmPXHWtTd7N4KureIkh4M4zyLjrzpLPjaSfqUrudPBmUNiPVIhIoYy9eGr2y1jB1fwEu
6t9q1t/50Ottk9gEoE/wnnwXGjxX4awbX9trungX2S74I/lMx/WvcvW88yaWLJu+MVQ3V9UZvBwR
OwD8asjbW0k1nrPvE3T0sl8onfloVIDkrHe4pIcF7UQEUW6OKy8MUMydTTrhhC47CrJv6DMdUaJN
fH1DMmLea5+t2z2+GJZAQWjEzJ0L5ZdtTdbZ9tpryAjylmOAN5h27T8AhERvro9e6ru1jh+P+gcy
ykKwBzrvOBpHvMScuFotSYKKcKGg8agarBLHM2GDuSwI/jNp4waDcuHDANEyGOVr/z0OB9I33C5H
ywGvw/l0eZmhLz8PLhrrYUOSLe+2Zrl7r18cyLAw3dbHbx2nVAMEX6AVXGi3c0T9+Mi9SwIlXakS
zk0s2+imEZac7XVeIocn2UjvOx8lDIcWxOJZJPeVU35FoRkRGhT4cZx2Ay4fyq4OFjq5c7y3N6N2
HbrkQhXCAUuMRlfHCz1iYIJMH6qQZNRg749dxSA1lYQDukFD6/p9a+TDRWrleiFNnFWMulffJm3+
lC/GlF9oNMA9j3Y=
`protect end_protected
