-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xV1iLktdF/92vYjv6WDkJCbZ4QWmOIKlRSrGfggDqoCwEZOy28tCmL0CKgi2bH8+Ptwkf6/Dz173
4ZYrHMVnRvhyaU9NqZO8+RqnYD8lQt89oWSTK914gzCSQHhONL4ZRC9Z2jdoiAlnM1K8QeuTylGC
FSNN0O+DJYbUBw6EOFzbDJMxOjmWLnwH3u9sR7OJdCbaNEFA8GZuezD/802JalcfCl3I26LW3UXM
EowdUWf0ltjiiAA4J6WzAqXfL3E67wl1igZPRqxzjP9XL/Ytuk5tHFWFXOYwC54sX4GhZLFMSVkB
MhbTnmUHgc4IS3cmV5GhqKrXh9+AvFHSo2rjhg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1680)
`protect data_block
yUtRBH8Gl7k5bTgUpd62XwOfLhjbvfolOFNTJDSNrDPJyW+bvfXvSnx1kiPzDT5M1kDdGD0apVby
Ta5TTdBNK2l7YRCBzIpJlADeTnnQUGn/AenDwcYsmCOpBi2B7EzV6f72gXkQNYeWo8O34n6hUUTj
YyB9UlEbubsiYV3l/YGHWdzK4kYiW5E4EGUOzQCLsGEdqmWsahORbYtHhbh2BXER7kVbpbJrlqy2
LH7OzkLEvsgBoXruWGIss3kmPKbBRid2wF56H1KpkhRkTvkuyJjDecSEjMo9vHKitt+qF5Zu6suq
vfyMoTkE42kxT1BEilX7ZgIYKaVdRMsPn4PxAgLC9VP8Y8HaVRauRJcMoUFxj3nkugJof70XAMs4
EXCZl/hsOLYqLbsp/7MP3n11wpFEeM7KW88r49nOpAKWY1yaCZ1LMY7L+axGhz1qV8gQEVep5OAR
r2xVQ3/dyNISBbS9k0hG182xd+kbpmR1gaa22mF+Ny8MdWc0BgGfDFGoUx/XYm4BFJlLyEOPcUPH
C9t5XFs7b/zns70xVhEOTN6q5iI61xqUXwiI81RNaXmekTVAL0krmSNxeed/rNNnfOtcjuXfvqex
BnVqum4mGLOfcxj0GholBnUWfWmbbRgdEbPJoEaq2Qn6GwGhb2s6JgoZEGuFrNAJ7nzYaMl2vlDG
QkRy+PqwfaQ/OyRfUk4ScXgUPFG7/+UU5nZnXXS7cfBlRqL5UjxODAuTNIXX7C7ircXAZb3rAJxY
h9sDRfV+7gaTWZ7Qr5lAHwj5eSSZSfndX83QfdtlozAnoHjMjJdZC/P20NffQtiXw7tF3BLwYzeH
yL4X2mi66smIrbqkP0YvaI41GoDm4XwomHCg9PQh2D2x1WKxgKJIP9ZfdgXrZsQEnG4x8gffKROY
gO9SHv14EsLyqwdN47fe0jpwUj8y1TK7vK4k2GVi0SZ+y0VI1dCsdgIxb4hkJLGi/o1Tr8hnd/0G
0IjlgetWvF6W0MCO/OQW16h983ytGUmr2TrjHcurKrR6Zl+Hv3VQEVvRgpTErttRsfBJ1hBOF1g1
jPcocCVklrQGXpVRNY8I9BJjUzS7/JRDk0EEsNUTPSqj1X1848UmPTlECLTc412vrFqqY7Tzwm4X
zHmRXrNFIx3LAtvWCw39S1cQmqC509WVaA/KQQ/7iEnHlw4PyMADG0bRGyg/KOPepX5Qby1W8Wd3
9d5Hxf+4ufiTRju+33SAiV0CHRPi8kPwufpXEYveT63+2eSz/XR0iPwA5CRR1E/X7Qy1u2jlJXX1
eaelkGFNFFFbjHs75AnxRjxRB49c/uB2Qk+jWzQpwumEabZw2P6bAvgSqXXB3NrtT7mGjeNF771t
zD7sWjdehIgMwWdLdoqUdcB4sclRV/cGnRRPaU2rpNu2QrlFuWSK7PR5wXtobhaEOtDyezDEkf89
TAzNCczXOM3nPsv97AEFQRx+w9PznL7kH5fM8GZ5B7wjsHonbAfopfCb/L73lvKRUjVfmB1Ji3Wc
o2J/xNiIaKPYhCG7kMcXPvxLQWhMC9sjiUqzog4ynx8ccFjc4WPMK2NZUIEgZTXB0zoIsMduoPAY
hFeMdGm7Sfw3es3cuyCs91gA4BIcPAUpcUe/1bXj1bOnsGS01FvyS8Bg7bVAQ9f8NszJDpBylS/D
WeDVGG201mRIBlJDAK47w1HU6ukPHUj4XFIYLJdfUUjG9fCO86LmaSGjVReKnlYunMSrt3o7CIzn
7JifJ0IPmr4z2+DlmMY0wtEkVOw1TzxSZS27nPE8fPQiqXuYR9xAGfz/VQJCQTPizFlCMyAUQKyI
HuTO9IFTXBTETjTrxlScmghS8hzA8av5Yxukf8jPChdgRH1f2qtzCgZVhhd0qiEup8Ov/fiPR1Ht
8qv8aTPsTVlhcenzNFdTiK1XYZeeyuZt1Fpm4qs+ZmEs5dKsLpIxquCD2tC6VZtndLhoo1LwVIMf
h9eqKN+nzO69/fMB9mPkT7n/AdqLg2G3ijLXK4FpyI1PhHgxVCz9DVeka2v9AEwH0FwPyRUQG0sG
/ubpCeq8YPqWlwCOLuaxKhKgAMo84p+UQiBtFgZGwOXE5Y43o0JVhL3g7yJN2P2bRvuodjDmSxYW
WW7ozprvT3F42PihTnDVcUqL4YPqvV8YrOYryJQzXzvX0bSOI4wQz4MQcdwojI0vdEFpC3G7pT5j
SKIHD9Wft3ZiHqJi88if5tU/3l1ie8m3T7EZ
`protect end_protected
