-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sH95hjKCUCnLeQhTM3ZaIfipfmKrIM/foNMlAr0bpdQ/BrpNe+3xdbudyCgsFsXz
zscItKiCwjtnKHBwGWE6q6mwBOY5rGDcZhf1BBeDfB1JTNLO8M2ezgyFk4NFD/bJ
bUcRyQEa6ESrgdud7AAjWiROKutrdSJXGsr7GmcQC5w=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 22640)
`protect data_block
g/ljVEZB0JMAB4XrtFvmRdD2dVZajcmnNeL7SFctkFPgkTLNcP8mw99VFIGTtain
kVFya/J3LXqvp7IeA4Q5Pi8nAqcYybn/mse/3W/3/W/y2wAa1TC4rkD9KpEBCilm
ndjIW9z7Mp5SgKpLlN0FOxleVMKOFXr371A1hpIwSMrd2sWNFVQFJIt9+ORcNGDc
tdxL++E+E4SCxKV1EX6zxsDd0k1demU49KpaxcKSGYB9ndXl4IdON+Ig5eAdiTdH
iN6uDJHmhPouds5WdFPIpWLVhSIJSEk99Tye6hfO/+1EGvpLPsuKuX8O+nrmMDW/
g1Xy+HbkntOQ0h+5pdfKWJDHIEXSc0/XmWscKAvR8Fm6DstskMKsqPl0Q3oVa3tB
oDfRyLGM4koCsRDehit1cu9xSOnzEEIA1HbtJOTKIT/s0f/adwWScDq0g+tKisUP
G5f41gKYT73ktLQpBwUN/pmv0BaPs5R5rA4e4KApuHQ8+EbysJFGYF0DEiWXbLhe
UaIEocasp4FivEqJXm2U5UiIdmXFuA+fna8Sz/Tspkwe/LVe52ea0W4JRHJCSxVU
TX1eP1+1hu+anYBSGnAbtaRYA3a2aYwPhmXxS0ndByJ9jBdDsVT/7OmSrIKWyIiJ
MMRQ7Hrq7ayj01q8UOPn0c7BsGeLbBxo7S4ZvAL7Mt+tVVyXoSQAOpiccrSEzlRq
ZslBpLDsI6vPykk2GLpzJd0N6dVt7chLw9kG54SnzX5rMNR4ldLWv7GFAomttpEs
HvVBAxpY3WAzHeSxgss7pBPRAHxC8qNJGW/kIThMHde70pSzRrlldthXAMZOycsY
4I8gjRRQfnDYvygpstUQluRt7YjF02yYNtISRTEZAKXOeDzwe8E2GHvU7qveiVFv
46gzU5PZtkU1H0My9B4ODV73WEiNW3imMiroOXp6sIE12yYNK4ukIQ3dHeIqsVu9
PLP/pWou4et8pUtQp3XWK0bu3lJEkXp0Hz0VsOl+BWvn8vri3Ma/70lA/H0rQLgf
fBEbBYSgSVQyjPeRe4fq+GXa8RuvpJkzy7NOXfbQL81bfTzsWMXATbVHm2ZT8zHa
layQBHpH3FIXVXQlnVbhkzsAgM3DCvN9bADcUwGetNMwrsb8JWmazJu01NZJ88uK
H5I3IxBCKakNZZdXy0boAPd5bTlRBabS7XN5V8+zo8ymfnDr9tTGJvgtQQD6Xfvf
VaP+lbFTGZAFjRGn6RccpniZZ3ewXTxjWio6ickzhCnH7Dr1VURa7DEKCAT7i/my
HYAKhtQ0ULv3F2v5o/lcMVhwr2M/6a4oGkUUU2TGG13f/QMoG3PVvghWb+hOCt5t
pkhjEij80PoJMJHcZQHwdvSYhOQOfPFeoGKKCRnH8BHkZYlCA1hs4r9imQRP46Z5
pTVz/82LKjf7RijTZQwBaUaETUEN/Y0sVKzBjmvcGC2ikK8HI32QEQDEuBi4xMt4
42BNLkahu7KQAR+aBqr9lzJ0KgTrsaSldtZRLak2zqUyjvZzI868o9JW6b58JuW7
EUgxeJMCnAmu771aW4iJRT7tD4iSkdxdbVv8aQ8AzKnw8oSts7D69g6YokHvPEvs
hsH6ejlR7tl7ERCEsOSW8yPv/+TA0lIy2uJaV+Nx9qjj/oorYEDLH9zjHMrWpLpb
+jIoO5IAYeGORl1699KkIlG4jqFzrEKSoex6OCql413s8p4R6oIJymqXLsUgbtpW
Avr+k9JfOf65WBP8J0J9hq0XVw98RXJ4+AFd1svKJQTneapXB9ln6JTU3jDm6C2q
4h20czQAscnSWbJM7FzFUvicyyy6Tx1CffGwBer7P3WZqYDyE11OmwSMO2hr3ajM
tgvnIBiQzbQcbJaTyoxXb5hpESjaiI4EDlZ/r1zfzeAoEiaQVJsjCjWL9PgGK9xS
7x7Y1xPIM0C30dH7hZlNQtns8BNwC2fhkFI21HclKXH7WGlZ3BnUAKVmheYEai0F
+LPgs8iT6yjkCLP8Jty65tYVJGPdcdMSuEwLvoTtK/NkY8gmGUwpFmA/dj8kTR0K
3vFsCBT73FbwjMl+uS8t24bsGf08bQuvb7I1ATv3Kgrpst1kmy1vjCajyJrO/6I0
qbsm7WhEnM9ERd6mA4PVxQM8FHbHvzFdQZygiHdgB8iA07F8HqccJf9LYh3XGij0
zfl0vCCDpVvA9JwrvfjzH2x0ABEKWVpny7O4LQRVuUvN0vJJh9j9vHD7z2vwi0hk
ftQ0zVaUk+j/r9zgSEc8X/v1SrvYxqLak/aJ21lofmtarHm+Zgf2WIc9PbH+nMkw
QV8Wo6J533zrtXsp0ak65E0bpNX/5Q/NdzRFio8BBkuOiYxe4Is9Nku2u/lIOP9j
bI3PBnlOFcAjDMUeZJRjpObNj6hoCDjCilLupJTZ6fkli0tj0uwNViYiQRazgopi
1bC6xBnKYGz4qhmILC9B+v5lhn+NPwnl54Z6WQededphnDSnCf+u5j4z+ubSHdiM
rJhf7NtgkqLM6o6HHMkHw3XyOLMRS/pOOVv2JMl8N7tUTHx9lEqjoBJMNHhjGWuO
pdnYDDN4JA1X4IIK7EJ4lv7QtKCk9Dy7C+v4Dpd/1rRUuvKkGP22eELFznSj1PWB
vLgdl+zSqrngGxE44kXl8J8l4KAzZHidMirZ0lz4ZKPjqQ+vZJtHblzdLH+YkJsZ
bTiRvsNbQwB78PjzvT6Tb6JukaqTAJbF1YjQ62oSe6fBbawK3HPBqK7M7jcoHQco
N07A7k/LXRzhT5jQRjtFc2OWnZklp30uxXDZzGfTo9cZeSX7udQeCL5Qk97mhucr
+qLX+iqAgX7W1IsaMSwil886bZ65OXSo4GugY0szt63V0bjqTGjQGUtAkCmMLisR
IcmV69KF3HmRi6cqgrSWmtk8gT8RZt5puxmrGlXxEtcbPTJSac0hzq3pwbxw7IfU
eLAG0Hk4bLm9wNpTaBtZjBcdRseF+qx2HN7IR+g+0QMyhTwHcwr4HTeJx4Yh9P1i
/72q5ArLxSE5u0mzEC0linasKJ+PQmwwd6BVeCboEtpAM8RnriBycXZUJSfboXQC
DhSxQOmnRyl74x9bluyDWpAnjcKl8k/rFprcSKvzX+3MKYbODjWZDwNg+RMPdbEV
1nK5njMdT1UGcvG9YbblJSRR2gqh0gADj15J/axYDhPS2NPddSYEaaeCcRKHSAit
z4iilNSyO/zYU3V358b1hrxp6m4Bfz4ldup3LC9emfePz3jWC1kvOlkBZ3jF2Zca
ZxFyi5jMVcVix+OEO8ACirioD1G0A7HoHYuz0YE0Dv5TEaZZP98n5MP7qkbEhVsg
NCiAC25Jjs49tHGkY9rIgVTUm6IQ0eGP+0GlFiMAeewWk9NNrsqoH+J8kZ+UUXpB
Fk9V1qRv1CTzlvaDrNmf6Hcur3oLbDKoV7bAQ1c1gJ1FMMPz7dOf9Zn6bsZZzV38
zKkxTzW/JwEtgYVURDi2xC4ot1VuYAIEMY8uMc+NQFT1r7FPeaFCpnUHULZi14uk
8f46n5b8QMjiypNkbEfyOuwUK+piaY0UfIjwMSvtuOk3X+/Jcv/2mRkMOB99jq8N
9StdMCm4Z0Odkg4EVLDsTVogA/03VC+duI91ggBOJ+liliHH0gZoOXQs5uAkAn4B
ENoRhUrnVUrYFwytgjW2GH80OepkOjECgbPS7Vlv/V9Y8aAdaIfmXin1Ja3MwdVR
2n+nHlJGgCh++mUWs8vBoqoju8FFgQ9qg/4x4pqu5YV9iJuQE7ljKFUZmKTsN5AK
8RWgJ+F/U+pa5OcEye1nqjF7IdMT8UXa3lyCFW7rnjSmsoAV34m06xFyBbohEUHT
/5/dAs8mHJHbIMdFmqkzQITgoJCa8gOutPew/OCOHJEq4dvyMkYio4f+frn/sYjQ
4NCPufRCyFTO171EA09vuguI44LR6NguBJKT97KpFFeR3R03YJTiV7qTjPcbunw/
HD2wvtjCpF521iRnCpx0nRg6BIKy1+hymdeBxeEnhMNrHS5A4XIzRLkyf0RfPEE+
JOEHnSmf77YWY/j+7SWPS13v8zn0ZwANSg7eZQkHHTC83UXx42w0CvHIN3f2zWFI
JbrmXinCprFwc+oB4ihPijj8M3H2OwnilOoFPwe8BNxz6iK8PlQVlNqLcsskriDI
eKWwyXtzGTg5zzScPBXopK4T1PexXsbWobbtroPhxSKKJY94QLuNEs+4QyqzBQzK
4sfGhaFtTnLLUONEtC2UNyZx9cBYv9+KGxmHF1HMrU3xDwUCGJFexQxm8QI8pFzN
XQTJb1+5aiF/aW93yTr49TdlwR/Ef1agUuO07FhuVv7uimJA5thMOysrVJAxf/It
bQdIitXWYqy0/mAVYhq+PdJHryRKXcAvxU0v/+Brf/7MTIznw3pvXCD+/Siqv1p9
cliymiBuYZB0QQGDpUmuS7ToPQnigAlV0vm+Zqpp6RZiYRn1O4Dtq/sAWo/yg+WM
IgK4UkP2IUL/OxgoWIgo6UezdywWUQTQ1gvuRMdHH4i5yb7aJYsqhVl3rt0nJROL
RfuLeay6Wj3d83OHG2Z9Mpw+G0d1F8v7Nmwjbh+oLLB6SyyMUkrV760mEEB3aMyi
21RDBPFCppgtMaE8rD5o+ILy27k7imBAu9I5y04hM63mjrNPzzgHjehqm0CFFjSi
cDKFHf5qkvYSX1UOOdhgzbf8l3L8rR2L+1ePHxJ7j6VkKluVpV8bIP8g+vaTK/7z
kf7HDSORehYEU9wHQUNf34qpIZup0RgcT4T5luHqDWa2CIAXSLKtlee7EuxZgCt0
1Ct1vu4ccZpythdlVFxiU7gx9JVx1LVrOenMghWyaySjj8ipmEtySOcm6I94Q65B
riCb6m3K+3EjsH/3ufT36PzDVybDIe2kjhT4LzD+2HTbuMO4V3Z0qn5nyNG0OwlF
WSDK8Ye27k6hm/3f1cLtTYLzfvlHtx2ZJIw/3AVyPznzrm7IiwhoAnwlRDLxK5yT
S+yjRy/z1NyFUO2Sq1dV/jJvC5vmGBP8dsWXJ/0DS+H0xIGjd8QHSDVXbRn+p/ba
Lykcsq6MfVIVy1EPy3nU8s9pRQNNvmvYht1ZHQJ9vEKkSWiw12wSbFicamGIrJ4D
VWB2ZfQ6OM6ybFtjKnTxtUCx7pFgNnoUfNygfxXcJw7IBfZAVYIrJwb0l4N6g7Kp
epwljI66McXh4yo99wZMAIgixx0qEGGTvokesaiBsy6JDKc0PlsR8i96ClSz8Ljk
6MO+/dBRuujNaXK3/f4ECHFXPl7H8wPtsVVV7ToQtS1WkH+dm9BDD5VlVn2kBzK0
dH7FvRaHi7W0nEOtVJKshtOCqM5P0I5fe93wcDZEITRj352yrSiEyzCDZ398jyWh
1FIwZeeUhpggZxc+q5FRDMa4cPLphPLz65cUmzDWuGe/IwbW1w96Zwn1YpQjwPCV
YYX6IxEWiUWStlYtNiVy9rViyVataUoWqi84RJQKvVxkJbaImhvfbMbS8BU5pNoB
YjCH7ESSAFMC6VITj9NfM3iYKfIRQW+iR9HiE6QdqrxqVfgP6IKsuAeEYf7NtdI3
VkTqT4Vgo9RyY98h5ZR+7yBzkllYduYYBBp6fPU9Rps+Qsw+oFi9fKSd1ZSXcY59
JDavGSZl7+3UtRL4ZnUAqO9miO2lLy4CrglimkHRB+lHCXFEOjCjqqQsYArPwoeL
LFetJ1kpowxqI6eDJCdYlMB++HboVBQVfwybkSJ0mGYanqmvkKn9M1sO53lRUOYG
+75FGj7FxYIC4J8t4y09CIhTTGFFL3C7zVe4U8Dtubfvw9PW5oD7gzKr136aO+Jq
twcjShGImeRRISUX6RHLIYSp2/kAVb6Wjspy9Ds2B+Kw5v+/u92n/WgYwwYDugP9
wTxj2Q/9eYHSbtzX7ZWFYOGuO/wuqaOYuFniCw91ZxUegobeV3sxcHWQ8pPzD00X
ZO9O5sbm0C8fq34ljqrGMuOTVsH8fbjjtOJvbYloMtIN5Z9oUF+HDR/DIccrDy/1
aDBx+TpafEOxD6qn2JC7UJuquNZ6rIgmUCjA2c4AtiVUsDoEGengIorLLA8HWpfn
YlHWqHny3uUQYh55anPmNQnuP7cH/4lS2PMRYQr0d7DycMAmPxrhnXErdF4aw3EF
iUu3shsQLxPFM7AVDJq5qDRbnQGGH+wwGHBBFxNtZTxiwLyudyNARKl5hidJ3442
lCjSUPECR7DcO51q+mOVlYqVPccGV2kjuou/Utxj8ZHzn6LWkILO36ACuQPMzqST
Jevl3gSMFwol52OOwx8/xjgxCm6eCNXOrDdRyZ5BNt+mq86sJITmXMDXPK8dEJhQ
fKewFD7p+CM8QniebR7biaGTd6D5oMy1myK2XrRaV9p9zufhI6qN9yJXYy+BZdlS
GtRGzFL8oXZQndRcqgCvbcbwtWjuA9r0RqUGJ68U7TBkIk06qDcFZOiKdS4gLjvR
5dn12Z0QUKEBMmECHPQAAv8cl2xO5AmkazYboLq/wo0ZNR+qPbdGZWJkmkWIp98K
xfx+JH4YlFMbYyTwds1QUTa4jtDCvtE91eu7LzNdjroWGmLs7so7lhIEFfk4tkbE
yc9fjXTmlDGkzl86I5SKr1q1D4M2BBER4N+oB5GhvJSF19qWnHtcZyYN9xv7isjX
Xsl4a68LNcFFfGEJ03wdgxt85Qfpzg1SLrUmiK2oH/UXA0Y05dtUde2LE5cbJdkg
5keqrh/1JJuklkTi2N0XXIguzcGX4kfo/SEbwB0213vYjpbuczuWYQq2OE8psBXh
mzeOoDEMGUw3LIsq4Ct9tSWhmiGdnMAUzovBWuk9N5AovBZDO/zHDRMVh378dPTJ
zKe5tDrf6Ftcwnr1yqydvMr9z4P4g8rKNqQyXB5x/M8jGKQ1/NIAlN+Od1+1UWfa
s9wAAbQYJzcaLOB2WTUKbPtmJn56iw22R94WnZPds8Ow6AHMLosSq5fIjR0/MKWe
vxruCpAN1tv2V/Eao/j56AMVS7ky4HWUlyb8K2nfk8kUhaAZzs4o5/dy1Q5TrLh3
O5+cSoOTOp7PRcq2y6cDRo8x/5ZIxlqg+paHHNiacAc5DucWeKSX/wOYY9Rn0l+V
IGY6QMIz8exUP6X1g8jMkbA8mcyI4U4lLYVUNMkan4Ihb+MNXklWy5+SkYUS+k6l
0iEv5PIRbk/Y3Td+A/Gwo5Aj3QyTHXPawrC+Sj9W5I8Izk8QOquHYhkTnk4CPnoX
ASUMCDGRAcmWEhS9lD4LS54gfqXrU3vOtFdKgGsln+FIsO3l5ukyg9SGA8o2c193
jGiApYwSbmjaalmEmeP2OJrcDmqCN4p6mRwzJ4glV+DgKQzzXdAmKdIVnGj15Zt+
P46kdBVCcO6IrFOsXn0JuoctxmLFPDcQzD446ER5gDQkNgm9TnEuDQboLNFtjG57
G2zbtGJdFaEPAna1R20Aq+CXAyVvri2+GlcQPxxf6IrqDsfkhLcox+UIGkWcSEfq
6XYDvoQdriG3iuFIvOsxa1exXHerIvHZogGgddpmxTIRGII1BU+fGok2d+fpLbGK
1XgzazmPQ+jSDNtHXxgtyUxCMGRe/JxU4e8rwg/CwnvLgQHOMcTcLRyEN28lY2YG
7m9D2NRY0cAuDhAmRYhzftoOjkkiJU4gKT3T5zZ15bKMxbX+3zH2nnvrnu2ioR0q
9XJ5iAzTj+wLL2FOd2znogKbCNPRJEv8BsAJ0VZc2JzZ1yMoz+dN8B1Fihwewqq1
pYFXSEfMg4+wDQigekUcwYZxMa6M4VuhtovZiZwKVvaLLP6sChFbRBDfiHR+vdW2
8/qApGfhLCbu2eEMjpsp5TAjPkwYVFICoyJRxouTo5fYow89R+GXORG5iIRW2AGa
ja6i8o0m14yLRMS4GVMtJ2bGb8Y1QbF3aYmB+0n416YU2YbfXR+eGbvdNPW6O2YF
6FxwUZBrA3W1vpCLG0ReAuY0XM6h5jJDCtKJb0bu2v9Odj7d6jo2kmLERYZumgYS
shbZqcWXaMzv8VUq5nFW1hns6Y+PIrdg3DKbJWfEakC6nJIUYIG3tAkSh6u7kU9E
tNcyLZVkBj6vnfrhPH9ZmYVpDAuAGwKPyZI3zXrqNSIBedrKgSFKujK/bA67RVRN
lMmW8RCGEVShYYMUvp7p0GuRUkdyVvhHXMvN4z7nCkS1crB141rYI0MWzuXWkPYj
CsppLbKZRU+MKrMdHeB3giEZRd5V/eOGe0fOonqmDWKn9P/2YTT1zE0A/qoI85Va
0CMnW1CPmQp6xsgQq28ou7zhcDA2M6UX+KVKdgUh71vQaZuooghdlC2vTysoiubs
ZE6aNbaKQAQZMuXxTlcXqgNd0TnbkF7mrFQVdMYVMpJsLE6d5mOP+L0JYvEpapxf
ccYVfVgrK85/pL4ylrTr5nmxUmFuf1KU9yqYoxSW/+zBSnu1yqqVzp6xJMDEcw2Y
0SUUv87hYbr6ZDELASBiBozgfek8HKDEl4HwpSd6DzDWWcA2GjJ4p0JIHdOylCJM
m73P+LLObuBdpswqXNmrKXO/VjXqy2zxUm718mFLcIfyKni6Nhp73/SC4wQwXMfk
ZOzg/0Nza57LaFmU33uLTdmeZYAt9OJuLQDlRb9Jxtu9nRiaVs1na1c4Lxjt8hXf
JYi9UGrF3eFd3oJuwHPNVm6eKj1Hj4LoWuxY2meY0APkJkk6cV0H5QuJ0t37OFBY
WR2qI+ZtQBzBC12rcWMY5WSMD2EU/hEsIzKUVaGRtvHGiwxdBAVVrxXjehBSADyI
JfCu4GAYvKjIbWm7fj2PiYkxZho9XblJCCOBDVKS5iporZ622C0Ys/ZY7/0ZlGtm
AZ/AAj+86cWIcHMLtYetyR+6zLX1d8JqGzAKiwPXqv5JBX6GtlXA73S0T7YvwRGw
jSqNk5NWW9xUcNpLkF3Gw5uaR2hBSJF7LRWpbHH9rkpuT4ughSCH60K1IyIJTK3H
Hd5YsgQDxxqPd5mRajhp0nl8gGPCPtnugcC8NLxvlDIKSV88sMrGEmybTJgKLlvN
571ihCwBdMwkOSDxzll2p5hzfv1GJyCQ9YsX/zZdk24/qqtOk9LvevMMYeyXiYgm
EbW8fiKMA3CSR6VGugVwjeK+3PxytxbBuyqP4ueJKMCpjVqe3H75su2zUCOaFKzD
o5JsmwLZtJTGu/8sdO1G4muwLQQzIXMQkWk3a3iQyHMeZFc/COd9hw9xI0OMYeIG
MDSIjPzYQC9gXqp4xzqVlJcNLzv7wDL8V1Wf0pv7p6tmQIXOcqocMKubqTT01tcN
22hd7oxHSx5r5CUlGfj6voRwVzy4LUEGP8ghXIrl1GeBJBOMGD8nbyaYEwjYaIZx
5iQrOincGg/pmtLftM3ci0olyQq49Y/k9IUV7dCE0Ts6uDezEcSHYPOUMX2y+7dO
KuDb+k0NQecSqd1eXdlwA0vA/8PhRpqNxT5OfGQjsNiLEkEnloKb5XSYM4h7aqcQ
bshGtErK8ow94sh9OxtYisplJ0HMmfkrmaNJZckH/wsH2d9jXLxvD7xE3iqaI21b
GZOk2H2Gz5fWWCvzWlHIATNqp4Cf5JRE5ppaxmRoNvlzFmFJwPenwwOJCK+xUt12
w6iJD2HdPyBeEM3yikjfNDbSLSDiMKeYzTCvBc0juHZWjUi4tmRT+cn65nwVF3Nm
lMMK0MQiD7eUxc9jDKYDRCu9Gd1vAPVAhlXYPgnhbG0NjtVF7Mg6Ui5Lk3kVShZo
03rOoLwyLrAoE1kDYsPU3pvqi/rWp9QmPqvjdG9ZnZj8GCOt8xQ+06AYJJeJEME9
wjkCPlATbU1LUyqU3gAgJK0ZxC5yLvvBxzsQtGdnBwnMM7k9JtyJR8KMTqOKOeMv
7s3mW3e/GscMuozv54WfWza6bM0HHIQKlHu0rvm6F+DnaX87CLRtZyXWATst6qHD
bObFA0b0sn/eSKG4qIjBbfG5pOy5kcpgrEe9m+E9CpWOydsvcz7M+uTmO/1GOCOK
hWfOCOeXe9a0an5L+6KH+K5V7Qg76J9i3ZMYeeS8RFBylYsMxqfI6L1jeKguedB4
ahyfIf3/oIcODfL+CCK6PCCXXFAB22mVJoj0HVruM71V8Zdrdlzf80QH53xqPdiR
EA2C0/l3eHILObOdegTM1kpBBkC5dVtN3LBxFpLTJXkbk1Dbb6lGK+AvZuSiWJpr
+mAI3IezhAEk1wTYgMHeVxd82y2Q3DixlRvX+WW+lp5GqU97pGtwSx5URV/SZpXx
OhKrY1Fl2If6A7JbAeW+fiM/FaxxE4+DCSxWv0jouQ8b9vJgtxidyYOeA9F1vND0
td5LCB2k2NHp2CZbQEFVJDS+h/YKFSDDNfgA6fLPgl7y3yQSmVKBk5t+h1guc3XF
DJOAsXCq/SypxoQ7QIBB4spJMkpOJCKKwk4aFJ3yxEMhIixyCk40q2x/s1LwRDH0
xUp4ha7y0dthoZAaCpFO+J+janEIK6pjcMJZpAd5aW5tctVktyX8QW2WSojCa47b
fdLpMTmXnawy4UGGOyNz9dQ/0cArfC5qRjtYYrgPscTNXs0JIKBv7Q7uHe4eGfZx
6vG+6+3rKCbMgXhwXXIlWoVcEMJONWXjtNA50LB8PnT3hX420GEaP8ExK36fhnoE
Gg0ktvexaCWQtzmwcgOobu2l2xL7avHtPbajbNQLwyj2fwcosZdwyZ2IwOB/2k/W
Uhhu+jVoaa/sT0J7n3oeShaPJifRcP320itNI/28VDeE64CANbwEmP0EOVEVPh8Q
pzZ/sbOmAt1zocfz1EnL85AVW8R9hlPgCE+mJa5RUzxSagLqiwm5OBEty4PyTZvC
T/CjFtMGaAL+at6oQi/f2HU9zDIsHh2BEaOdJXI4wslw8E6kis1C18068YQk7JhV
9DwXDitG4xma7R/I+XZIrzElhfOLp8vyeF3rsAUQGLkzafPztQgqHHh55O53MHp+
T4RPO+WD9Srm96CEJsIGpe6hzjLOUh7NVzvC0SU2yCH8nHGBH1odYZptNavdRGwr
yZCY+WW6gWokARg1QVfr539i0HOmmo03pUtvgva1Z2Wcf8MQ7YjEWjiKf5TOVm1y
pj5sH/2cPMO8N2sT9GUu4hiXZ1Q8LvH3SSMryZSzK/qbicgIu0QS5GQ31qzKcpI7
ZIG5hgo3bEv3SDjx/6e92wZxOr5KfAoxV33X2NYKdZ22KDr3d64iQF/QeyLDAAbE
vSiWf7528yd1MzW806xf0MaSA2y/HIOI134DUNW3/z2lRijuOEpd3rnhpXCnrDe5
JbbEZ3lJwfbJNC+h+u8vtyJNxc2Q5rSKMj83+9OsIef9I/+7r27Xs/DgRkVcqhz7
lH0o8EYocbHMF0c9wPSWn8WbcJAqYw6SKeIDpDBqkDweeQkYIAAduzS2qLRuWRKD
aA9jw1Y4yTS1aTF1fyW98bzw1ecAUIERd5/QL6Hu0RWpxjeBoUS4PahtU5EyCj07
oScPCgbUUUyyUx8c+5c7/vHEIUsQ02goAe8lnCbL56ZiDWQ93HbhNG8CXzHp7yXa
dLlVSwBH1I0K1ZMVOT4Pd4KX/FHbJ5T+CeFwvKfmgTlv2WXU7Vls8bxadO2G/8fg
L/pyMJgxcG3uWWGJWgOijKTNTzhjs0LJwbIDKAlOLo66FIJI01O+/2RGliwz/MXx
A7qMYmVm/hGkwqBzWsc7ZYO6C3O7T2vai/DVQxM44l+jJtC/5vkf+QGOI5uNXlRd
lo2T3iy4kiCDwumgC9ghEubb0nig2gDuc+JkXwTN1CO3mE4ISceJADT7yadsazSS
7QON+pBoEx+DgVfzJX9gX182lBN9+oPbdD6uq+FjJUSbdMVO92CMFTtGdHp4Kzpg
Ty6iquTT3R+7RBvw0nJbqxT3qD59CgCOBEoIwgesgcPe8A8dUucL2avJsuDjeoab
rdNVP5Ymycnf1CLaCz7mHgMq6ULzdIE2bLTOvbZ0e7pdNxuD5Q5TbMsy8UBPC/j1
sZcVKlUSKOaoFtalla/oLtrUBqes5GQH6HsOPO5JLnYqtb9Adz8jYuUzF1sBKecw
guxJSGQ+QdtRvEqBbXhpVCJWsVc05WqK1WczsJAgGSfOGbqHHRjVb6/HSy1vsu76
6NBhxghIwq5uwCdeuy3s0toxDOTO4B+3IGzXYfdr+eQnISYohPvJ/BL+viBlVfQ0
4HrWQBAY7/mZm2h1AqlLuyu0/ina9OJWzXk4wVSQX0E5lTDtvwM6ilD6aCm+9gKv
pBjj+vlFQFHIIFqwhYhUI3JgXHg0xgxyPpgS+1ig+Z3X2opDXuSHUyRZxWM//qeD
bsvPdlqo8eRYpRJwS0EmZvtdgSCGub60CcuFrGhI2QkngaNGCvW4uvSMljx+yKhj
L6y5A9WG2lE1bPzlx+eb2NzuTXL5XrDGphVUh0rBq5ggJRMfOi5Ejmqyq5tKvrwW
pGEXgIAX9GgHeaVxbTIKMv2Ifn7LzO1cOd5a5ilQivrO6jMDf3bnlOjkcTqH4+5H
L4wF8o3kDxzdvn1EG4OEz2pVXSuz0Xr96qimXpZ5uX1tw0XqevlVVY+f9bM44kv6
/IjslwoURIOaIYC8e8EOK7I+xDMZGzwlT+OUjvpzcTaIcM+h9Iw1fql3YCElxv3l
fwq4hSFUmZCX6Z0LEwymdKIqkZJpIzL4soY/dRYVbGagWTg1wSBbw8bgbSsqE51S
ihYFaXenG3o9xHDknElFd90GxSI6alntiXrTa0lVLwoNkHVj5FqQRDlox2sfOKrE
NFXcICG/pfc6cVsUyGqb0d0hL34Bbzs5TxxEvpxPYAx13JpNJ8PCs9c5HsyOV26s
pBluBUNWolwSdt3r+zoytUVPrVQwVolC6VXjOFGbcath3ojck8nayhVo8aa3BOHq
aLXBwi3xX1wiAU56EOZIPDmDg1/jhV5DHuYTWYe2bqIKcOKVL0p+Q8rnl/XZsO4k
Gvwp5sWrpc9O6wUcsktXzv9Nj4KO1aukxv1whQ9iSlxD/mfH9rUJ6rYW/4rZIEIZ
WDUGnzkrcabdRCaHnoagYDvY0DhlcGlFUC3et83FQQ3dHM4I8/Q/7DnwYB43yHIR
fj3yC/KnIkhHbRNUjuo3iHjGytfpp0l5zUJG8nE+EtRtNtitTe001Vqx3qYBNYlF
MZgllio2QIE4yZVS2/0GUDEUH5rIGHmL8x6Y14XG+vxMdLv7AqjysAoIh2qeJsDf
Ppw4L/3jM0kpG/OFDuFe4dTTT9Fod7mixi8Gcw2ZUMusA6ZG9TfTtuj+FmekSVjo
nqH/FmNxiFCHeVL6mfZdb0PfGGjBc5XcRfv5yDjlpdOLQ2wSkD3tBIqL/hLB8ZYB
6fEqznOxsifKiP8CVFX84Ay0i57OqNo+bhS3bWWVwXxZcyJemRsmc1dh0fbr8EFF
LcrJqB5vPj0iy5HicPFBmS/O4hmHgV4L6WqxZTVKnYcn8mSKd3drB5ikl48lGxLZ
ZoyCAXnL1fS/8xOSCtZ1FUo75Xl8ECBN3FcIsDGFPty2YKhyRRMf6d9IwOrQG7s1
U1i3L/nXltda4sITH00rw2ZOggWKIvv+mJTHcJ9qaoHIU1sKRr2XPQcPj1O04zR2
igFqcRpChF5SYpLfMPsaIQxyIiz+Dt47Z1QNEjy4b5FaNGY3E5bXXLh7woo2m/tD
5ctZ4qF3cAniXw8VCKAaOyv+E1yNn1cjaNtSPnGv6Q729td7aDSv/INCprNoLvhi
oV/zbNDrvhdf5IbpTy04SCK/6AnUxeWo75WNkmpZuxJnEeB0g1ysxImiD8pQJF0W
AajuNXWzWPsSgKOw3xIknRyuwsgEtl8xcJ8q3qQgD2VCRux6/uopG+Uz8Zu+bvE6
ARmmtB/uhD2hrzXD+83b4KdJBHtA83o5rXt9YbD+XHN6DhBec/7+wwVYESDphp/D
0+3ih3dZ+kvOFVwLQGkxfrkdAuv/GNvwVuUBK55RzURkvmvDJSEibvBiZdull6jm
F5jIJv6oaF61BWPw3NvKspzByvITFbjnMkW1qwO2wBS8W/KcWBIspqOIyg4rlVCQ
949b2ea+Ag5uqMf/lbxMJFIQiXhitu8z9/Y5/EW5e27K8B6GlSXzWWVKqcHBYgEW
0WCLBSOaIUDxiFr8sr+cgibIKPwVoVtRH//HejakwBIKFaODAed710O0/551N+CC
hlEYVT1WmZpKif5kGrZbOS7QZ45ln2yoKwWFveis01QFpeX868QRkizQCK8xM89C
NSKaHfOwQFXJyRhapq7GbiavyLPYdXzxCsYDAx+h2gpN7LCPXVb3lKUZtWfc+4gU
FIIKvdtxXd9WS+M/0LnwGpImEih4iU4B1o5tUNBlHn5UsoZ/a2TyOMPA1WcOqarK
OJe6sMuLLWGZtSM9c4UmdXve0TSJUG5g/kBY4HZifAGOjuZUxJr2uya4V+plj5I4
6faElvzWdtRuuXhM+JwtQ5AoRAyP0CRIR4KmGvYCYGx/vkY/6KwIwjzTnREq/mNf
SO6akPeACw4io7h+9FIpBeBLCS+ak72GiaGhk0VOXiyRrlpgJsQnYRXYBsj8VXCr
8nhl7lO3ssiX4N7UEGtHHD2zs/sNoasMOAw7umMDnL/v6WYOf/EdRPFlBsGH8zGA
7ExZwKILaVqvWoyJQTWqROzA7vbXkDMkg8lvpFTpK5iRLuogbC3/9kaswe2dJVkp
MyMtdvIeU8GDuXPEmkIwftufiESSeklPfwmRUvdM0Gm5yYcIeT4Vf201F1t29Baa
0xi98A70hRO4rz8KNWQjKMCe3oDPAZ2q30J3a/4UELd6RrDPPMmcLql+61ko32g7
vP8GkbRKy14PApYuk4TStnqPMqqfxnFt4iWfGsdVcZbsOvWtQXLYYHR/Slv5XcQS
xBHEWS9TeyB094PnnXC9GWNJKtpr8jxLhFfTcZpnonlwUXPACQ1tlUyNHMcl7QR+
EPuMGGPul3y2IB1F1hFDyA8sbZbMtXvIk8lHUctUDPWUEx9MVpvnbOeav4QAwp/b
f+DmgKnwalncj0mTcA/Kwz6FjWT/QzLzcl3tQPyztvk+cyhaPL110WysPvBWXOZg
vAaoeWqkkpbIaP5STVb74li/o9LEf8VX5xh/W1zjupOUH7FNRDVND7YxMyjGN5Ru
MNhS7D/gWfPQOS8ql5Wnhv/C3Ib8BigeSnMUQGUamGsW17ApjbMmcWNaf1Md60Me
aUcjHrre1Du1uVfkVz7AGZGXRWChGoFlzZ91kl3/J63neNRjayOZgMRAYutAHvqJ
TtbUUUPCGinHf8o0yevXkIq9thjC2cOy9N40GSE1OAbzACf4O1k79r95OL8Svd5+
CSaW1Lj5CYBonLkrnb5AN3+H69EwKVovTxD60EHme0ZTIa4eGoUuaoeAn7+pb8z3
Y2ZXm4Ji0chz+ekDulMwj1t8D66O+4uFEgc8YiAR+Kl1tuNnvImwiTlvUK/PG8NB
wtv1GaVVz7H922/uegYnih/YUfsv4bAKsKRX3+F4c3GYA4WFyBwbD/uzw6YVKJS5
jyZNMoaJaXhZ1tjcX3KJKVjRMw4GGFBfaisRmITmK8f5amIEPVmGBuk3nEOV40Bi
/hCoaOL6NEqvqjEa+ocMk0i5ExymVSj6k1XKIt/NvEF5JwOFVLiBsbFs93fHPtCx
zjOOab5Z/MKf35VapBBI06alq7bEdqBfnQGrXTno1cphw0/5vAnO+XPpgGLoP5I9
Rh/Lh70Qo526PGMCWqSpfvJTdwohuVOaYunUptjnJ2qvodxIkRJ0dkBLEgyEfalA
HWn2L/d2rUTS92g9KvyJU20rIGo4xIPEM4S0XWbKOEYv0dZCxmffqwnlHw742CGn
9MHZimMWwI5aMDVnDS6LaKVQxeTiaxr8OFQyqbX/c9T7Xs/ChQUK68CivNbLRtrc
HcFJBQmIUTtvYAHqmwTCXgbhAiW2vpkaETkEIeHsOiZBm8rHPqHaCxOB3Fd4Nlzk
GZVR1Ei6feqSueS7CvAuYYJavShECE/wakuggVlohtPt1nLCsAkjCvNSHQU93xE7
zSp9dm4STefId7/y+mV7NSIy2fl3dY3F3pB5jq4lJaQ2OHCmgs4kgthv293Dp+88
FiWKI8CJGqO2+Sls17a3EQMJrtq8CYqX/DbyxaT1wfJ8dADDBryQ0jnqExMAV9fJ
Uvey5qV+ovr1n1Bwm1G4Wvc9yR5G5yUHdFARxL7qcFJqSnyIuHSvTZeUoIvcUPC9
te2Fu5VjOAs3eWOiDFYyatRRsKMd5ctJZNx5Pep1flArIPvI++hOHXIh7tATS5o2
d4GKIC57uNbTGcv4IkrCOpGoeJyfqt/LtWwaI/p9C82l3D94kdvTt4IarFPBWfFU
WnGZgpZv8sVeq6uZM/pBEe4WFZxQzDksRpzB5tf7kxhz9UvPSYD/mCm13n6YD7Ys
IerIOTmV6P/8s4DQLNQgfBJ4hSoGk694B14eLMUAibn7fd+HlZIEBKNpd/G+vY0d
viNH4paggxlSB3WfWugptdZtw6XtJzN6GogTJ9uulC/j3Cwng3Y1BEyNnQ8soRHh
97uwiHunvSp9ZO+T1gdxvw5cbeIEW0N1uL800OGczfh3wWzXD7UG5vgUQTS/J/Lp
yuvZM1lfgnnKYSxh40PNqpxNeCerDB+ux1eQzMrU/vLRdqfE0shW42xom1/LoB91
CQpGzFLVK190HMmEKOx75EEqbIDlcJEL9gDYkaS3EWx4QZ7g2k1Mjx18iXw3Bdmi
GJkPzLQ2BIffYuDZ5d3foUrBFYSrp8qgbinzxmH8GbXy7yuDhVr4Tm1Mpw6Hqby4
dPMOH4ct2VDvPPE0Ty5pcemNabmZcH6iU1UM+sd2SmYDHyk/ScT7gPRcyJpdj3X5
KrtHIchjvEcv/bGvvGQEr8/7UFF6AE8EYEifQMp/Qoj59wUfdYT76TcL1aOx2Wpe
IxVDVy/+o9PbLeqsWK++HWxqR3oEHJwhalynHUZHlm836vXaAXm9R22UyXa3kOpq
HB8BGQ3Tne6pRy5HIxdmtdi5vyX7wFs7S3LW7GNTmejKItz++U5LjkiZ2vNUDVVv
1HWVwXSR23zik2BXsBsby9aCfiK45SCdLW5fpG5MtibsTDih87oBirPFLGU2lewi
tG4HnNlrcfzs7xNfZCkIj0cbXlDWdLFkApTr6XtAPERa9SMncMh7Mx+pE7ejeRx6
AQDcCvGk2FIxwMDWrzZFnPwdA10hyfuOO3f8sD8dqRtwYt37twULhs/QppRBtDjy
bMRlYcYZgnAHBn31j7rgQGdv6RMYg9IEmqUDNx7Qf5Owz3PjcnHUeDVaD/cIwH8x
aEPQbWbNd9YP+rAwOrdtKwHwglSPY6+bXYX5hSXbPS2ss8eeZM04FGbS9WgPEfI1
BmTQ5w+ka2qBaUZh0Ofc6fiNJHRzEnl2yWMEocmJeXJrSF7QXO+x1IJby/VwxvFy
mhMLvwTfiBUsOm9Ws3vtHVi2cbeMlK8NQMNBKVxBKbNAg/bhM140kV75iaq3Ip/S
xXVErEFg/a18EpbAa2YKSW9XrfpcZ59iKFVPokEIVY2JJrCiXfCCV2hPArvEpg8d
26fqbTYGuaDg9UygKlHIZmjO6zyLI709FrFmbzPnTjbTnBWFS3NrL0MAKb/y1N4A
nozO1Bfz0/f/lbF4hbBgMdbphYCcL5TRCWXymHZPa4z0WLXm2kHk4GdT6mSvDc2q
6oK6Typ5uvRFd5y4pDWrBsBsk+w5BQ1mf7fP39Fer59Cv0E5tT22/c8jk0CMPHeU
dEcVzHUhwjfYVBnprbZKrRw5pAOLixmvTTugoQmb6PYoMfvegAOVEcrWqAwJTfMZ
WEJ7OwJUlRYgQ7je8zRUrXOOO80zbGUQKyfZNVz29d6PoCKwT6Xn8hWHuIzxOdL+
MIU7aLHzfTq1VOK7PBg+1VT1iG7BQ3RhOdElVh1oanAuV2gZu3sRFWP7/61wMeD5
Uf5WexNOgCfGoWB/yzexZ6Pl/FqWipgkU8/alNT/QYv45OXJW5qFG0ZsW6hZmmKs
b0OuH1TGxSETfvIZrsKFTH/HijsB4qhYq2WAlIBENb2SlSfySyCGrUmO2J7Z9bjH
k/iM68WX42tnNbwwYttCoES4EsXc2rFzIzwHdlZHAQtrgkyHcv7OUfDBzXuvX8No
qgBmiztSmMSnDucXEw0Uut18WrXXbhT2Lw8VAGBo4m6V4dn2AP9oFJ5yusUF79Js
3G1jz2Lv7rbO1eD99wk/Bp+Oh5F3munC1A+ZRA9nIFYDDmoTh3cIybXd5fVcdKrA
S8pG6u9JPffU58nMQEgej14OisF+3tt1QLDSj1jWoT55cBEzHgfJgsVJa9DeFg5j
3vBVECRITCE54bDI6AhfnXgMNCC2c/t7FT4NL8MILODafFzYQXXbNKMXorQck8LM
u/5od1wPtWSab76KPffWBSH7LS3hVWlwbzBWYOZQnoZHfzmjzvrBQd2rlNfikht/
Zi1LYzRfGObS3+LNiR6RRPKFBA29MBLmm5pTcv+BgZpFbllHbOvs+3lxszb1AS7Z
bkOHcpV6j20OwjZO34NZCuKWUDgd2hz/S/odRmLHYuRABD3vKNXYBvK/wdP8YUWH
YLk+vVdy40yGJcVLXBj8+iMY1enF6ll5k+Wmpif70hFEr9z6lxrT14kgpdd2qfb8
HjRD/MLdWQnMznpKgVoAPTveH/jzEqOo1SMBRUi9IKb2K29FJxuBsr2oMCBXmAkl
/7awTNhkKhUgwTFXnScO2qT5XgYtEJ/p75VEUlpjMWS1jynB3GkP0kOBgLhvs9ju
S46577GpmNhAMaVmMWc3R2yklrNHT46Whu+cNqEG9DZAUuAcK4J4Bry0IFQflfpH
4Kes8zoFR8V1Gn3qO8IgWTMh1DKYA/M1jPq+HWnA33oXf+HMI3rhjDi6ZyZRUcmX
PTfZWS+qFLISKQoVNwBLqkwtT/NB/Myz3HT8Iyxn8AUTNjgIOkLWufMaKPXLynst
GEAncD2nHEwN6s5Ub8X87KVtFVkEbaonojF3/n4ftmZVTwdzY35fCSAvL6BIzJTk
wronjmIaNPsAyEPtj+EFCvUVkwdPrtUZOwh6iT5NPLPsyG8qtDTw2D5MfuCBOSJS
wotOTrpZZbFU0H9pAS1JNlvoAMvvgQuf0N9M/JPfTYzc1w90iEQNTcpxSgXufqXc
6hfgoxpMYjSQiqTY1jnK2H013boivQONaoBc2eZq513d2lcCNWEPtt5HPd7J7OH0
fviewY0Q14HSzzvpZv2KPP1My9ezkoSb8jWkUH3hn1oJkq5p88XjeKaf5w7l60Hq
8WJQDHGCalti7hq0oGkkCG1xE/8B7sullL5d1cIdKI2C95Wow0A/NO43BH4qJSiI
OLqz/4IqK7Q6MMSh1uQi9/rX2WAkkf6rd8SUOawLxNN5NcdJA/2QrCdXSB7vrvlj
LfyYfOc+aCwrQZfplAM3gy38d8oYS04QWAb7SDKuM9RPa1decbP5S0FPcncpg2Ns
5Iz4HXS4v7VTdaQ4I4NUHLoGQB+Prt6S6D4GjljtRyjHk85V4Bb+bGnPeo7J1eaZ
lw2GnmcysQbjHJGGZEp1ykNyLickPCRNvdEhTblI4fg9qaXy84lCBCCr+5npwoH4
p6YAv0aB3NbugXr4WKMrXH2r87YgqZr1NaCUUSz2JCte6kTnTkNmA2dfquTLh86s
kRxG1qjLJbAqD73E0NnMbnlLtVRbFV7NkpnlKZQKlMeHJIGYC6tfBxHXwmPTjm4+
mc6orVUxTI8dIzUtrL5l9W4cg+rYigspJeio+5VyIGLgVzqfqNlVR9cuNPyB8G7D
ZbM3Qlp6zokIkZWNvS+hdpiANAMX6Ot2Gv8cMfnAv3PTI8xXdNmQql/CqNXdDipA
Zb8K55+o6HeHrElXXUMT9Py4M4Wo8o9R/4DBx2YQU2Iv0W/i1FEyl/XV+V6NMbtd
UOiuqGf84WGqwoPH66/YlFFjS37SjQP1OdMs4FnuwxAlcZnv4DC0AHQID/0eQxAX
NxG7RMjECI2QMYE1Ba+v0Q3bIJexCmePbM2VBKkcU8FT3X8mameM/9sxHlTzolpR
lKVO23w5qlycM/Km6GU6hb+pzZBQrOoyAvT65rZfmctMfK+SLk11v6o2i+3GL5ft
24QP7GWG8mUzmRm42B7EKgSOZTym8+bIn05DmgX77t3jkbarhtFt7uMGYuTQfO1a
qx5EpNr0+U1OzftDFI7hiYT9BA66/6lwwzElLTYUb52+qfeYc4uDW81WHCGxZmln
wwJ0qGSVbZf6uD5bgx3zHqu+VuTgNzNlhwz+hC/NuvptKnkEkOjU2iOfKZq1L1NO
j61uT4GOMiyt9hwIskFxU24jfR3GgMOybY0b2F9cVoUBa7g++zE7XlWPw8AWsqcs
oSirARxse64OAFpHDUD06e66ARM6gE0ss2sDcsZia0M8VGqAfrbhYrFBW+G79uhB
JiKVAV54T1GJl9kLE09rWdVgpBYzo8Doa6228P4032HzuWC7hsktZaIrtj3S5R16
q+ZVAxdaPHwrCfBbElibEStVfkNquQylyvihD4o+ExYJQL6wuO6OjjztwxFfNIV/
b9B7XDrH1C2jAv0emtaDM/EUCF0Y5SkttZ7PJ8eLh3ZtqzaB/CtzMqOPjkCPCjUI
3YSu3p0pj2LeEFiXOOynjYVcHOC0UGgaOCbWgTEcqY+iBjV94zmm50GilQgqLVU5
RLaiMwFZTIARiF/FLq/T9SgN3L/pPLN19xYEy+3T/i5IxO2htw07QbWRS8ke3+UF
jBp28EPCWGhmXUUoKXJ2HUd87BvoFXQloRCKN/zSlrNJCSy4YrKTsIpc5RRTB+wh
qcoYdLlVIQLog9GhtDBLBWKiRXTVDL00cskNZKqW1l9beLjfvI74uWpBjXY5QfZd
cn5HvQX3X+vuwQnRxJVeBynCwdcMTC+Kr6LjuqGn9W8zBWoDqroFPQYTIpJey/vE
72WpkseFGB0bw6g2q70bf3xSyPzMMQoEgTBvYhxtLyAQlaX+mnGIIcXPqtsq6MAc
hbn/HHF7xQ6uKPFp22DB/HvEVHVelsufBVUNqX8cjIjDnqJ8WRaYU07aDU505WRy
DpmxWpC+1c6xdU2zuwnGTO9uB2xtPVx+SwZAEiqMb+V60Ezi/cxej6F88Qi4Dh5o
jG+uxnTbYxCQOxdKg7vN0LzbaXzOl2XKLdrkxkpQALv5rNR6w1r4OH7tQSPj8Hb9
SPA6jAMK9D0K2tEBUN8m/LjnG5azgOU+vlbcPzCnrkugmxryGki05C2DPcYS7Ucs
7gyUBazXMNdpAVN7qrXV2a3/L41pWMaACG9VDhnZzSe15VMpHKJyCRzwiu8l7yRA
4bDepjvK9nMk19CT1M/pBWNbX103dpKkB4RP9In7MElx4vFarXUE8yYyTexHKfeg
bejnVh14Yh4QIQEoonrg6NZOpPOajvanITz2m4DvTdkXgeO1nCIs8XIOzogWZgat
L34qtruXn/3Nn3XZcrLMUHFXyW8/hCHBgdBlAC+HixP3lv3kbweeDzW1KgwBTwFJ
AhqihYdag7GqUhMe0kN47A26F1IDN21SbgnW9Y/kTGzg595ZTmM9wgagLk9z/ZYY
RoVjcm7EXA285Q/V2zqz6loecHjXOu+rkpXr25d2nn8PirZi+rCHjPCZqgzB3GmB
GjZ++PyM4TTO+/cxvxIdu4Ae+tYyEvbwfIDPcwk8qZBoqcyDiLE1+HRxbcjptubb
IwChhcCYyaxwbitvMrGs/G7o44nD8TW/tkmUW9fJ2Tnio31Fl3SCaW2HFySo1GyT
cVTZfycuDcWbXX6QCunMKA1R1+BoRmwMBva+JG+dgu0zF3MAZztsx3noe3NdcMEy
v0vM6uNwPn+jTDXUpqJroNft0yh/Sb0hjnx9P8JUE0VAYa7XChNakBfycrLMWpi8
mWONhuTrXS2FJ3/OIbNGEmbFdIGrDYF/LvfzUZz8xpOmcpvnjCE/uDiRHCn8hZGL
E1ERsVQkv1T7uxZNTyV6wC40POLT9H7CB+9NLrvSrgOr6AsIg+n9pR4vPDPBp80p
JGnADOXBsihR5G6Kn+T4c2/YQX5SjpEQoIDrHljjH9pU0iEGa9JWaJH7TtwFYrv4
CIEX7l9QmR4o7IkiwvIjlj8RIyj+5doO2jF4ID6Fi/m3/NfXTDtcagZfWk0GvNGa
/FdRa1ojAUcQeJnwM/UInPJWjEqc2MPkCkwg7IXuUG+8G1cwkzyjxIj0Zq+A3AWJ
6BtHN5JtVfNJCMgUHGUl1b4ooPI70qGjMKJUVRDRe5CxnFce4a/iWLE+Myttez5l
PtQA44AaEUsgXadHiv1JMVnHjW+i/4UrZC/Z5vKftLqi2gDLbOmw93ip91SpOPyp
tEJG7NSWSIn4z1niRNIyrDBxaZtFvis/7T50fZvSYDRjl9mN5G5yvY+t3TM5AyUb
WDUxX0L4iuM00yjImWL2LOCowDr1md6GSIb9blvXAk+kopWRc90Yygz7KU/kqUgq
YpxircRvwcIQfhQbeWBIJrCf8Gqjs2rtN2GPW2OILEyR8st54z5egSaoF7YDkVyr
6fRbzYtDU+iz/VoZoBPtPb7jI4ChrLyveXMUSb2BsblLEsYzAxeqr9NNPqlZ9Ys6
xmLWIto9W319k5Q+/JAdEoXmK/oAy7dLpq/1yyaeMkHtIP8hdNaGocp6HpayhTuJ
vfrItyK7NBsuiYGRivruJfrTasYLOLKZxt/pcJpz0zth0tBu3WReBUCzt2iUx3Pb
ocTWL+mb7JHMZH9UjSBOQtpmPwCpUurkM3RBktnHgAqgDqcZs5qzC47TqYn/NDUN
7cz8IxsiYV8IvNZLiDSFdAKV8BR9rnr2KZzSg+tBLUoJSj+NSkSDGvFQ+7x05NHR
WA5trk9Ol83SuzoGqa1frdypD7sWvZLkk8Ny/3wLJtsXlKvu+gGsibAMuR3wKhNU
OtWNP1MicXUelxdiKg7jT0sLueB0N6/q8RdQBZfGzL8judgC8JBUiJBykS1e1ZRd
s3EBtgyt/BAEEqfGbTCx178Rz7ailqonhVZj1rYCmaF7nxD7M47+6qCB+16kacpu
smhUld0QHVVOhmxMnUMNx9DxwCoZvXnSNy0DyfKRvMuPAEANXx5JA18juUlnrdRM
nYsmdzGl4K80VQSehPzVKweA7Gs1RvrQOG/c+PSXZIDDTjDEQv6tqvmHgALEQfJL
52tZ767Ssbt8bAxsoyHhYre7YCuGOPhJhy7Z/AzX1TLKJVReeO5tnnEBBNxKC7C2
Ug/q+xLpROdU0jAPx+xP2CtFkOmvVgx8eo/KwV7DE8bQUTETXw0w7hy7UvouSpqO
12vFtFQqiq+nvRTiAMRx/AWBU4JTglZMXr9wS8QjyNPhl/evrJ7OMqTPy7I8DbhB
XYOQLYvJft7908wyux3Ub5gN1J37yCQMryUEpcbZpe13IeJMhO3JvpcwgElw5P8a
2H2jdia24hVZGunMYkkedlwPubfx3z/eSsPJfBfptCAFBbjOYRSx1skV8zAlnCK6
iMz/lj4SnAnQ/TUr9ct6YVy418Tza21Sv4IICc85FXkVVGO+RSgHNeX9keRqqrFs
fyFjBN6XSr+bsHgpvcvqdSreIRKlIl3SM3Ta/EwardxYAA7SUu0/tWFUwNJuAuaJ
zeNt0FWjkGz42+OdPIqS7+mpnsEEJs0m4V9aSl3GcX9RVXa+iMcD/+HYlweOnsLl
EAvtOU9Qi4dOfAGhUIobeglJQIlLjfseQ4sYEpCmBfxfmlOsZTx0UZx77FRLzt0w
3gawsYtBlDjTroHC0ucaRv3oIn7GSlnp+dZ15XpK/8ffuZCJYhehKhIfKwq1MXm1
YXdhZXLTLCvdGE5JyQCKeC0oCVppR+pKr1MiBOFzipiGwMjsNeT3ScPZoiANWNGE
OxyxrQttb1rZYbaLXPOkdppG3E2QLaYxelPaQlwljLj/QH8skJ1GUgU6yoX+Gp1S
jWRIySOQzCx8h+UIN9IdYWwKJzPKaMm5BJknn1f5D/O1DpMr0BDLg4No1+u9S92e
WLLQEnK1zRzKxydDh6vnsAijBE76IB0V9icQBKCTBNLJB1WfyjFXONApmel5TNwj
ZBkcpyunHggqoszNnZCx8erl20/1lovsUgEVsulW0COkK2Y9mPT5N0AWIFMBiZb3
olZLpB5utGxv1lymWyq7EVnNr0OQ+VNhvnBroWqUUN8aqsfifk3kCXfVp48nlQsw
vSGkU02UnDvIti+hMTqQ7v/FEu048rGczFD6lbjkZVrcUnBtVfDvlGHN+ybPhV93
WbftQqjTrGb39erUUe/QFQMFpYnpCimf0TkcZ75vjBjRzsuYR64t1/wmEvQS0F7N
syJRpV/E4vUuD+uWR/Z6FRT0dsmgQWBl+85AiXVE+k0fyP/WE+OdVTq0NoUsLTuI
w0iJKNC74z8gsB4MQYGV7a5joXDrnhXXiRFWYsqasjAhFa/V4XNZobKZqy6lLJnV
p8RTuL2HH1KMMvEGvOQCrQRpqcSM/0DLH3DLu5uO/AWi0R6iLfKdyl1aNqTRCfDu
jwBN93KW+BXgGm4tcEy/STKtLXwignpy3RWsrWOprUvVKT/NPNnCSK9jr9XDDxSN
hAo8qfAk2oM/63feDomYKjv7ffopAkNAEngkMkrV8p0bCBZO4pt/k0eLNjIhtet+
0d8PmzxZWwF0UXokK2J95Qv+96puXcXg9EpNwNGz6dExtZiJmcgsYYlwL8VHIMjM
5xLEY6oIKCsFZUHv9ibAtwsgM7fNr81QBfm+pBvb2n82k8ooX0iVjDu7JyaS2Dsz
w8kmYGQuYdwiKXnqFIy3mu8kqfZ5ZWyy+Zu/lKhwznDCUdZq/ABfsQUCZ8c158Z0
CJo2FKsbe3w73hQsJ89QEQxLb9zXu7KIxyRh0RnwVFKPwYp91g0DH5GiZ3n+IazV
PK3yB55VWsdo8Rbv/pNsMfPEoWvkNAYbkSSf2O3OifxJd0GlTBNKeaaigZXFJe+Y
pnEGUlgYr2we4OdNZ1XWiQ8Q4IYA6wKeXvmJY1X5C1WsZ4alXpkk6DW6Ucftjuye
dWVgXMMD9lEDyheHy4Pb3svCA5EXgGjjmhIzGt32upfRJI7lYavpWVTBU0MxTukh
9HXdx4QzNTDX1sGE+zYzHBnbxdjBiLjTWY4m8jXaTOrtgglQazdRQeYx/1/JqrEK
fGbraWmrPVSDmC2RhAGam9ayliWtzkyFyTjk7Ix+TYeiGAbqLgBn2ELhQR1eJC5S
Yud0J5edf7jKE28+F2RTHgHg/pWFVDoourc7o7ajRSx8ejLhw+DKSk0j6VBx+skS
KVc3cOpb9CLBrL99PfQOar3B+KfquBem2iBhdl4vov3+f+LAzGX2oF4aq1gWsYeM
M8AcHQmQwwJqmNG5znqVQgP5QnU+Kux2g3XApbwWO8y2FyRpb5eKs9MyUZ7HMOok
vzIbUFlw5SVmPjWJt3hGSBA5t3ydi1goXrWwzKM35Zy+11e7LtUo9MeB13WzgRPY
ZcBvfoRvxk4Y94VKFw8Drtpnc6USeAyOsPBGy/hiWlXnHGEKW1vHQYPR7QOJxnEg
BXX1kabLKcmP2enGhlYmigp+hUTYkOut44iQ374G4a8a6sOFaVnY/7AgXdlFmP0p
a3OSfP7K4Ef27KFb5IQ2k92NVyrM1hZrMFfvYFGMF0jJSvi1BAIoKEDo8s7xwgEu
FSEhZNHnicsUL+5nfJX9g9YcWAELGcNznSbaOeumhZR190nCwO/8hfkCXZJcrSnu
KsBsrDGeRYiGUiYFWJ0+Kx4sGxWukyKgpaPLQectWkVz/VODdUZQRU/8/r5miWqi
E8eFxgTdq844ZOFdDl7Nf2cpSb17wzm5CyzWsWgEqF1Izg7xBfQZ/NsFxT1hmZ+i
mBH3ABC2SmXPJwJ45HynF3DnVB1rrZ90ICw8/2ddflwBIbhH5EGSI4viSkbjerto
3dpWUz5gHV5A8LhVneIJLS6xpfJLL/hlKlECUxxRn8GyBnwdsT1ld8ifWMCephjE
LBI2kHbUcUKNUdDpaqBlRPmXRZbbJZeR2awVcgnvt/8uF+2Ri4Re5SdNJ8X5hc5I
zo1qqtkudMZuAPmVGs4N5gRXkUB/ybdZzIJGh0/Mh9HEkh8Ngroax9rgebFGZGKa
mWD8b1F8Kgx0DFxYVkZ8J/H2vW8x11TZGpmTU3gQvXk3Ff6QrVTKdoMbis1rZ0LV
dPT4utPSJifAVz+ekSGByDrvUXFXgmhx+s/HxIDEYei+BaFz8Qq0tUOS73aKSJ6S
LmjHH4uGDy87XBR0ONWE8b7vMgcHZoXYIF2p38WUmxjSsKsQ42uiukxB0NLgtzJJ
9p8KA3cOs1MV0K4DU8vhrTwnjVqAF6l2F/6K/mQ+D5cIu5lXI6yZd5OGLGWxKyzL
hlGX6uH2UzyjK0LOSz267L6yoe243PShxPx78TCBVw7081sq5chVum9Fj8QmRYy3
XS+oYzcmB7T/79UYS6Qq3qckVN7WIVxDFIqEoT4Mkdty7p7hxGZWD5itZ/07OFPw
83bvxB4NZ91rfVyzZBqqE81RhgYEd+0mOZF8yp3/4dzMbzpWSl/0oYlyAZRtZR5F
GCH5dSF0kW5JvoKA2r/0qptw0B2YCflvp2Ci3gG6weyz6a/vyODjSqvvLpKq03xm
NSTrX2R8A605qIpc/igdZQdEOfItywLA01Ye6lzAANm7Sxw+M7WJwZGgWLHaKeDu
GbtywjlPSQzjxv72HbPFwL8aJ6XyL8pI5GABFMiU1oc1T8ShCDW+gEwDRU1LzaGk
oQ3DbdhFUdNn1RXTCkgubt782dMLmIqcqKByn36kR5Q+rNxLuEsDQow/CRQaXetL
95IeAXuRv5uA2ObgUKQ/C8XkX2zXqamd0n/2SJU2R/aJQavVGfDFqFNC7UCACpBk
LItL1YleGzAzB4Ysfx2OBgPYwEeio5rpV9oNB2GTxJPkbEzgaViQex7ToVbQc11/
4Qz2xlawAbvzM7h37lMi4yEt5OxsmULFrBEJuNI4X2Vn+h/K6x33yMY/DKMGlz7q
mBPg/i2MOomFJu7lviBDKkR+tdqfhMsnglELCaqhVcjhTqretlPPibLO3p9h90Jx
TdhtUZMRnlBiqB+O7AwIkWtww5eteQuOYAvOBHL0KIecOg1AePMzIcHq8AJWzVAh
g8jd6mgkQvU2BTPJmoaYq9JKwIKQczTPOYnx3XQYNf0rXdcCCCarXDtdeWmdpgm6
8vazSJzVfxr19ob+0N8a/0RIoZBQQY8aerWBWVMxLoL/AhB56s58MknpH6exKL/8
j7u6PlmGqF5VVBfy57TMNaJXCVW7yQmhBI1XsrpB1sTe+5az3NkPM8pHvdmpll8R
ZH8Rs1Ukg8OnfT723Js+t0qOgKCSX2S1PP1HVXTENRNv3oLOfnIcxbnbbfHNKi3r
xYmGSewxilSorEejdzZJEVKTbML0ee6XnzrFmSUepg6B8nBEIzle3Xui1lpgORJT
XE77Ieql17UMfa+ytgYvwhvjd2kWD4zyLBzHKleiJJE6/C0cO5KHNqd9vdG3oYZf
WXPYROk8xcEDV3z3/yoZHMgfbYVGy26Db20LW56TMUhCBduO9zYx3qggnE0JVVyo
Jy87xBTHeC8vSX2+hvEbPmz0wFMehiKH2J1T6di/CZa5aL+YvxYROITElLJDdl27
ZMJ2fdBLxVTrvZTKEgEZfRYGQ9dqJsTR9QuVf3GL1iUVhW3U8+leMLVxBrEL+xSd
vu7lx7cMNSNFmF7fVxqdF9fTTvj4vRnq8ip3I/y2Y9l494AVuetehdPIcDldcJny
T3rS4+ZmOqHpudPPymP46ZBIp+jWP3DZvf/iNwUdU7/Tb4injsskfyu/p/HTbTFb
tffvNKPJNrg3JNPInLpdmRMPbNjj9PSWAoBtV13jqfPu8H85YkgMVQAyqru+S4OF
PTi7bbHFZZEG5kQELc5Y1mdxKKIk12wyQ2w17d2io3T1ox/4cxNcv610PuJeLzXt
3hkcpbniY5IpsDhCq3Vey99j1hoVNWKt1lMXsKmpiEBCjwq4Yocz5YsX9pr0fOnu
AV3N6IJW08hpAjDDGwb3e9MEdt0jWw3G0FP4a7BJvH0oPdOF8/DEadH64eKZosD0
zmR9wHoIh8jLHPlnycl9H7esaHXNop3gfGekBG7zrbbe6MJhNT7kOxTrdgcLCBAi
dPI4I87OQ41wE/uvq/NRSgl1/hTtcNeQIc2qN+X+hOupxriKyaHWduUJUDpScI/4
b/y8LRVbztynJjOkdtkZ7ZkQy/NaSHuK7dhri+VpaYBTAiLFPXhRzPs6PSnA+3/Q
34kL1LNsvvnSJ7pZb82uHXAgBZvH5WW9L2jP7hTWzpBxrI9K8YJ/OHx9LcvTHRYt
SioNdCc0ODPzdof3wc5LdLBqVrbgtRM3PFh27ibaXTOCSTmwxNBjDhSP6TwgMrjG
HpDAQZqS4hPoN+BKrgnFldLvDxEjdeIpNS3bx84tIOokaQbLzUhEsHXb27e+nz+I
1+yMQ6ng7mj85+UJKlYw8p2efisSXOGDmaKay9RdYpjxSdcwnYcqrAJKFbKbZmn0
TKWkJrss+gEAxLwEWqmg2yLBxEjh7mky+51Yd0BsPOBs/aR2EKSZGx9zbCN9FXzs
cp5kAvayLD8pXl8sZHKkpPghTZ0XHMHmidg/ZZpJrTFUcWnoi26dCT8bce5keyF+
Kdco+HKbl4sclVWG/yy0ZZpGyhubs+M9ktoqQIFnUP4AfLC58cLKfppF1KKHH2wF
fCZJMnZBOO/pU38azdzgZ9aUrMSbP+O3XHaYUQNtVLP4S17TJIlDPCGIwQdjrrD2
arwi9a0jC7FdZ36nbGYplka/SLGglCuLM/XJlDcv1G487zoXTZgttv36yRMr1L/T
lVWpT/fvi86K2tHuSPaIMLK3DhXOKvxQUwpTk0HGlHgkAxubM80ucoFCiXLyWuLR
KRXK8iEKNu2REgQWAG8+M4aakvhPqVZzb+Ww3BrwLEhrDUSDgJObLpC0yKfRCqV2
rQ4UR5JN8SN3eX3ji1ImP3TtdsfnYQGasGa+jFfVzhNNKnWZ/I8tcTm4pEs91DY0
MUSy3MCETwIPrGwg3d9sw2sD+Au7HVOm9TKPtftIDUKrwwQFEqjuhStAXvKA/6NM
nqDgf2IwPotdtYsa/7OTaG/EGfW3VKxPjlwSHI4rQ6QG+Fc2oOx7oTUY9sbOC/VZ
cYSWPOAtGcb9zVTOFP/LL26QntxNpepzb+/ASXrQzg+aMfonlqtj/gny/cBt02pa
qbhWlUDRPckAe28NUqdSLScy6ilrDdoIR4hZ1RuO3Ruy1vl+5xUxqbROWEoXWbwx
ltz1Tvqp0sbOmvOM9dJgXaNZYuufxWAA7YzTPeGRn3H7Hf4nsEfLj4P5zN4drzRc
WpEnPtzIYw3l1eaqCB/j2hNpImY2Lub20jdXtEAQGW648grj9nVJk5AbHwuRwcAs
H3g91w6+YOdWwXBH7qmLHfvxdJNG63DcbbNFt36BxoVyEocRQ9Bpyvg1+UFi2ig3
ZchTxN5Jj9r/jLWzdlevie/7iCP9QlEkd0rh7Ffye3p2bJenORD832h4b6TdQuuI
e853iRVsLMeDOLNa9iVdGCZyITsznL+GErL52gZMAcRia2qRyi21rma+zA0EizqB
XWWF5oS5JafRlHNfymbZ0UViZKN9SrteVyj0RNn2848c+TtPF7Tvz3PJCBje4ddM
WnUNEeCLKcM1lnQPVBOb1+EDUQmaazldcjnCAoeRaRAeoH+JhRSHkXd0AKQIIk8q
TYPQCm8LuglXugfIG5FeWL0fodfaWY7oMSSun/007Hji7kXk9GC4+Y0LEskF7Eua
AOossXWPqarnh43lwn4Ldr0ottiNZVKJCi13hAbPpFr+w4H6e4SHfo+G2uCg91oR
6S9z1WP6GzNDp+ycY0ZlEb5q83sDnOE5oNKWnTIlPOTA1GeTco/ivDpzOZ9iaMUN
O25MRw8pbqWwx3Wa8cy6k9o335xDcdIepfitAxDT3KA7UNUonB6HR81j5ZyeLSp7
DPpuFsPtiDzqhHxbz9EWDdCr1+Y2Y3u/IL9m1y/2q9exTPlhxANVBH6XI8REK1pM
l/6bv+qOGlryu5xNfkzG/kB1tIB2HY/z3IoINtw17EY6H54QoYHaYnI+9YbPmlvp
HpT501baTc20oCHg4nH6Qkqa4PJmaX70v1avN1rsUEk=
`protect end_protected
