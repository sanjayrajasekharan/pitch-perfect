-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
g5lCyH1oNrwqlc0Si6VH/jDjO89yImVJbS16B/JmB/KhiyJFvnv7+p1ctPuQsTnr
x1w1Vcqwav5+SFzckkWffTdjHB+CeXcIZodJWd0+lfKKm0zWgsaKZFQCq4fIMgvy
bPgrbvbKVh9Ba6zO9v3s9LYR5euCwuP29hrXE4JVezQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1012)

`protect DATA_BLOCK
Uqor+TgalqRrvsrEdADiHQ4l37H9dYmt1a4+iV2zkb6KrPJEI+gQJO7o0BD7Alnx
h/e652smWMHTCPUf+4bQkMOfQal/nD2TErQXc0NZyJvq0DOi/KxUpnBBX4jt9zal
bBU8tZBPffu+xcBYKmutIAWiJ8dlg9yh4T2ftXMjEu61OyxsB/yQvKqgeROXPbMc
oxyYUWN9dVSf0xNCAxw3Pxo4pY8vc/y+Juv7gaYf0ylGvlfmR99DPfvZazdcpnzi
p0LnC9lyd8bjOngY0oRUqc8Rpz9LmvmfM3LTS/8hDTXb+dzeds9MaMvBNP3VXdgU
QcnV/QeiX/kXXUd8j4Bh+o0wjHKMQ+M5YlxnKnpKwylgs4GCH6MUDKwJjgO0M7Yf
8ok0NPB28xrqdcDdr7yNC9iPd7qklwcBD+VA9bqaARdPJXsS+Dx25EnqGSylXuus
MY+daZzlZ+GU/uBAS4eFs3BwbBaQGJdNebkolJo0sCEU9NrMXoZuB3LEv6k362Cq
5KYOexAuplj9NxWpmSZS0B7UMzS2H4SQpBn4S3/R6YcWC8GsJAnyVBgrge+xiJX5
dtgVo9MXY3MRiccdqLqQuAErXEZLxB3EGFRN3gM239mfsTHbUK2nLsMac2c9IpCL
a/QoQdKxkl5L9g8Boq2lOOT5ALDk8GAgUj+dEPbaJamiiuE1obzqTVIleo4zQge6
TzPsuJOx/d+NqdSlAcixr2KXf8i+IR7YEyEbag6IEpmAW5/fTwq4JZbUV4z6hDxH
YyDyo6t8J4FSC+SO7SZ207CDmsLFnNFDoB4UEh35yHzssRIqvm1tdNWkPd6qV7sL
0IFOLIMnDqjeUm4Fke2/mKUXFP788FgL3fBtIOBhAFd5cKVY+G2R8HSUJk22Tpl3
tdlNikCTlRJ8wASUMmgtgMWyGmYz23NTeITnzTw9JpqGQtzTkpndNPdEf6s+6rGm
7WH19oQ2ksf+TmDpWMg9Rpt2dCrFYQzc5i166WdHP24WknWTPjfSutzXkQUCsuZw
WLHaTuVhpxD75YrNOhkVlWyBC9vH4Gh5FHK+SnCD8fAYmY9yZMnJNHx6Z/oCK7Vy
QWwZxdc58HoB3ubtz9jl8sy4+RB3YVgVh9vv97X3UHrGfs6z1ACHDDW52JnL5Usk
6JwbH//Wliu0PbvQcZhchDcFttYVL8sskIrlbQvDB/hWQGFY6nmb4QAGjaMGDP3Q
XGewoSG6O9WhdDr5rsbTvLh+ONh0Y8iSvkBKpmlqmQHvxI0akCauQ28T0u+0jwki
+DgQ/3mJfvpeGQTQTCWtL6ZcdAdxcT3TdDmx8ZoPj/OsD/VW6EHuLxjViAoCye6L
xkgQZNVXlldLu07MbhIxj+0lHJswIQiqCu58ykkjNp4=
`protect END_PROTECTED