-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vDSOxzPDRDcTvt17izv8rT9Xh196MnfK2px3bOyWaX2ZxySgyMJDtkGRP9rvWf2l
buPkOxqQEBC1u7bxJVkfjMgnpjlTDdSoNnqcl+ahwlbjpNS4inIfiIm7bd5tDO7g
bSrb8nXJPb4Ds2mAGy53siS/tVaLjYTKtm41LnZMWSxWWpw1kykHJw==
--pragma protect end_key_block
--pragma protect digest_block
E/DLBVsp4pdOUvNMC+uYrYwmYoE=
--pragma protect end_digest_block
--pragma protect data_block
m8nVlM/WSDbhgt+JgaJpP82Ov1l2lmrlHUELts8eR9lzlQex11h2LSqWZjjNwHwk
DnqxrrgvUemjYWcwUqqIF/UZmlQwCihIZXFQGLkTSGkGKPyx4yTKROjxITZCXrtR
dufzWwKyIjXxyCEraOa7ogd4PD85bOTDWfWLYWFcdbLjqAF9DyjVxtBJ8+BJQ6Wx
cMiRsSecQYNRgCdjkgY37HfE1Rit3+l7sDsEI2/3cQ0lSdpElUhmuc5znsOFDH3j
dcZfz0X1K6G+Zf0SOyw0RsRL67uB55vyZlsApplQN4L1e/Zpu8J+DgY4MSjDC8s1
mGiZ2fek8BxSvl1REmTWYuUwxWBMseM7OGnlR/D+Gsib+7MtDgGQOkxsa59QnDjU
mDFIibqam5svC5JT5B6dkJ/lXo4T+Dr96Ge7Y0Zakz0MBs6abpTH5yZhCDO6CcH2
8p7sEKrajFxXvQCqGGEvk0OvBzYXJ13vb5CcUegovgcWAMD7NPCb0VsmF8wwXNoN
/b0INBGvsyvR3ZtD/VXRRNKwqnX5OWYZUTKt/YRdb7syXETbcZcl0JGnxFTm3aUA
shxRCBpcWworS04YQu08wCIoE1MKyV2qcaDPGaETxuUv+/7OUxrWGfWwCbHvvoSj
1ujjZp7WICWTiwkSFtmaKLmg3F0xUaPhf6AuVxmSnUd2Wf9gFbaQMiZDpAN7JLzH
/qLLfQyT9gWXkOFnF2dlLJXHfWuQn1hAS4FFxVdVj17+CG43JV+7Ul0sldQ8ll2H
AsqvHCQTf7iV1OTiLCvrDYrKet+Ddhe0KGUuI8HcLBWwnp6VU3LhiOWPmsQETELa
6rIA8i1WKGIcLoAvJbV4U0OaGCrszhCBXNw3FW41sIKrbk0YNVFIJD1I3yMsojdf
b6t87yE5TSUvaUJw402VAJhYcigj8Dv7QrGOLfzslorVc6RbJ7VIz/McdeYE2PwA
xfkwV3iaZryn4FvCA85WELChC6Z8EaT+52mCccFy33w8PBDsMXr5ehxPntioxVJD
u27OVhwKvn9eUK+gLAztQTordG2d3caRUxsL3yYLrNPO/AGmKfa3vWUBU9sLeJMP
6gAJ2AsCpl5dF2Hx/mCbgKjJgjKqhxaXcX6QW/tPU835PwAV2czBR4HCLEWOX1ue
AF8dL/Fz19enxjmkDbbTX2LHTdkwHo3oFTcva0A1/DDBBsOuK0LezwnOgpza+tuL
w310grg1uLkJywYtGn5CDcXXmmLtcaZ6ukK/t49XvF7vaYv0KyfjlRx+40nQ/Mr9
T1MMrNyh9AnFVqR9iQMYd2XHQu6LZTicjCIvCy19UApgZd1KHZk8ju/SZK1o+Q4a
Pyyp2yf4YRUQ5pYFK6XSiFkXJbGkAqg6iXnwYHDLVtBmDTXB+8SmD2GYEYtg6+9x
1G8uSBsbKWfTJRp7nxZKMiLBbnVfdtqgvoYScnZ5aRCd5L1zcCz+LNO1Bsbq1eA/
qgF/vK/08K8YFNBvBXKoyCflNDyUxKDUYecUWdsVrfR6LbXNeY/FjYleHs06XA3b
jVXSlgKq7rrALOLpzqvFxlEa0E3DhUdrD8RzEJVOjtp7w1vSyA4GNOcjkmbSH0Aw
owzwnapLTnEX1ZRfE+2oyqhhp45wqP5scgKA0tQNhagmy7ipbnG5Gdc2ZctnovuR
JO9voFaZCNxW7cV78Syd4MYRLqwc+l51ZNBVg6qwZP6c83STXSzXi1hDyacSj60D
ThEoANUGSxdT4lJX2SzBSwz821Ymqt6UEOaQSZyN5gf1oxKyjcmSiaIynxWtA/1P
K5eYeO1Kfey8N/NhduJWCbxW9GA4cSkBipKHjhvYE7X0uBE4lMQigS52SBzRxCPH
lEQFafULjaUugaYxC95ZuuOXuEYrYPwZebLmm5PKg0LHwx17E4gWY26sqgsDwYOV
IiEcgrPDbf28+wlw+ZPNvrPmsMSg1jdgfO1fG6SDKsu4b8YoWfl04JmjSAwYsaj4
ICHfNw9YfYY6B0TQrvX4vO9WjYGMqsrFzqI7haTvaIFjcIxj1CS7Mno154gL+EXF
mBI27P5w5bc+hC1lQdqZecdiBjmXA5a6ZI/zKH8Jehyo4IaHZAgZtUkMdfquzCfs
r+Oo32UpGh6esOd0ligsh2d9puvnZJf/GdAPF5VY6Ufam4iB4xVgFYKep7S0vekN
QMICmUDXhmYviHr92RyqiVGXHsALLZrC9k2AEbFrddJNetVlNMjNNXJSkWnY0FD/
isFgq/WSyeuEmyiYhJ2uYiqAT66zCopOQZSCUHmTXhYepKcaAKNPOiO20qG20J36
5BN6AWRJI+aF4IANvPQby5zeMATtS1wCQafU3wTJScDQC5/N/NMVM7V5ADb7z2S0
22aUtBmz4xM/Fqm18NGe11gC6LCvzmru3YpYnUxT5kBxce29yXUwTcriRkrBSxEQ
lOY2UVFvX356J87e5n3i+VnAtNpA9LJehWBaFxEJiJ+4zD4f+uKGTGhhK7OkKFXr
hOiASp8k5wvk4KLSTNPaIf1GQwhidC72tkZXn0UcYB8E1vW/l1XZqwLICHyqmGPY
6YJ1W4bkwq418VbR2VCaqGyzRt3uSKqKS0N+2zNL9AzA7KUyoiMKVCtEd6rdmh6q
Xw0D8xGVuqoE+4pbjTlQ/XHFXhq9vesJY//FoO/vZTwOt6Mb1s2iQAFrKkCE5U2s
rw3F0Sas3oz7Upr4AY2UmbE9uXwa8Sv111zmv3aMHAYgUP3DYyq6gkj1M+qLwcSe
f1W3k6lgQySrveOkefFpgQREy962fp8QklX9CG75R+vwAW9kNWZ6E+kz/Z2Q6X95
Fvxa/X9mchUrvHKiPVpzKTkeOyIixFnb3pFNiWhLjMkq62U5x/rUgDETVsoVsNtB
FozMlnALQszCeoMkoUOLWJbceNbU/R6OxFRWDnBIXiMctOXJFvN4nDciaEUu9nOG
GfhazMQ6jRhq9n1Yej7jRV05AVlnZUaRtx8FuJfHxcN6pbBPmOr4w2YdSgxMUWS3
2zWqXUOk4lyz5UZDnQDxkg2k4vx1jyoMSSDrqbTt/kgW7TYC7MPTx8623V2P8nNo
7jzbydoM8BWkZzzwO82MVi7r3Xm6JF5yWi4XNs+hFVZGjEHmdmMKCh4LaNLrIv7s
3tYf+LIk714oDl6CJ6+fjCcFY/aYsCk+923VaPlgaLF/CErEJZtRpoWOadSUu0hN
5rH2w8n6vwEWQSyDmoU1zwxxvb4QIknswKCYiOY45dgG3A9CsGnbgYf+eXVMwGr5
bvuHGAHB6yKI3ofpkaiFASrO/sBcfJ2B2s9ffXjFKojLQdOS3/DvmP0fXfr9O50c
XwkJGF9RhmG+9qjAau9yM2W8sWT76P2SL44oSq52EBaevyCmze0UCRlaXqYik4jN
BOp5wiYx+Rn7Pk8QZUeNMGJmi0X2fG6/WQKZ0a/ZQ15kwrPRxDhz8ayG6IcTjiyw
ShelJyWAkgeNt3t4tKs5/QfDN1j55wtInhA+G4gJEEYW2EEzZj6HJF6Rs5xZHbY/
odbY0ofYQtbLznghFr4QsRct0SwfsXqz/tmQnZDgFvciDmng40QZFwodLuHnQO+N
/A8NxL1jmoKW7JKFhgAsdaVUW69WJkJ74ptIjtCWY1DAuxRJ8//kvkXYBOKcdPSm
cBlUkF3jU7M3KW5LMJu4chWbH0L0/wPAX7ux4j5DqnBp9XnP5NLuk1EzEle89DTB
S5SLL14vD3/+7izA4CAbgFu/gH5zCt5mGm0P3FDPc9fvWVT4v6BJ9PU726KwCIMH
yhA56JdYJWC9+CDZUPNcP5bPOyY35onW99i4E5YhajAyZ1gMkVMvA4/KPtY7FayV
DkUx2vgykEjs5OiCgnhbRkCXK975n03JFi8W46zcyy1K8HE9gJT3LQ/Sxrji6Sny
Y9wYfQrrAqzsxCWC3dKm8Jdtq7Y/dXccxc2oX3nPMoL0eQiZrXXfKQLEu6ua9Fv+
mDSW4F/7I9XlI+6sbx6lYWxBbWkzbQj1rsMwTSXxfxam2EzsM4jdPbMNvGx0TqzQ
8q7bBdBT2aKH87eHiISs49RPaihFX4tO0QZNVYT3ejYsLTeOULDAOeoG8CgK2isv
PEMwiMIJi3+i06rYYSVvdCWGvqKB8XnCMoRlI6ibVRszHrr2QAbGuRIUKW+6xTLW
S8Ez5s0aSVwoWQZisCLpTcHTU7Yo0lYSVhz5nAGDsNSESA5pQyJtANHUEgYQU7lN
ejm9h46Ah//6kpimGUUHmVx3lZJ2UMEKU1sOb6MmQXadAnsP7Q7rIfo2pFgZl3nX
fo6MnfR9A7dUr8/La/SxCbZHPisOcafwkqSxeWueSzHcxVvNelTta9bY7LPgX1bj
wGPYJrtmKMk/Tuf8f0fmtNLGk1NYGCuzUNHU1GKDXiOmXBOQmgDCZgcy/RmksCA7
rSKE7pj3sKmG3XM7jMF8F4nkDnLYKIOmiLVkuOHDCnVFLxp9xVfufoTRe2D+8Yao
j1Ph2OVhAWS6i0Ay+oaEoahbVG3GsgD2nBhP+C/qUjA6GgD+dtPymoer1j/WulMK
1KNZzcdFC1IrDFI3WTEwTJL+zA3UJxue9z+z1Uc1GIrqjRwiw/T1/RYfdXskJ31K
ndHJVeM4SgiXBV1f6tILaK4X4JKwcRsQRML+zELeQCuy71YiOZMzZ9mUUywTS6dA
g0QMNJDZJsAKtaDmO2jmdeeuzvIjbwU3ePvnQ3RBzHoEdEyzWbFBwXzjIfpclaRk
6SkdD8qe38WN4lc0Mb7PCubQUp8h5WnrZRJ+A3D/kHkX7bCYfGPW3JbznXYLPsNh
WRA1hcoDDex1MJ3TsgkQDItFL2pbJtSGTrlgcw6ed8YRSbntNQ26LWZXUsniC1jM
ckE+QQ9N1PMBlhoNZHSWYzkJbwdgjVE0X0jH3SFtkCQQYAw9kOKpa3nTfjrO2pvR
CL3ogYRholoc6OOauocBlEPvQT8eJjE5PITtPBAy7OAd4AcZErsv2l5XqxfJCerE
B1EGtZE9HJRlzLTvADsTamu4LAPlrqUI61/BFfvHd8A2NgpIsRVQks+YjdB46rom
5r6dfoPmh4TowIdZilo7lECSeIlCg/I0g0QwBd/fTh9m9DrPzTI6TwTzXkdVwejz
aqGNNJZVwci0UL4T/HSZOTolrn1Oo5ViII7QqeHoScIW2HM1tjOYgZp8NPlW+k6I
4KGF0+yGt+HZPhiJPHM+ocKVk9iD2PhShNVls7nRSg56gVO9L4yHJ+dEKCKYLSCB
72JhuxHiUtLBq2Ldvw0j5ZoMf3kW85LWN422Rj1x2OTjnLWaQeoA7uF77nEOf5f/
m3Tu6IYW1jy6Skwcsb8ZLAxsqbw3mPyvc8ZIp5XTA1T0PrxhgL195NJu/OIdvUuY
R5gm7iWgsyiZ1YFqqa4r5jJZRWZ+mblbKXzmcS+onL4BrZQH7At5qETuGHIq44CY
+VTu4bz+DeIsImDKZiU1YVk8GV79CMLnNVYPX7+3Bye+IrnxXuCLFM66bAfuk3TC
6EqZItfMzNn7l/1HRTp0wljNbm6+2pMWXfuCbvQzewDGRnPZXJWT4+JV0mE+JZ7K
rGPPUsLD9Ybam3cXVeDqOsK5fLYc40nAdEv78Briqneko37I8/l6JRaU+ulOqqNL
MNMEI9xZGExPEUInY6kR5MSWvgQCj+YJas7SEUlO7HGlvgOYXCClSYqyLXuECg4R
uh9HjJlXQL/Lkyd3CJRAES/34ekxOPzC23nS1HT3n3Ok1kGIZzPxgLuoTyKgDzC5
dDjUoUO3MktDlbRN9N/3x4NnOZx6yVVehODNWBcO/lL8lR8b2mZNp9rjjFrkK9ZW
TkGEHeCMZeVHl6iD/R2r7JyX1J/Rv5KCGMPtTVZw+T0KNLpmkCOWTBDP3CW1Mh5x
mxi7XOOsxT3eg6xJ6vCHULUF7y/1j4guViYm8ITBN+Y69JSMUd061/v3kZIyCgB5
qmX1fVO+8/aE1y1UT9qMwObG+cyVGmHbGOPBYFjIXrmhUKl+3ZzlQQnRjZZMrCqw
eCwUgA43nSYKbE1lGhSu1sZG5NgaBEOCFhoUz1tJConGaYpCWZrxccVK1l2XDoR7
sEHwzWAecZiw+RobwwABhtcGNL3qpOyb7k5CVh/k+kNi8u6777friQzfRkqZURwi
vQipX701dIkYGlXBrtvWMYHnw2NGIPjEtUxrWAeVl/v3WEnMcRzet9jaGPMwKW3k
ihJhchaNffLmIU0/ByKZKt2SLwDFSW39JyvsdovLlS35muXt8/2u4netHIwfmT2S
eLu3c3j37aL/CUtzCG2Y6L82a6gksjkdVpFvC81nORBwUpDUGoiBzCsQ/VheiI4U
MVxSzupwizkW3OGhdIE+Z5w6PpbIKxsLoYALGBy0KUen+p84slkSDv4f1U6PI998
RCBSk4AZ/1PJm15Azlqn9E41bIDs3189tk6SwPxr8nUiwZPWJrX6FyRTxZpEBqJ1
7tse4U8vK9tptuIHDhLCqA3N+tiJ6mNsX+CVqJlH1OSQ3Gv4tOW5o9m4IRZug+nk
nCo6z7S6VX7ANvJlAz2O5xE7INnhpu6Z5pxmEJLq+F5TIKjZJPdszd7//2UIoYNV
hr8c+uQmWX38SBJu9O4iRXB5ES2g/s7fYq2G+VkmHBj5OmJcNBTPWlDpvjt41ONc
DXC5yqqv06ZhyikW5o0UEKSi/1hyDil+YaNaawOX/ukA6nHNN1gtXCGEv9OpclIP
sgvXf+nLkoJV/27+n5fLxS7oQ3Z2T77OCbQex8Is1KCDDGNFNcVwsTjyUaDG9Tr9
56qF3sB8a507/94wpzwmgQViwBhSSqngwIpHkeRTWbmkXlF5qpFIhu8BM3k4LNSx
cPtAJDrDoj2NLss9U0mqvz4myCd9igd3Km55Bnm1ZLpFLUv+56YVbLLq7ccG7xmA
yj54eQ7b3wJ59Dmf/Utb/jGPNquwgpiMfsktx7EH9nn5lTbpYkd0rUN1tU65S3Jy
6Z1gp6oalj7N15VLmw32X7E9ffRrJ3x5GJ8mtPZG9M9CfF7ddx1ksTnkRLRFQvAH
ts3vQmc+QjIXwJH234GOexEj3+4FnTBlQztTNqnsLiBrfhfft7qRQWjmH01RYYAy
p1EkJ1M+6P1z0u7Qe4W+PnN1Z0Uyvd7jicc2QKXLsG+q+AF0a99+QCyQLCCQ1pWr
iajDdkXibpBD05442hZsTiZPiqcApmeEwu71kC8SeL42M3siRK8FaHGwHeIBC0fn
c+Me/KQf7HMRwNXmwQfuTiXYR/KGnZ1LeSlcTHXvFtV47z5m/WE5okgoh7IltWwH
YXtq0GCPZ80DJ1ec/Dqc+RQC9KYCgm7MQDHeY+hMw4kLRY1d8k4ZAZ1lsR/Zcbcs
Q84FK+FStrTqPv61Fb3Vhai4qWG7kE/Y+dtMvkD6VZbt9soFGnots+y6GiwSvlAI
hLjWkT3puUbGzeXtc+QVuFMyXPBkkDnMdfvlvE0sepei/LAmL3eWTiP/N/NfgbTF
GMBeQyiyAyIjPYxmYg1kQJmYd7N3H5FMNpFjvAYmK9qeFnzQaLxQbGlIkecFFRvD
hNxTSYKiyIvTOTdVZoYcpUt7Rtf8jZXIRfxa44p2eNi46R4izGf+xtUC8Wqt+rEG
MMPouPghI38rRVgreFf66EV3B6kqe/uA89FaGxTMxXQTuZS6pBKFsY1WZqF8zZy5
DCWn4c5ccVFpwar/VLkIUPSz3IuVxH1ihWXaM5kbSWg48NhBQeaQFB7zYiT5Rpf4
9/GV97znJp44sbACsgB/9eyQbMPNvZZFuPhuKzZ55Kt0nvFowC1LGpDgaKfqv0+3
AK2vByRnC3mW4pEH6lICgfwEw3wdA8knbvHs8PKfnsAHDNXejFDiEGbwxBZfF1PI
bPDwp8lTS/KHZIWmgU9++sKazEq+HNHJxwLPCFDQpZs7D3Ee1P0nhAb0oVvW4jrO
XwuJ1bKS0mnaRKSlkydP6e3S+3UHYYcwLme8gO3jZwiiXlvcfgQkS5l2DuObleh5
0N/C2C/e5GryraJnThxUVOALQ5fOzQ6AOwrUY9R4RuREGjbpYphjzMhdXM0Or/MA
gdfiHU2aIX9aWUV/TWAFyXhRvNRaU7okbIVTAJfcFGwqvs0pTuMBoX5QYs1raL+E
2cFji7eNUPdbe+UrsDVWj9TrpnF4ourWJF5BNpeNcGCskFxYfc2/xQ2krIIPBoXf
GM8aNWpHhBIynZ5SZc6uyCSkBbdhkfdl2GIRZTiSiA1b0Vl9u5eAboMCjIj5Et5y
3zxW3qWZibx4h76fO9uXjDSWzdrlh13WIlt52WnaH/0AqJLbLuG8ckZcys9uP68i
bRiOBxE232vpCE/gtKc+XJf3vgPCTq5DnqcizrV44dmavBcbGcHuckWEcA9Ks4bK
DmXCHcH2G0X7H6fIOpaTVYw5wtfP7AzEvbCJuca2/Ik=
--pragma protect end_data_block
--pragma protect digest_block
rvoks879OJbRJzrctwkML5pFdc0=
--pragma protect end_digest_block
--pragma protect end_protected
