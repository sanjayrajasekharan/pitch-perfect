��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki��Ы�T���NDm9�x22*z�*���Nٮ#�;%�ֱ����n�D�����o���F�	z�2-S˝���D4�I�f��b�r�e݌�f�H,�,`9q�&�?���w~�j(;���9�$�(�%�,�\��w�=�z��K:__:��4IN@hVe���?�s��랳�#,#��j4��b  ���\_pl3����i�Q	_;�M�p}ĸo���w�R�V�d{#<���!��7�a���R�'�Lƃ,�hr5���i@g��-<��V�C�WF`f7���883��9yo�f��h��;���>�l���=�(6�ӣ�<
�An���9�Ga|�r�J�R�U��Z��m�u??���w�~��a���#-%�՝��=	���Ob����o�#*���
AJ�4-�1q,��v]
t7M�S�f��jq�_�W�^V��T�]}��� ���'�r���������߀�~H���	9�5�m��+�O�y����Xd�M֬�����F��)��Z�\�%��+|��ipC9
�����O�� �bm� �߆D��!�R �Y�d/�����9$|��<7����꣚@~d7Xk}�U�;�0c� W+d�Yr�$�{�<[���.�Q$�A��a������$��6L�ߝ�cS�*��X�/i�8k��QA���&���Rt�P�f���eZ�;����Y��,٨��L�63��2������TH��-��഼`�� 8���V/�!s��ڞz��[*�Fm��x��Q��z�Y��q2��J�?�>μ�z�
����n�7����� �Z�?�>��|��D�N�` E�Y��ѳG��щ��?��샘`���'R_A9솨I���3c.��F���cD<<�����=��o3�.K�G��@3��|��tN�._��7g!��t��}�>��vNn�ۃUI��q�Q�h���Z+X� ��7��(a���b�L�:ŏ�($~��>4擧b\�G�d6ݙ�L��I���ԡ��1���Y�]�;&��{��[���2�;�{BWڨ�zt��f��1��غh,"��m��<W�53��#}��W�̨O�m^��ϭ��~�xb~P�}�uN+�⟹d^9�Il���u6p�������^g1b�0f��I������D�qJLWg�O@&?�W���p��r��<�Mf��N��N?�ok�{�N�CB���-�v\���4t���
�!qܞWW����Ĵe��ٿ2�Y^>��_�$��+�]���hu�)�9G���AG��c'����
����/�?����i���� ŵO��UΩݶc�)X�
����Y��k��)�3�=�wM�������؍8����Ñ�A�U��7�-�~�j_ԹQfH�\˵�>�z���!�ðݳ#]{׋g�,*'3*�
=mT9�@4()���C�9���r�th0迾Y۞�< �����/�`aW�Br�HOL�I:'��#����jn[��(|���y��E��4���b�zRf�x>/����t `��ӆ�Ұ�:!q*B���@�3{>�ی��:ʏ�_ݹ����A�hl:��F\n�Z��F�Cmf&z��ɒ"��le���W�7��������fPm��IYt�Lɤ�V�yG�?5�*�%�S��x���	#�bM��e6W(��$%8��gn��Lq�����Ȩm6��-k�ٓ-�g1A������n����k,�0��3��Ca�ږ���XQ�V�o���
�3�눓���t���M�M�:;6_ϧu�|�¡�`a]1T��N��
*��+���^x�:�Va����g}�D������}� �
��G���B�V1[�eA��nZ�ԍ��U��붑��W� �^X��4*�#���mV����/��}��>��C����q���O�i�:�*��r�x.G�V��M�DM��ä� <�/���N���cZ�ΰ�6��)�̃S���(�v�n�L�0�.0P1��Zu}UH��UB��G�Sf�����q�YnIs��V����m�ͅ�R��W*��ܪR��EC'7���S)���l6�a�E����o��ua�ԵߑU@�G����{O�{��(�z��;�e7GX|��o#j���#%��y̮�՚
Q\i����Ic���x`}BoVޠ���[��7XҮ�c'·C�s�<Ɉ+O����p��G�6k���Xː�ƻ&�j(����@g%��#������ZA{Pꏬ���*L)�N��dRg�l�M>P���Fg�"�� ��ߣ:�_�z���Xi���R����,l�QU�a^����-��|���3���kSCҟm6���!>Ҿ�-4x9?J����.�7�d�;�>J��==��N)S=�&+��tZ88��F�Db:t����ioK�g�e@ḕ�cE�^k�m\����6���t�`�e@pI�Õ�2(�Qf`�6nw�KjS��2g%\^G^\/1T��Y&�B�'Ej��3�C��y1�Yh2w��T� ,r��(ȬAiUbw����$��$��}$	��6~�	_�%y�2�7����ڭg��/�c�2ğ#d�ٙ��<��-�c���C׹���
��o֞�J9�Q��P<��8�T�l5����2R��@����Z
�7���%��\����e]��/(t`!<
A�,���z�b5F��- }JK���7~��Q�=�����j�������j��LI�wz|��f>m4QR�
e���#�����߶q.���p��DH��;*+��xr�o��e�z�D�	�7��.�2���8�On���IsjOhY}��N�[�>�	_�Z2�\�`ך��Ǚk�$�eb���h#��FSTl�ybp�_AnH�{��L���!ނ*��q�����bm��a��'������nUֵ�'#�]��6�Ȕ}{��䖭��QP����^�m���e��F�ʣ�ΥO���DB�19���.�$9�~���ʑ*7H�l`@�__��d�x2��B�#�� �"���$Hj��<xd����~L}"c7�U��:��C���x�2�g�IG8gĿ��i�9mߓؽl1m���#����<��kښ�"�����o��3��4�T�"��ꋾ���"����`�.�C\�<�^����7�!:����?�o�kkM]/��6���/�iY
�s�n�%?.������1>�D���>��&:a��23�͡������m�m`d�����]��ڍ?G7d��]�|p+��$�~�:���-���V�{�N�׈�C޳�m�k������$����
�F_k���v�S�`�x�@[~�E��l)Ǎ��G�y+�R
��#Y<��s|"OY��~�zh�~\�*����H����=5׵]N�!���ZU>\5��-<�me���)�-P�ݿ�	�p�э�4&���j�,��q�R��Y[�<
�%�_�?�as��=���ْ)�\��ُ��21)��c�a=z ��N�� !]t/b��g�
��{�Ki���*a�Qש��s��+�i#ϜdR��A�6���>�ы$g��P%��4�%F�&�v5�A��u����~\ ��;}eإ䵫��D��b��k&D�@6�Li������Ge���5w�W�H|��y�=`����js��*�����t�<K�Wߛa�Ȱi0�fz_%���%���Э6�U(M���sq�aì�&��RuR�4���_V(_�p[����Bj�x*׋�z��ZBM�Lo�W����Ȳꑞ��&�5�و|���:6�C3���^M�����=��D�����(�)��ؗ ���d	�Qq�G{��6��~L�w)���U�<�plR�o-e�  I� �.3�[���I{�K(�Eu�g�{:]��AS[�ve�wĝm|=.%&1@��Y�=CL"3y��@�~��ȉ���0G~���6KwUviӝNtxvD�t���q$�ٸ�:�7�n�����,k1^^�}��W��Hq�����ȹ���c����.�&AG~nnz'�le����d�&ڞ��f�@��s�ԡon�U��ӭ��r�Y���_"�b>[c@喌-T�1ƚ����%tj���\��E2�e�����Gu�i;~P��/�H[���af�l�k3����|��7�QB�Z�T�Y��q�:�kQ�d��)��2�D�4KN�|��	w��"n�����=򙠐�A" m�GD�q��!Z�i2���D	�c`�E@� ��I�O�M�jQ��/���s�3�?���`��k����Q��6s�թ�h�I�G�3�h4�m��fb��[�g�0.\�$|d����m��A����F��c�?��\�N�����;[D��%�1�\�:-;!Oc(�|F=b���QI���Bڼ�q�6(�?b�n� � ��#�:���&�[�C�չ����4Q�XZ�!�P��T�H�Se��};6#�����HT��n��u"Z(�����g�cqf26���F�
)�+�v~fZS���ŝ��˫/��1[�2D���L-L�lh���>$M�|�x
/G�E�y��C3I��]_�B��G����D�X��'�+2h�R͑[�hVH��xf����m�U+������d�4�'�����.d��qR:f����:>��@($K�v�T��o+KKwP�����X�tU����g�_�X�KH�k\�`�����RE�מ���p��̰/��x��+�?
�0|����2��m}w���E�฼�������U���_��f������R���0��M�~��>#kiZ<Syo%�3���h��T\Y@=����Rb���L�ZH/E
g�zĪS?A�5��-�E� ����UE��G�rt������I%5R�lu������+��ih�1D}2��7Or6~�}}Z��	�#�R�1@F<07{�}�%�C��n�Bк��l�@�AU�	9!r��2���β�n_��t�E��W�������Y�g�d9ڸ�zz�/�5h��p���:��\�v������O�r��P��:�u(��wn����< ��#���9)/m(�Q%L?�#{�����R���.�` �D�;T9��B�����+�d��Hbg�3�h�Uyf���'E�����-l��/�f���OK��c��O�H�)�����sCa�W^�Cf�ӺuqT�j���w^�g���n$�H�XB-4��u���:SL�u�l�0BiR�		7OR����5{����EǙ��xb�L+~`�Z?�lg���3c��N��ͼ�F��-�[�ţ��W�"Zv�S��}�K	Qc{[m=~�����Q!õ��F,^�Ac�%�u3^1�&̱�������3��`�qg�؟�y�RXlXN���=�>J����9`�Z�!�:.�eZ˛��T{&[+�O;Sڥ��㊹�\q sM�xgEP�Q4�+��݀1QeZ���]݊�'9��#����o����ݥ�F�Wjh�{�!&�����m�@/,�%*�� �L��+'�u:�Q���i�L�8%����>�6SU�r�^s�A�i����:?r�tO�7UZ۟�+��.Mc��ö�D���ա�@����_��u��Fa���xP���uh��l�|�>���pM���#�&Pq��L��1���9Vu�65E
WײַW�֡�RNB��)^���	��{2��I�2���f{b���Yfۂ ��jb9��FX���zLAn�F��g�of��d�6�����s-ۋr��/.OJ
x@��E$SF��nr̩�n��������sQ�c0@�=�P��|��-T�c+�eX+���V^�����tzy��^�46�H����H�J�����|�Z�iz~�R�=Is�Z"&<	0A�,$#�	� o��|�?~uDz�A(:���>�2.\x8�>(�M��tmF�7����l*d�on���<�~�us�`L_m{��)�@s:������~w�[FEkݻydT���ёjϻ�1�"�(U5y�6͕��L0T��t�2�5icg}: m3���������к����&�$e$vj �\8]�`:e�
-�U�!�t��X�B;�*��u~f�	ǑEGHB�n�,�g=��*?a�䣏��,g�Ej�r'P:�Ľ��PX��k�m��y��<�ޞ�߇`�	Y�N�>4���/l��1��bw�7ݖ�̛�F]Y����n9g�S�i�����B<C:$b��h��%��9���00�T��@s�ר˾�^6��t��J������ha쯓F�:���[�� �wz�����a�W1_Y�A��C|�C��%�����a���ML�}TЃ�Oa��/�����a}�|�?Ǿ"�r�������/H~�������pr��0{*`i����X@!�aZO���w=�e��F��Nt�tH�)�k���JY��z[A��R�_�����k�.!��!d���·4h�K�S{�����>��t��q���q�ɋʨ��fD����X�.�9���"K��V���Z�ZQ�x�P�N��s�XxƜ�6�M�'�e����{q��mwz���+ĘJ%���e���T/�T6�.�oU@���]p���I	;��7j�E�?���WA1j�O`t Q�x(��R�P������&o���5�ކ�B5[�2����,<]�x�x����� M��\A���;EF�$�чN�ƻV>U��ko�x��6���rH���"�Z]�4�mQ�؝m���~����v5 u�a8T�v�HoI� ^�@v�!:}�H��D`�������ԝ���=`C
)Avo�����}�i��	z�[�g̅�y"J����&)k5�%�SM/�&�@*�/�e��Qd����A�ԁ��}�������͉h�G�/�d���G�UǸ#���S>�E��7bۢF����n P���$�]M=�vVƫ���@�_�^e7�E������2��<Z5�}�?��p�%^W4��'Y��|�1"H��Z"��=w��J��M׋O�0"|6�q�qX�6��.fp)ɺ�N�ـ��ﶽdhBϪ����K��b��H��yL��]i[��X��B��Q�@!��?m7#K�������?���$�c�7�Ku���,�����t�y�����f��g�O�y*�Oh�e�����IO=%A�z�x��=oK? ���v�rꊋ����??����ߨ�n<�O�C"QA�B�8׼��Aƽ��.�ef�)�cr���흇8�e
zi��?����4��-���b�^�����]߻�������A�:W4�-�s�8��Hf���K�{� ,K�P�>Z�X*�p���W��Z��7kP�2pu귞+=զpWnN�w��>�b�H槐�4�$!��"��&FBpt��MP�E3qq� ����HV���Dj'��T�i��#T���d���+k���ln6�MW��X�5���������Rxj�Eǔ��J��� `x$уi��;��9+YP���T��B;х^x5b1�Nj�!��Zu�r�f
!� >-�sk
��wU3#�͑)x��������?��mۗ+q�6�/�j�*`�T�\uq
?��=x_.;C2����"8nQ�cy�N#����2�JW�����oJ+�}n�}��\�H���|Mg���ĉ�NP�1�R���*a�ViZ�1` 0�$}3�>�.C�T�y�v��j���~6��V��E�:_��~g�u�6����-y�I4�%��c�O5�S�;���Sb���J�Ն�{'�k�]8~ȃ�����i���eym9�W�f�OO�=Y�7�*�J.�%;+PT���*�	�M|�ͦŬ�e��I��) �ޖ֢l!�wd�G�� ��l�V�@d
�Iݓ%�q+{�:��dRQ^��6je���4��S���?�������M�FFz�u�lt��?��#�����oo�V����7}l0�`nlkD4��<�*���I���b˦�jye�替p�U���ɀ�!��I�>��Qb�_�-_��%��\zO���z���S�NVJ%�d3a�OꯋD:��gL^mM�_�"�ˢ���Ґ�!�M��o�P^����Α1�<��mrtd���]E���I�9l�7�uj̻d�`�S��6�~(�q=�;m��D�h��L�B��!M>Y�B��q��|��&nG;w�%�|��1�N-�=�J���X�r�T%�S��d�s�������m��2<-�ԙջz�&֤e=L7� "ᅝr$v:4�^��4�a�q<C��܎�t��5�E��56�J}(�4����cESK��rtEX@XF�9e��wzϋ_��X
&�����ҽ�}�vsGY������%J���WΌ5�/,�s�b �*u��J�TxG�	���\d��@�&��1����d�=w�jD|t��yqO���6�|{7�.�������B`�p%�-πs�ڲ�ϴ��v{L	>��]}R�v��Q=�0^	�S:�µ��	��Et�~]���x��t�yi��-4�;�坏��m>=�����2g'�� ���z&q��ԓ�|�n�1����BN'��
��)�-yb�8x�Gځ���r��%��@B\Y.��gu��H"'=3��!�E��F&�v��U�]���H�&���<>��,˅�x��d�������FZ=��I�F��ڢ��V����%F�,R���7�i�RM+��g ��'��Σ�7M�@H�c�m\�wd��C�{�� ܇�:H��*�]�o9*'����JI6�H~��K�c���Ȥ�&��<��H˳�/���=֞��PTH��پ}�F����bc!��^��\��ﱟ� �����r��I�{��>�T���J5(7�7G�����`l�3
��� 1�G �]&���+׭���d���}�0H�n��jh3[�f}ߵlʂi\��_�vD���B1sگ����AV�@����ݾ�nKK�C�Ob��ﳁj�X��Z �s�9��s�5�����Պ�lbt.��O���';=5�#�0�	E�b��_�����Ԙ�v��z�1Kd��X�y��0A�����0D�&�GUܙ'Rrܞ�2���݀t�� ��(���~}w��<����93ȩ9��A�n�8-��`�Nzs�4E1^T
^�����fZ�7:�Y�-�y֯J[�Xk�)&�x�"�� $�^��T	���/����y�&fK7�@eDZa���SdrǨ����Pe�΋���H�-���V��A����a�I:V�҅�b7����:~'��$����P�}�p�CA�c��g�hIVy[�i�	+��yr�T�Ȱ��۪ qj�K�2Bͯ�k�a���n�;�TJ:|�F�ԥ\p{ٸ� (����a�ᒎ��3��q�����݃��"�W������f�)'x�u��z��&���[U����{��hT���%ŀ�z��f�u��d��~�iF��m���������Z�Ns�� <���l����������|�y��*�?�X�`���>��z6�<er��rX�%Uþ��g��"=�5:<1��������<2� �x��c�hw�L��翴�֎�z�h��e@~�,۵�d�|�윂5��>է�s�h��q��ߧ�C4؇���dYR�"��O񝑼�sY�Yp��Y�(��բQ��/��8�.�dc�H���%�g�3���o�GTߛ7 <���y���Gc��K���t9�z�"Z�ڹ�Q���#d�������4R��H�y��-0h"�L(�>Vذ#z�hV����n���ӔAL�1ӌ���Ƭ��XP�P�O(_u
���������J<@���ġ^?
Y�_ՍF�C[�{�@�d#������|i�a���1}�uc�%�->~�lS�9w*��{��ؤ_�0<-!���~M<����̬�z�y�<p��Ak0��D��������v֢�z��<�����pAi��,<V�:�u�\�{T���4���2����E�b��~þ�&n ��.5ғ+���&';�:x��D[�2���ьKļ)]�i�zv����3;Ä{g��x�q����3��ד��Zi��!��C�	!-ś�
��8X=<^1���PG�!s��sX�ل�*�|�73��׃kwzt�Һ�1O$\iB�#.�uSa���3k�z� ���X�.|��kca
e�q%�Rt� v�����Y3_$xYg��}2�D�g��[w�w�*�1��=3�Қ���s ���!e��5����Ad�C<1i��ݡ�1b�Ղ��J(^\+OZ/FG)��%�w�AC<T�+�"��V����^��Y��C�o��*�k7�3*Q��sx�Ι����F�nl)�|�Ħ�+Ǐ	s��c)ѺBR��S��1��78A;J$�4G���b�]�=7y^��Os��<}�Z��3��`箽b�*I�J�?�� ��P��kxpI����Ϛ��V�[��'��W���߹y��r�[�S�H{Ɖ���$S���¨��R\ �l�ya���*NZ�$�h���OD�P2���L��WC�4�����,dRJ�NΙ�c?�����I���&�4��O�֤���p�諦���7�(O`h7G�Pw__�BFEl'�S���l�{���s���_@�.��L�X�ʺh��`�خ��od�?wO����Y�RD ��]@�z?����#�6�Yy	��d� ݱ��)�ޣӔb��hOa����M�b3� 3�M>^Ҕa�?��o��ԗI�9?��i`��bDr��2�>��Ϛ�	e�`]N��	�y?��6z��#D�g�H�Co�~ail=�%[�'J��I�k���Ud���P���F
�?�%"rT��%K>�w#tᡕ�c�ʙB�HW� p_Z��s#�Ŷ\��O����������8�⿻�*b,�ؒ�;Dx��box����;��!�2�NbŇ*H����?L�h��	WN�O�a���Q��Q�D��hd�I�!lsް�����f�ٱ��a��nՏg�aqW]N(���.��#��<�%o�8��-�ڙ��.)S�Z���� � r&a5Тx�6�@�[آ���LJ��|;B���㇀ʽ��㒷@Bh� EZ�A*q�.l���_�I����=6��$�n}���3DF�%�pCbm�b���eT����'���׎��n�B=��މ0�m�'�5�.E;sS;�2I$ͫ}�r��`�ω%:�#3�x�"�E��������yu�����'�p��Đ+@���9��/�}��:_(L&��%�vqg�&�r���N����ịf16B9�O'-�[����E��e��4�]���8�?�K�Q �l6}~�_�i���5,E����~�]�񢫧*�UP���~��QD�^���Q�Y�h�W�	֬�KG��Ӥ؅��4�M~�X��-�>������t@�'(�3�`oG�%�(?��L�M��-��J�c˕�G�P��U.3����Vy�ڷ
\�[�90ճ��ⷺq�& �!��W@ܺy������qw},�-v�f�"���=&1�w��`���l�TU�����"���嗳)I�^@�ITy-h1�g��l�6U<I�9P^x��z�|RG�:�N��W*���;_���\#�&� z�\(���hV@2Ѓp2�t�?X���û����-�ɵ�Zq'ʖ����z�>��1�>�F�9�_g�s�v �]_��r�Mc�<���t�]+��H���bY�w��kM��8	�VT��ѫ�3�	+���X���#��0'Y0��ok��
��Y78�fw��bލ(V���v��k��Ի ��"���[>Z�c��8���ͳYj��\S����Lɷ��-6�6�Ƈ-��*�t�:9ѝ���og~S�b�W�F�93٭���_o���2�:��Ν4c�j��8��o���S�P���_�j�q�	�p�T���D��I�(�	�<&@n���L*ȴm�ǀ{%ƴ��Z���}~��R��?������ۻ5ct��x�g���KCf~�%����:r\�Ǘis�dV��aKt�� �B�atCY5ΞM<�u�k^8^>� r�*��#oqG�!�D%GD��5X�W�����R��)��^�r/N�}�Xzmpg~�y��D6�����������H#�����M<~�Y�M%�������,梶�5b��m�>��G����Tg,�J�`�n[����E۞p�3k�W<�C!�����Y}�	����K�b���a�bk
2��S�7.��֜E�۪,αgSL<n2g���h�N����i���G���J�`�Ph؄���[�~Y�z�>�R�������e�/�G�����~��98���M﶑�	�[���m�F�����3T�jD��J�,0!O�� ŭ{��U��"pQ(��r����eyo�*ُ&p����u8 np�_ܓ���:Rٶ|�#���R�������=3~���u�k������JX��!p����Ӕ��I~|��C��G[4�W`^�w)}l����Y�uq/�*_	��X��hхH�_�!�]�z��)�)AJ���Mb?��Z)*�,Y77Y��sP�7�#B�A<V+sCň��
���~Z��{��XZ��A9�HF�\ܬ�kT��Co�lpP��ͻ �<:��@1��9�:�!Ѥ�<�<����� �?&��>�~� ׶��L���\��1"��0�5�퍑-&ڰ��x���ߔ��n�(����t��q�q��fb9�1���:��fK&�;f��D�S[Jˠ9���L��ކ�2�*(�����\��T�����#+�2��{���Cc�tD�m:�O�s�ۃ�aїD1����ܞ�b��[���񶱲���1Z�9��4ܠ�
%i�ٜV���*��AxH�k[7�oT�6�45�0�ݗ�H�i���w-tw��+���A�Q,(����§��D�oZl֜h��I�����R�n��L�5�浡"���� �$p�|�zV/�R�c��$^BS9���"\zb�K!�Mc�m	��(;z}�,T r��%�j��<����G֛[��$N�vcV�XGͯW�v��Uv�I�8��vl#��]��:�ȱ��1��'�7��ii2f����|��E ���u��cUt
�1d|w��,[�ߴv�֢�����"���5�z2� �t�/��r�������87$��P�9&шZЯ���ۮ�{��ɞ�����r�|	>X.4��� ��z�ߤ��-���3�Z��	|��ZN�˂k6����ߋ,�0�*����;����Nq�!�d��8 Y rZ�Z���l;N��j���ǉ�bq8�b�["H<d��6����:�^P@�X�=?�o�G��[��5��M>`ݍ�P�?CFn�jJ��%��ђΊ{p��ڗ����#�GK"-���5$n�,��32�����^eE�k5S
|��7�`��Z�a:/~�?�G�������ׇQ�]TH���u�塯�� <�?����O_s�y�R���_!cj\���d���:C-�!T�)��`N�<G�S�xî*������oT�*"�aߣVs�6�z����J�09���Z8�f���F������l(s!e���X��_�T�C��1���y���}f�4�0�'�[�����opB߭�H<'h}�?i��'I�z���y���'J]l諲qv�z��M����`���Ȏ�x�����C1���Oڲ���M7��W�j�oN�N�E!?g�?����0�F��eMb~�O��K'H���;����B�*�6�Y�-���lx�?�TU\L��9^�Nj��GJ_��#~jm�W�b'lhͱ�q�=$�jY�v�7�n��g���xWN(� d���L��ǒ�u n������\%��u!����QЧ�1?�rw�aI���?f%o��7&�@��q(��{~h��t� 3�������sY�;/�'y�(c��,;�Y* ?�/QCCb����We�;�fs��w�s�Rq�;��?r�9+�]B0Og�W4�Z���p�B<��ׄ>խ��>��(պ��=��4d�·��[�pO�@�@!�=J�-�5aY���]I�l��J��NW�[�)�弡/x��C�d	���k�V[ q�~D���s��t�C�Km�b�W[ W�����V�{A���{Zi�u��O����"`��ܻaA�Ɂ� ��uT�D��-�ص}f���QVҁ)����U�}_���'�â�V�ߜ�yԶ\�"������"�=@�u�]��)�̻�{���+��=�R]��U��s�z�3#���z=�&@��*i)��Z����Rt���P#�]�� �cS�H��8i��g^�ƪ���m9ɞ��_��^�9��|E�;v�ן|̿�P�/u�ʋs�d���'��*�T�)��-T�D��F�j�㷌o�wz�ݔEp�8����ԉ��-V�q���D.d�-]b�z���T��(.�Q7`���"��f��q=J�	8�����������m6�+�0=�oȕ=��'��K�g����\?�4h��s�t�A�re�̎H-N�rS����p�BHb(���8X�y<:�M�����Q 9�����sn������$����a�喿n����4Ah{x��1g&m��������._h:�X��1$���N|C⨱8�k��/gY&�R^���_W(44�p3nV	�%��r�h���jc/@z�}�c�.�Ē�wh�w��M�A�y�_�J5�h�����D��^������"��M��*<�0��]�\���F>`�440��s| x�,}J�����m�zP+Ry�xVA))����S>��c���y�lG�k��2�F����<s-��w���޺��ҍ�t�(v�/a�J�`{��"$a�`6cN���K]3CFH&W�a��8�R������T�OS�4dK/9�ﾥ�Rfx<��>	�H�#����s*��`\nH-�U��/���Ò�8����0#H�=�H���`��{+|�ȸ�BX�c�a�fo����e2����y`�hX�WPr�:+���l× AE�,�H!���&/�k�j��T�7ٽ�,��P�~��;�28=D�BO��#���d("�H?��=��/n�6�C�(�j�؇^�xN
^&5O~�ء��ng#v�>Y�/�����Ϙ������I�Ǫz�����]w��lb�s���[ݓj�u�_O�'1A��C��~�$���1*��\iD<V[�q�a���Y�)�gzh�q�õ<w�oTh����Oƪ�0k��_HRz���E��_�rZg+��6�{]o#VB�Bw3#U^D��^I�~FG/".!��9���eb�$<ZHs� m���}�vG��k�[�õ40���C6*-tY�p�h�~ч3,�$���Z��y
(�$׾Q<�հ���e&2�����������T�� ��=���ح"}����r�Ƭr�j�:>{|��~��P �KY�>�wBÈ����k�P&ȣ���pu�V6y���9$����F��bM��ѓ[O��I(4��[���H�g�����(@a>���"OQDw=�|A��g˕Ԛb���}r�[5��l���2Ce��g��U	�ac�kb��F��-s�i�a%��_�f[���`in!�PRt��?��Δ�<��oNA�~��o8@n�O�� Ax���1P\��̾��v���#�~���߻�ѣ�D_��)�Ɩ������k�.��@"'��$�~�yV)^�������-�ɔZa\^@7�FJL����ad��t�}O!�I�8+��Nߔb��U7�`f�>X��q�$���{�k���h
c������f~�
ﳳ����"�çn*��O���w$���=�ջ��[�mlPJ��-��#_z��S��8�g��Q*��@��%����R��uhP%��Zq�ϫ��T9 *��.k�~@�����ׁ�L8�&^�{}��&�L���|*+�N�{���ҕg
���v}I�:�����z�W�0��O*?^n����l��{+<�E;7��=�;�?W������3�5XVc2R�zل��H��>���h�~�P����6�ڐE��Q��iv��$�x�*e@c
���.�}^3<]�č�Vx�!�@��b<����7(�Z}�I֔�;�b�&����7K�8�~�7��Z��~�*�/FO%8�G�A�-e��4+��.��6�\f����\�E���&y�t�.�������Q�q��*!ʲ$a�w�������\�R�C�\�㍼	u�����P�;��򫝒#4��թ�a-ȹ�tԶ!�[�O�k�V�h�19�́�*¥T�ǥ������A��������I�呍J�Ӗ�ڲ��z	�E>�w��"��.����ű�q#MHR�%�J�ǉ2t	b�� bq�\��$XU+o����o��$s�|�`��58�y(.7QzO�N��5���ޥ9�冦�:YN��̠��HAy�w���e�z�=�ItqW�e����?�q+8�\����.Cj�:�A���s�Y���>0��\�U ���W-e|i"J#Y�Ou�
YMP>:��7�h/Lx�Ti5DP.�q��Wuʴ���Ѽڇ����p��=;�f��A�ԉf���3�m5phS�/OT�M#R����`����oRj�EJ]'#�/h � ��n�\ݠ��������c0^���_�����X����;�_�'�Ǡ	M��p�'��&�RWr6������12��3O�3�� K�DcI�|��Q��	l:��G�-İV����'�3c�[a������y����s^���OZ��HFY��L�vZ�(��3�1�@.��:!-l��e&��<���tơ3�]Ǧ~3�.��}ԅ�óʲI�nJ��E��f�ԙcE��9�#Pp�2?��k#�wfM�j��IhU?���6��رإ 6@ jT����
"�@�I���#K++��� ^G{AB���f�a��C� � \ A���ho�Ry��*�	m�w$0C�����~�
�[v�\�����~�)��m9.Ń�}B�aA�N�h�$6xdNy\���0�s'C
VY����q�}h]����[{u?Sg�2I��9	1�lW�lS�gu��>����A��Sv�B[�۔KT�J����_Q~�G��3^��ӭ���@s!|�\^���PQ�y��X���.�(A��Y�r��ꛆ(c4pݜ|����餒�k��[�d\Ƒ��<"�D��S�m��{O��˦˰,�C�ߊVO�T��·w�cl�� �ޔ%^�:X�	_�o�
��!}�3W�Z�P�o'fS����6'��ݎZc+�-3�=�7��r�F"���-(W��ڹ���S���� d3��X�� U�8�KN��_�J(J��K=ue7:鰅!�CΠ�&WY�����VB�o{�[��?�ͳ����}Q�eW?�rڇɱ��;���ę����ԼI8؍�׆�q\B�Sk�Lٹ������C�R�m�`��V�$߈���Mx�0�b���=j��X��<��,ᢗ���>�Ͻ�����*���џ��� ��/.�l�ꜵC�|��p���{��N��ܥ��p6��G��v�w�=��� 	+8���W�9&�g�^V-����Ad��)�����b��Du�Ş���/?�yo;�;�g��uX#�I�\�2cq.�;��͏��&E��d��~"d?w����[HB�����K�q����.�Z�$|%�����7����{����*)!���k<W�cΥ$3���J�M���f�����>Ռ7W�@�B��Hw�K�,b��	��� no�K:cn|�R�}�X��V'�D���&&*U�����m9?[��_����p�W}Au�L� ��Z�;ģ��u���pPm�4��Y��CE�nanIB_ A��ml��O���*��f`zǳ��+���!�b,l��x�dNv��*UQ��7�l��������A/���.p5e�U�-/ז)��D�.%n�47�Pk�p"������~O�����<��TS��1)�H:�
P0����Qx�J���pG��|�!� $�m����M�7P�wM�W���,ANg����5b�&7�?�	��4����M0j3�w=VP&��L�����^A�$Q���`�_�W�w��;C��x��n�2�~�x��{��a}>���UL���F���`���E
^�͉V�fn�g.������v���4���&�� vxO&H�����'+�r �Bv�x�f�$k���^�����ί7zH�*�f��-87~�C��r���������GZ���N9Vq>�.����n�܍%T�;蕉;xR�7�ڂ%AѢˢ�X��B�-4��&�qmQ�e:.3�=N�����*�`Z
��^���3IH|�W�+������0CAOg٥!��"z����5��ٓ�o-� .5Ϣ��l�ELZ�̧���_D��L?�/K&�Ef1QN�)�Y>�A��o��9��l'm��3�W �d�g���C0�
n!-��1U)��$��Q��g�τZ��$Ϋj'21!�,������(O�@vK��b� ��SUyع ��*h;M�y4��]� ������IQ�j D!��*����K��I�t�ӘmN�$����h�{MrC�1V��T������T��k�[���c���<Ղ���H@qa�H��\m�I6�R�e���#�l�	�s�Ջ��R/�Ԫ$S��C4�kN?� ��L��	�ko�7����gHݸ���GER���ƿ=�g.c�)�y͠�/t������A��m�@���v�f�i��BVf׊��`_��֬�g�\�'�� S�?x�F?ěڔs)�)1����M�-J����mC'�}3�S�;�,<����� �]cZ�mj�W�<�(���3�LC[YO6j�;�C�[�m�<4;��4?N�n���EUn�o.P;ǈ�7m�o��T�.P����mp��E�AڿL��eG�0����I���-*���7�y�h�>JKʋ���eEqq�q�>�{�s7/��� ���eh�+H�)E)H��A��W_|7̠�S��£�X���5~ZjШޖ��I�#}�1fN��&� �tlB���"U�ʉ~µp�b�3ưי�`\����RT_�̠=��t�;#��#��O^RP(�}���+M��@?��@��hO+�7O*Pg���.�4H^��#���� ��:o�}��py�,��A�$W���+P�RJF.�qS�\UQD�?�=�
DŔ�����Y���2�{�
O�o=����x䫷�N�;9w�U�?7�>��>om��_�g�,韄K%]E{��I��j���d��8 ��B�:^`Fs�lG��kr�4Q@�O]���C����;v�8��?��IZ��6�hD�R6*��u+cD.(� WOl��З�?��D��;h��n:@�v*�o#e�$Pn����'��
r�B�i��M��P��C�t�^��ԟ�4��N)��/3�O����qU�j@���沛/��w�Dr�}�j�����a]��M�Bon/c t@*���u�Z�x�Q#6�Tw�2���dִ'���D��Z43J���Dm��Os:O��A���c��db"h,`��@!=�[�K��8�Q���	���bb�=���\4z}n�7��T��yx2�K��mj(�*�4���z-u���~����h�����SgSը�GŲb�A��]k�A��5%�S��A�;݇�T'���C>�덍$�ѿ�5	��?%�Pʿ����NnF4Wg�Aʮ(�d��p�!������H�/�˘ذv�o��Ȯ2ާ�2�[����c�<��*�v>������*��)p(Z��2sm�3�W���"���)��䤨�����쀘S���ܹ�� �(B���ʠb�A�\z �zU�%<��d�a�iLȹ��ԭ��"��*:���J��8��;�����y \.[���<�qr��_s���Hu.'<J�!3�ΝX�=�q��U�_����8%����T�l��Ե��k@�)��'�3�.R�l�q^^O,�Ҷ�-(����3W �,�IQ"4�v���<Z�e���;�<U�6n�R��Q��X[}&l:�B�Ca�^�x+U��Tu�._�����%9�C?�o5��aC�e�s<gܼ�t�8��k�6O����ێi�����ix�+H�9P�5p��'���*:|	�u1�|���9�LP��%K�I��R�ǪqoC�,�c�Z��X�x�nsgP�Pky.��T�)����I=2I9:�^���EѸ1�7�=���fx"�y{ǰć�N���g�!ф]�.��.p<g���o�e�f����H��B#(ή4DH��3l���oK�I
�+ΰ.#�:'������.�s�S&�rq��� �/p q�:�ڭRT��<�e(S��v�����-�ϱ�K&e�ȗD��ً
g��k��E,mV�:g*Y��)�3J�\R�F�bi�䉞|؎e{�8@ū�w���n�8��4��E�-���<k�����b�ʸi�鋷\��	�u�Ai�0�>�I�M�d2�-��C�����u�:X�����5�%��=�������c�j�3�:��D���y���L�@o�-��F���:M���&A���4Wg�!�6-���::,]�[�O~@÷ľ�_aҭԼ�٫��-��p��/��YT�G���Y��y[�`��a��.��R�<5�{
B�5mƯ��j�@��djt�4'�tԥ]:��@}0��(��3-�C�<Y@l�җV������������i�=I�8�pZ>��F��;s��
� "�O�
�
b������`�TX#�s`<�(:��	^�K������L������z* GTIP�\��i���v�֯⋶Qex���Wi�I8 B����d2�&Ձ2�.�3f��$��j����cH3��S&�ʏ�|N��1���:�"um�ʻ6o�?�H�E~�d�����d_����=�2_�A�'�ƘG���Vf��F�R�.(�͕��q��znD�;���}�c<�'�n�i����	W�ȇ=w�GE)��y~�8�Z�Qm���.� ��[C�Ƕ��d�������ϋ���莦d�x|.)Ab+�<��TS�z���t�]�^?�I!BU������'7��O�y���;S_p;��f�%��td8{Y��4��Fsj<�i6ُy�~Xo��8�;���Rr/��ݰ�b�"������li�ό�ۚ��=�G�;�`� 0�� $�Yn���C�_��ыJޤT�=�fhb涑@���|�TOZ@��:K��񄮮��"U ?�C6ps:���7� ��OW���\;Р�um�@��|�'��1�,R�nL<��#8|����9:�
k����N������eF)wr��O����>�ӔRF��W��{���"u�L�����ٞcͅu&��J�#,M�1�L�ij�9X���5�`xj���j���6�]k`!�-�6�Ͳ(�	q�}�8x�HSn��-�߸��d:�'��(^���j�U���Q4�۩�܏�`��Ɲ�@B@�>�\�r�`�s�Yů��TҾ�yC��f+OkxA:{�}P�kr��*�GOy� {�ل�HqG�I<��S��6��r���n��np�|��{d���#���+Fw�2�'�U��A8v�:�01��h����g������G(��;t#�|�fŋ�]37�tǽ���0� ���$3u�T���� �ĕ�;Ý�&��d$
:�\�mA��"8�}�^I�����C�b�X�qFm����ۨ�GN�����l�<�\�Ƨ/�K����O��'��qby�ځ)�����xc�[�N�\��ݕ!�Yk҂�J�
�c?%�|g+� ��^i>�k��P��!��,끆KV	�ֆ��������:E/����  ��|Bv��1E6��^j��U��د4��(o��X�WE�GI�[�O�%%-�RI~��3�0z� 0W��FU��oTooe�c����1�ZH:�Ooe���o��p���XIK�b?���7���#:M���y��6~�?���7X륱��$�T*lU=̚��
;Je�2bZY���BK���'2f�X^�f��3��C�_(�0�Y>炩l� a��Ba�����T1��"٪��s�GΞOx)�z8��V���G�01?����8���웠������F"���V�`�bX�+��7�HZ1Il_(�,��� D�~YZcӊ�{M��y��q5]Q|��ȫ��-�ճ/�O�ܓ}M�{_�^�~�TDV���[y���P�����u�JRkh�*���D���F	�5�	�I���Y7��Y��{�>�[y�b ��������^��b+�XuQ*������ޭ�1 )I�`o.tmN���b��,�$w��,�^L)<n'������b�����	Z�.H�A8�S��7�th"��v���!pصC�9m`�?�o	��sg�{,� �Ț��l���۶p��M��C\�f.H8�����ȱB���bT�ْ��"�&�JPuF?�3|
>m�r(�/W��3�*��p7>P�b*�]�W��Y,F��͐��V��7I��[⺡w�Q+:Ū�<�;"� Qn)��L���6�!��rٳo�lI�����Q�z�;�G#���E�=�}�S~f�"�@�r����eoY�J&�oy@ics��`�b�);�F�)2��o�K炙\���Փ+dh�{���,̨M�z?q`��g\Կ�9J���a&'����Y}q�L�Pf85��M�m*���W�NY[wQ2�7��C+�MgqYm��)��b���Oy� JE�/mZ�	F�B@�0���R�[�	贙|�w�ҝ��~O��7�)��pb�2uf�9E�<=Ët0��CY/SG����O��=F�D�&�}4"�d�-g�:5��6�n ����a�vuH���EB=�_k��4��/��Ǵ}5���xt���j�N�@�'`��W�1:���7c"D� �K���rod���p"R��[a�j^����az|gٍ���@�_ +���a�7�⷗b�I�أ�2o;,o�C����`��d��H9�r�� ��#����<;2s4x���_�ܡ�W��D��O\�����[!�4�HO��UO�bB��Я����	N��t���&���H���r�I�^����3�>1{S����aw�<ػ�J�WM<���^�8}Q�X=;!�ji`.:+ '�ʌ�VTu��c�SZ�0���Z��fK��o�$�B\?���;"ӛV5��I!���3'-��Y��L���
30�h]�6�G ��1u	��)�םD2��ksAD��A1������d�\3�>�`�l�r�=�5���_ݘ�w>}��SA �7��s{��{��˟P���QS��%�B���wKs�2���� *#e�6@���ܟ$�����5q�_o�����w���(�$��o��D�NM%l�{�e���"B���MHCq�ا/q �8���%�w�e�S0�Eb�_9������G>��j��e�ȫ#N���*h'�`i�Z�gp�*��`�x[�f���{�+I�3y3�����`������ 8h��D�����.ϸ"�Q�z;��*е�wp�k N7>��|�J�S����	����SӢ0����%I�ѱG_��n�i�帧W��P���gא�N��.�{�K'>ϑ�}C�whm����<��k����_��u>�
�Ћ���y���tI�Ъ3��o��������������&ا&_g�ʁ�x魭�6���>��߈17]��N͖����C�`GaA�L�lO�Us_ebM��ke I��Ƴ��$h��H���/���f�t�������E�WUl��r��i�G�m%�m	�h+S�:d�*$��px��Y�������ԝ%���I:9@N�Qr��ުO���;��p�[F]Ӎ@�4��WB+:_h��� ��D�r�,O��������/H籆y$F�"ƽ1`x�B�=��ǂ�x���un�����&�@;�I���!�\��flG�7т
�VE<������q����]��3�&�
Ͱ��5��L����=w�j&��V��C�wr� �5��b~��U������A����@̵��~�BU�s)�F��r�ֳypMr�+0;�LS��<�o��B��-���8&��fkp�m&�`D���a��QA�h����"�hVa�b)`�$�O���ߍ.�G���&u��i[����E|`*m�����C��{�D��)��uϾh��\�>�p?&'��%��O��i��QU�éK�oS�>.�i�}0���$(Άߣ �;�y�p�� hgf�b��C����a`��pR%�3M�ą�.2�1�̜zڙ]w��S{7)��/D�>���WwbkX��psj�X��R�����'&tL���ÚCqh��J[��_0|.�"Zo�Ԯ����������p�#�_@/�����\5Q@��'�RC���i-��Sj�U�r�C�<�??��\��-p�k��u�\��GQR��$�}�Q����cF��{�����D��P$h�"$ri���tn� ���HxD|��,櫬{�^�a	^LT�N:�ִ�b��{�����歖p��ǒT�t�=�		���e���/2�2�汒��1�ѽu02"M�+�.`�Do�qE0"nx���Pkp�R�)Nf:�>�U����F��*��9������ч\?�	�����`E^�ߥn� 2���<
�y#28T��/p�b9z)u����$1� q�=4�y����ĭ{�x��O��iV*zō�9X�A�T��8Ս�i)p�1��EibS���az�Mj�QAVI�ޗ�#x<�S6a�ZZ��(��@\����&FK������q��HA���Їs���^Bjp-��z⬼(oϩ��n��/k!Ô�|��E'	�$�I�s��;�z���u~�\=_%�{�%��z�M����y%jc�c��q�:�<=�2�[���$�b~^��r��&���U��JY;GV�­�Ag"��+��E����s�&X��U��P
���X?�9�꼈��|�V��\�)�K1�3�6��s�>�Hw��+0L{�5��o���S\�L,���yL�Ǔo~S�dk�9���-�њ�`����A���A5����|lF>ХG j)�`�N��y���G��R�W�ޯ��%���-U�����6��b%���� o��l�7Y��72���g�?��G��x�l3r�j7��8�z�d8G�<�W�D�>�
���N��<5 m'���Z�/V?�rö�'�b
����u���0qT��w �Ĩ;��U�=׻��4�uE������j6_�}#�/�cb��g�.�%!�(ܪM���k%�Fl4ʣ�ma�]�\�ƺ+�:?��_���I���e:���U:O��@o�����\a2z��vc�8<80s���D�\�u|O<IB���)l�.@�E��V���.��r"�C�Y?���`:��AG����4�/����aO��^��q�#����0�1F��[��-I��P�eU�ᤄZ�2�ez�+���ȦτJ�l�CW+x&��w�s�st�Oal� XA,���wc��a9�`m)�B�&�m�`���u����s���/�����3BQ�������s &$�C�vs�Wrј���MWY�iZ�,�N�Ʉ��v�=���
��(���K�b��a�Hx���I	�Xpߠ�����4%�_����X�o�]�#���.{J�Ȼ��vʄ�db�����;�H�@	���L��D/f����G$��K歃�i`�/!�iP"�*N.~������9�c.C�+u=�u
�t��(�F'�OA� ���Z��bRu�l� �"�(}�%y�Pyk;��-ad��q��T~�w���D�!U�	!)��9 ���4 I��YeVM�֘�?��:�"t.�w#�_��W��'�Y�-�j��vġ�.	� ��tQN;�/�E��/�\�;�p��Iv,���8G�k?���Yu��F�c� �oq�{2T"� ��ͦ�c�<(��|��"�ů��	[���ު,�Wgdþs��O�Ȼ7�?K�}E�:i=`�8�+s�N٥��!swШEW!���2��1���:��E�K)Em�(�'{(������.�*+A�R	ԩ�ޭlH�Cl�$�j� ,��2l2��B����5�Q9��g���o�[pQt����O���hQ�Gh���r��(������*i��� B��ҭK|���_b,�q�Ā-ǔb�3e�T�I������hAR����|�%}�)��zg�����i����ن��)��� �p�ޓg�s��
ɽ#����r�:��w�2��|�
#�uJ��a�{AS
�c��j)�4���*��z��$Z>�S�h�JVmmb&)@:]]����w�s���G,�"q��������
%�ϥ�}F�ϝ�j�I��겳n�U.���N�Gn�$��\�$�?��q6w��������/��j�x��k����� ��:���q�ߡ;4���嬎�[���N�1�u
�J]����o����x��0t&�e��:���?�~XfJ�/G���D�]��;��W�9�&����<��%���B��  ;]	��r(�K��=���	%�7��L�>b)Df:oʁ�O"Cp2m#E���&������,}�����$���bŸ��c��as<:��X��"�y׵�p ��>�ka|j>�{�/�Co<oh�KЮ�Uc��5ʅ���&U�z�!�f�V��e� v<ꈽh�.?n��<�T�]��M>��߫H6�o�H+����q`.䓝��L��R�ۓe������Zbڇ��$0�&P�Gh�"W=|�\䚄�ֶh���s���\Rne�\e��eʙ���_d�o��/�]P`xWޝ����7"˧9^�%�g2>�i�
+Xͺz��
s�G��4��z����e��U����z�-y{Z�NMGy� 4��m�q ��E u}(���)�u�Ѡ�}�&wJlQ��r�=�i��I�ўi��Q?"	�N�I�F/�Om���Rv���7�1
��� )��H�K�*
&��LĖ��©���{w�|�J���������{u�xR}�5U~N~D�@s��~�;��ѧ�բK��T��\-�-�ƙ�b��j��g����kǀA���W<Q�ֺF��*���2&�0e�%�a�5����N��
�G8��Q;U�c�S�>�P���~7�q.��g�Gp�ۅ-3�:Sj�%����Q=��xc���&0�our~*EL0^~A+��ɗ����?�6� (p_�������ɉ�33'��U1� K��.�H�:��R�Z��c*��b��6>�s�pލ��W�`Y-�3��W5����dfI9h����eTȞ�t*� )9}�44��D�C`{l��$�?Ā�^�m���AIM��;L�$چ��k�?��SF��Η�cĜ+���D�����~<a���DfŴjaE#��ޚ�eP�A�C#��bʤ�mL�d�L���8E2.�G���c^(X͸����?{^sa.�+۱��[���z�'�+'��(a}�4�K���8w���4R���b{d��n#��*+�'�M���}A2����!���7�^_(6�<�T�����e'���$�1[��M�����_����k�N�N���w�7�9�w�)��_�ʰ�����jI\rLym.�������.�u:������~��9��!�C�u;��,�nlD�*�?d~�]����rs����:h��H�>aT�g���q�j��Ñ�e-�S���:H��\/���Ba�\��x��e�)L��<�9�xf��_�di��*���Z?�ޢ���C�& �=�"��M�E����ެ��u�wf8p�[)Hf8�?h徳����1wކ��IhTymϔQh2C)��s5�	+���7�u����{R+�01X#^����c���� U�+ɭ����Y�(��1W�0�/+n+-��g��O�Y��;�g�	+	��\�S��u�R������V�wc7�A�q@�!%�5}(q��zG��FV"(���ҕ�
����^WCD�m�q��m�U�<�2Ȋ�L5(�$���K�|Ny=���ɭ8�b�9���]e��6z3at��`� 8;�� Nm�
m�_�1���`���?٩���K����޿e�#��"�L7�9(u%xq;"�F�ح�r @r�G�$ s��h�ff��ԟ���II��̔'�=�n�������i��(~���)����)�S�Ҝ�>��lbF_���`+N._!w46�CWS&ϴb���Hjg���8�A4�L�����9w�v��2� ,[��Z.�O��X��u��јJ�EtM��#Ĕ�z4���b�;r���ye&p4���������A���o���A��֠�{y|�ya�ؾ}eP.;�mp���_�^�?���FR����@���f(l A������.<q��ajq�T1!=_������~��vY��Vz��Vc����ą�8���Q�ml]%��UZ!{R;��z�D@��"����\ۄ+����gN��[Ie�Dh�$��K��l�J
�NI���<�(ݹ:��L+5�'JPC�tU<w�J�D�W��|��E�Ǻ#��F��%\�--���1�jy���.t/'s7{����2b_�|6ge����}?kG�x���^��H�ow��8f)�M����3雷��MT��.� �����xw�?	��ۿ;h�r�d��F�~��ė���4ݜ��VSu�S���HU^8���O[Ԝc��?�X7hI �T��kx��X��BJ�|�\��d��ڐ/DNX��ń�*���cI�ٞ���p���_���@�1��o��Ӕ7����_���JNf�+c�l��0}'���d�:����v��}a7,���$�Z�(V[�>d�Me�@/�yo�O��B�p��,�6,���a��e&��X��7���4O,�7��!�U��@Ht=r�'�Ar\&s�\�1���������zȀ�-��O�P�����l�"$:iR6պ�_w�b.����̤\e)n~{1�u����m���J5d�oݣ� c�QI�)f�H�a3�<|��1��h�h�������d��N�Y��d�"��;��[h��7k��
Ə��j�2$ݛ!#��(��-�G.b�,�0�>���FB���Wa��K{�����=��x��c�IA���ý&��9�%� �h�+L:&��Dg_oo����?+��CH��{�A���Q��\?vu*:(:@'�vP[Dw�<��|��-�>F��?��і;���A a����K��Ӄ�Q����I�^��x���k�����\c�d���<���_�\��N�+���m�:�J���o7u�v��xce��"�Զ��qX�@%�+�Tpq�k�(����:
&"��^pv�5�[��HT�
%]��_�D����t9 }pXo�6����y�dhXk���Vcs���M�*>I�k�c���2�Ws�|@K 6nb�u��\�n�{��w��=�$�;7�������B����'0���CR��P�7eV��rhJ����p�:F��7���?�MD2���M��	QyY*�j�`Sk�!��u�9\=���k\}�V��}��f�gSO!���^���$!�iS<��VC91K���k��.�C@JY{B��c��90&t���_;��n�b�*z�r~�/	ک��0t1���/�$R��~
VN+BB<��Gnju�]�}Lۮ.�`�N��>#,M���-�u�h����E��f(�cS=�Z���U9e7��b�7ɻ�Za٧|k���N��eo�i)��oT�gu�ep���NPRx-��2r<��N�G�g�s�ݱ�ol��aN%8:�P���v��h;W����;:7�cS�O�CMK8ǯm"�����J7����E����<�~G����{7�:�6��X���������-!��c���!ͦ��P�̐�MOU�asZ.;�yzdZ,նN:�n�a��m7ü�,7���U�G {ԛ!���>�(z�]�$wc6b�N#�!�q�^��qm�Jmu��g#�7M�7���Bɸ�����#B�
$P4$l�G7��~����:�v��#B�Z�!���'!/��넮��zD�UzoË������ru��i���)8e�F1���(��C���jgS���ʷ;�^�K��wқJd+f�4(�p��q������ܪ>��=Ù�~�y!��1��(>�ʂg�=�#���j�X�X{�[��	y韯M#�Z9l��N��*��F_����.}Vɸ��=#j�����3��"|�>�y�W ��0H�����mض�t��&�_۷��>,Q��8�&�XBdrӖ�'�X՟~Í"��c�Z%ï/��/�+�
UԨ�.6'O���Eg*�>#^Q=Rς�;<�����g�P�NCUxN��ܛ��C7
�	��V�M��'�@����9k�`*+b{S_ܿ�Q�l���������6�ߝ�,�V��+a��@撪�u�w�®Lq4\��&�ڶ��p��w�2�IC���T�U��k���Z��hg�wJGp���[�y7y���.tKQ�gv� #�VSL��k֝�z�܅�6د�w��ΐ�Z���/�2DV�ͫ�9m>��РJ@<{,�d���"���?)�Cz�� M%vf�0�\-X���3Q�F(O���/;\���^u�]ZW�C���4K=��m,�ð1����~�fl{�d�!>��ys�9igU����ݩ��'	�%��3����G�E�6��ip���mBR{�PWֶ��r5*��Nnb0��6��[�Y7���U4X�vV���]�{��7ek%J[�\l%��(I��%�^�T�!>U*!��'��U�tz�ת>��<�#���뫦ZRL	��)���햑 `bS'���Y��G�w�i������=yn�r��o�eஇ�*%���$�����:8�cTs2��9�&���4����u0.�4,�$cDc�N�8��=��=�5Yr!g�M¤!����!�c2ԝ������'��/���� ��cUq7�õ�0�V�nȅ�A��<��J���Z��1�4���͍��Cmq0�h����٨.'<-�ןˈ�r���(:~�n����t蜺	��>�F����I/8�r�� �Èv�
e�0/=�=ϭ��u?�h�L��Z�'��C/�s�F-��/�g��F3T0x\-�,GM���В�*��o��LD�]:��s�"�xmM�H�iH����P��☱ Ƕ��C;�j��{2� S�ŗ67GcHu���5�����`�T���ᡲ�d�C�`�N�G)(�'$m{�|�Q����(��uwy�ӽ�2�ï�&���:ѥS�Ԅ�V�S����F�1��Ig F���R'��d0H�=؎e[?��DG���#>��U��ɀgh1h��c��% ��z-��6[�)�+�ګ���Y�{�� ,�hD싨�XtǬb�+�/��-�����sR�G�G�LM� ��&h����ž1M	?��CU��ënJq���X��X0��Y2�z��[��m�S:�y�Q+$V��M�B�+�Ru\iaZ�4��Y��3���w�nT��M�(�4ǫ�T���h�7�2�6ʔ�u������Y���|� R�:��N�֖�NYX-�C�7�פ#d�(�K���V�8gʤ��'^�3�{����{�;)���f�>�/�y'���BL����%��8ϯUƌ�d����@[����i��������/?<sK˱D���G���׬�dr��;^3��HW�x�����w1`o�b����������!5�|�%V?��S1֕�}ە�xr�z�����5��@��9b�X]�ؐE���'y2<�'���a� �*��|�'�0��
!��P->������|+6ty��6�p�S���\G̓�
�� vk��(���:	��$_�c�	Z�/LT	T �}�����
�1Ȼ�3�j,��|V ��*zo6�� ��6:A������M,½���n�A����B�Ҷ���u7�`�:���&Ϧ�rG�p�݃jM@IV���'u�&��I���8��	�(5�o"��e�yUF����3ݨJ���D���u�"�7��t72��jm���1jY�1�_�C���>1\�u
�Fa?�3سwc��u<L��j`�*����N��x�����/��h��.݊�n�rŔ`*��W��r�q��x%>xF9E�d�����>�_�A��q�V��;X<�#�n]ε�uKn=u�7fbOBM=���p����\�5�4)����u�A��d����׻⊞8N/�D�zi	���t8q����vij���4>)6#M؀)����4�,_��ؓ��"˔��]�"��M��ݫ�ش�H��K#WQ/��m�0Y�ȕ�4��]W��"�1a�=+d)��5��<)h&�l{$�yG�����|� ֛o��7�W��ᇆ?��Et|љO��xԵW�kJd���m�@j���[���N2��)��Π*���k�1+��l릺�]ߌ�T�q�ZT�.����S �y�N�R-}�����	n(r�uHw�E����DX�E�)���'A_v�6ai?d����>?��C�B��6�m�˫о�̧NP�W?{�'M�i��2Ӑ&��=�H�������W���]�=�.�i�[u�h��%�0���o���V�i�~ְ��A��THD�?�L?��3e	�%VKs`i(�<m��xk8���S�K`�B }]�ΒG�>ed���������H�tj���\�U�w;�����V{�p�M26M�S,�f�ۮ҃��5��1~���3���| ���y�� ������l��0/�w�=���P����,��2L>I�#�b�>+�� ���L��i�=�F����E;�D���3+d��0�%��Z�8� ��ߴ��t�Y�/tB ���$��"��d���5�!�-h�o���v'rK ��`���S�&��"n�؜`�o�LOLf�4̭}Y�/GL-zt�s��
���8�`��2[0���S�xH��9�?��5��[5����k.�y{�.o�@�#��/;MJO}G�Om|��8V���}޸�]1< �)�M�ޟ�W�/��0դ��(��߁Ì��Y�_�CY�P2bJ�	�������s��9�R���S�<Ca�n��2� ��6�a��}8�X��]����e�L7�'"��V@{-��;̵A��m�d6,��S�� O����Uvwvu�a�6D��l�%��'�'����`qY(��7 ���O.L:�ҕ�~��B�py�3��&�Vڟ��l����-;6;-i᷑�������A�b�zK��U��=���q":�PîtpB4��t��H#�,��ǥYX{ڵmz1b��h�Ud�7^��_����(:�h�?�ݢ���da�Q4b��Y�Cҡ5pRٽ2�8�tۈ5��3ſ�)���j�)N>�*Gl8�����~�vŞ���>�\�ن�~I�+"ý� /�lqd>)`��;5�(�gT���=�vȫ��X�N<��)�c۹��s[�%���j�Lk ��傸�a6g��{u�4��v<"R@H�t�]������(E͓��&c��G�Atb��|���L��CU���Ξ �@.f�4�j�00�F-#Q���q
�����vd�/g�N���E��/[ R}XU��qhM���8r�g���[���xR�C��͟���#8��0�� .����&C�}�!W]="�����l۫�>�F�`8Aʦu�M����:�ʃ���8g�U�U%82䏥I!B7������ٽ�HA�$}#�(x��I��#M԰;�M:�ٽa��?�Ru|�ި*/"*��G�J�l��"�S�|H��g��%h1[x�ץ��e�lW̸�G
�v���m��[.q	��H����ώ�,7`�m�*���ͽ܋ԓ�(A���%�������T��띷�J;�Z�k�(m�L��S>�v�lh�R�����|��:�`���L��$����1D��"��M�t��bx�cF�Fˮ���Z�&�*|3+�����ۏ���-�9��h�N��r�S�| Y���(��Q��.�a�)�r�Ol�hN$�\��=�[����cg���� ?��8s���].����J��gհ@��Gt'�?��kŧ�P��F��$N�*�.o)�P�m�w�>�<��M*r����j������� C�l�$����}qi����.I�� �/��/����N�Qj�5z�Su���27����M �&��ڸQ��IAW����٤~m�p�I�M��R�j��~���n��J�21�BO��f����o�0�����zjlt� �����bq%~�11���/�'�����4�������4f���C>��i�]����\����%o���w}ﾢ$d�Q& �s �t�56��ᏉFo9?�{7�"~�n�F43���Cp��>ȧ�1������.e*�~jh^�7�-�ڡ����d�߾���-Rꈣi��M��UJ�/A���5�� �}ߴ�hT�O���u�	�j_� �;7};ě}e�b\. 61J��L��A|y��E���30�_�m���5њ=�{A�Ũ��U�����)w+L. ۲w�(bz����\��'űs&�6�A����)Ԗ�2"�4� FY�d�Qi+�jJ��A��c���:7w��L������ۦZ���^�B����4ћW�E
��J����h��(H����D���3zі�E�(�X52��3�]���*o6�ao�K9>�l\];Ʀ��ޔ�yD��� P���I��&}RϷxH�?�'FW1'�Z�o
*�:�u� U6�d@�S�U�`\�T�&`]�1��i9<�~v^�ȫm5��c�-{4#���#Te�ax���W��[Le䨶4�4�g�s���:Č3n���!�r�`�Ky��٠�%c͉��I�˄8�Ϩ�##��vQEʿ���/��i	�Y�����H!�����O��E T'�a콉yδ�M�c���'�<c�dB90���>��`s��@n�5��A8�=p�?q\ت���u�2p��Ea�L���pV
c��+@	Ë����?
A��k����P��jÏ�o�2?� ��y�?����� �>3�����ue�Z���Ta�������U���JR��3H�f����(c1�u#/��2���?0�'��ǽ����I�y�b=�?g;r!P�J��0���ZE�nj����?�q��>�u�_껍:N��u�XQ�xe�gcs+���D��p���"��KB ^�]/G ���ͤ��>�<�ꉴ���F1��~���9�ƨ� �
��ǹZ��L%��I���'�n��̀�j�[�y<��ss횡�\2
�B7	�f9�Zr�ʾ�;q?�F�N�x+˚_fc%t�tn'�Uw�Y�����1V�"a&~茛��8���;;_M�b&
/Q۲��Ե����7�@\�Z;⊛��@Wv^`fΉ�$8El��O�Nz�2(tT�L��.7�9�BgE�p%Z�6�z��ƌ=��Hw?x}&d�ϋ�(tR(X���
��DA�/>|^���Q4� q5?��OsRGьI@�1,�m��/Z���=+S���H0T�X�rU^���~~0�o�	z&�?_Pg|�8�)�ō땗\��S7���"���G4Zl�:��������/�:���;�{�Ɗ���l��T�j�����E3T(G}Ծ�]�	S��->�d ���K��6vU,�;��q�s�{���z���4"��ߕ���Y�3�.�ח[����	��7�ᑓ\b��)�
�{:��]oKl#�}���7e�C��OWs��H{f�t=o;�� ]�����\���`WVg�O$�ߥ��au�y���0<��Z�}�'�|s�j ��#G�+���ܼRľ�O������#xlgx�
�<C�,����ӁtE�>�����">�žg�~��T7��SX.����-F�'�����JL���v��,$���렽ܗj_T�
;��g'¢�%��C0��~�W�����Dt;?��~�P��=� ���]e��O����Co���
������B
7�m�	�y��aOE\�aJ���rA�<<�f�pRBs�/qD��4|�����66�~2v��p(�O�J���K�"����Σ����7ũ|��PＲ�x��x]�pU(Q� $!Fؠ*��AZ�!q�S��H�c���gT3ią�/f��y+ե�h��9��t��t� 8;E�-���9�+�>�2�E���af�˛�i���|��6�C�ߎ�yV�@Υ�ڇ'@�Ǽ�0�^�%�+ic��o�GV܇:����A�E7/�ݨ��C��������6 �J沺P���{Rp��τK��b�ۃ����%f�MطS߫���{BM`�>���5�m�Ck��6�4�c�b7�+��wʱ���SG4�}�=XT���uc�� e��a�B�n֐�f��V�B��%C�;Y!P�es���#�<�����0~��	:�Ƈ,� �1I��>2�;����.�K, �uۋkE�W�T�^�D?�n@9�!��0Z!~���vtһ�3�%4�e"VTPw�yy@kw�fX,<��|f	A�P����n�^rO��wG��AOoo5��M�|x�}vU^o�8c<̘�d�S5��@�Jp����k�8��Yڞ�n�5f%]H;�1��Y��R�=l�EҜ�%j��ojl*I�;sCzd�$#b�Z�@���x,�F�>��E��=�1O�\��w�괜uĞԌ���S�
��l����
�o�a,<�|�Thx���[)�`�����=�#������'��!o������.\���5�z�n�Vk�!s�cX�|8 ��Gi���q ���˖�D�s�gb�W�N`KA�F�D�a2�N&N#p�~���Y�<Luw��ky�Ap���IqȒ����(TDth�(]	�f���yFs�6d�P㶈�-�I�����t�T�Y*��e�E�->Fzuۉ�O�"�y�4 ���$Njm3�,M��i�.��q��t����1��k�"j^כ֢�v���h� �>�h��Q�w�>̕�&~�F�>s9�>[�U���Qt���=�a	^���1v;Dtyg�t`��%�`�C
TA�c8�´�Tt�#F䲖��[F�.���a��:���~��wivO�/��N����d?�f ����E���2�ɵZ-cm���0���� r-��234쌕�ۉY�i��a=p\� kl���^ݍ<�s���C��sG����C��y�Z�t�.N~����+�R���VD�Q���%fk�-��˸�#�f��h��Jf�e�2	�)��x`�ܬ��J�~��߲�c�.��^���ʡ�Z�--��I$��hQ�"�|0Vͣ��D�n��uZov�O�9ҙ2`w�(;&��`���E6OL��R��UFh�'�-Q�9�Ȥ���-��th��E�H ��X��	>�Kd�qe�p����ON?��	�n�"�1�G��.����*�e��>�{%^�\��(ORY,"��j\�[)�:��.�f��~!��c���29se�@sx���t��`�l����ߔ����S@a3X�� }��Eƅ�N�X7}q��\O;�!O��D�N�ye�<��$�p�;�-�@��W�(��}���Qe���m<� �B`2�(@=�Z;;P�����d+�í�;������^E����6�$������̯���#ь�qxF,=�.f4:HM�9����<�VUc rH�LA���:U~���T��iR�i��S�ݒﴼ�Z���Y�H�mDUC>����tz�\6�p	�7�I�8R��	$���{F��?;�+*�S�j�`Wģ���G9�GW6�5�����4����vg��-�h���Pu+�o��:Y�E��i���s�u�'��Su	Q�6�ī��bsэ;L�'� �F#s�չ������1�g�jX�uZ��zx�;
w�t�f�ǖ.Q�D�m�*r5׫k�ϗ��Q}�Q�]4o�B�6*g����)+�0_FI^�J��L*��eo/��~�[Yq�1���v$O9�����$�Y�	�FG�k��"�#Q^�ҝ�7N���}iyS���H��wl�<��PA�z����&�;ң�y���[*�Xܦ����������ӳ�BbۉޗzG�X(�]�2!R�J�=WķC�e�̷wq_�����/�?��������9� �Űc�u��0���U�o���t��i�]��t�Q�{M����'7'Y=�G��yi�kԦ�Bn�;��"���2�)�ב���rM1��0�H�/���R��k�
��3/2���b�y�Bѵ����l���$�Q�T���G<�u��.���&�og��Gg)3����VQ�w=�
# ��K!U�����T=F�%�޸w�X�/�4Z@�/��|ݡ�tY.MG����W9�}�dǺ���Q&_,��*��E����kŖ]��]���N��hn��0�����&=k�^��*&Sm�Q\���l���'\���=�>B�y�s�s���������b�f;��C־3;��Y���Y@.仦[76�l�Y8�hv��F�Dx��3�t�$_4C4���ZQ9����(�/�� �¦��n��U���G�ZS��_����@�4Qs�{��I�VK������Rh���IK5�>>�"��2�H�xfd{j�2,}w�m�
����nT�%<��
�U,mJ�.oح�WH�Jl��=�� [NB�|{���J�7"�˞������2�LYR0d�u�!¸�;�4p8>���Ҧ�����x���S��p�r13Xg��"*��K�@vH�ud��@.��n꡵�WYg\L����b�
���ə�俫VGia��~I "�P��x2NF�MV����t��SX��]�r�pi�0�x�Ve��$Lᣂ��/ͅA����!��D�Ugm�9Ґ �]��*�ψ��+�� ���Qy�_~�����3��@T�ǖ���q˦��G�T���e��
�#;��<�$?��P���s�8jh@R��\�P�3ŏ�fl)�*+vp.m��k|�b�mV�� ���6��!�91}._��Y����:4���P�@<Ȕ|\[0 ��a���c�����[W[�9�S�
���ܦ1�eOϢM`��)R�y�иSo�$���}�]��=;�&x�1�Z�y�Όj�!Xy�e�n�b���9�~P�E@��f���C�v#7ױ'9�y�D0���0��D	
�+�p��Ƃ��XBG�b�,&@�B��3�k
�%e�r-��|l�+��z\ب��դ��Uԧ�A2��<����4��!z� n/�5�oĈ�A���;&�`�ǟV�s���j�S�F�}&�|�"x���)��kn�}�OWWe���n����i��Um��|��\�8���R�ɓ�)�_��잭�"�^mi����3�. Ʊ��)���9�U�7�J6l���3)9�=j������>����\ՠWA]s.��GK��c��4}��H|�)!	h�٥�M4���y�t���c�hչ�~zN>�\z�$�%�i�Ho0�an�������y�ڮ�=ʩ�H=��M3�H>�h5��x�*A	���=GQ��1)��fi/�X�(Lc�8/D�z�Fb�_;�T�7I$v����؇}2ISm���_ٻ[1���a��Ct�Z�S/_b�zN8�G�1͚��P�
���;]u�ty_��Q�۬+�Ø��n��+$���h'��c܁x�ݤ8�X��C�I���(��z������F`)����w?�aY�����:^�.Q�K�쎐ќP��1Y�6*;�أ̞N<�w��_�A�$N��t��W�š*��{+� ����)�F �-b�2Gv�:h+=�6AY�2��@gkv��$���Z�EP�u�df��A1[|�/Ԩ��E���9�s��~6 �폚� f����4���p�)�E�/2
�٢A���(� O��e���N���:7�Ò^*���l�	�w�Je\�� ��� �U�F�t���B(�=����nIl���/�!*���V�q�b�[K�T�1W�ZHcA���T� Z���ܘj<�%�3�'�\�/�8�����Ō]��[�(Ee�n�ࡢ@a�r���KO�RO+x{��V�q{�UQ�����gw!��/^���<�������o�큧l����q�[�V�~�u�N~��6�>q�{,sؿg�	T٘�Y&Je3T޸T��8A�E�8�H�������B�6 ����u��~��ޑۉW�P�:�#��������?Q�fs&��>��&�څ��*|Y��5�'�k�����{�c傎MX�)��Tr�D~�
��6=��n��'��,p�V2�d��~�tX6�<:f&P�A�0h��0c%����nV�"����Sǫ�Qj��;겖��u��x�9σ�^�6���s�P�����w����nIv,3Ø��M�=y��/n�ρ�w�g)O�+��2�US���</��E1����.��m7ܦ����OM(��x7s��S����ƥ�w��Bsd������8bJ���S2��R�^5~Қ���	��ԀDTz���=�P��\׫,؈(Cݏl���g�(!�ǘ�pU���`7s	�R�4��eW�	�n�0)Sי�υ_;�ja"�z���;�?"A9���g�� h�3�K�-���=������Q�����+�/�$��е�w�����e�KAX�*��0�%��p̴5q6:'IֿވI��^�cv�k,nṣ�`C�,*�Է>r�s�L8�/]��͕bi@s�8s<Ҿ�'�cӎ6�09�|:з��?��c�7d�
�+b�F��y�j�}4�`nY����A�1�<�ֱ�I2,�Z���m���c+���h�𡓊̣�V+[���<�i_�GC������u��r�Íz�>�*���Ԟ�������7g���p�*��]��#�+���_�8gA��)b��or�����]�$U��_�U��� Ç��\"��$K�e�)��Ψ�NE��F!�2b�b�y7�����L�"�ͥ�<�>��(īVh���$i��ΣdP/'�z"�WV)�,
|\�w�h��u �zn��Cɾ_ڠ�g��l�aց�����R������g	��8/SM_
75$:fk��`�����������;+�$ׯ�x0�-d��.�V��W]���a��_L�Xn)7�B`1��Dp���
�
�d�S<�#�f5���zB�t�%9�Zo;�;���>@ޕ��(��=�O3ݘ�1��B@���b�1���e�%�������5|�Q����2f�筚����B%;��"�5����*L����H�v�������*������/hj�rҀ�B��+T��@�F��'�?�LG4vۓ��P�di9��Y�ԣ�S�,��&����`�#�۳@��8ez�\�5G1�t ��a�4��^D�=|���6#d8
����5��A��5���7K&Sa�WG�+Y���We��ƺz�F�!p�:����)+G�[��b�P��+������6�" �w�3tc��	����|�S�]5u�=2��ƭ`���.�S�ZQ�2����e����`�閶����rsP��_�����@t$^s�3Ј�M�?�E���߰}���E�|�c��k>�6�����
�To#���4E
%���x��$tUiI]�����e�I{+�&9�q��^�>0�8xemK<@5�]z&��#�Ƴ��6T,Tw	�t�G�"<��n�K�ȷ�^]	������4�YJ�K��2�1wT(-�`���f�~�(�=*;��F�v���>����V*�a��qi��Ug�Q������ʹp/��5 ��A��U4!��3t�z߯����l(T������1���u���zCͻ^��|񆝿J^���D"�}�D�3���n<�q�:w��S�`8v���� �U8�x�h�X��fX���F�Q��ZB�R���>/K{S�Ɔ���m�e�%���U1���PX�ү=���m(\m���:����xQ8>E��{��NÒY�9`�t��]�l�̗!� r��S�C-*���[�6����Ձ��΄�^�!�<��R�l�������E�tET��������^�\�^W;����C��1�թ��-v�z_���SN���6�n4�x���}��c����x�:X�Ft]�[�r�3o/�f4`8���e�[��h����su���(2��.�]��g�`�V�|E�eI��=裟���ᖯ,� א|j܄���ȭ'�FK'�⼒T��ͫ���8��t�U]~������� y���{���L+X�,g�����:��>��rį��&����|U&����70B>O�K�K6�Qj�6�TJh6Z���J�pf��=�y���zyW;ff^ӏ�;{���w)����m�!�����~a�eǣvt�:�?:��-u�Q�:��ތ����o���R���������e�>O�1]H�)���WkY�/w^^6�J?e#�ݬ����@�F23�W]AE
�쇹\`\���W<��i��L@:�jv��w5,�|n�:D�Jm~
Q�HvK ����/.�F��.��b%g�+�%���d��}�P�ׯ5Y:�J'.:��:���v~Օ�_m�h�ྍ?AzH��"��b��� ��@�|)�*���y ���H��⸼Ѱ�qB(M����۲���:�я��5W��k+ d�a��j68��^ �U�)�M,8�g&"�r����t��* 6�`2�w�L @$�}��VN�#�)��oKa I~3�$���DO~i��F?�}k�Ћl�?��JSvP3������On�����;�G�
A�[�������a�ա�a@�2��"�(`�.�-���@r>M׃���E�"|z�jXz�5[YҔ�8)W��i��c���9�$�z_���� �y��B�LG�M��5�?��e�^��p<:p����u�i�pŉ{;��E�נMhX��Wrm��E��c��8O,�5؍�|W���N=�B��"�ue�G%~b�*�#�@:ֳ4@r���r�ŪA�:� �'��㐏Y���M�J�UV����,�p��?�^�Ŧ��D��C�w�j���i�rR5����'�o!&�p.�q��" �Cg�F�#0\pC�G3^MP\_nHZ���s�%�k�"�k*�U��	¸	�@�gu4��T�Ovh�$<]Yy��;�(Z
��t@`�I��,�u���)�;�����pU��~�N�4dH��F�d���ۣ�K7J �������=��h8Q�ne���9�+��ZdRJlq�oJh���wr��Z<�Zg�*?3�7���(&T��dej����6�m`mI�t����+�k�v<�Н&M^��A
3n�{]��ގ?�d}����4E�J�����Gpcy�$B�n��g���v��K�ⴵ�'�T7R^����?�ZW=���\E(�k�Eu�u��l�Ѡu'�n*��/�E��:R�V�8�xA�u��� T��]1��Ǟ�}����!�P�8���B���U��M%A�����x���׶��y���!�1����Husi=�i�k���-�W5������A]����\k؂�P&79�i�>�i
��oSE�j�5>3hY�����y��9�.�*ҷ@�q^O	S�:V�Z&�@�����TG��&�����I�O���s��C{��%9A'�X���>w?�%��7��5х3(��'9�٨��EqZ'R�Ie:h�i�3q;���f-�9x��#:�$���bp��͗��4P:���4kH��ȷ�j������[��@�]�tWNzCj��>��1��IR����2o��[�O^Z(�e�H+��Ē���� �=h��g�Q�@��8�=H��1��F��@�[���)a����������NH����iq�GԈt��IY�Z�>��*H�$ƨ�~����]���daD��,���]��K�~�k�"��IP�2�;ZW�h�k��K	g*#�{���ת��������Ph�NU3�=��V	���a��䑻F�ɓ�����3p�]A�3)� �������xf�2ʪ&�;�[�g'���
��� �h�Z���(�����,&��[���fH�3�zM骿u�T�V�=@.���&���p�,A��w[yL%�] ���8��6l�&���f)��I2���g�h�:�!;������Z�
������3�!�����X�����&��S�1�߇�\#n��P!6��Ә�щ胛����}]�m���9����|U�ܵV4М�/{�Ͱ��
��k��ڠ�c�0���,�.O_2�y\`)��a���m����N�/�vs�&���*a���<�e�$M���w�S�Q��r3��*�|;��oQB�"���+�4'��n��e��k#�j��`�ֹ�ִ}m��纃�3��#ӹY{2]9B�9�w��N�О��<���;.�w_}n��\4�7gޢ��
ܾ�p��1 �њ�l��d����
^�Y���� ��i�0��Z�Ws�t4M���x���a����j<!)�ܼ>@��K5jt��F����L��yu��Y�O�����H�_,Pa��"�[�Y���,�*�q8�0ܬ�z��O�*��՝ˌX�4Q����e��Y�?1F4�Z�58��K��l5��� F`2���M��G�!R��v�D陸�r��bʙ7�_���{ו����谧fԁY��i���fr7p�=�0�#�y
 $6dtyǖ�Ѐm�P[p+�0�5�w�_Ƥn��ayک�BW�t�)_���qʬ�E��ڝ�t�Q{��M^��I���g�L��`m
t����P�M�����v07	O��;M��0k-�w �f+��/�a@�����y]T��
���"ׂ��*��!ڜ'*� �e�A.ja+�1芷�b�������j�[V#u�#��\p��S�e#�]���W����v��r&BCJw3��� ZN���+�t�{g����-�'�1��(q��E��y^|�X��Z����)�#_]/&�� ǂ��.�PNGSD��^S���?���.Nk���3�G�ƥ�e³�P}pk�2���%	x�'�B�J�
-wZ%��7X�r������Ѕ��LZ�a���9���8�9n��"��N�.���TyCQ��?V���l4��#҂��k��9��TB2Y<o.\�P��a����䲍8]Ng!����O����sƲ�`%c-�Z$ټ T���?v��")p�y��<��	�+�W�/7��6~=.���K[J�)��� ��د�����Ђ�J"��':�-��y���8����]F��C2tAJpa�T�Y��F��Y�Z,�C�I�
i�"��_���K1p�g�����)�b(W��㞴�?!���_F���룶���õ��?V�#��\������s���ו�'�]��X���o��Qt�If�Fa;��j�u9���#F�E,��w+ ¡u��	�>��l���u�����T�rӴ͊��L0��v�\����>������M3ȼ����	�^|��j�fe��oGjy�2_�p�˴9�v?!��N̿:�q"↍k�Ƨy\1��̃�Mv+�q]��/��5-p�x5�����Y�����!�^��_Lm�J��<�C���R�*Z�`��p[v��A�)z:���I�������#܄eg��W�^�]���Vtb�80�:3?@���J��E�����O��>m�|J�s?�r��J>y�+Wp:V�ac�9�^W8��T8K����4Ǵˉ�i4xAONf��+���ܯA"��R�$���Q-�pαJE����
$<C�|���S���j$(W������B��2�8�xw(}�J�K����C���m���� Ԁ�V�U�x�QNh�X�!���/�4K�VQ���l㉏CC�5}<�!��J���M��͐RXcKE��GJ�����~u�H�����^;J�*Jz�T�>�'�lcUK�RNz�b��(9�|�~��7��f9pM�^~D�\�؁�⊋��E���o�g�gl��̷�j\�c��N�;[�a�/at���ٯ�Y�*���59-��v�y� �2��Vc�,pXPh�Wr�	!����]+�3�gn�1!*��Xl���؟X�W����*�T����lɶ��Жi���i	,��ێ�-�U1�,�>�_�D9���T������F0�e%c�J�so�k02���s��pwqg!�w+VwIs�0N�tv:�_uY%܅���{)�5��I�N�@3�f b�Y�V��JX��{��@D;���e�B��ӋUe:� fU�H�m%��rH�'a�!��[���U,�%�>����[��0��/�20�3�C�."�� �t|�,��r�N�!��-��[�-sQL�f�8��1:~ys��?�_��OL2��w�wX�?(N�����d���W��R����A6�Hw��
zɫ*�"[����[Jpm1������ޗ�W����g"�w,�2@��L���׉V�� ��Ke��V����o<�����o�J6���Zr5颚��Aɰ�]��IC cJ�('�p��.�7�}�0��ाJ��%��h:=�C�sA�`�#�ߚ�f�����7~����?�2HFXt��=Ma�9*_S)A�E���,���C$:��%C�^����0!������~ĀrhMȖ���������7x��ڛ��������UEGe�%n@�W�+vE����#�* �G��`�xīo�5݅b$c"4~r�r�W���`�' ��ok1�/^�8\�Y�����J����U4���C�~�9����Hq=<S콈
Rh�@)��v*՛߅�W���K�Aï�\$"���Vp���/O�Xsp�\Ɂ����Q(]C��Ml�/Ѫ=��N�7�ې$|�옹�2��4��{���_V1��_:�'��bRVW���p1��/a7z��D]R:�|s���^a��d��}���о����ո{�iw`88���M#�Fď'��Vd�~��/����y�$b�m{P�W�Q�4�v��kþd>\'.ʰ�
	�w�&ދ��1�-������H�fҙ�Q� �۟!�]���9!�-�0�_"`���X�?O��;�v5�a�=�� 0J�f�6C��)CB�k5�;��8Q~@���DO�h_ڜ~���!+Q
6^=}����	��Qi���,�t��cݲq�GDc��ۉ��I������P$�WKc؊~O�f۠�]���bi��Ђ��sV�g�q����<��Z�z�t�(�[B`���WF���Op$������'x~�JТ�\�n|��b�|f�VN��y�i��.�-��)�Kq-��ح��/D,6Ͱ��Hh]��o㊕.���;�Dl�%,����^�8�m�N�J�����<�S(Dtk��ɢ'���y�^O�`1�����r��XŰxol��#���X�F�=��-o([O�A]�?6�8�۬P�3���̊��<�9����k9�n�1���0����dK��K�k1����=�2���{"g�ϗ�daD7�	ܒ����NjY�*�Q���`�l���J ��f��"(��/�yż+��
[䚞S����p13oF=��V�s-���Z�v�IՃX�V�:��j�e��'����.zJ�E�Y�R�e#�t���,p��ͺdxm�I;�J�,�%t�䡙A��b]� \�Er���	�ǭ�׺VB䁎�N�c�c���E��n��9�w�JѬ��l�R�8Nb���X���"��@D]Y�Y�:�[���B��RFʌu
q�J��V��cc�S�NjTw&T��E��⡦�2��y��烇,B�[��T0��Ug":~GŊ���i��N��Qn5v����v��Ot�WN�����-s�R?��2Q*�"�(�Z�%�af�C���Q�Y��_.C��&���g���n7ԁt톧=ltX�n*th1V�`+x�s5��N�Swgs�)J��r�C���P���,K�e��.�����>���6��#ή�;���3��A������K���p������D�Th�y
\���P�fi=���S��0Uˆ��-y�ۨͰh�6jqMi@C�^d�z�6���y~�����4V��-�����ƪL� |�A!Rۙ�<x��d��@JE�ɴi�Ԇt%�7�1���
@��7��P��/�$����$�F��K
��V'�tM��#~�����<�`�y�wr�4W�%��=�D4�6�H����Zv��BP=Z��|�~,Ӧ��,�Y��� ��{�񭀩���-K�/�~�4� ����&����w�1�-���R*\*�n��u��]8�+�����2K7d�W�x�!Jm���$w+,���w�}S�W�v����)/E�ޚ��'(����c�^��_��UQ�����qڈ��04�ۖ�ޒ4���BB��|L.���wٺ��\�gQѳh���8�H�4�fE�"�5��d��+ܠ$ݎ��%U�������C�-�d��,�QlH!�3� a���Mnr�>�����X8�-����%���!+}a��K}l��ZQ���~|����g)��g�J�s��bf���܋d���.����L�
!�Vу�v�����{���L*�j����3�q�n�O��:槏��b\�)!|�;����N����+�`����ߩ���a	��U������IR��KMEM�4��?*e�p/{P#���m2�=��ƃ��o>\B�m�1�=^����y5L3��V.]D�$�� a��:�[1�$���)�n�����i����p�z&fK;hiw��q$X���-�����i$xiu4X���D���R�U�T���A��n���&�4�,���������S�:pH~���Z��s���DEW��6�ҙoet���Փ�!^���S#a�I��-���J}��q�J��$-C�0��6U�����Y��R�k��������˿��aLM�`�U��u���Ӧ��]9�珺U0��rL�Mdjr�r���qe��8O�b���$�_����mݕ�_E�l���${��1�v�bVB�HY�6���	�Ĵ��2�rb����:,�O�V�Y^!P9��	��1���i�6Z��d����b��;�x�o��[Z:�5�`3v��|�dP-��չ�}���Xo.b5L+���_�'��7�:u5Hu�Κ��z+��a��K���ȱ��|pU��3�I�����U?Z�	�A�Z��c�'V�m�eJ�e	���(�񈆵��7�"�-Z1���Z���(����ee(ɲ/'\Թ7%�d �ԍ������H�g�m��l|�~�]p���ڴ�0��dKD��!xi��9d����,��C�B.KN�Z3(N��a�Q�`��'PtQJ8z^���c���5��g��ڒ�<���!P韛�r����PI�5Qw(l�+�z2��(���U�ݞ��8����� Rـ�_Qi�ǘNS=f\�X�T��'�9̑O�p�/{P���"�u0ێ��u���������y[�Q��'+3F�#��k��}{�J�)"%
M�����;��;�asֹ]�wm�V�t*�m���s����P|A���\KÔ.�O3Y��!?�����΄�H�+h|���~`�Z1�>۠3ק�:54��\.���K�1l�`XN�E�IF﻾it��n�,ny.��%�ǳ�wB(��{B��$95EX� �! �)��ۅ��e%�i�ImS��|�`���.1aS�(���j���1�c��y~�5��J�Yf��M�ƈ�P1���-�\�Ct���Wv0��̕-�p�WG�����������ZG�	r��N���Y3��?'N2Ϡ^+����9ɰs��2����H�}�&�>!�V�gS�]��)wj�jȧ-�/���������9-����1�����8Ǆ�6�@-��G҅�*!e�7�Xh�k�p��.[ͽ-�P-�Ӡ,?3���Z)��HS�M7�-�J��=�*�����ly��0y�JS͵�}�#$�
�fB�Y�G��];̩$��٩�kNŽ������h�@"�d� ˀã��Ј���� �4��>�9ugX�=o�������;�i�{^�Ys�3
{~g�O�m;e(���1Ϯ�A��~�τf9g���3ފۑ�Ͽ�!�����ʕ%͵5� |�g�E3�t6I����!���ԤR�F�C�ImZ�|Q��=Oy�EC�c�t��}�A�[@cv��LgS/9T�HE�Cc�\����~4bkCG�Ns0����Z*k,g@�jC6n�{����#�?�8��z9�p2=[BÒ{�P��5���*`�~y�`Mc��^cH�|j��P��]  ���!	-Њ6;�W{ܠ�q��痕8�f9�cRg@� ��vy'�	��l`o��B�9�T��`���[[@)�b,_���BOΪ��W���%ȕM�#o7�*q=��V��*?���v��d�G��ᬈo��4�<~��J
@���߿��!4��ȷ�!e��2"�l< *���v��U����Gwc���D�)��x�X��湐M���-id���j��ei�:4b�;����7d�(gdR8��2v\�_���F�2����O=~!���!e�ſ�Wn�qB��O8��D�##3i�qI]4R��o4L��C��(*���%���H �a/�]s�x3dn��F'n��K@�؟#2���Z�L�d7������F�1��>�����_��%���ko�W�_� 7�����8U[IRj�	�I*����}�� �n��\	��~��N���)���\f���f��M�lnl�٤�%��>�^��M|�hˈ��ʿE/~��b'r�:,~�O�0�&�[k&�)7�A��Xl�� Hɵ9��[�z* �Y�U����
~T�_��ͻ6(��($��i
Z2��|\��|,|�듣������{%�y{�n�7Vܚa���3�.���v�,p;e��e��<�Q���?���]\p�����1t�a#PQ���٥&)F8l� ��B�~l�`�Й�����8�e���{�P�s��nlE׋.����
J7^�Rw;�\�B�Ӈ�e��P�jUͱ�R�Y��\�ɜ�'�E�c��2A@��b'ME>JQ!�$�k������2����;gO��H�p�H��_6�"!��&Q%-�3�O,��� �L�h<.�גA��V<\�/�t�Fn�k��<3�>�l��w�d�\�������K
<�2q������h�����K��H�8	#��'?��㘸��g��#�2�������,f��ݕ��˧��q_W[Xb��bK��j�GvI���S]�kV��d�:�^�P4�0r�E�{3ܻ����Q�d���7	�b�3}n��m��c=���+��irɠ�����s����͕�Tmp?:E��W��"1���bi�&�Ь;x�X����4z5�c;���*K��|�d���� �Z#2�3�S���S����������x�AT���t.m���gf���M@�"r~E%�!Z�6��J��N�<�a�����v����]�ǲ:�G���A���<��������<#�D�/2Jq#>T��|�;���-Y�ʜ �nj�e�1�L����^�|��{�t~J�K�d\�&>z�C�k�:���r����8�^9h�\yG�Ǥ�V���˨�C�G���;�7��m��3Z�4F���;!kDJl�80�д�ן��W]���G����w!� Wz1�b���'Y��q���Ls�������CS1��r�$O��	%��=F���5�I�͜0)uxW���J�������Ϟj̋��r�f֞�.ieA7������ ��:���)�Q�v�1��7�����]��u��W�����ᣏQI+�9����2�u^��<�%q+0^��g�z	��
g	�-GȖ-x���t���Iy ���;ċ���؎D�()��ZB���Ѱ����׭�6u,�ӾH��@f�_8֮���N
:kB�X�`3�B$��jy��i=���A�i���>�"(�$1��*�y9^fۆ���w��p��l�Ä�DzD7f�o \yT����ύXo'<��n�l_P� JLܭ�^��Ȍ�N&A�ND�X1Q^R7|�7�L6���G=�43�S��T9����I��s��d���唳;`���\1� �r�hzAb�E@،�'�q���h�F��N�J��6~Dn��C�H��}����!>��$�;;� ��\~w`Bh�Ǽ�MҚ&�y������&AR���i��v�b=m7s+��{KIjvb�s>����x��'d�:�>Ƈس�Ǒk��WE2�c��tڟqP6h��0Pj�g������kY�d�7���۸d&V?Z!Ū1�|*��\m	�W����P8�]�۷7��A�	�8yۿ����$����,�����&0ҩ1x-�U��5]�A<�n�_���b���kcқ�<���H҉�����l�N�b�F�{��kr1�8�ͨ�,���oy/� c~$��P�tX��0��2�m�QX�6�h�w�y���<��qN�`|0!�*z�V�,$A���n��	{ն�d(gC�e�� �1�x�j���1|N��� 	��D�K���?J�vD�bx�:�h�I��M����$ua�Q�� E��*�N�A7#ڡG�}�n�i�q�e;�5�Dʅ�����cE6y\-е���1(ZT��?�;��'�8��.��N\ yPY�#�<��Yчm;߇�6+�(���4����j��7��?J��
�h�W��]{I�g��U�ˬ�ROh|s����%�n��a��Bg|_��|�.��s���aϦF�?_�*��3��o|���Լq���V%g�p�U�dF�ZA(M���	��;5wR����M������/���۞�[g҄`xH�g9�:�2�x��_�h� ���� i0�����{L~}��)ʱ<"��)a����g$k��W䤽�Sܬ�&�� p	����2A�����B4���cK����K�׏Ť�w����lcK�7*۵�+�$v�]6��y�0��g7���
R�Y?�����[�<�|���F��[+�؍1�p��~^c1R0��tْ�p�Y��ف�WU�d�!J"� �8FMpQ6���#����iD]Gڋ��쁖!q���9#�}߯9�u���φ��*���Z�dw�i�ק�5� S+U7���d���9��OC��<���C�n�`�@߀ﬔ���7� ���Ѯ}���^E_xQ4U'5�w���(3��-f.`g��cH�,7�mu1��Τ�VMTzLK+Cb���(�V�s��7
E�)�k�t�7��������1���T�f��PV!)�v/A�eCn[�e�{0��1�/b���W�� �{�(�u�l��o�+�,�ƋR��P6����<�G�?7j�wS��$���5�� �g�x��:����L�1ql�l�f$�� �8&?�1(����N'ѕ�z�[�*!Le�Vg���W����|���-�a���N����P�Z90�܄�`��ѴH%�"UPl���8�xٙ���ſ�jM!l�m�.�M$�^���;�� %͵ɹ�Q�Mr&���Љ���`��$ȋO`�U�,�(LWg�֔��$��_ �0F�\���ī���x��p�6���n��&�����g�����^��ax0U
��k���vS)��0�>3�9�ξ�ӱk�$�_*�����SyڱnIT9��I@�p�
J�6
�V>g��F�����#��' �<�/ x*�o�0zn׀	a���u��uى� �=����o���
jwýE `�'�2���F�����E�h<�
I�A��bH	�Q�%��)9���t��ͦt��=��Xx�]����1�x(�z��
B����*̯D���Q�޽O3��U�y�$�����J�Z|����2��4v�8('��2_gJ����K����bC�1V;��Z����Wzg�|#�f���v���$O8Q�����&��𸘢C᪭Vs:��[Q���� ��\�;�o�kA����|y�w�>�:�R2�P��a^w�J�c{DE�1v���^�b�T#&w}ϝ8���r)U߈��#i��V��/�C��q���,+��H�f{c�H}��OA���f՛��1V� �\G��sEJ�8����J���nX3r���Q��@CD���p��Y��&>@*="iG�M��0�<g�
"�V�Ld\�օ��Ξ��28?Rw�i�՘y�*�5�w����(�Kjxד��cMu���0�-f[Ei��f*�yk�Y���[Di���5���Q2���a�r��Q�m��O`7�Q���&n�A�7�͊��ɥzj�{ǂ�>`}L)�5���I���q�b�uMAGM�����T���''D� ���,B��G��D�����{H�K�/�|]R��%q�4>�qM�a�r���8����]㣂�;�1/��k ��*�q����'&��`b�@�nC_�i9
�p��j�/�ӌُ��y��Aʯm�XkF��>0/�	0�JǤC��P:��k6�����гȔ��w908�:Nmٖ.�|^���S$������T���ЊGJ�q�^���E��J=.ZN&|�J�OP0v1�p�=d�)��Y�'ߥ)B�v�����h���1bi�C��㷓clM��F � �YcMn�I"�
~��?Π?�����"�	��I��_�A�iM�Ӈ3�c�8�����;�e|�Z�C�y��߸T���4�;�ܢ��jdi�ZƤT��g��K�m�ݗn]��Z�Mв��)B�d6���bUR싍o�j���$S��
��D&�擅��(�o
�^��d���5�$��Yq�E��o'A8��{u�@}���<�;�6*��{��19%} �'��+J�ﭺ���B�3-��Yb�J�Q�mD��� � `7���ɐ�JW�W�ņD��?R���,�DTӴn��BY�Y؃�q�j�;20��)oM�4������"Uqd,�go=�
���6(@~+y(ș�@��P�`�8�^��8W;YM�Z�N�Հ8@�0b�Q�Yx	f�2@.3C(�u�8�N.������Gr�#�-[yy�!������pu�!��/��T��>7����U`��ԏ�>��gǁ����Q��ԅ?SZ���&�`&�Ñz�T�p�e&�����)�����n���O�=-�ؽ�Mc���.�e��JHw~�s������R�b���w޻4.%u�#���p>Uj�I�2EAq7p�n���)	^����I��L6�.�/���B.OŶ/���#��k�%�4Fs<Su��4��r1&\�js�%�Rip�ek��t(~鹔q���}�m�
"������>\�S���e%V��M�kyg�Tu?n��WH�g�+r|�8�@����~�ƻC(������M��\��n�/�a׸=@$�e�	98V�1���h<Q����Ȱ.��|��5Z%�C���H&R���X▍�f�%��H�?����-3�R��k����S������߄����I��/0|�єS�/������2x�(�ٵˈ�`L�]
M!9�zp�R4R��o�FTk8}���Tp�:![ږ��ȅ/�?�F�{oi�)y�{&w"su��sYC��p�e�M��;�V�knP���>�FT��S!�jq�N�PD�&Y�f�iY�P<9:2�yg`r(��&����'�Gw<�5^c1�+*0ʧ��=�� �Ŋ��������ח7C��D�1�$���`�|���U��Π S�Y�#��a��Q:s��9M	Ӹ��L��?�=Qus�D�Ri#y�<��I>x-�4� ��.X�@S�h[N��0z9��G�kA���J�s���U��7���z��Gs���0&�*�Q�,y�\t|?_�8�q��F`�6����/gA�V8�����{�v�&�ZS g֨�݌,�����kT�����`޵c��3�]=���Q��s���_#���nI[P9Ӧ����^(�����AuX�e�����!���&��d��uY,�:�5YYsxM�Ml
�Ҋ�:lO��-�M��m7�.n���� pZ%Ω�X��L͛,����G���zߔe����?o�*o�^=E� b����G��Qd]��6	�T��Α��r4�ڔ[y��ϓ��\^�ak���YY�
/D��wt�Bx+_����3J9v�Wo{��zU{Ͳ��#,����`���^�������AWI���z�k./�e���H#~+`\��6�殖<բ�0���?N�9d���J�ə�b��Ώõ��>�`���lX"�X�0��.�jOQ����}xz�fY��	��K�NjuW\�D�%؊'5�?[C������(<J��E�� /AEc�&IO�_#=�0I�6��"�؁�z��/���ؐ��%��<�ե��E���̵�}]'SF���m<�&kn�b��ݢ�^�0�'�=�	^��5\j��t�~�Yo䭓J雸	�c�Z���e����#Қ�j3�MY�P����K-����a4�)�y-�E�Q�!i���&R������QٕN.nd/�?�ŘG����),�s3O�n�a(C���ֹ9J�B�t������)�v����oo�6I;ob�<Vl�Y��W;)UX>���y5��{c�W���lx��?(��o�J�62溰Ɠ��	��>Z���U��^������R��c=:�e�C���)�J��\QÞ�'Ū'������rsUG�{��O�X�f�_ު\Z�|(t>}�QV� 6/ݺx�"���Y�	>S�R�}O�6��9�c�b0��ht��ǯtVx���~/����)VrP	a�W��{8����Өw8��3��0��%F���Y���tA��}�9�i��T�np�1�����@]i>e(Ĺ�GT����;<Q𯔵a�#(|������'�W���_�����o���BQ�,�y�7�n@�QZ�/Zx�)���&RT>}I�g	F�Sr�u�A��)c[=��v<u���T�W4y��~Ҹ���S�;��]Mf��$��̖�osF������N/E�è�t��NU�� �����(�����$mZ��Ɵ����B��:J��	*HW[.uқ^C�>F/�XTgT�ʌ4��z�Y�sӓ
��}��*���J�������a�e��k�UvH�D爆[�7�G�!A�%��B�Ԡ�g�(���m֐�ƨxs�L�n��d����#�`v�0���"���w�����>�R0A�׷�0 eAzq:���H55K�ب�0Bxŝ���/' M�L�3�6��a5�����
o3G6��߆��U)�ѿ�rI�|H[V ��Ė���Q׽�%�~R���A{O�NGY���Ml����fg8Y<xi&#ކ�;D����E'`������G�;CA,"$��Dm���-�l�rc*����i��5^�e `���t���o�)��k��W=�w\!�ݶ�i��a A�����T	�s�dM�NafHU�XXT��o���MZzXW�-j�S��WvA��\[����m�5]�B��ci<�����i�	j�a��^�m\��V�1w�kB:'b÷n�懋�޷>�S�zI��N�Ew�Un�~Bߗ�e!�D��
���!̯&:;��yy3���3�'&S��E(]�8=t&l����[�`,>���l�&���'8���f[3�_�x�%7��H���)_����ï��<B�����Q��<'e1� R��JY��£H��o)���F�t�+��G���A��Sܚt���܌�i?�<�m� �>�-G�zހ��\�-	#�?��
)8K���j"H`��R�B"|3u������-`jQ>�/C-۬�O�8�॰�&�I`&8Z�k��>�
�m����j}��|�N���!�+�D��@֧�������ͽY��[>!�]ץ�2�����g��u���dp�!H����^^+����ꘅ�74��Z/�@��D����ϗ�k1�&R�=��V�ੴ�N~ߜ���w���%K]��5~jk����8��i>�]�L��bM,�{Nã"g:�48:�17jN1h�2���U~���(�ȷ�̹�	�7Rj�W�v��pJ����=.�7�.�dD��%�����f�+�>���	6de����I �����Ĵ�x���*�}��LU%u��E6��&��iВI��k֒�"^�))Wdr�|�5]��kWͽ��nT��^�,�Q��
I>��\l�;��ʢy
�覍�ŝXU���!�K%,s������W�yv�uț��L�.f�HVr[ɉ�ň*��L����`��&��b�n�m\J�f�M
5{�NIk�����XO.�F��i�.µ9NC�u��R
�*���D�L-�Z�\�`��I�t�U�\	�����{�/�@b�mk�\q��c9�{*�$��Ώ�$!�Y2���&
ȱ�<�� [�#6�5L��
�6�o>�6�ɋ��!j�܈�l�j��x���&�{��vo�������	T��H�I)�)��XE�#�=r�.��p�my�Ő�NQ�T-U�Ǔn��6��^()�;爸ɮRQr�/,����6��7�l+�Ф����@�Au޽8p���Oj%����!c��@���nzd��93Y�'���^�*�F�)o�r�Uz�q�W���k��/��lj\���7�B�#��x�MY��@sd�Q��:�P�H�G�Q���D�Y���� +��tgphN?�9Gx�h�y��nr��ߤ�A,� �8�/��Y����i�T@��ԅ4�!P6��#�)��4|$�@H�|5��|-�6S�0(Z�ֳ�kWR6��}��g��-Ue�P�C���6���!C�����>�bf$2I�n��?S���/
��G|��'�������d��mV,���X'�bNG|��df墶�����x0^K	盵 �oA�`pD�sR� ���8VuA��y���K�U�k9��,�����C^�_�6!9eث_�h�������\�`<�٬%ʰ��U��`�t��4��+~���f���_)�rUY�b�A��w��.7d���}�y�l!��/𔟳�U-�.���`�ĹKA�ޮ����I�n6�@�յM�}��2����Q!��:�.�w��A����w��*I����R����oZ$��e�o�#���=7��^{��t�:>����p�$������h24�9�J-y��qty�7��?J_d� �c@\ސ`)����3+a]�����i�~�給ɕk�(�k��*L�*�]����e�r���~�\8�\)h�Gn�\8|RU�5T��Lw�gCd�&�I��� �����e%�?�|����F�͂\j�^��'إ4e���"���o@z��2m��|�M�6{�fۉG�[Rd���
�wō��쭋��/���Huì^��LL�V.Sh hRP�%�}!�&C�ôyya訏{��9�-wg�dϮ��������X���9'儼�O�2'd]{�@hlz�k�0ʈ3}v���+�$r>aa<0W��~JTWB��d��r��L�)����$J��k�O�',3$����}Av:`;Y�G����Ei����f��0Wߙ�e����	�ڌR�LoR���m[+V:��x�5Ξ�)��&<K.5��A�K=�}�r�'%#��A�4�I�n��l.ge��w3��L7Ψ�-�D����±K�ё�j|?��|�8��XL��̄�;{����)��ע�?g�Q2�t`�1|Q���Ο�sOI#���Mr��]��Ǻ���W+ϚYړ��K>�q�=M:�{-�	��v��Lru{:;��UG�~���
X�k�<_zX@�N�kY�� O�5�`��C�<4���h���J��g��\+�[
�s^�36/�\'� ;r�����Y�
��d;�r�����]㞇ua?l�g�D�kV[��Z����s�V�č�릕
t�]5L![�D��y�~(����*�[*�7E����u�B���p�Ok�m�a�制�h(r�xt,�u�1����6�����\��7Dвt��zj�$Ws�GS��$�D�J��W,�%G��%�VK�q�|�SL*v T��
L��
�t�_�v?T<��}��n�^%w��|�w�����ȅ��su���}8 2�� ���Q�4��P^^'nc7j�Y��[̣	���� d�M�S���ǂ��K��[��Se�����q1mRF����v���		-)��2A���[\S�O��EW�ѯ#�(+x�����[º?�m��VÇ��J4P�p�r�t/�쮲Ȟ;?�h��61���j�P�ٲt�\�P��
X];�n},(^���k@������󧴖XB��d����(��+-!��yQ�A��?@H<��b��J.6�߾��q�����2u���򋃽����O"j5zj�J���*�6�!Gq����,K#V*�"��Ӗ����y�"S�f��p���su��N��-�y4\�1�Q3(`$E�gOή#a`ል��3/:�\Xwu��L��3�E�^BM��:ީ0k�,<S�U��+b���<�T���L����%�!aE7�z�~r�&��wk��!vt+�U�C7��ۄ��̽pwa=�m	��ܰ�~��r _ �c��qF����S�ح������H����_�'�x�1\�	��p��W�q���5.�u>'!�^��� 6?M���q�Or[������	m���e8�#ځ�	�~*.q���wM��~e+�i�;����N(���uci]�qq��-�ӽ
7��̦�H�,!$�3w��S�1>����;C!��"�h+b{��Eo�	��ków<�F����6�+��a���D@T�!�.,�.m�P�����g�%�,��<��>AD�I�VaK0�$|�CN࿳�@¸GlK�G��3Br�� J�վA����5�����׾�7�cd6��jwj����"��{�
�<6=4�89�E�����h�;�'u�6^��х�m�x�k&)��� F�{�g�x����rEmC_q�^Q��)v}3I�.��M�˗}YR��B���l������h&�	Ѷ�I2�`R�6������\sHC��+n�f��ß!�"���Ֆl���@���AN��+KS��U2{��Q1`vWX"=����:W��u�b�����R��6$L�����YM�{����Y��9W��*�@�&��=&,�P�97vF�g��ǟ���6;�,~]��;Ѹ �SY�[:��w��e���#�-�����I�:�0*ֿ�/�4�R�~<PÞ��sS�� ߿v�U?��p�H��&V�	O�qiԄ�¾�o ׵$�o˖��u�0��@������3r����y��+[�	W��d���4c�/�0��J6�^ͧ����݂T��0�����S���)�1�S-�U�҄Y	�5����A{�G�~͕��+ME�ۡ!G:xXD�Yvq��,��us���W����&`�7�
���^ߌ�,��8��*�r=�ƧT��,[��\y�
ug}FT��r�ā�*%�w` p���=�"k���t��wp������,���Oz逝y�ar�M/#�=coe;��	|\q\$�3�^��L��݄�/(}8��2!���R��ʎ�v��$�rHo���g����>�����c���G�n��r3�ɘ�ϰ�>lIF�>[R�$̻}<��j'�t�2Nef��Ƃ9�(�.J����i����I�(�F"@� ЁΘ�J�g�$aM���x��ć<�:t�R���'�=x�$66� ��Q�R���}J��w���M��c�7N�=�\E���1Z�Uǒ�Q�,��>�\�3�hK̩�YD�� ��g9A�!���E�dT�y���ۿ`<m+��`���d,�O1�"p�Ɏ)���pn}��g����l0r]=��ɠ2]��ҥ@,,~�T"#�Aq#`c!������p(o�� f�k}�+:<,���������q�ǡrP��i+$�0!��*%��I���+��K�5s
W6n�3�ū����a9�.��
�J�O�&���V���bE�~��B�0�M��닲�1uC+��LN�v��l"�V�O=��_�}+�ñ�9���M���ZUn� ���Bs�
	��;4]�4u�t�-��bNaS�ǈ���S3��zEtf~F��}5�k���Ͱ�Q�O�ƭ�X�F3c�s�X��!Ѐ?.�*]#&W-�4�{*𤛣T��4�91R^�5z��Q`���z��)g"�tZ	|�}�k�.�����5ji���:��I�oҗ	&��d��)�՘��޸�U��1=���@G��Z=2���s?�C�K��;����Ye���M������=z�� �*#�Kj6�h�`%_W��2[(>0m��j��Gsb2�@�Ft�s�d,-b�.5݅�ER��{ ɾ�ܡ��A��!'.�:����Aϟy6��O��NM���3r�
��wGn$A�M7)�g�i�&Hf��/wXQܾ���0�v9�.�m��A諾Y/s�L趕����{����4ubND"2�Β��"�����yjԝyZk��'���bP�"��
t����4ϴu�{�?�T85w�G�l�2ڄxC5�ݗЌ�� �x�I�A9i��8��1L-�
{�]2��K�j�����RN:� VM�6�6�����A4��+�^j�j��0g�(X������_�k�'u�W���F�m�LMH�����.�V71$�E���?���,�ވZ�\e�T�d�o��f�T�dj �jh�R�c?=Y����*� <> ^Od��h������&*���-ĸ��<B�e�0YJ��-��ަӻd�)"W����a��yC�� J�'L(%vݎ�n��oO_�S�T����X�t���b��BǢ�����~ƻ��@`j�������ցj��N�лq��V���Rg�H����uV��gO$����DH1,��OM�d-�\�XA�\XE��V2�f�$㧾k"1�%Fcu���a�e��}2�a+�9��e�Nk�4�����O2=x�ἄU�2�3z^-���tA�UʳZ����%p� �W�/�7��`2aOa*N���� �ۨ���k�i�MnA��Nx"ҖIi��1 ��~�#��I�r����8X2՞L���ܽH����TcVD��-9٠&�������ڹy��4g�F�?B���ּ�=W&�ו�E��>�i��2u�g{/�3��rU,����Յa9�*�Z��	�1�]���57���2�Iq�ۖ�[���E5�q��Pt`���j�Q��d��/�^o�DH��\�0^���Y����Z�|�wQ�	��ҵ�O_$34ƥ��6��0.�̾i��$ ��@q�JJ��#�+ <!@��u�R]ĸ���
�x��z���]��%J��>�ȧ+�h>�1��x���p���mt�_c�w�k�6�W�������3Ě��q3�$̓TX��D���[3t˧s�;����N�
6�:���JH�����ӎ^d�?�OZ���WB��̌A�U�܅N@h�mK���Es����-�������d��I��d�#�g4���m	��G��9�=���<��D:�	Dz��I����x�(�����^iN���[�����x���
flX��)�;]��!jsm�Ϡ�á����ek����sG��07zw���ʾL^S�v�t����|m�2x�C�Z�Bz��G8���fX塽�tWrjt�dB7�v�e�q5tӻ��eqa�֬H�/�\�N	��?�X�b�^f�E�c�%���xXs$~-<9f�1�A�B���'uU]!�pk �,�BX
�����	]R_�-�d,�dĮ���['�k���Cď�5����p��,�	�㥏���~��$`(-��?Tv 0�`��/M2��a��|x����[�j�E	� W%���������O��*d~
Di�K-�ܹ��
�} /i$��m����T�W2�:�#����k�m#sѧh
�U##�}ޭq��1��T�����Ntu3��K�!a�P�0�1��3��m�.6>k�5{={Tj�\��)86��/�mوI'J��x�?�T��Mt;�r�m�Vj��k!�V���=�C��V]!�f��𘨐�X[ɫ�yF��c%>�jӑ�����+
�ŝ������+ijlt�����W	2���,�UM��	T��iCŻ׬����lx��?�����M����Q�N'4_�h�ɆawwO�Z<%s]�q^I�&�U���#$�3ƛ����+���N���?���>�6����B����W�<|5R�~1yw�XsFP�3�	?��Y�"�L)T�
6��ER>�D�w����+�-.�n��К�jD�4��h���I�,L�v�%�}��I�J�,c��L�-i�䟱��0��+o#	��4:�� ;�/�@�F�� �aR�HN��y��=J+]�2i.�Zs�ak��w��vk1�*d�n6�t�{�j��Np�M��|�b�l���){���,�`r�j�t$�gu��Զq�]����K>����0K^k��vр���e� Ά�ߋ� :�g	C����oIλ�/�D��F#���h�^�;��N��3Wъ���DN5 �W�ٌ�'S�^�7D�E�\���Fs~�tt��H%96n��CK�n"?6��ҁd�C����籥2e�VM*$;�w�y�������5x�	S%*��Rr���rO&.���������K�]=T4C�&9GI�l٠��+�>o���>�<h�őJ��&E�g@D���&i�\O��jj\	&��V�	�%����O�y��$��zM��)n�o����{!��)��D}��� ��Bs_P��.2p9l*r��i+��7y������"���?ͤx��V�n�����]s[s�:�	e��r�K�� }�E���@.�b}	�~$�>�/�*f�B���/ͣ~"R2TA��?l�j���O��U��f�G2%"	�F�|�JhFP��e����Ba=9>�_ :�Z;FpPͻ�ż]Z�[��������67������hEe-����a�d~oxq��B"���)B�b��	L�Z��H`��-�x�EwFa'69h}K���XiV�;҄M>*9#��I�2���ɘ�H��~=�s��_!Q�{~���iV�w��Y�V�̪���{3	t/����6V�hG�N��J�����>���u�&��ƈ/�����*���<���d�8C��+�������յ�&���\�A�1�ӭ�
a��SN'���_���o�8|��b�E�1/%^���Q�ON�E��F��m�G�A��8�"�"
S��V��#+�����R���a�=7ټ�e�	'ѐk��%��Rh�҄�dH��u��2M�(�$"K�=3�m���d�����{�֥�Ũ ���>��<�bNH��-��;������1�۸�v�&�X'�TPHf�������_阼��-�ĳ��a�A��Ã�:���$Fa;�]ɣ�+T>J'�u������þ-�l��+��u�ڍ�ᣝ�`�S���+<�y�qWc�g1���Z�����ݥ[o�رA"���XB�On'�⨧����s�a9'I��o�k#\yL�l���7����[~9`�u]>y��ܚ�	jΔN�Jj0� ��%�3�FqZK��ӿiI��G1��O��sn������(���B>7�;�^���Ix��s}�Q�#5iEz��Ԯ�7S�@��r�r�߈���Z0 ����kBp��X�� �V�E�V��\m����خ�������C#�p#�X�%���Я�ėn���^��!�d���!�x(8��+�A[=��f��ͳ���`�y�؅59w�Н����,&��(����� 
��D�üb||<�-�DU�ӿ�T�4���@B�m;T�h#�Q����>-���t�G�i�6�â�Mi����u���\�k��s����9�J�Yx���E:S ��<�Ut�l`W�j-���7���xlr�^�ρ�1��Ӣ�:��땇� ����`Q�5��!G�m���n�~��Y0J
���hv��9�D�QQ�fQ ��z@�:ۆ�]��H<�u�r�A^�"\�/��C)���sumF�%dXي�1�[_:\�j��1�@5ߴ"��W;@�Ԃ�X���� ��g�1��fb.�E�E:�_��0Ց\��@	�b���%"�=oBR�*x�\��`h�?�}=��ޅ�H�/q��X&Jg��������묥�?N�n5�����Ũ���� ѫu�k�0�š1��G	��S~V&��ʽ(w���?�	=6�b W����-�����7�Z~5��`����LI�p>��2@���8}�7��.(~S����3���QR�X��p�����^�]����ۮ^Mo}2;�Q�ܘB��Vx���v�t�O ��ˠ���w�֟�����	���	}1�f�e��!iK��pVL�S��!F�,&W')�.i(Jm�
q>E�1�� ��T)�scf�:A @���W�'�4?BbV�'��w�$7첂U�y{	i�����r���`
Vm�q�6��ʘ���/�����|"��^M?�bE���Z���D��t�����`pf���\ ��e !����>��e�2�H�dx.������A�N�
��g��g���o����2�5�+���K��L4J�d'��%F�D(��b7�p��m�:kt$^�������*�肈k�N:�D�E��76�l��>���gD�(
�Q��������Y�W��(���}�M�7|�$�|∑PB=�Jv�r�֖Қ�=c���!t����V a0u���xܓ��F�הR�KS��_���׼���~���<[��'��C��D#䞴3�!g�hЭa���E��Q]V�x6Z!\_W7x@��H�������>4�]'�rw�/��R.�ȕ2������^��:<�Y�ڐ�Hl��b�"�F~��O�D��޿)�FT�HF��sy�l�M����1��\�(6� �f0�I{�8 �$k?5�VN�n�z� "�bh�H�p��2�B��07�qԢ�r��w��k����n���̿;��t	_��`�˞����;�2"o�+� }n�H���+�3/;L�|�q}Sa�"z���!�~����DǤ5�N�n_]G����pڡ�V(�g��pl>��"�'�R=%�_�
�[�q!�#����R�j�1��,i%�&۴�a0n� �1��Fѕ֙v���5��>A,sJ�S�
�%A5( �/��<����W��BO��,}J��A5�{2�8[�
�\ X��L�9�}�Dt�\r�W�&�mȼ�6�\���Qf,	���>z���yFVL/�z�7������H�nUS��t�8
��@�J��uC�U�6��{q
,���_O
G���� A���3�S�9A�ҵi�$�3L
��睟�F�P{���̬ϻ�7n��Bo�ꚃg�F	�ַ�%f>VS�?e�s�r}� �Q�̡'IF�ò�\Nlz~�))@,X��ŧ�GRq�����(�)�b�=���Y1����e�}�5��t_��χ�~�1�Jz�_٨�����'v���>��������9I�_1�2?+�K��"��ͮpoo��@W����#�<}!i.��q�Ϗ��g��}����z�=��IiC����j����D��3=��>���H�K�%D4N���=ZIM\k�� Va�̚�p��]����^��@� ��Mo  z�f�uu��|�Lq=�����`bZ�C6H��=�v�a}]��1 �g�������	���뗶*<�%�]yW�9(�⡜{�k�U�J���Ųn���&N�-y��n��#� [��7{�M�bs����}��H��e��ta�H��\�\�jܬC��X�ق���Y�i,O�^&O�)?�4l[(���v4�ҩ����	��;���2������{R�)��_M2Q|A�l��z��WŦh���I�-��i�kԱE�Z��,`�0����64x}�P�?ܒ{*Yb����&���ꌝ¬��l�!�(�Aa�v�n����4ͫ�a��&��y2���9���2��C>2����(p�ua�NelXi��~���W.c��D�A ��x�6��[(�~�t���C~? /�BjH�YM����}]����?Tһ~>��M�x?�b�j�Ti�R���N{�Ֆ��5�gI��?�r��2�%�͇|�=�?XW�
�7U>sG"�Cu��-J��
Y�e���@�ȝ8�7�"�M��%q񶒢�D�g$�`p^˹\�<��|�;�)N[i�N�k����vo<��%^��c�A	p0XV#>Ĩ���оz/�T�[���2�ilTӴ	�|�*:暧�zG!���Ԙ�ܫm2��
%�R���S�Ens�i#okt:�6:��D[�R�k�[�QyZeΛ\x+�����I,p��k;�-[W�JY^S.�{9ʸ"N,��/�&V�'�vv��VP����2hc�o�?cN�1�]V.)����\ڮ2>��ύ�����[oaali�Ȼ���ܢ\�j��<.�M<�W��Ӽ$�i$�6�娤{�޾�1Mxs�J U��B��K�~��⥏��׃�bZPaj[?~ɻ���K�$���+��-2�I?c�6��(�G4qv��&M�mt6Ɲ��Y�mt��8�#�3T��1�Z��k%t�c'GЉ�+L�q3zV�j�xu�<��Ev*X�!#yzUS��GI�籽n�}�Y�N��̹�G��zE�
���+�e
P�Y�غ��R�ST;�b��ELU�"�J�v����!7ߖ�~��P�^��s���V���4�'�	���p�
�A��#�m�{��\�p_��*"� z����9����+�s<6�T�[������
���v]��͗W,�ꢳD�Wu���dK��9h���\ъ+��~Y��̸K�ɖ�<�������G�u�$�t�Ⱥ�j�U���o*�P�O�}OP �a��E��N�"�6>�������� �iz<"�^�=6���_��s�P�6zQ��0��,o.8KA[c�����6�E�#h��s�7	�IE���t���1�n��:��H��.�æF���se��;�fiR��5y�����_
�>\�]��S�~h���/�g�	�<�ᚧ�S[5�g>I������Ȃ���b"a#-k�u���)C!
���N�� ���e�XTz���KuN��L���Һ�`h�`�sy�_�t�M�Ү	�``2��`��*}h���D����<��R�~ۂA�P�$�g#*g-S�����[& [�}�S08N��YƑ���Zb5��h��*Y[6�3�oP��X@��+K>���S� ��,����Cs�f��@�4Fo7�Wˀ$Q�sfۧ'�l��{?�p9��#�SޤZ|�P��/�{�0�M�X�*�Xx�a8�D$�u��%�)�E[7CS�]
@�S�܁�EgA��_L��8����|/~���w�8�Dc�tZ>=8��~ �(t*M})�S0�
�J���n�����f�u��N���?��3�VEM�²,�_*W�u��]&��(����js�e���L]������w�>Sۺy����W��b�]���W��&ѲF(q���4,G��dD��(3�[�p�A@���w��:ױ�1�a�N0�>�[u�~��l�΅��Y\{��xQc4<G��襊tj�lBk�	4݁'��TMq��_���;��<*)�,ޗ^���)��Y�h��wqW�������~��Ĥ�-f�zw;����TA F�	����̒��a�FR�zc���:n�2HG�ec`I��v��B�����E0����N�	�:�Qۅ��IP,�J]!�o����ppVb4C�w�/�d8nX`xw��H.$>������p�m$�"�t��6�r�7'�v(�6��_���ܨ }�5韹��yu�*�)�L��"!��B�(NO��73�d��f�ĭי�����4��^9V�I0�ZA���#�1e���P[�Q?�� �n���	��%�n��B��/�e�F�<8G�Iȑ��
�eL�Zs��Kα׼��ZH�pE�i�S�.: �� �`v59�s���v�&��/�<�.�|��L�����Q5�:�~x�!5N�3P�������:79p_���]�I��
#�|���0rxtԨ���z���j��1�&��ˣ��aƯm�G}���l��wM�W~@�N<�wa[|��^�k�����~?���n���E^�u��R��x�؊�.����#��$ ��L��퓜�/_H�Ft*���Y�>������6g���	���"��|���f��ʲG)��i�ZI�م��u�����b�7rO����k��.&�f���m��y:(�E�D��%EK����$zs��S�0)��N���iV�>7ַ�[�F5'5�����
k�E��0?����^�����H�xK��oZD�@�L���0\���k\i�D����6��Hh��:�"�j�(�^[��-��yq�Y�]�B�Nfc����»��^8X�V�9�\Gw�+�CzM[We��	�+�*q)
#����4��kT��@(�\����mА� S_�a�I:��}0�Y�8d�F��x��<�q��Oi~D�XdnT�Xm��l<�r��e�ٖuO`��&`�?�W�5�F�6������X:v���iR��^,�`@g�&����_L�P����SU��<5U���	;�H6��᣶~�C��O�s`g���)����#�{��b�rz��54m~BRʚ�����ӷ~�|��=at�p�i�@q�#n�]so�wl� �_�*(��!��ȟݺqhiڳ9�4닯��
�~�"�]���z���s$`5f�O#��.uEH��'b�2I\��e�5q2��r3N� V%�N�gԯ�� �������������ъ�m5~�	�]'�1N�m\�2L��������݉�C�\'�6�� `ϑ�h�#;�Q�"MMK�O2�*�g�m_�Kz�����T*@2���UC��G���T �X^/.��sj�9r[�?�6�~�q�A54V��g5ҡ=/`��l�+���_UC�vaj�[79�'�/Q)b�It��T,n(^��pO�:�i�͙�m�
�QE����_���kA[[�L&\�d/�P��oqf>��GZh�K�"Ԩ�!��&�)��.t�2AAY!Q�º��o�E���<^�ᑻ�K���>Z��D��AE7^��f8\�Ҝ@]#���qD�b6�&+Hv���+��Mp1���� ������l�P�#�Lyx3���v�,r\�Π����[%��{�,��vr֤���ɁZ!�kXA]���#�p2;��,bS��Ώ����Z�O�@Ƶ��l0�$�7}pD�n~�;:�+~b�O�j���gմxv� \<���=?� �l�U3#g�#sh�ަӻ�y��[Z��A��ݿ�I�r$�?��Q1�C��ܮ�/Q�I��C�h��E�)��<X�K�����p��$;�q����X̐i����_z"��ǭa�#�+ڸ
�M.~�O�!I�E��.^ٰ~�� |O,�D��5�_�Z�3l�$Dn�dp�\S��[�z����]]�� ���������y�ybgKQEi��^Z_���h;ȗZ�n:4T_���9���T�h*���jFq��R�g���xE�1������̦/pc�g��v���,�"�ԏ�j�~q@%�(��-$`$�\?,�-m[�=�P�Z�6��(g�C=��>6���(����{7��]N��w�ah`	�ҰТ����Z�1� ��lݻ�8��N���@��Uײ��'�D�ImZ�4�!����c�X������t��<S�
�^9�d�`b�e�}�Y�v#�Xpą8fHݡ7n��(�[�95[�szU}�����Ș��}P����Z����B��c8Sh�]�Q�vow����S1��7*i2+č��:�~o��[zjU�Y5�nQU�K8�ƚ]jt �)(8�ŀ�kX�(�qe�si��-�cV"B��
�
��kN�aJ}Bq\xZ�ػ�G~��6��S���*��e�e=���U�:�Db+��J��$�����&%��u3�.�dv.��]!� �_6�f�S@Cu���y{�����cS��\�g��d��O�T�޷��2��f-��&�l�q�5��ݭ��%�33�`!�wF!��HM�k�Cळ���e�A��	W��!�}�o$�P	��E��D��^��r�A�/J�ݶ�)�[:ݙ45"��GƴM��d��:~X��	g��%�B�OF��0
�n
oN�xL'yK
��RDf3�+�4��!D��ڎx�K����$���m���؅s�,�B sn�rc��CX�*��=��Y#H\�V+O�eVM=����1��8M�2TW��PF������[Ɍ�`��|�kR��!�3�YCݩW��p�>�Q$C��
�5yĒ��;]�4E��;��-�X��8˪�C#�(��L��]h�:)fB��P`�vO���^��T�¾����~U�ְ���D���o��U�ț��V	�ݡ�13�D�L�n����%Co��[����٦�L��h�]��-���ˏ9�M�&���=Db��8���l����q��g��1�tyf��:�c���gW�<�Aɒ��Zofm�'g(�H���܃�~"�F�w��7À�clYm�|1̩Wdn_ ������q*�z�k8���%ְ��ax��ڠ�3�)2�t�K�z=��`�����9���GO7�'n�`��^,���^oяq��^��)&T�H�]�N����
|�7P,P�ѳ���Zo�eȓjX';���t�4�- �^$绊��'*8�Ϣ�y�2��G�'�S��¥�_�w,��z�pX��u���qW`3�C ��'Y0��š,4��C�I������w�}���c�^����ܠM��8��i��c������S�LM�l���1�[ݓ���&:�>�!yL	h*O�� `�ЗQZ��l\V&���q�>C���|��<B���E׾BB"��|G�ys�c��j c7 +W: OCO��2Բ��9�����̀D�/c��1�vs��	EǗ�t���,�u��2�XEf�0A�rtB\<�"Kq�ާ< \;@�޲Q:�L�Y�V�,�b����qu�~�h1}N���M���*��[|~�xJT<�@��sS,�m���G"V+�W��ڀ�N��4o�+�TΕ��i��?�9�D��á�L��R����̇_����8ݑ5%�X��O�)���|]dN�u �O���<O�ϐ��mׅ�ٚ&��]d�����
�ܚ[3��4RH���Í�ӤB��=��v�	� �.%�q�{�%>�P�e�3.cAs����U�S~� �+�ϛBu�(��Ҏ���]�~��Li]��!\���ž�t5�f��q���߳�c��4���B�ݴ����6O� ؇"��#��Ч���A��Iq�������Eg1���!���{%�����Ш�)
�YW�eM�%d�[fs��d�A�2�AP�/q"9��u�.���q�v8L�/�s���q΋mD�B���k���>��]����������g�}#>Q�F7�O%�Q!|�&]Ue�1�/��u���{4�1/g���h<6Ζ1��  䭾]��o���j�\�T�S�}m����3p�2-��$��x���	ƜӿK	�I�o��іx�l���z��9Q�t2����/X<�3��4�9�o�>T��/�V��P�Zwo�8��&�^w C���|P���ݥΞ{B�*EG2K'g9�z�nƔ��kxN%c��)Ѥ�3�v���P	�*��	U�
| �$$���U.�	0���pBT��Y�!K�Hd��)��I�ؘ J�/(<nP�Ö~��K^�E�NB��N��Dw��>:�Yʞ�q����
���G����8װ7�Ի��=��ǳ~�^���G����`�_�%nő�[��ӵ|��b19Z�> �xGWWLG�qP�bZ�&��{�V�E&�	������8!ﱦn�R�����<e̘�S1�. ��D���v�:Zc�����e���5�AqMw�g���n�ٲ;`�cP3��E�_�P���7-ӭB�_4d];�swp�I�[?����!�s�y�!��ҏƵQ��8܇n?c�`�R�`�e�Ѿj�\�g>���A�C��]lt)/�HE��lV�7v�`4�o�և�.����~�Af��wy��� �3\����x�E߃�BDN(I�^��S����} ���8笷X�D����'�>7}�
	�����cP��Uc:4�\
�_Kqp�$�R	��i5D�'$A����\���lGjK��4q�x�\O9ϫj��H�� �|������ '�Z�mտ5%J��?,�8s�����+��
$���A�|l�\�=x���,+�+����a��5�#�G�A��P	�B��iV��3�!:{��v+�V\js�����jOwE�'.�ֽ�݆��N��ۡ�\���M����xԈ���n�H���ֈ��,�[�B����C�:b��]Xv��l,�;A��1��P�=�>p�h�6�7��8}-���`��s%Y�?�`z&� c���k�3*�j�b���p)+��tx��7|.I�:!2mG�'1C�X
>_[{r{9�T��瀷��A�����5O��$��x�c���~��(\�?�C0��J4e���R�>�>ȭ�5��6�'�h�y����z��lrP��,���,�
�yHn�)��?��'��Z��jlP�-чv��C�"W�蛛>��d_�#f���:���W4l����@���|h\�*�:�d���TO�TPT9���q�2z��x�	o)�j^� \�$wԠw�Ǎ���+�>ӿq_�/iZ��Lu�"Sw����]������1��l8��/�Y�?�ɪ�6�j��G�C}JB�ܠ6Liw:��P�F�K3O޲p��=�ݓ�'I�:uj�dLs䒥|�V
�T4�_MU���¼�"��(�|�FXJ˶�<m�Kũ\ǣ���9�����h���Q���	�}3�A�
V�Te�J�"���[��1���hL!������6��gX|�����U��-�%H�&��0�Ny�-��r������"�l�@%gNf�����ٹ�vP/�\Fz���/�h-}��f#"�Pd��hw�
����z����Qs�0Za���h ���w�Y�r�$�i���!	4�1M��G�hg�i��LHgO��Ty�y�^��1U��Y�A��)�i�B�&����Ӫp��k?�q�:Ā�<F,`��T����5�)b%��I>��#X:�h��1ؾ��O���rjC�0�E�!I��ͷ�m�l�y�2�W�pi�'?�41�^*����\��6�����gg�c��?ӱ�'�Uz���&7ɿ�t�+e��dG]�%l~�W� g�r�e���[#��V����U���U�z��� �K��I� �t߮��\��$�M�}1D&Q�i����J�CI9�D��R���6���_���M�a�������;�_�
6"�ñ�I�.J���@��x�T(Y�K�H8�'�
l�).�v �O�����ulA,�|�2>B�����
����NDi�ԂS�A�	�~W}-6�e�Q��l�g_��(W��""Y���1��4|��%7�V��C�R��P���^��*ڻP�ЯKh8��HRTN#�����4�B�Sh�fm�*8Y!�(V��)7�_
��,��sHq!yʸ��8�]׺4j�e7Ec
h�=V�C����g����J���CP�\ X�l j�5�Ӥ#&�!��nC�\��-$��W8S:B����Y�].)m�i>{�Ng�K���N�?�,ԹÙ�����,�͝9�#L����Pla�5t�f��ܗAU��h�j{���IJ(T���ʃ�״~��;������H�4��Z?�rh�Lu�Nn
!�di��x z���9n�y���y)9A�k��,��L�i�F��ᠭ�}���_��ϻi7���T��qme��uӵ:ϼTYo_��j��`��M��n��I��`��{��ڊY�+(�nv�b=�[<���n�%��ڙP�APv�����<L�$�0�$	Į�wvw�x뾓
m�?�+#G"-��X�&��d|��2р?ෳ�2�y�8�ZK҆���a5^�>	$�eQ�{U�� �����pAU���޶Ҵ�`%��'�>�Y#�^����+U�I�Uc��8/�]x13��(����%���	��ݟ#V��4�#�pҤ��a� /���,NMq(���f�0 b�:>�(_yU'�8�lC���j�)�zk�ƴIu�hr��|Ж4�f\G��?��>]�b�u�Q6�e�n�,ģ��%��x���jq(J�4h��G���'~��D�j(�T5����L۵�K�6��k��ߧ�,��M�t����D�2�rq ��V�U�<�y-�Ov�n�D�#!eV���
�l-�|9l��P��g��J�L��ۍ�p0K�/��/��kW�DQ��)B�XqF�퍆�|����I�S�W��L�{�Ռ����B���04Rg�N�	�+\|��#�g �S�!�']��-��(�U��X�|�c�/Ty�O��D8N9h�98)˰�݋��p��~�ʪa�qa5a�U��vɿJ:����V(�q���CH i4�0�Bg7�j̵�Sm�6�qg�k8aơ�h�4	����r�Nv���f�����*Ǽɱb���ܗ�*��-)ek�r֓�}J��-~��ɖ���mؙ1=]n&���6|�i�Zyj����;k6���;���d0���wh�.�O :B���*�b*�mv�����-�22��-�(g��}?�qܽ��]�U�1��_�G���@T�r�F����ָ�>	�h��G��ZMI��� �vlvi��K�����i8	2��/.�;PL�2[y=�x�h���t��~_qG���r��Z<�<Ś�8�n2����+~y`gOA1�0�n���<�P�JN��<k?�_.Gw�ASʶΫ�H\f�G����1�%��+`�%phb߯�*� 0�>8Q[��.l߷�O�K�yt�E���|�r�T��w)6�[�ԣSaA؉��t�P�J!+�A e��΢���w��뼪���9f��7@Jj�K��j��~�72�����}�)4���׋�3T����J`3r�U�jJ�t_͝NP�	IP>R�c��>L]�g�s�YMݠ����넔���sz�GOK���Z4x^r��Vh����Ђc�bQ�Ƒ�w5�*�S�1˽߳��ꨈ���	!�r�mx��[��EI�{����"��쨺�}���5=M�|f��u��T=$5�4@!�>�W�z�e��+%7�*�*
�	݈�sR#��Wk�F��[�M��j����txY�6���l�q*wK�g9G?4kN�.s�T��3Tu�4-��h��#Ҥ�b: @���V窉Y���(���scQx�iJ�H�pꋩb���dB_�%��K���H��Sd�
��G%&�a"kɯꮑJF����ǡ#�aW�Ow�"�۝�	Pټ��s�?�����^��t������%E�
��bΦ�n�ms7�>��{Ɲ���WFW'U�L��� w^Lj<EN��ڐ��Y�-~���}�?�-j���nG#ZR�tV���G9j��1�@�[�K»���ăft//�
1IE��2��]��s��CjW�BLGk�t�P�hI� ����Dd�[p(�2j@I�{���s��f�إ���͟�����xM�b�R��;��L���@;�o=�<�����Y#b;Gr��󩌥ȥ#���U���=M�#܇�gEQ�ޭ$-7}6�t?���(��r�p���.�5��̢ĥ�=E�`'��zW[�wK���KUCON��׷#z-��1e��YE�ޠ�:J�Wňl4�o�Rt���m1ҙ�>�
 ��̓c�D�p��+��8���	"������5#Q�/)o3�1����	��V_uW���c���ў~��gV�NU.��F�xFl$���R:=�_+��v \M����t	r_�}y�IC[��P%ͩ�Q�~�$��ay)�V����]�с���r�/���`o��_�&�?���`��^�׭��4�gx�34�5���ЕDs"��7ԐpI�Yjk��[�)Em	
����ҁŲ�N��!�B��Q@�"��Eí[!������Ím�_�Ö�b��F%G��ҶJ`.�!]8�哫��]�y�k�.�h������d*��dŭE48�l]sg�R�I�Df����j���MeP?O�qyQ��	�-;��"w�I�-���H�izo�>6v��},1+�6�H�
0�}(���!E�q	)�8�����-!W���)J{��	d��#���zv`p?l�Ey#��M��3�t���Y Z�%jA��W�4�C���n��6@�܅�K��r�ñ�s�9���?�7���T� ���$YdC=(�XCƎ��g<~�t�OT/�C>�V�ٻ�rJŖř��u�M��^1�ټ1dE�ik��G�w��8��&⩫{�磣�ܗ&�R:�#wGDx���%���"i"��1�����kn��%�U��B�%�?B����ӮK��w`hl��߰`n��3��k�1W�LE��o;�o �EV�t�O{�u4˸�?i	k��3C�����&W�Y��#':o��ꂺx�xVE��-�]�(�83����p��d|.잟�K��r�����V
o��x�9<��z��"��qx
'˖Y���q��)��Bh?r*i�-��VZ��2��kLh�R߼�@��D������]R�.���:��w�qN�` z�ll�Ix�ʐmo$��>=�x�j��ko�0LK?�znf/ԝخ�,Fu��A�Sʕ�����0��A*��H�ta�#B}�`JN����0nq�8�T�.�;:��?�jp���nzx��%�e�\j[&�Bd�-#!�!C�b|^~{���S!AT�R��)��ˆ�_�M���u��{-uwA2�Z i��"Ж�9j(g�ୢ5�L0�/��wCVc,��������CjB+M�����K�S��T�s���ݵև�;�/��S0q�dC��&���x[�ʰ��<�>�8������?����q�_лO�k����7�<Q��>�C����⽲`KQf`��s0��Z���ɍ8�Te%Ne���a��B������!�
w�^�(�6��$��͟��-�W^^yј���Yt�q;S�{���Nw��w=~ۨ��.�|9�q�a���;i��?�y�4�c��}�#�tM?������@nX�׳P��BsÖ���G��Άw��mr;�#Lѩ��@�I0�����V��<������e�{*�WK̐�R�P���'6��v��tE�݂9��Ϩ�.9�BhC��#� @��3�&%���/	�I�����x���^o't�2j��{�L�����PaWsfH��o1����Lֽj�.��o1�ؤӽ���2r��ف5Բܨ�V4�3�EB~I�f�k�
ЩDQ��=��^IS%6���'?"���(ǎ�2u�s��>�j@��q��}@��p��a���J�������
@?��	��\Z{�ZsOH<ؼh�v��U� ��M�-��J
`�1�0�.����� Z��sU���a�%#��d�_�}��^�T6P�����ھ�H�E~vF7�	��^(�����+�`�%+4v{U��#��Z
T53R��jn��#?Q����� �ʪ/ڊ�3�˦�9͞�����T6�F2*Y<I8�vm|�^�G�tV�"��2��v�P;X��@�U�ɐ W�L6$k�L��`�_��3��pH}����%=�~���Fi��V(��`O�Ŕ�K�Һw�碌��TJ;���b�҆��9da��27��Y��f�4w��>��deR 8����{�����fcH���wۂcۆڊ�Q�:�*R}��2al�"]�'��^�0�kP���zR^���y�r-Ht�i��={��;RX�"*N�����Ĳ���{�2*�[�ehzt�H��a���O�P�W\�+�$:J@�9¶��5h�j��s�Ŵo[n�r���ޣJ�\Q)9K����a:e��7a��$�� �Pb������m�$p�q:�e�|�q�<���aȒ����%�i��򚻻?D��Az&S%0���R�J���
y�u�o�EFv�L��5�=�QF9qI�	t��+��3�n����g�$߈OW,�r or�nh��toQ�2 I ��*Hk��\gK����}�)g��s1��nɒ���jO4|��u�Z����H�c{�d�h~0�H�����e�pD]�C�����+7\�-a�,M\�t��L�)�$��^����5�����k��.����.b0e9��ȼ��̺��%��MN���僵 ��_�ߦ�!t�UMU ��S:�x���(�r��s?��3]$i���V���z����ض��,�՗1���s��
>bc�j,HP�\�[^eA4E�M ʷ�G����8WU�_;=��\L}���}"�;�S�H/B�%Ynnb2Jy}���=�)ȟ10Ȑ�v�qS��*[�˔��H\�r�uo��w~�~�O�������D�a���`]n,�V��V[ ���(�Ɍ���V`����a�_Bha���Dw�G(`�.h���n�Pi��I��ǀ�F�v��J��|�`M�9J㶏r��ѐ�JY���.��sw�v�yS��7�N�+S�#J��dnuz�z����+Yu�1�{h�i&�	��Ȯ���#���Ai��D�3^O#H����v��;� ��"�_A��m��XȺ�\�ʡ��U̝A����~_I�����aq�O��g-*��V��Ǔ��=����[�E��&����<�� ��T�?���ccك�~��NUn�!���V��g=����T4&Ӄ�oNI���Ӵ>h���(ļ�ξj9C�^ ?�Kw{6$;��9�2��jJ����zj���)`����fN��*� :��~.�;���UxLl^M(��ח�|1�����e�d)Ae���t�3��QU�srZ���P	�J&��9X6�2M]���1�Fn=K��o�
�m�P��F� @2}}ڑ�6z��ӆ���Ri�R�/�Z�����3��jP���1����s���I�H�	�g1oKJ!; �"��O=��_T\nd"�*)�Qų�G{1\�����z�v'�A��_J]U�z�*E��pr$��e6�B�
k"
�%�&��i�~�ёY�ꀊ���t�8�V�b	��L(��>���@4���6y:��Kd��]���z]ʥATb@��e�ݡ>�iҶ%�G��a�1 �|@zo�<)�`�HUh+�q\�7�C���r�g�dŤc.RF�fA�Q@SN�󵤧���rC��K��=s�K��|+Y\��~�*,�<q�ob�zТ�+�z.��	z��i�1ܦ6��㓇"��A�����2��B3��x���W��X����A�	��m�rN�^�i;@���{���j�1.JTY�L!��;čG9Mrq�C��z�\Lv�t�y���f�xV��e���{���I@a�����J��ts%+}�jȼb���}V�%�<98�*`S��@��[�xl��{3X��#����u�{�t��=��BvaJ�A;[ ��b������E�m��2��Ǻ�RS6�(��GH%�L]��"b��L�j�v��O�:���gn\���[}"BI]�g*��|��m��,P���NK�^�RP��z�"k%X�'Vi1N�������Z�u�?��'�5�>����o'u|vit�����aS��sQ^��2��>��'��Z�0M�~v��O\{�]l-P�-��"fyp����_F(S>��se+?�u�UY��WJJ�S�	qm�5�oa��֤V�Z
��*o"�H�;��-?mKѩK`��ꅛ}Ŕ�c6�Y�a�=�3��/u����y�o`�~�ߺo�=b'�ƕNy3��Ϯ{=ܜ�,��������\O�D�#T�%�����E=&S����_yC��Q����=o�k��~0[�� ��/S$J5�Tk�<w��rP,�L����pVh1��15sh�V?��� ��EԹJCT"�U��I~������y����z��5͜f8��n0zk��]��VǪг5ho3ʡ*[d� ��6�1�h)���>��tj�jS�4Y	'��!��a���hA_��5���WC����y�سHʬ�s���k0�W�Ýp�ʭNY�����lqJ��r���u�������týK���Ȣ:�M$y��Ԉ�9%����H?��/.��80�u|>���{*�]y65P�t�lf�A�яnk���1�����T����^@*�i"x�˴�)�S�����T�)����B��hl+����â3q���䈺�dX�-��*\��������X�"��h�J�H��Gb���t�ܳ���7�̨�U�jY0>R�W8�y��v�өS��`�����^r)�	n��>�?���Lz��\�'���Ք������� ] �P�����X�6.�Ǻ0�'��<�d��"c�惆)aX"��,3�n/[wNIM�O����0�p�k�9:�('��~][�"���-�6j~s������t~��{kOW�K��'<�t+���>z#L~���h�aªbz��K���E����ff�����lN>�au6���&Z`���fQ����JF�JYE���l���
⹤����ޏ!�a���z�W�Rl�h�a��w�GxTg�]}An���A�U$���������2�zʹ����{R�F��D�6X�������9���A��Zg�e��%q��( û=�p������n�J�v��}��x�Wd�Ŭ�2^�#|���j�z����	�*�P4�%no���b�J@��r³ڈ�3q��4��ͤuxH�]�v�t�iHYс�4��&��.�֛�0��q�p[PE��3h��a]e�I����8-�!��r{��mŌ�a{ �d>�u�}o�}�'�XX���������d�{�ΐ��[�cP�y�&�*c�g�ZgΡE�,����Q�4�n<^���_#�,N�)��F85s�LQ����/e|;Wl
a����h�Rk�Є���yt@U�B����7�B���'�0�|,�7����@2��f��a���L+MZu��o��R�
��JU���P��?!?��)kҤ��;���|�����M9@�V~#�ُ�]��;)Z�Qdn+��L��ry �X2��H\�B�i�S����� gDm���q��8���1'-�����+]��U�b�e@����&~��4���[4�Z�b˪��b�]�uӭ�R���{ٶ�PŔpX��;���U!��ϋ�gPA��75�����:-	LD�;9�3eK��&kb�ǧf9����p��!�)�gۨ>R�,
�G��1�~֢e��i�����'��ڝ�z]L���-_��Ė���Oب�E��%�E�8RG(JBaT��l�|]�Ԋ�{�H��z�,^�o���q�+��7��@z�(�	���}�b���z�K�5Cs�0=��-W��M�J�^�쥗��W�ƪb2y�ӯ��}���"�����3�=<Si�kn�I���h��jG�'r*Q}�8j��j�^M��X������4���/�]��$y��Q֌���Q����tu��K��2��`{�|�o']%Ip��r6ʹ�{������L�0��9��zU{۞����+�Z��:���ؾ��L�G j0\ ,iZ��]h��K��ڛ��c#�I$��1�\UV�M��Y��i��w~-�Z�#�I�`��R; v��  U��Ⱜ-/K�g�?y�x.Wpp>���`��	k��-slI�"�}@��6��pku�DE+=������E�i�=��VO����#�D�k,�2?���>��^��}Ԯ8;�:��M�sP�G���+<���c
Mŧz`Ϫ���7P\��2`o����8�7o#� X�K����K�� %�S�|%��X��,��`�ʒ�mW�5-��%�}���u\ʻ�C�F� %L��W�Q��+�|��%˗`�!��ޜ��v�n�8l�yH���R�m�&����_��	\��9!�Ī����fv��ФAe���͎��׼ʭ.���h߽��?���o� �_{�O!F��ɶ�b�*7���7����	���'&S���w��<q#1�ȃ��m���Q'S�?��<�ʋ���d��_~�"
p2'������3t��ܢ5����$F���H%6�F��d�␔)�yѹ�u�X�GS�Š���@����Y�L��WS}CN�ݤ�Ƅ�7������ё}��� )=2�.���ô18bNU������V�>��R2W�c�ճ�T�qY�A�����\�)W#���D搭9�ANŚ|��?*Il�ш[R��y�i�S��*qg¼�V�m@j~"�f.���4�N�� ���"j�ó�@��X{�9���4
��|:y���\�RR�/4�CV�D��b�N˲��4X�au���n��BI�T�orf��L��7r�|͟�+�"�H�ͬ���G⟒84�1jgYX�C:"�f&v(3�O�A�Q��sN���?��Ҝ}��	�1�T��Y�X)n��VD��"�l�fس�.h��o�o��f~=����*U4n[��D�rq.�կ
]��^LE^����=�#���v )�%nw��盧n '�V=�oE�,�"	�~�NP�݃6:S���O��}��7&w�i����臀�#;V��W�� �Y�E�e�a-�g�(�9褄�����7S9�3��~)w�1��^C'�8�bs�%��>S���B��d�ΏC��$���m?�k�?��6�Eiw�K�t<}/�>M�&P�$oK(��k�}�NVΆNs�s��Um��v�K��\�y���!�H�F4�R�M���D�k&��r�	��0 -�� ��0vپ��٢�������;��O"�P��	ZK�Ь�UtK�O%I���q�QTn�QpG]�]m�i�d��D�+�V�^�L�{�7�EY�ǹ@heY�'�PC~e�UN�P�e�s�w�귇��)nc��Ar%du,/?>����'�@i��#�x�J�n��ѳ�)`�U���a�6%L8�?`ZV�&}�����cI�%*c�Vs:tH���;���>#�R���:�K�H��Qδ.�q6�扢�``��¦tb��C*�l1��mm�q�1�����{� K�\�&�P쇚L'!ohWi:E��
3����MSEK���> �S����l�
��E����e�{+fm2�$�X�=��o�0�^
$�x{q!���)�Á���<��̧s��RÓO��W��\�i�T�7��; &'`(@�pkwE�ص��r"
�CLh���7׃kǴ��G��1xA���7���6��՟��'p�(I�$.P7�/c-3~[���k7�Vэ���ZCw�&d�9���N�K�*Q��_�,��ǖK%��
��f�Ō+Ʉq�z�̰�K��Q`b�͕.�t&�ushjI�R/j4�۽�+��:Z���J�D�i�qJÐ��{�4L#p��r����k��[9���owvm�D-��:��^���������q7[4J�w�G.��,e��0[s��<bGe�tkT�
�v��B����U/����d�D�7�Gy�hrG���gs�(0#�����Ň�5ʂ��;9��g����~���j1�u3~H���l�s��P_,�q:�W�z�a�J������T�����$��Tp@J-G��e�1�j��V���Һ%�2��!�Zx�=U��Ho��-��ʣ.�>�w~�ux(�g�DZ�\ࣆ�)�o�sȟ�@"�c��$z桹B�@�X!\�!�������z��zʽɲ��V�
�R�k�l�V��V���U�	a?\����r���� 机'�2���<(~��y�ѭ�ٟ^cX��E��S�I��3X�[Fۍ5C6��c�2���Ӣ���㽜�� "�|XN&'E��M�a�Y֣9�gq�֏铤���&�%�bܷ���Y���f.��mJ������f�Mu^ށ�.�ͽ��𞌱GpG��yB||1W:�Y��)�D�ɬ��	Mۚ�H�!����j�WJ�;I�����a����-��cz),Q^{�·~��o�)<��x�*֠������\x0�J���>�-��1���jdŔ2��5]�"P}��c,yN�����꬛���n﵇۟O�f�������w@`�����mW5�Z1J?ƛ=b����$ٛ����[AH.��NR����˹���e��Bf4�9T�i�����q��r"���8�_��g�^?�o*cV-k^�6��� X�k�f	���	N�.�sG<@���������\
�΂~1�W"����W����B��+WB�q�rf6��� {��"��A��Oݠ5=䰆�s_�H�(�y>=�^B�9>j���~`�0Q�֚�R�~�ơ�w��~"��32�(���w�!)w���ᅚ��+e�&\=���6�Xv�Fְ��sU8�.)�J��\8p=��Q���y3��_=hܱa|����/Y(	��xJ�I���5�m��D2!�<�Œv�$�0t�s�҃/f09!40�k9��m�1 �	Ě�Y`C<;��_�x#���eo�z,{2-}���]lɑUA�F��������e#i�Ty/�?$�^!q��3O�s�����gp��d���]b��u^�2��(�x]g�}e5�R~5YoL��MƯ]D�#�-�Zg�'c�5�Ē�W��f6�#c\)|��6+���d/_�F�'6��Be;G.ʙ�g�|��)�Uf:%���awB9���F�i���Ѝ����r������s�s��q��gA��h�a�W�0��g��\����%{���T��W�v�å^��U�EWofU�9ދ��خ.�5�m�9��VQ�l'P�����P+�=Z�w�R�}p�B�e.L�7^�a�D�O���m����<� �4j�󪑴��,�K��B�H/6YchzF�����d^���xsf�b�_�Nч>ߟ~0ꏴ����>���O���e~j�_f��T�zv4�]\�� ��n2W}��`�|>$
�ja.rt.�Roo�;��A��	@N�g���Y�� ���0��,]�D�9L��7X����l�!�����͉B��5���ﮌ�(rI���`@ ����4-M�:[�Lu]L��w��H!�zOៀ0�"_^���aT�n����mQ���G%V�VZ��δq�� ٴ�iBDƩL�U~�aW��%;���b�����[ʠ�=��up�c�w��q68�I������z��~O]1ޘ�ז,�1ЭlyK�L!�D�tH�N�$���]���<� ������01��#��ɕ`�nD1>�K��Vuh#��'d����x�<�`��y��7�����n{��w�D?7��p͓?�i�V��/#nk��J'b��IKٹY��O�;�S��?�L��_U�G��m�V��� R����#dDG(zY���83y$�7�I��u
��?^b�Q���8`8���{�[�WJ�����o�����) �����xe� i�
&�4�,�H]���|�jv��X�j�uG#�@�>���J&�0���k�g�A~A(v�ڏ&���� C<��6�u!�8l
�Bnc�I�157��h�ɼ�}�vL��F�-O��)
X­\���
u��l�X��B؍�}1��+W�7�ލ���-X��uǙdc���� P��C~�}��j�p��١.�j��g� u��+�	�A�b�^�]�����S͙0	�����T�����h��ϊE�|�p�S�X���KH�"o��F8�����K_��k��6(�y�aJöI��Fڊ���X8u���n� 	P+�pr���a��)�*���(bkvoF��#��:�2�Ia�CΩ݃k:*9�ޟ,��O�G�AV�>��R��]�{��|��	���|I/{b�na6�e�%�N�k����kĞ�hۨd�pǄ�O9q7�	���*طwk�nkx᫿�m���(##<ɳ��@������r�Z�-w8#+W`*��/���j{u$S\:������H��'v��1룋�O�g�Dӿ�H"� B�\�����{��8-�dy��DG�;������8(�&���B���pb��B#>�chXj���=4Ǖť���SfYY���3��x��4*	�����nA,0��5���� �O��WG�х.t!� �D�e�?ީ�=Z;����ɱ��J����Z>d�:F��!!���1H�l��_��z�x&�ڹ��V��Dҩ(6{��'�ŧ�o0?�IƧ19�ѭ1�����3�a�>��a'��uq)7m�#��bc�x�����pD�Ll,V_��W�-4` �ӣ���7��
��"�@莱��&�La��-��#��R����b8����l�}�G�=&*�&%�4����-ob�S�
 M���˒�S}�[�F!̢d�� ����PoX�J�x��	���W�q�RB�1��2����(�����S6�����)h"��Rzd���R�/k��X�Q���L���ؽ	t�'���j&��#=�D;[W�U9����ɤ>��(6��Ez��!`e�8!kv��:�9VS�ɽ�l�v�h�&N��҃}�4��脿7�eb��e	�IOP�CA�<�8�#0��a%��R�~���T`{�x���&��G��Z�v����WJ�
@�p�\�+�4��HU��'�]�T;,tVd�vF��B�-���Q�g>k��j�j>�x0��.�Z�{ۡ!�*�q]T�) WC���k䄞�����R{�Oy�N��N�g�&��O�p	ܬp�9�o�*[_MG|7�ˁ��\0�o&�Z���\��]Ah�~��L,Z�Ѐ�iȉ=�f��{�^��i�so��v34ˉ~`}�<B�_�����iV2$J]I1��[�ZE���ܬ�T��2�"s��2z=��L�1|/O��d)�
m�t���6m�Ϊ:^���������+��Җ{��q���d�x��0'1���>���6I'�#;	�	��M+����6��?=��S.r}�q���B=Y=���s�l��fR\��z$���-�W5�����!l�߸�V{ݷPZ�t0B���Tr%�<V�3��ɒ�L�);�]X�.��.��y���v�ak�24$ƧKEU>��/�ca��Cf_��?/�L��DD�	S��n���oRTdU.C�S��@ϭL/͸-?�׍���䴾+��3X��Y�3l��	҇=��ĳ��@�4�gl�$����1��$2����.O[%	��P�Ba�Sn���0���הx�@Q��:I��n;+����]�H?H�&�sV���7E�_���y<�x'Z|�8��x��H�"C�2%�]�Ø�S$��� rR`67w�=Wās��5�j�Å��� ^g��ڻX�L��$���령�";unT`���џ{nB���擐���1B}IE8�5����a.h���C׌�L۾?2tB�Vo��@��$�l��lgZ	ЭܷG�X�a5Id�|�ǫJ����x�Ѳ�
烦�����(Η�/u�f����gu�nћ��̝ �m8�M8�Bا+��M���*����5��!��Cul�c��
P=�R����Z:;t4	+�Co�Jog�j�����[�6�:��wˑX8����WAWo��Z��[ڊ�{k�G$)��.��,���Q���k	ׯ1�
X�c<H�B5�~_����\�q���H��^�y!w���\[nfpˈ�\�MK��=����Y�=�V����j��oyx�i>�6�Z��j�7$$+�g��S�{E�F/:��ò��J�$\��.	AN�E�b<�[���:��N���@E��3ʋ��BWa���r��yR���*��<��E�s�5U���3��#��3�/Ds���6L/�l�߿ޛ充�PF�vcW��:g�?vV�L��}� G#S���W&��l��#�J��j��!��ԡ�������v7�4���/�Csy����F�&.k�\�3=6���|cJz a�C�g@����"�5Fr]~�q�z���n��7�����Q�0]
	Qכ�E�]^�S�N ����	Ou�y��|z�`� r�5��]�0xzB�F��Y&�"B��bA*&)�)kw>�{�ں�>h���Z���RI����j�F`�m2��{�t�0%�J?`џץ[�/����݅�^)|�G�p����{x�l����	k�7�n26&MH�l�m������?�l��$y�*���&��	���R������̬�[�V"fg�b_[�Z��5զK��Zdz�4�1�Ϭ�f���-��$=df��fy4�7���q�렊A��v��誒���Il��������]�4�FgU�Z���`�C�����1��6-5TҘ(!h�=562V���wg����єx� uR�H�m_�BY��~3s���1���/�Dڄ��Wٴ������rƛL&8=����ooK�#����0>��,m�ZA~�]32�9��QB���"嵱}.=j���3U���!��۱�3z���sG!;� ���~O
b�}?A��N�'�e13��y2�/"��S+�Efl~P#�Aq����8�*�"'���1�R����߂E���k+���c�����&d�Q����Sɛ:��VhY����>e��9����N)l���'��Z#�8���T�k<w#��o������ٖAq���Ĵ����}h�R�)#����h��dn��!�Aљ�j�r	'H�-�O捦T�%0(����P]��jy��nfNn(�rQ�5b��bE���ٗ�.m|&�*Y�9�����
�UY��-��ɱ�`���u'�YL��˓��%=���K@Ud�Y�An;��#C�U�]I�u��N����gY��Z��A�U�0 ��M��_�8L̂�����Nq�6Gj7��m�Tr
�8��a�׳&¸��ǃ�z֗"DX���9�5�88m����"}�gZ���M��Z(���޹�F���˼&o�3?�����v�P9.�WB�6a�wnTg��𜕲SL3P���E9]��w:���B��I�!�]��)�Ws�BYTq�v��f3�ꚅ&�-�ړ)�!5�/�$5$v�A���l��9ͤ8��6���!J�f�$C�
��r��D���5�+>�y��f]��K��zH pyUw
���>?O��Aͣ���4��/X�ǁ�{�1+}�wiWP�)�3@;߃a�BY��z�.k{~/M�����M��
���g�{�zv����|��8�6�vh���@݃�d��������.��8����i�-Ax9��6���(��r�~%�_�V��y����U_è@������V+�X�l����
#B����F{�$z�j�P����7;�چ�opfLϷ���a�K�ڻ}?��z�8#K�,�)�v��i�č�M��^ˆ��*ԩ�=H�Gn]e�#Q�N�gFʘ��O��p�����@�d���v��Z��~o�+p�nN>� L:'�C	��]�"���Ã`����:�̥�Z�ɝ�ZjY%z��P��	s���0�B�h�e#�W���S-Q+ٍ���aU����n����u�|z��|�$���>�v�@�7�AD�vk�f��q�p�T|����+2B ��6������[�7��O�/�!�������Ȍ��\�>]�Y@@�9�I�*�b�z�`w�|�䀌*�$��'�h�S�]���5��L,U�PñX3���-�*&fh��(�"��D�`�16w�����Vl�D���f#������{c.�@���df*rI��}�:?���T��e��sV:�VBCq��q5���9gޏ)�&o���%���s��dR�`��0~��
���D���=�I�9!M4��\�5�UpNQK�87��/Q����!��`��Qg?��>X%���ڈ�����=�	I5B���Z�܁�rB��q]�U��&�HX�_����B�*lD��{�k*i�w&��Q�>��|�Q�~��#�b~�� }d���P������x�5�ws����j�e��;( �)驪�Fõ(�>O87b�ד�=�[�DSH|�V�i1��x[X։�/P	�,n�܍�5}���}'I�,�Y��0�tJl��X�:�й�e`s���m�>�.��7!/�2�j�H� (B����))|ir�W5^�,L���x����/��"���{E9yX�ڕBd�"�}iX,��nA��|�p����@y�/&��6��Fd�)�	�8��8F�1�Rx9�����N��߄�WU�\��o2�@��L/��]��+nB�Z"*y����s%��mi�����xh��Cj���W�����ǵ�aZ 21��Z4	�j`m_�<ID�p��8�m���E����y����N�ld��>h]J��r���,�*e�gX�L/��^�Y��*�%�/��җ����B�+��vA��lE,8B3���y�YW��<��7�h�M��W�7R�p���hyɡ�ɮ��wB��M��5W���jF}��*"3�SfYk�$���Wr��:��Kf��-����6��&Z1�ߋ��%�=n��ߨUjMZ3����A�К�n�ڌ������g�f=�Ӂ�]?
�+�+���ǆS��Ǡ�0Ei��n7~d������(T9S�b�|���JпҘ�W��8����\�#��4dtx?G�N���x���UJ^��ӚK�ʑ�C[wǑ����"9��)ʝ�
;�������v^��| +�- �V�� �m\
��?U5=q�ab��㲾M�gu]�*i�j�}����T��F�n�Ny|�H�DUHVE,�4׉~��"N�]ٰ�5��4YU�j�!��n��l,?>[S9c��1�T�݅����t�,������%���9p���Q=a~�/]�rǯ��h<�FhK�R-�f� pc%�J�sM�ًmKd������m���$:��be�_3��7��XNڜj�Yf�u����oiX�Yꢅ���X�;2���4��i]�	� �ۗ�T�.���Wj�rhS<��&����D��7�����ֿ�)J��"�Wꈔ��f�����A�Hc��wRJo��X_��	��V\w]���#�Zn�4`���ӫH�yKwD���B�k���m)��5���gQe��\7����Rqf��{��QvM����sH�ѫφ��-3�" fF��w��Ƌs;��$`��i�?Ac$$m��c+�s�Of��@�,/��y��'��c����=O�)��`�������V������u
-1c����c�dr�n�X*��Z�l�;X���y��۝�%�֠���9G�|�ͱ�4DB`'A�k�ȟ3����AxP������>A:R�#�:f�����,���q��M��:{���̀j6�[���R�3�<�/����OSQ�������z�������"u,y�@b�#]ۙ#�����c�(ϭ��3��;P$e%[Nl�*8���.l�36T���0�r����`������;A������x�&t����×��ov߈��p*	z{�Zs*�����0 �� �$���Ks'�W�Ý�Wq�,[�~��ӅyoY�A�)�{{�7��'h�<��ڒ�<�X�5����NXL�0��"����^����"���3��K_6@A�y4)׃���E���t4yZmI��p�f]jm'��:�@�?X/�u�΢���tf�[ہ��v�,D$��jb}��jֳܶK�h�#�B!@߸ux^[�9��dԪlD�roOO]d�����Oe��&a��-e	;��@��G���34$�)�����߯7�(�c�$�©��&�F�\*4��p�3Q�W꒸���.{gH�t�9ߠ��`�jG�f�\�5Y,�d�rA�7�;c��~mv.B.���ؑ=cIG�7�m�ӎ*�p����K���$��39n���:�<TT���$U�����r����a�`�RX�bD��Yty+jK=����E��h:�*�]����A���*>��mt._9by�&�T�� x0Z>.{8�]�b���*��:E�`�`����>��<)w�2J!+��L	��l�(�ͺ�����|�0b��G*"�������]�ъwsQ��HD��;*�|�N��`Hi��(,Rc���Xv�Z��y�E)5� �@i�&6�$�:�q�}h	�w��=��O�}B�$Z�����:���W{�ȈR�%~3��!�[o5l|]��Mm��N��U#f��K&|5.�Ԏ��ͦ~��O�7����ʼ�5.���;��0��(�k+WǱE�ٚ���-��/Am��L���eюTK!GV�e���y�"]6W� ��S�H�\��#�t�Ȏ<2Ļ�Z�''�J|F�}/�ݠI��A�ܮQ#B�|G����i^�Xڭ&C�z��z��3�dכCb_o�K�8�w��p�,�7����U���$E���@��Zl6�S�J�f��7r���[ڛ�����ZN?����(�Fir���]��H�ܣ\��Ư?���B���^~Ϛ�4��e��R�b��f����:�4~5��b6Q騴�D�'%а�	�JzE�3l �����O��E�{IA��c7��`�;J��6?d�꿲i��q���;�+��z�\�:O�5�)��(�c9������jߪ�esTa���E�:xJ�e6QX���K�ofײ��QPs^>��\A�p5Gn�6�ɘ~S�,f�<0�j�!7ؖы٨�O���a��Z�8�c�<p?,�TW��q��Hڒy&���9Q�{q��lS+��E����m�� �l=0! ����έ���P��Wѹ��z�$pB�s%:��2FW� �b�+x�x�7���=�:-�ߞ����c�ذ/�H�O!xڛ����M�������%�(g"�3|�]5D�B�מP�Œ�VO�����>w�[����OR�7t��U3���֖zڡ��KZ��ksfE��h��z ����ʑa���u���7��{��?I}�G���M�f�S�*��'І|¨��M��m�-�7(�C�_w��xY�߇ؘF�ݥ,8�u- ���q��Qu0n�����MTHW4��g�ؠ-�՞4~��m"{�E����c�'��Z�A�\E�Rv<�E�q#�?A��v�Q7Ҝ_�I\�� ��S�g��K&�;�s�$9-KW�"��&W*,���g�7��k�Iy���)`zgQ�_Qm��������/}L�v�!�X�î|t�y�=�.l}��y����j���/�M�i��+�P�:ۗ���*�D��c۠I�(W��ѹS�������	5�g�_�I��5'���J�.��`�m��x/̿��ʛ���t���k4^���3I�c��*�igguhD��:,F���������F���T��)��n�N�d+ꑤSn����4�@�%􏤤-~h���K�����1���z7�j_Q��M�Y���x��0_��&	ǡ�����A~�v@uE����
N���;:]��)'����mA��$�P�����̔� ��AF$4x��Av �M^Z���([dqnS{Ut�cd�r©�X�A�̰���0����;G��-|��������d|֨�vbk4�M��\p"�
_c���B��[�qH�q��~��N�2��>Ј=�	V�I����/�k�&n`x����G{��"�D�i\>J�B�["�_�t�5�˻f��uo����0s��^�~�S>�w��+����"-(Âc�A�X�$�@8suv��(Dx�Q�!&V�s��[���?�@T���+��F(G�qh���A����X�OM����E|׮�R��ł�&��0ˊK�A�:�#'��A ��QO�$6qs�π�[tQ��@F�v���@��9�����A�,c��)x�:&����bJ��aڢ�� �3e���߾h�R*'3D�ҳ�J�SEd�SO�1�瑅�׎�2��|Ob��\�z[���szn��=1�U�����QV2��Qj�o�E�����dh�2� 2�
_���O7!@��6P	򭨉/H<�c2�ǂH��/N����W�n�W��������]W˱+�S;ӑ�3�)�P���f��H�眵f)C���e�d�]��W�q~/�8�a�4U��[�m��Ӑ[_C*��p�����T9�/1���ūf�e�����a�e�2��V]���͆�t?F���i�e(o��ralՉ�0�k��#ʨ&���˸�a�K�|u��@zLq(�bte�(���W D��]�M����	+Ee�,��Lz�,6K��_mb��h�{}�/K�Mr��(*�c��Ml:�Mtc�4��X��%���<�$�5e�3x�n<MGg�/6��&
��`Z����/��v�)�`(%s���W|�G�����l��^�l���� ~�i
F�a�\"���>u�*������:��
"
��!u�tL�3r06�)$ϙѓ�D��Rp����.��	Lq���J��A˴�����4۝���%YAG���uR���D��]���nu�ޗyn��؈P���|.jJ��ckc*Dk3c�{�:�>�)@�h
x�s3CLݏ�ķg��76�]����=SC�&�2�n �wu��M��J{��s#(��{�8�K�o`Qe2{�s��#cA���33yG��SA���[�ڎώk��	[�S�p�,x�R~k�D
ζ�Hz
�r<�gg*� 4�\�J�tB�2�}���#����ס��՚L�������٭>I���ӯ���6m�P5�ݮp �	��Y��	{�k��h�D3�H|�
��R� ��{R�Z%��Dx����B���)X,� 5�N���0)�@"���K����CD;^m���
>�a�
���̃�Z��s@uf�i&�ų	�
&��Z�xؾc�Vc]]˧�VL�t`�jVr55_�x�t��O:�<)߳S�@��Zv����/�${^1�n��:(�ָ#�D>*�A��Z�Z�K�#_ҧ����[��o�2>�1���K�j�jH��[ʷ����r�XfJ5�9T��z���/�lO�A��2�Y����ó,�/;aQ=�ز*���/|/�-����,# k�� e")qI�)����OC���+5�I	��	;Nda�d��y�(����d8���k���'�?K8wB�Ӗ�!�@������OǄ��_�_b��p�@Я!"���<��ܧ1���y�E؛s�A?4����	^�g�.tf���8���λ�����5�9�ܧ��q�L���q���,
�RJ��������y=N��G�����l��W�I�G�t�-�Eg3����bS0�b��_���(��O���Ni�6�շ,��Gy��P�O���\��H5���lt�o�^F�Ts��p��u�n���ж��?��!�7�#j��KiZ^��SX�fX�"��L$V�(+A���I�$͓��>
����qQ��q�����2��=��֚-!d���]�n[��E]��Q��(�8���օ�E�����=Q�w`m膡؃*�2��]�D3�^9�W��B�u47����d �=�i��8��D`��b)I�9qJ��2!���c��X0�˰d��LNńō��}yJ[	!މ+Z�V�o��Q[��s�.|	�6��H��nu*~ةu %H*ek��v5m1�k7:��� A�N��,�>>�����%J�t���������}�"7`^&���
"/�I�A/;�=��x�l��Q�����Fbf�n�6z/�*�kN@%`�nZ�ў����5w��ɇ5�-fٓ���it��?��) �?/�'��s�J��w'��nxP��ԈA}#\Y��/	�$�>�ihB>n�\���&�.o���V�/D�D���h]�g�su'����g�!�>qq� 
��?��Q�`\'�����N@�����D�n����F��;cd93���i��}�QL|���BY�Wug��{�̖��M+���}uGFZ,v�E��c�ABH3I"�(Q��eU����´�~̲U�	�q���qq. E����l?nz:2��m�ڑ���g:Ӗ�ԣ:6 },f�4�Yx�	{��mt�H1-4�����^F`��&�e��+��f�����@��r��ε���`z���?�����\ ��#��2)���ߏ-�Ϥ��r��up)&n�n�0V ��ZC`�+W��tD�F���F9 ��%��]ol��o�����iލ�������ToP���5M�I�l�]"O�3<?��59��{���.0X�P���&/Ό�a␬�ŕ�﨏�nWW�7Y��_�����{��.f3�MAc�$|l����^y���Ι�ok��&:�\�:���Q[�E|k�7��^����G*�*| �Z�Q=�tR ��&�,�$�@I bĒ�<��B��ֿm8����7w^a�?���Ҕ�T%a���9�ře#��{O��J���!��fc�竹Ŵq��1]�A*�4$��)�h	�;��w���'�nn�Xm����IG��{A�g���ѵ��m�v1�:Wn� V�&��`4U^���n��zL5!���#�>�Xp�:�a���Tf1�kii�����0�t�Wfa�"����X��0E�r��H� r��,�_QzmRx'.w��#㘆�o浧�>x|��Y��W��ۥ��d)�-},�R��T';�ȑ�h��ޝ��#0��t>Z�����P�.��DQ����)�����IO"��1�|�,h����O��DStֈG]�ʓ�l,)Q>��)D��bn����C����]h���=�6�`�U�ЂR�rn��"�Y�#�����C�ב���7O���q�)�4[��I��.#�h������^~l�(Lė�R)���jUS����>�/��C��k���k��'{Ay�A�p_�g�;�d���a�&2Ω�9�����Z.}d�Q;9����uݒ����ݨ+�RLǃ'��K��8{)�]*�(n�-����B8��3Gޜ��]O��\����}*������G[o�R���_y�Ϝ}�B��݅V�߂"A�;AW�M��9���&`c�b3�	|�.`a��_���9D�ж���!�L>olZ�nq�����+�_=�J���Y��ۙY���׿fR���f���@M� mi��:��S�5�]Z+)lG��;2"��H�̧����6���@̅jx=�z������R�[d~cQ�__";' K�崾�ZS�8<�mS+j��p}���-�B��fw�@� ��?�<U�ؿ�q��hq_����ŏ�z��Z�r_����L%�;&b�а�j���y%&�&���lv�W�i)�i6]YxJ�^�ش1+;<�Km�M��uO��մ��-.�GcK�ea��h�x��]w2-SiN�c�Sb;��j�����w+�ra.&�vpuc�(�ء��A_����\�R�I��a�\0���0|\߂���;C�,�hH�����w���.U�9�$������=H��{Amw�I����Ab3~�Je���8¢!I�J�>1�,ΗkI��u�x� ���p{y�K�����{����g�9�Ҫ�QѓNQ��l�W[��CR��x��`2�K*j�(@���u�� �q?��j��QEq>�Q��m��0��(�����jT`A�����|.P����4$P�=q��;P�UK�G�9^im�Zٚ�f9l�-�thdu�4�C�`�~Bc>�'��HreO�>�8�|V�2�5��z��4���5�����C��l쨽
z�G_i�G+π�H5g�KbV�sԎ��~R�~j4U�S�E�r<d�^gT[�M����%�y �z �+,�e����ט�*4$��Z��k\�i��y���L��z5$��_��YI���+��t��c��<��؛z��-l��-�M��UOj�px�ݫ���+n'��g�v�C��D����E�J�V܄��;K�w�]h���z(
��R����i���X�cj1��ns�f{D$�r\�X��7�g�ln6(a��*�_h:5F�;-_�������-�"���	)^��x'6��7���*D|�OL���X�K�u4�ת�O�F[�6S5��f������
��n5��!5�>��?�8�9lb�a%Z���Ջ_�?𼋕��.K*5
a������/#G���Ym't�`>> r������V5x�-��*�La�����τ�!�#���K-s��8}+THf� �%
�{S�U�y�<��)�������y��<�_��6�H<=k��Rk4����7)�̊��zHn���A�Hȩ�qB��El��W��m����g�P���N��q�md?:X��6oQ��;�Z�6�ɛ�{���v��&�(bC�<�)@��q/[dX�5��@�s'���]ٯ@EzF��jHR>�Hu`-GR���N�,sU��:J�.O8�Y``r�~E<�pप���re�\�q��:�K:L�6áP���u/.�������"ų�|S�p�c�OB�+4u�.>X��h�d��	�t}*;���SB���a���O���V���4�rCr����9=c�9�m��ݙ�jw1fу	/��>�>��0������q�C��	p��������"���>�!~nPj��[�!���gEDw�ذ�rrK�"��Z��~}̬���Ҿ�Y���c}c}�ٓ�S�B�j�Oa l;���i�PD u�g��e��� !UJ�\%���.hp�h/�����٣�*;�W_J�� .�W�Mj<�����ia����������`��謜���r���,��4�5"�#X��-_�tN��q��tձ�k�*���6�12�B8�yDVΪP�q������^�.�~�ƪ9���-�s}f#�:rCIY���#Lupysa�WN��Մ��wn,�n�柷w�2c17�նW6��hJ&���&'j^�3c Ax�I�s��j�����`"a�w]���b�Ipdyo� ;ⲱ�')�3��S�,�z{�B�D�C�H���<��߉�f���0ZPZ\���?SL>�;���,i���,.=h��.y�ʸ�����Z�O����o�_��mڡ%�m�����iH�Իm��6�1�I6ɹi-��R�;� ��V�Ŋ�
��J�)�@�����y���,y�4��f:V���2��,-�F��{�Ŷ�Ҕ���r���o�����22�����(�҂�8cD�W�xX+���
�#�&#P҃)�WA���-I�\��s9O%$�V�0��:�@N+?n��������%�w�:3�k�|%�����@,<-��f���f��8���� �Gz2S�� ��>l���Wl
���\"&�[�A�^)��R,�WpG�Rb�=�?m��6��[-�jhL��k�uʺ�*���l~ne�2�!��H=�p�	��Z����y���}�n�Fo��W�O��7�}�^?�
c�m8�1Q�]�X�^���)�h����$�Z�,���k�Ȼ� ��D�m��-�1�_��]�n��5'.N�MA]�x�+�f�H�Ľޙ�Y0���,[���r�ٶ��J¥��/�;9�� �$ߢ&[�kR6�Sa���Bh5	�נ�;'�Rn��Ԥ�o�~.M֕-�|���6B����W?��4u�,���`���f�~�>w��������.Cv5�l��X���/꬇~y�)�f��}����������@�c���	� e��,���~�z�H�Ծ�e�Ce�hwr�L���7{%�z"ˇB~�����T��U����i?�^�yu�߅���[`L�3�|.
��T�z��'�B]�De��5��f��x��R�+l��26�u�F&�]����X�}?2��H����� �!���y���L�5m��۳��,���#	��@xJW6�x�l1}���O|����TvR��8� ���w� ��u���I��OW)8@�Nz`ӓ
Yd�i�ph#}ܱ�j�peO[eX,"oF'�O^�#��YW�w"J�i������*^B����PD�͋b�z����E�#��'�H�n'S�0͙��{� �H����%�(%�>� �ϚVg�ѶM��
tNb9����R.�ьaז��7�q�߻����m���Uc���"�[�7����]`�t�F�9=�r�aD��<"
���I��U��[��9
�v�	����:Lu���F5��!	�q���@�1��}A�����ՊZ96���u�eq�?eM�bd迩���nb�eCguA�'���8�	�?5�fF]IhU:�9��$'���L2~�����
��T��/"i�
�,y��������z ��L���hkj١S�B�2��ז�����F��!��Y�$�i|�q�O����ʅ}÷bgI��n�ɦ0�c@=�\�q�:�i4N޾~Ec&܂�o�W�#J	i�S]X��*���N�� �,���*)�/~�������
����Fz�D�k����a�8�c�n����7��������V�y�w}f�����oz��B2��0�|����2m9�C�1�/W�N��tI�2��} aν�!�����M�'��;�>9u�:��?I�ڠ��ED�ʱ^�˥	(�esH���: �j�J�ͨ`�S.oD�� w�^?-WPK&}��=��6}B���f^,��旈 �xI��N�b��{%����Wv]gr췿�Ok���.�D��Bpʫ��0Q�L9,�ח@dJ��������ZC��$���W��(�P��ư*,C?��G�o�-�gՕ����j0�i���Ob1B��>pa@n�B������]��|-���]�x�џ�`�Uq=n��^��TΉ7�]�xX�,s�!X�s-���;�2lͲ�&lxbM,�z��n�4I}�0��cP�%m(�7W-^�:���d�Y@��?���
w�Uܱ�-�ؙy�2ס]�(1c$u�_�-�D�!!�8m�������#�f�k��Ix�`�m�䤚�2�F)�*Oμ��z֑��[b�؃�4Y�hu@�g�3����=���}�R�>�R"����5��g��tF�R�
Ȁ���x�"�K��P�io�A��,�_�L����*cC`3�f�ɦ	�+�O��,�:�I�����<����m�ŋ��w��i��_i���N�ɲZ5<rX�0#��;�ܤ����r�]a�[����}�r'zn�M���+,���V��V���Rh�Gx�u@
�R!�T����$���T[7�6<NP�j���S15��Ȭ����$6P�S�I;&�Yo����.���Eh�x
�*)͒���,�8���M	�ض�.M�����])���)��,��Fa��>;�j.
�{~����9T�ȭp:$UǎJ���d�l�:(�ԉ�Kk'�I\i�+����^9W��?~m%\��F�6�~�)Hs���z�=�Fꂱ#�t����j�\G���ǘ���!y��zڴ=ܮ{��cY�D����h�BӞ0��*����ߒ���A[\̈́#,�k]"��::��Q��8�j�D�o�b��Y��l�_�ë�C�����0�l4,|�E�6r��\�y^_�a��Bf�w؞��q+c.3����U���'m{X�y��J��*��|�$ n�Y�w/�T�s׆2'�`��)�8���*��h�P�D:&m֡K':�KHq�ql-q\A�K.Ut��R���K����������.�A�[�����DH�zM��ĶrD7�6�M���է��c���f�~� �-��e�NӨ7�l����[A��S���Պ&|��,�)i��l ��BmJ��b�^��KFD�5�NA�4������'{rf��������
�\��̘����&=��V��Yl�2�쐐������r�#�B�I��LKu��0/AQ�5o�e��X�=�l�F���6^����;(�0���!&6�X�c�ӎ3�bu)[��]c#h��,9,mΪE`C ��&~,�[�����E�&�K�u�k�L�����l�����TV�꽗�(�o�]r�̐�Gy�7Z��[C����KN-¨���v�O�m"�+"�'�������o��9邕�����b)�*�U�tI+�G��9�"���oTvWB Z2�[�HK���d��]c����TU��$�ۺL�U[�m6-§ p����oE����G\���]��s��ã� J�O���gx�f3�X����2�`[�)�e�0��l|o��yo���z[K2s|������<�A1��7���"�_�3�Z�t�$}u�D��I{q���'R�j�U�=~7�0{�6
s�Y}��+Ӈ���R�����ЫD��D�dW��)�	CIqo�.�d���^���V�d��MazW��ĉ`7]W�#1��V~�����1'�,#�V�!��U���t��*I���x�𫏉���X�e����˷�q9&�3���xs$Y���?!��o�0:�q�\9/�]P�2
�*f?�f�!�x�)��&�v8�s1%����el��j&���]5�赪*���E�쳡M�o�����OD�V�t\y-�eE�P�>�ᵑS��V�k[���Zn�b9�L����Ǵ��������`H}^�"���|�6U3FG����נ�@|�R��{�M�gV���_�Ӄp��]t.�
ALM [ՂѨ�vo\�����g���r�3<�����pr�j�.gB�!KN.`��_Eܛ]y��d�_Γr����>����e�W�}��?���TZ屣���*���<:h��~��R˨kj� �o��34���&� �7j�m,-���Z)�M�<R`�W����^aN�#G�v&��O6sA��s����0/��Gp���oW$~�b��l۠�>5̋�����!��paa���i��KF��>QZsuWg�����M���Y�:�e�6��pf����
5��G��mx����o	H�7���v��G���DS	
C!:��%frɍ���܁�"y#�XK���Q��}�)qkz'@����҃W̗�YH�ī�?���y
(�g9f}r-f4�Fl0��<|ޱ�����dS���7&)���ŇY�[��(�s��.�{����mr/��O��&�-�g�)o~'����������{�2�����b�a4�w7J�)C�n�L_�Q�ހ�:��=ua*��x�%S̿�
�9��g����2�F�RGj�*Kz����&�:m-҆���$�� `G�4�%�N�h� �]�f��L̶Z#���5C]���#!X���q��Y�<�Hu���?"��$d�����X�p�US���c��L:*�gz#����L�n��J����Mtkc)'�8 ,?ؓ�'�6�Z�)m��]�a��Ы�D�5�B�N�m�r��_t��c�fkrA�E��g�F4G���4�����}uZc|��t���"o��(&&>x~��15s�-�ה��B�էѼڇ�v�(������lW�?*6T�+S�tB�]ŵϻh��gKH�e���������'� ~��^2�u`�z�9OA9�n�m�^]�ϭ �-�$����V�1��?�W��b�R��� �WԿ�h; ��Cs.�񎉞���N����ǻ};S���d�������
�=Wa���yP��I1�>��<�.�
�����=�����Y�?�?*ǁ��H�i�J��}\Nf������o�J@���@����&��KXE.Gߪcr\�3�]@���n�!��v�v>�T�g㖊>�Z��G�NJm#���
>��.����la��{���U84B��,1"2N�VjOCTSTy�b������֩6��<��l�;3
\C/Wfnj�jlJ�6Nt�q�����o�0Kh�_m��ąU��V�W� A[X�����=)\�pHL.��ܿ@��D]��EhP�#��'�]b�Z��-u�W��Zsj~m�3�m�%���f��B87(�]�.֞'�I��_���?�b<��u� �Ư��IP�چP���I�h(XG��_��/6��� �q��_z��4wC_h�w��9!����j����$M2�Md�h:��;ݬ&�_�W�Z$�����J��B��� z@}��ӠCs8�.Ov3Ny���$u�7%3���x��c졅v��v���fc�+���������WW���T�$���~?.��7�ZW���0�E-u�v_g��[ݧ���Oƶ,�F��ۆ0ݑ� �����p��	�e � �����mk+�fa��7s߇C{ LR��TT\�K��}��(�-ʅyl�0�!�L[1j�����2�W��'o}E!W\x`0���to �u1�=��]��������>������ j:$bY}��w�d��f��	�<Qx���{�,\TۙPn��s��۞N.6>�K;��#��8?_˞B`�̘^>ב����t�^�-�~ڐo��k� 1�J�O��LJ£�#���ZQ�M����jG�C��y� 剃ï�7�}�.)�P�,��/H'�q�4X�n]'�D.���n��Ѥ��h�]�K&����;���G~,�Ϧ��E�A]�X��x����\�����P�i�~���+۰&�ZE.;����O�W�>d��"-�i��&N�I�a�f�P�!�ˍ�j�W87v��u���F��brT�_|7���î����?Vˡ|\4l)��B+ڧ�iԡC
�%c�a�W�y�qKdA�8�/\ ?�z�r%���$�kSU�@&�����������Y��(҃9��U־7'��xi�jQ$���VC�~�6BI��@jk����vE�ZlY�z\ _f�X�1�xH�G@_�qRȢ�WЪCEOY�	��:8`d������T38@����xc��za��o�?D6!��cW�!/�A���7,6�%l�e����\|
��=��\�Og�ׅ_k�$��A�1��|O^���(�M����!BZ���+��}����w�F�No��ns[�h�:V�:HQ�6A5$�%�}����	)��q���O���;І�*��*��dh�X����qQ�iA�dv��&M'��g��9;�Oe�%�
Y߫��.pea�w+l����`n����>.��:�ը��
bJ͏%���;�kn�oP`�v���=u�db��\�6�M@�a�m�,�2l����aj�~���8�f5���a~ĥ���Q���1b��f�2Hq���X�=XJ׃6)�	'����U� �68���e��m:
��0�t͵�8�N�R5տ\Z6�@̒uƹ�Լ
c �
"]�.��^0V�z=��QpK��#�pX�A�wE&���]pb}�X� X�����_"{�=*� e��!Wl��݁v	����g����}���b��]��]�G�r���C9K���Y�<Z�Mۂ�d����ai�/#��_�*0����%=q���쨻y��m�;���il��6r	!��-���^=$�\ ���pw6>i�̣�{jR�*�"fN^�]�#S����p�{��t�2�ס���+=S�<7�775m�8Pd�Խؓ�V�OX�� =�/
)S����L�}�T"/�v��������JE?M��8W�@�W���h��fT�Xj��|\X"�q�������CP�GgS�����X/�j���� �e睭�L�B�.��b%�JX�&����
W�
|*�G<��]�Н֡W�*��+&擳����ML2��e�`�IJB����qAW��&���ܓ���L8y\v��g�K��]�a�F��;۞�����K__!4���r$�m)��9fϴ� �)���7�z	,�?�o��nSS�A�ϔ�ׇ/��Y./�,� �Z44Ƹ.�`k���`|�T}6V�����������t=��� TMs>g���3 o�i�s����9�{1���a�L����b��}}�|�Zf�>	�C���c��;��]�uoow_;��fM��$8O�;Ѐ�d��u(je����7�?|�K4i�-�OO*k��AX�W�e�]9��Y��E�`� ��c��:��B�����ݦE�_�2 s�
�0kw4͈�����"�6
�i�nJsW�&N���J��%���V����%h^�!��5ý�JFI-.(���<��7���r�z�)D�dt���#����،�3�T$&lX�F�#�����bX9?�]";�