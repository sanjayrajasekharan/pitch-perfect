��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q���17���B�I]L��٩{�|���e����F���˅��L~#�|�f�
��������%����U��M`�>StB9N�P���t���H����B�ԊeI�_k:���
Xݤ/��R��B���C�[��U�	��j��~��7.���qy}ov��yJ�r�E�|�H&��k����~��k�@ԺL�!9����S�6y7�Y��s<h<��o�<�(���z>���=3蔫�'~m~d_�i�{c���!�H�	#�i��t�h������F�I�q��޿�m���ՂF���T
Z �R�n���@��$#h�t���S5���<�:(���%s۪��2�s-�I���&pԉeD������4��W锐��-��z4�)^�	7r4[4�����, kJ����F.�gh.�xNݬy�������~x���T�I��aL��`��ï��_��pk��{�b��s��s;�U��+�%fB��[�����'=/B�� ��@�>:*ͭ���#��`��]���9�OξtԱB0u�U�k] �k'�.̌��!���&�[��L�]����F���N�i�:��)a�����1m���_z���qwԀt���	��M#��;)��"�T��Zu�5���'�d_!.:� �x�-�һ��m�i�So�@ �����Qa�" ��b����g|�e��X��ӏ���&����n�U>T<�8fӟ��
h�Q8�����6yX1\�#�g8��I��y��) �^o�Ʀ������2��|��:l�AnސtbF�g~���c����b�N8��p�����z�;i��&f�=�㏠