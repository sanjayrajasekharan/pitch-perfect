-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Hp/tJ9gndSjxl3+fNsNXH4cAncR/wKGAhOY6g6US8WuuzDdQA4INyhObnBHsA3wC
hYcFNYHbmVeTOsJR3kZndsAaQH0xmZs4dnzOywvIc+Eot58GN7stFkUCWp+w337A
4AbaeWlp7yKMRBXNsn46BbFcuGWQGaop43XN1GHhEqA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7984)
`protect data_block
htZ5svqyAKm7TlPV0gSWpuQ0WBhp8QqNf8yXLf1pLOKYv4bDsCtGnYpC50A0fgya
Ni9Uh5aybvuNyfCwiBsBEwRg1dRmcdhcyI/HSHAHKx2KrcylWpj44bz3TyFME8tm
nzvDVYF2nukcLEXxp3CApDz5iNml7y20Za4sHOUQJ7z7ac2u6kzlESC/aDxW0VbF
Go9fWEosONNYdpX9iJmF3Fd5vDcwlg/SPfW6RnwwWJrZ8xhIlxal9eE8z6A0vedH
aWl9mUFp3vgYYzo1EHabg40UnlXKOmhF1Khf+YANsWFxnGSav76zkX+qbvrAel4J
8qlnVlPoWA0nRaIzNDKk2Y01KlMZltDz+2h/bVt+lNFtvGWtbEGNT+4IqncAFqNA
cPdJt7Ztzc3u2J4a/G3N1M64WcPtSIK1p4Q/bZMOOw0hCtrVJTtItYPPjhcFqFyV
jdrVEHHWJqmgeZcDt7Da8ET0g2gqxRLjbvz3ge1fVRDBrZpM5p1rnjBZVRsC5BJL
PUD7zwQ2nq3MzoAw6fHbf3tuqpoVTAZlWvqgqq54tfPxoX4IvPQaqMgyiXqefGVJ
GR9M4anD5a+tcv75dnhJrAvGYNTElOC/zx1HmZF9wIPQakkiRYCyLK/rIkPxwaYn
jJDP4iJLQF3mhnvsRn5MWViwZVqocpIfbmhNOoRPPsLiKODYJGkxhSbuS0Cl8WOl
wMz2LeU5SaaLkiYlYMZY6KWogYWPiNezhtbj4kehhfhhYIrgrPKZ1HgeEy6EBtbw
447m7mVOavOLwnHXRtmk3+GtKdgNQiHtBAD7QvX3y0aF+aaB2Xeta0O++CAsGYI5
KVwiuEu5VJ+FYZL34jHlK0VgMDWLmAWN2uOHWMZY3pL7O8DRZaBdXbt/lagC3zkG
J6fOJTavGqPz4hwLXFwfV32h3gIuJWRO6sghK9+SoLwONteQzM830pWRbgCiVQ+4
EjnByg/P5dz/EtxriFMJw7QNK8JBDoRqf9rZqSReQAk3joJzQafh+TkZkJf2n3wK
5tBL4Q70z/vPYbgwvyEzMTV32ChNOV0svVoJ6QIFi/s7fIfSakR326V18KumtK/F
VmnoEKCkKQFabAJYwZlARs9TVrZ56YM4bu3DdRxSfL9m4lcMSfPHZEU29zLSfYa1
9XuUobkFTQ+GyiknMXlIlcY+Z13n/IqRlwRdlrwVAGX8AVhgAYrRIKUsWUEIykTN
b3eVHig7R76T3e3EPHHw33c0F30T3Y46i3F8uUaN3qdJYBg+3Ma37BkrBcz6sqwh
zgCFhCu/xd9CZBu6xRAGtUMM/40Q9F9uMb7vomyMhERHT03sNdOcnbQo/v+eFoRe
L6PrnST4peRZHD9i4Cc26sTzEIqkrDrB3AXkhu804vu9fQeewc0vAd7w2+2X4fEk
ylg0MIF+VApmjQwpx7bb/bBvvc5nyAwZGFXBAPxtCY8WXN5y6AUkL14OccK585vT
u9G00IuXbKRVDD08YwAdUhFplRlP9ChneZfiAfsRLI1BqzajE1FwkP3qh9k+wY8f
XUqA6+5AVY0KGcnozyo2bsOovprPs0fwop+qIhft4fPUp6pGFgAPpPd5zEVUkpJP
iJwf0Fu3vrKeKAQwkRv34GI+akLzqy3CvAyEtGDCJyGg4oPbHzHjvd6wCk3TLsif
lR7bc8n/utjB0l2gRbu4X84cweF7TqTOqtAMHK8WU9ZLMYVtqbW7dT2SO88kMjvX
pQwCuwZr6RRFJpjQ6piutdzmyZZwnI1sgaSl+GX15+CPae+Uqgmnhq04CTI8nc12
ebbNqEqDSQdZYW9T2nDWgr5ZgZSt7ikE4dTTV6V1UXfLePs1BeBHdGFI2/phG9Ab
a+mKsr7Vmw2AymkmqJmrucxDvW0GLACn90BYWLmW3FBDf1ukvP8hr+E+yZrnzLUT
JMmiN0vlrUKFWSHqYxpu9/2bSII8UW/K2XUvcD/NjkGYb+Fcgwy4GPsSUGyUPBso
kjwObwV7scGHALSENw+nUX4LNkCEy3SfBfoseDFrawEMHXJzPMcwoNTTwToR5wSF
2jAzOgFn8YlaZXA0fYan08bsNZwkBjY2fHp8vQKm3cpSwNFRzwVOqbnt13/UNoTd
axrEg0eXnUIJiaYmIsOzcPf06Fzg28R0/mUWsZMazHeTraS6bHaEd2+RpE2QFVLL
bJ7TtI84vj2CVd/lvHO7j4A8YnrU6+QXKN2HQLHgDX5ZsgyXIwt4UBZiKvFePmzZ
BPZPfJBdhUJ/rUxq9+e9Pt/DNXdLOQGnv3JAkCg0kUXQTqScvJqrwhRlRkkjbO6t
YyKU6Gydu6Kdg9tpLobbWp41etrWj8+8B2jCHlt1U+5iEHCvIAta+NNESWmxdTeL
hFBkkcVx5bm+WydXHMeeT0lrDfVZNtd/jVKEHeUmaveajV7Bo0NYyYOG07tFo8Qs
4Wif9WNVjYjxdxt4+2X7FXsPHzLzfr1uVrBo8igpSqkrDuvJRv2z5KxWwhHGsh9W
lRFPxOUrT8luIMTJ8pWx3QY5OT4BYdVOVx4IUNOP1/3d+7zE6mFL7YVh0sphaJZq
yj6bTkBRI3uI3tWKvc8dE1viZ1L/+CHqtm+7j6QY6+UMTW/bLg0So1LPpJp6SrqR
u1osrmA0VG7dW8FqcpPaogklo8wa3vhdNgqD++p/L/iCQd4akloJIOKruW6CPBK6
/D2ee0RLBotsBVSOQ25LiM4nBpkkdGfu9yzjfZSZawIXOOcxQBS3s9oQc2SW1AQ3
1zELYB1Qg/O9Va5mDB/ST3YYReiO3xgaYTxpbtAKkWFGR5H2vLllsUttjAVFkR/X
BuI1YVT5iydhattLsLJqI2W7DojtJASlUGwDLzk/n61imHXnu3KmFZQ4Tpp3VTJ9
lmppivQwLnTl5Y1u67EdXK5oJc2fn8H5+vL8BDhsMF30tVbuIQVUkJqjRYeeQC+0
dc4S/zpRJLph+Zj7dKG1te26i64WHMDoD6Oddn5E9ZtpNGvQWCwaVvRHCkPGcmmI
VdKqf8p/KioDyTD/96BTtBNd58BYBpQ361WnriRZoVWena/coRhz6olLAcsSPqMr
+/lsrJlwQHgoZqG6D55QnxuGoTKiwQ0dGvBHzgwjbKZckWX44TTT6LEATgQxnayc
Zk5wV+0p9z0UrnF41gl5OHWbyiUUs/ra7+6hQs1uy8kI4qxP0AHLS2xQqin1xq38
pegojCi1uADUJ1RAwmse3zTNaB5094ByafZv7J9X1OQGzUXh9LhA+THvFZGZSEul
54mCEHsq02KPMEQGOiCe3ahIckC5hh2jrb1UDO4OrWzid3S6AMAQiUqecX/t9TZm
j6SZ/2eJ016M5ngv3RPZYLHXQXWZKlxKPNVZuIY+ELWD27gPZlItH246ukS/NOZ6
22DDtvFmtXs0k1abHmqV8ap27umGRiEDr9cqSjG6mJBJ+sOY8705hoNoE1+SDxNL
qTFNNPbwprB64/iaXuAkeP6iPHRZAQX8p10Nz4Wj4Ack7Axe1LaC+DJkyzMDcN7J
hZeZGe9TKM+Fibu8/d9Zt5XpoWxeyei41BDuKfm48/M4XCCiPJZPk5ighXfntNr2
p0acTQufv7+qjixLOOOoOvX6PK9rhWSfBoY3FI3fJNV7pXoB9Gm9I+hoQ55OyWEG
z+ZdEsX/FvGPmBTbDMAVCC7n4ORkxBGmttgtrt/dPZnAtIIghl3GJTNBjmudcnHE
heCNfQc5Qbzdx5H2TNVpXnNZ+zwfT/x9TlzAWn1Uv7hyWDgbPm1GOBa6WhC5Zoc3
IIaMQxMaXYIZHgeQwY0oQV7iOmoQoca2/D+yQwXzCGpeqLPIiR2vJ6hD0xPlY2s5
3sKRu1u0XYWEttV7LWsDqwELS1JQMQ5XuYHIsY5m6WLDRcgCgro/y2XIZNSssG0J
iT7JaukF5O1Y2wxPG/JC8CKd8BUnxcaM39DBCtSAe7Of9JRwLomA2epBjRDHwYG6
piSq/Y+3SYp1INXO2EQSW+oUns9HC56/rtzQIbFqjK5XYQP6pGdcTha5WDPJ2EEa
jhqLSpZsdKJRlPzY24eQr8SNV8ftZI/0WcFWR2n3v9KRD2nmjfDXTi2Gtd08WvaB
cWhr6t54Io1doYVB+1udrfIw8eJWwXweD7zKNVo4FOOERQwzS4tgsmPyfx1LENXn
vRfL4wEgqoqiym3WfWsD+m8MHpbf9ZDQTBzKlYIaqiRDox0Ay7d3tk0jTRlSPDb9
IHIH+lonnmIMD4j+UGnGFRFTNpNFPjnfH0jcDN86zXCnvHqOVyB5PQN91DHsM8ib
oLSe4wjJxx0FnBbzqDlqH9PlepjhAyPlmoYC7kdEZvf+uMh8W7AocV3NdFSuEWXT
fc0io+6Z69096ZaOZmxC+yiFWHi2sVn0QC8pS2AVoUzTuu9ybRBHv3h4AiF6gGFO
mczdOjZUAuWoQpamaO0DRiPwGitPmeKUIZcH5d8+Zu7Ii+HX3D96ryD+Xm1CVqbU
JzGy7U1E7OG3u1XErGD8AcOd4x5D28MJ3xPz3YJ+OF2ULjuG60/eBq6198w4apWq
ZdZF+1gLjDQXuMdIBCsV13BhFCVjjCsvEFsHRiZ+R6Z9e2jZzdiZtqKvEv83erpw
ulSfNhK+chInYP8lw/VO81yhA0YxVDiYC0w4LMcx5IsLqBQNJ07gOuginl80Svfo
eVB7XenLouH0LsZ6XBSBsoXpzXO6dNU5jU2t7XEVreiCOPCreWARaWYDQDuO5v4A
0FnX5uI8Lj8CqhCgombqjOFg1Kyw3yTOjOXv9IXGlZlBQ4FfLzxkg9gWH3msRNk3
3BSeVrr7e2X1vYtRrz5wT7SxVreHfDp9WrriIm8Q0QgnukZFARJRZWlvbhR4HEz4
1QzXv/tmPk4NPNVdFkl8N7OSHPMnIY6PQHy9cY4c5HslbG3JWWtNkT985CjUsP+E
s+oJ/55aCjTXGCyfRw1oed2CX5UEv53tJTtFpoXQinXZJDLR+nSmGwJmvygEF85u
eCyrVs8N4X8dZk4oncMiYhJBKKsFLcCUZhsnfpDdeATWKzU/MTwusN7cZPc/nl4p
PCStTIxqtPXXyNjT/wOv4nTwNgVRz4tT9OU5vfWPKD9WbIq3zf8Qu3hF67uC/cX5
yKKWSlADArklWoj6yeqWyzHdUYc6w3nTrHZfDNLidiE+TY2HQrn9a61cxX4YRIxl
aTJOvL7qPxRBRtgvO3TSBBS+x76NESzuz7iOq1lhUg+Kvx+1FKjjJKdQ7QOFgl5D
wjFltEnX2BZKqsSe89zmw9owUGC93CSHce64TGi7qMa6S3+k11pLb7ixLri0hAme
Krrt1IGGQeg0OAqJkKJTFPNkAyeT318HB7bwKy3jqkEWypkyUhKUSthKhI8ojKEO
bvfOcl6G+o6gqmN0qS73SXsV9hZfa4T45POSX6DOkjbLX+hyXQ7KWUzDvTVptnit
hADh8gdShCW9YEOmZMBpVkl9tO4Vod5tHV6aU3IKokdtn3DKB2q264PM4g1MaGPO
R86mctaMmJafD07bXVP2BShEb8hD4YdaoyIXqMCMW2egVXO0SsBNbx57zQna47dh
7R4nw4pIkv1JglV1WZ3XYbEXdcZQqx5icRCvu0IMRr2xBIN0ZN/zNKEU74akuTJH
08+2fESaU0pTidlUn7CHI7zkbqE8gaTeLeXeDx7xMsn8zgwdM5yzuvRLafPpyEro
5dkAS5QGBtW6ewSYnpuY+jRYN4KBqjxhJyouTkt+6IaLTXaSYrGfez2ekkMau3lB
0AF7k3Kv0AbkpWXYBR09FXkMfUv3BEjxw0cMFBhjPhsvUmGGzlVgZsOhGsOXVKy7
xtZQo6OCje4a9j+0Ki8zqyaisCcrI/YHWD1n19MbAR1bGAXTHvUCxUxuse84JBiv
tc8jfxuJHbIrKwJrH84WFRLR2+HwH3J45Tukr/p+5TVprb1bOnKTmriOKW+HvlZk
PJP2d1B/JRysNbsw5T7ukgMD+kA3DU5TniRpiVpBU2NcGEIwG0W+PZyn/qKMJJPK
oikrD+B8jQdyYTqOILkYmuRs6KHw0k77DnQlXoWOP2VAiA0z80YHrzoG4ho+sYIX
DJL9MgColmYpkf7oACtb1w0E5/8+86vebBzW9F3zhUOY3URSxgzU/qLEG0cYPBLs
Fca7y0Em9ASXf9k4MhtPtqupZ4mkKvAdnHrNI67ddD59xcL8fYws0TY2nKHF+NRI
NvGxO9cYlIWF7+UQDNXEbT/O3F7iVZ/IbIVVpZ6bxLZietkpYxNbbKWIMA1N3CDK
DnmWS2xbqrFzHjGbBB9PyBA5YwJd6VSZA4wVnA/WfmD3Gs1U63D8wZzz/7bnojkL
03ACzT9F0LYtS7G7vNvlJsTBP2k8gTvTj5y3Q1BaVQfB5W0okW5v+V6C5HYNixEI
XO2uz1ZBGGuT3fx9aQaVfSSQkzJOTI1ikIXo09kZBkU1G5CF2uOQCLpboY4qDiDN
/2NRCtTgagr8goLMEiPYbVpsqClKF1Yjl8FJTcHrymZon7qazb++0C7u44v6Ies9
TsWJtdfhkm1QzB9nWohrtWwECEriatVXt6+N5LTLno7K6kH1WXNXkkq8E+qjDPRq
8ORTR27BIPSCvTSTbfVsl2Tz9zg2V916sWdO00E8JC1/xf2yp5sNZJ0h/o9nA0ro
swIR26ytKckHoTrR9ctSKtbq+HsC9DNsHp8WCXUZxBuMKRSDIO0OJanwNGBbmg0K
P2j3zQmGQ09e813pvdT1E6MlV6P7TKAbd+sSW+JzQY2xnMdy2yH97oW6bGvR8b57
x1gn30GGbt7Awh4JSQ1f29AXpn+eUSpgWB7smpyjr5lnwbNOlCTT+3TrKQl0JBEH
P4cT+ZM5ZmAP34CaoyQF1u2VtsgZrbam1cmr5oR8/nwbunKAWRCbWaTADT4JfY0u
xNUt/sySLIdyZODw2mbEekABKqVc5BYP/2ZTRP7GeX/mjR3j7lcaN8Sf1qt5Qohn
jlusZMqQy/C2tj27LZuvzd713pMglUEOLLdeEs4sojimmbYmTLpPmzElE9navtPw
lxLBjrWYZRL9hRXJ7xSuOMgUdvbUe6MvOHbzJoi35QVjpkEUx1PcUPGKPDWnVZNW
j2DHYOUZO9Z/1ChP1fwVss7rozCit4dwirpCjwcxii0W25CsOWgG37+HsWacVoXq
I3RRDm572xeoLaCZwmdOsN0ZB2Kmjl60Y/WKbl/ERxjhd1oK4NYDCHAn1tZhqNri
gpoz2IK4FC41nJeTsWAtneKXxmXtOGf0QLwcJZSciq7/YJgTc5yCThiNvyj/VThh
aMukvjkBmtturkK/2529cQ9MydU+2Ffq58H/QKpfr6XHx4JKVTNXoiBXQh5W0FyM
M1r9MvbtKJFCyLYv7Igmcup8SAQAUUuo5BlUuGqeb9xTgRfTpCLgFUA1hyvAk+z2
pqTO/l5tqv1ay0AXCOtRvYdDP/GyU4aMDHOLsaOiR8roAzKfR4GHn3RubKlg6N+V
sPXxV+zGPUcTyZvvHVYqVWvAm+gHG38U3XEUZ6+QYxRx+eNiSu7wstJyyUc9gAVl
Tqf5XUX1iAa4cTTjo4e8M2NkL2GhLa9k6KNfpN6H/kbdBZm1BLEv9lT0aH9Q58xi
nMpitQWFo0vvGqHnNpCMn9GbHHbm4/9Uf0eCLogc2H9E/sa6EhIal/c1SXCJDy0K
uqMyu2p1TYu7sz5+JWizQKOrf0BRwz6RInIbGbreTBLn2EtadjFotL5ru9JL/qfZ
/WUzPUfQVfgrgSvin+RHbcA6dyeJxQRb9uSSHYkGcduQk3ZSR+LvlwbmgyCHs7nJ
kvKAPJLBQDX3Ion2i3+sJ41GScu9WqzbLrSpcqbXDY+OmoeMUD1Ei8/FyISVcQ9n
gW937+gLE2AwITwyHHld3duGC80bszl/wDpFNu0l/IaPFLjVqeAmDGhRhZfc2dXs
LK1/drq0dorLJ7tJbMxlLwc4XgE7+ud8kHO1J/Li/wMDVUcae1OOYbSCsMplRRPU
mXXJoUOPik8Y8WRcEfzLa7j5O4Iqd6FRA90+dRoGVz985CczLtACQzDU4W9izpaO
/HkEOk6EQj0Kh6lMeeqLCrUCLo4nGcOiGXNVWPdfktrSU+cE1kTsblhj+SpV4syn
6qra3q4m43ygaphaKLwEoy6l/VDj7UrGWawB0lo+SNUM7bIKfALpqbzKDsevka0A
6IvrwlXqYpWwWIYIBGOZp0AiMQNzawmjztmNFBt6V5JugOFXQJnI27kIRwGwZCqZ
3DO45H7onYufb8gg9jj6NUoDxs1kBll6H3Trotule1spiKS55z+R8gUkfTu5ZBt+
+VkeFIq1vvSla9qrjmFKwrCby/9RH7lAAIfa+4RRQLArETjOyuzvz5FWKoS76s++
jwe9YNTYs6cZ/PtzlYXwIr+DV9PSNd5h0bZm7CTQzggHlvAJgglmiMig4x8nlvTP
HiVPYkWXdaJlo9kxbj59sd4C4uxVr9XB+XvEFDB8/zia3Bd1wja83X289GjqiUem
oqvaT30SVTNM2kJD3GpbClhpXurT1HjmHO+A8AmRNjg93Z8QMA+9Vzy7N7A21W4Z
7KkKa54EERJ9a7sX97jGlsLSNFlm7E/l/mVzcmT6hfDcrN0OVk18/HuvyIa93Ls9
DSApDH9jE+pMSeol7KqiR15eKG1KZyLwqukNwZE96K0Xdori77Iz19amWi71LeD3
PiSd7v/adNPIuon1AlPd23dZzVIBi8Y57KAva6FsawYUQ7MF0ZA0oZA7Q9lYZCHa
zQ0iPJFk/b1I2RJ4w/J/W2fGz9AFSpsuEUwxwmL5wHkucDX7eva6KyYyrZVjWIvL
f8J4ZRs/lJ36/NBAa3WOD/qf7RrqB2l+jN2d+ydjPJGrwK/OdaFdB6uKkQNNdop/
0d9zKhZspkDR9KXxySrmHGZAsK3QHR5sbAA1RTIha3aw5x3lib5L1WN522uabU40
N3UOl7VERjJ1TKiA6nB0jUfD/OIwga2p35wp7cdW/DTU7QB2xopfJf946pcdLKUM
GL3yJbrM7WcNkZhzinRKB3C1iU54wbVmHkX0N2Htr2NCsOFhUQQMatdyxECKVVt+
i0kQ/q4ibjLJn3CUgX98I2TW8pFF5G3aSSUPf6o+AHunqfTlVBUzjQ9pS7sPbaTh
loJmy5WMV57Hj7o9lgsdWHwKRYyhWuK/OdgNhAt66MK3ngRC/HnBYXP2orj3Xnqm
7yE/qJplnTt2VHj5Fsv1L2eu+9GPoqgDDJ0Vi3BEKk1fRJ+mUctXapATpdKCmASx
/9kXN2EiqTBc+tlMWJ1ak31OGtTzGwAE2LJtwjR6NmNLoOmC1Hh1skqWQDqIr0rM
YFMoUunSVPJyUyCm8/EeKFhgKkbF3xXF8v9nTO5V9nbT+uV2jJa/Ya+p5ca2Cz8W
6AGaVVIXtwqTpKPE1PfT5m3DnEJY8NvWLkI75fIccW4b4kBG6xMx/gWWXDIDKjop
hMe0CQSUgPl58IeMxy5OfQmFNGoN0t0o8F27JG1ii2jh81VlOoDFx0QrpxMf3GHd
nsU4/uqX0qsW7+WK/gq+Jb78prv1GhK2xD6r5mnt7L9Fv7YfBr8gGur8CW1nv3SG
bPz9SizTcFZrtF56fCQhKRl2xdyDB5wct4QaAGL5TA4T3UfDCZpBTKclHNgQAWnB
iIIPKc3gCVxOQiBf0Z5UNQaJlIyyR0D1WoE7ONxsdFEiyUxhbyQ0FxLDFBo7Guet
kbv8V5Rhda1mt36prveogE3//Y7/ZZwsGNqSAuzEBzHqBRB4PJjku+D3cjBoBccx
UDDU7sbsDK/BK4EEJ+nSenXFIOXVKDkFYVARw5sfbMkW0OAi84dtkL3qmf+UtCrr
XgiidIADSgWkGujAKZ2onokvV4OUOSOnsmznh+DtcLPOa+pKureg9c1saYF/ylPu
/qcXBrxQa03ttVPg4mNnNmDp0AbOE0r2tX++gERMkJgaBXMgNDrHyr+GYC7+BgGp
c6zYbKP5FvVAuZF8WdaxwbRWK/99fKSQiMo85sv936FTzDPFJC4AfyiG5OvXA8xL
ARRKkjFKRDvfQzMGGvv9TFu7dE+21GBpNQOBmUCVWAXizZKVO4jeXUd7Hs03gOkH
d95Cjg9ohYuKO0uptz33Z4cJyKj1aU8xf4lgSeZmvH67eoUgCdwRgv+JAWeh9PWy
AjYFeLtq1ai0Px7FU5z4+GeGDAgPZubDtsbdZYeZ8HfjulrV2EN9/hByIbeoiFQ3
32bBPeJKZXXHEIKbG+/k9Cdndc2A5yJSyJXhAWi9fr0pyJAFoW3Kx0W8lHbS1oKR
JK7OIV5J8nq0XK1M90rEJBM5+MumWT2tcb6tBkhJat02XezCT4leRFM3RCSZLO4P
Nua/1QXSKMeYX3ecbdgloDaqIfMZw1jVCWeISi93wsk2B38MzWk3khg6ytOfbeRw
OIBXbzUXvdImcqaCY+jIibiXGfnhckIUkpY2qjYA8CXfAYLc9CRTeJrY2Wvy+UW+
PXojiG9joOYuDuRYQohhuropUNwsfNPwYkZS0ssz5KvcfzMkt0ixyzdedIwftbIf
+fVWh/g1q903QcBG1Ir3K5SkMAHh3sg0fbpA63psFXIZ6RdfoRcMVd3HTtUbTe5v
KboPsQXe/gbTmzzq/hAbdQ==
`protect end_protected
