// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H@L#+;WB?9T'B@%XN#Y0(TC*KQ/[?5+2X\^ZB$<N]N01->C_CYL2=10  
H#>9:.6L!>VDA>S_>VP#A0:DGB\HNO'>)!<07!*,X*F])8FG36J_\50  
H</[E/BF,@(N.;:KA\T#706]1)^T&&2@7*>G"CKGS-1IA_ZV%,I:U0   
H7CW50)&>O];K(H@VT)Y2-,N-W\^]'>?ZC]V4!KF,&!K*R)$U#A[/?   
H3%AJ_#J!=0&*$RZHQ/S(5FQ?!M.K0P33>@+P4N$JM.>-V07.69MMXP  
`pragma protect encoding=(enctype="uuencode",bytes=7696        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@P!EL/7D0O9F3Q(DP,91+4^E4MO$AK/4!&UU!,!14X\X 
@5E0-+6I>^U"N@K;/?J7M7FO!*W;,C"Q2KPA<SF(L%90 
@*$2"<FN]<3J9L1I2@>0-]GDUON1^U[O_#_V P-&[V*\ 
@S!<=Y'8RPX4U%!)L:CC&D<9L4%)L)&@ZYCJ94#Z78>( 
@\-A9QTHGO_->3)P(C-1KZ^ILQ3^'CR^!X1+:T4QE4*8 
@4A'<Q+(P'U5'H4+,<,)"'P$(YK53]&S]&N@=%@09 W< 
@GA+,LKA>9*ED!Q6HKFAJTCP_ ?&KHGC 2M;X3;&8D!4 
@+ X1OMX3/!CU#0P11A!HIPO =,..N1\3#?=/.I! #6X 
@!E?V@JL1 )Z(G%*ML<)T@B%50E'P\/)=IJVBL'[BK-0 
@F.7(HA:>>M<Q>![JC*^%$'K6P^1QQ5['YDPPI>F"N/\ 
@:W ^ASV/^.UVJILWM+4=7=PQ @LF23L@..NM,9&A)Z, 
@<!?[Z2S87G-8>3VGF"5.1>?4#X_E*?*?Z:2"!H/0?P@ 
@";AVU"Z@)]G2;B$C^&J.;IGD785N<#WE:5ZJX#Y-2$\ 
@8.Y#-!8$E410(C:-\?B/T#SWMG (CWMGS]H^4/:0KT< 
@F/[V+_!>ZF.8Q"YR1A8:4X5<+/R(?=1H3=1/,PY4F$8 
@H'/]^V\YNT(JLI:%[3!2A*[QDR/R2OWW%"6/(8KJ*U8 
@)<Y;ZL<%2Y"P5O 46A.3R27K&QX^3#/]6KHM$G>9Y[\ 
@&S!SJ/D+3 #)P:#G"E=S9&X_91%K5P"OX$""X_+&!KH 
@UXG9=\!GP25%1ML=^V(BBN9SE:)TP)HW[&F8#3F=D>8 
@O=+6@CGC)B=[MOL]SL^"J0Z/WS(1PMB? 2\^ZD%+!)< 
@],('SW*8&B#8I$/PKL+5U$D.*>&;A [=EX%'BQDI6_0 
@G]JU*_4>7'X#H4)9'M"FU9^/T--AR087$"(TS3]&3Q8 
@'6>MICVD@NS  +0Y3=,4-EV<',C4W&/1P5UP,OU^R-@ 
@QBO_/>47;!*)19L@-@B4G]6K"M#SX-[ZCWZ'.7G[M1T 
@4,R5*VK\NF[%+U3?"3R4WB\AI4$+?<V?*O7LIX= V-@ 
@M%)&S-L0)$RG!Q,^=R46U5S;]^X.[P<+\EGHS/NQ9LP 
@@:UUR=.^8[Q;1K3QJR@@UA)'^I_X_G0!!@I$,N=>_V( 
@GVRRU-:3(#WGFC8S__TC#'C>WMS_T_L&"UXU>;D86DH 
@RT^K7)]-/M^2*76771PQJ@;C[[<"YZB\.VK?+C"[\;( 
@$,>Y.2P9B#:>(,4.KCN9=PH'5'GG8O8[F&OC2R8H$5D 
@)$>F;(>DLG>0&EJ\Q<G1[CW95V*6B5$R$R]1?!P1?'P 
@PJ-/F8&@?KR -%33FR][^Z;0W11 >-9,='(VKEPX-(< 
@5N>F8J8*&!3#3P^=[V?RP(H=TPG6"Z7RTK7+98?A@>L 
@0O=, :6FCPH@=XQ(5'%)P=[)00YT9!GEY#BXXKM10%L 
@-WPR,$4TGB$2#7HRDLQ]VW5-::K/3-@<##]3=0PEJMT 
@CKKR%RE(Q#&R5>9=T1X6PO(UF)UH&BRNUL:+#R]F*L$ 
@9]VPLN; S^/^!FJ-<C3L',F 7G&0G5\YCS,YW% .;J$ 
@O5*L1UL%F<,*Q8N0+PX/=I%7/K1I:#SKGPUP[G3.\N4 
@@*(T5,8Y/)=-KX%L>VC2/YDK-#CNMR[]2EIR'ZISH#X 
@FU OGDE25H]N9N$N>73Z,(<PV3:^+ R?3&JZZW]-R(( 
@:ZNJ*VN8PTF?P@#>JC$;[-EQ@$^#5<<.D0CI4Q8*#$H 
@/99SD)?C7=+!_V,7E=DV0!9<.%6N 3B3B))_$K9 9BT 
@5<G(NPKF#%(.S)#L0W1A(JVP3HH+^^7,[92?:/_M;?0 
@?H2]+A[2$O<ZY+T^K33<TVRTX#EK0LCBK;$Q(F1@$10 
@[6"TWUM#&';,ZZO*2&@I^6_L/ L &(R Q*Q?*?9G(%L 
@4_BKB]B9F^BZ57$-[5UWHU2>-!82N.H0Z".8#?DHEOX 
@>WU\OUISNIY2%' &.Y^7V%O);=IAP24W6+ZKF3+JW!( 
@J[9450R+DPK@2XBXWV\I;N;:-_C>_A4*+D;"N0UMC:  
@']G4K#5X.3*L3CA#_O*1PHJHL$O<4?4#E!99@497P", 
@GH9)O\2C+JO4(J^M]Y7*+\N\UZ .QE&P1[ UX9>)_F, 
@6V7G 5P'+5&5W[,H<R *76OD2F+K5M3^&+KG9D?)<SD 
@]/!6GHE.?\;SWT&'(S7S,;+FI%RJRL$J#MG( 6T%2&T 
@2)'29Q4?B?C0YC>2H!.!%6I#BO=GMB$15'/Q"=)+<(P 
@L4#FD.*J1Z:/:P#V)5E^X+47S!1&Z5MJTK80F8B5%40 
@8PRW_ C7LTX,;#WS# ?3-+TQ9\ 0]P6 +ZD5;B";^S( 
@,NN&LT\NY&PIS'X_U)_P!^D8M!.XH(^#^5&I7S!XH$L 
@3.OZ\D7@_3<QJ<!5 &4V!+CQBDNIF&F5.[M-'C[I)0@ 
@L!7*KP\Y*=O#PI*?URG&CR2<N.F4MYS5\#]A)U>I?&X 
@"?(O$FLV>]#2,+BP"4' ?B>T?6]Q]Z/MAM#SEL$C,38 
@&T/6H2>::S(]U4;2VNA#/L)\;$$2<*K F3\H_].1J"H 
@"NV)GH@S_:P?G!IAL_,YD1O;^48E'!QE.">B*R@JMU( 
@U'N>LPU+X@PA'*F"JGAR9Q7F KQ3KS1V,\ZY:QIRQ8, 
@2:/_F59'GX+=H>E5(#C8#?:'7)>*>0[*/D1Z(*GV0T8 
@]X%C[)((HB;B?UA'>5/\% L+-H^YT1GR_%$F$[%>&L, 
@UG;N[1A6%.!H!6#M\[O/LE$"A(&7EA,_ONP\O\"9 40 
@0:FHG2&$KLB\=G%&4=IHJ8:[>E:LT(?>E9&%IL56T*T 
@<0OV7EDQ_ 7Y>K%T_55Q^%-P)0D3XJ%A3Y1 B3]O,-8 
@0N!['H @2H<F,A<HO-5>V9&U+:[+JK[9!'4\EF8=:P$ 
@S0EN:V0HYY_[9LBJTUT"Q?L=A(BCA=.M;P,].\18Q&H 
@S!:WX8^6O]L:/E^B!9&=(<*.A7,EG^'/QA9IAXU5 N  
@XF==XBOL*IL^D,,FK8(Z:(/0AM3I50<5-Y4:>";6$R8 
@_[4N;)\H#D%*XP#9Y-L>-?,J7Y&J7(#,8'\?,J::EJ  
@]V) N99/!P/+P3'1YM"#4:Y-%/FL&2ES9"$9C=!OL;, 
@8O!/E1(CA2YC79T$F,[EM>A@,0'SNZ,P;."! [?N/'T 
@; IA)?O\?E$4U:##0^ 5YT\;(DT)>JTL[X3B0]4@SM$ 
@OO'RR6V!R+V<D&Q5]>/C;J%%&>A[-0N @?-\68O?ZI  
@E7K[!6S-QQUTX3&97Y4;2 R_]EOJ\E1G;JF#[$ +7H, 
@[GOX4Q6C@JT7]! VMZ:W0U<J3*^R%=([Z.7*?I'E,\H 
@Z>#$H)/>T);&!^7UFO.&:E#%JNB75_D!?1%Y8$,=!>P 
@N 63*5Q)KNXH&/J5MX+&!Q$VID[GX_R<_"YUHP["8$P 
@#EK7T1<.W+@&T>'DE-/GOHCUE.0+QA4VSBR5"ZA0PX@ 
@KJ.Y,1=Y\X+]:9-%,A-M6-S!26\TZGO$:CV!H V'3XD 
@'K+\P&8'#V6 J?0HWNG:7QJ;Y[N,DUX.?(Q8:'9GV4$ 
@G5!)F<Z9R]-E;'QYL,=US5PO\0L+U-'X6468MALG(:< 
@2QPV:':E!=?SZ+P*]LM>],!0B0]U=]M-A[X.XOY]]9X 
@E!3YPZKH]35>_7>;6&][3</F6Y6'IVADL(1QA! P:*< 
@\X4I9J;458"CF??KV&OZ2EV0I<NZ<GD6..%#\"%7>U8 
@E13./%AW-N39OA!7I#*7OFM;) :!GL!R3OPY#E_%.EH 
@]KR, F:H;"#['65J<Q\&:#]^EK5IKD:9G7<LE@S[_(, 
@U6S @#,WATX64CR+MS-T$ZL5V([=*,:R\Y1(5Y[$4.0 
@;$"W4H^K-C38B, 66-*UBA"Q,@-0]'DJ?@'Q7 ]>[KL 
@QUT7WL>+S>?J[^?2_)2X75QAX_3VO+ZV_S.T21-ZPNT 
@1]]75P5$*G<>FS@--_DI,[4LUM0<@#[FPPEK8FJ#Y6  
@)2<$<2)1,!=D\E7+ZQ/9 T'+^*21>,M)6OD!5LOY3"T 
@F2A:+6UB]L*?H0"0U(U./BO52/BH8XP(:FZ\J"S/L14 
@3#PHNA[2;Q<$%E=#2AB3B1$) IR>#Z;T6$@ &=3M"^, 
@%\?F]S+ V57&/O8CLA$']YO\8!AXD^\:&SI1VK(!6O$ 
@ICC&O=7#YX_?P:#?*M3]*,<Z@B6\7H%\7[R%A_8QOR\ 
@N0UGAVK*!<W(MX>R69_BCGI=J5 -R9DA\=87'R_G1S@ 
@%)92!KM"PX_K=WU!Q A(0N=5KKY[2]J^9S2,6\/',+( 
@XX(D9$Q-Q8T:!J'0\X),U1BP,K.08PE6X7PSWOD*&[@ 
@"!)2AT5$BI,@')NQ?D.I:>MT-1&MK7$IHIKC-CN&H;L 
@3Z9+0L1R9Z RL!8R69 <J3MXS/A[D$S9_/GQ%EV.>?@ 
@U FI*GXG1.)$8W(&_-@=F&W1R5Z(B-@Q3HK<#OY>X)D 
@CX'6]\QF4_TZ3;*=('7;>ODY Y2Z.2$$^( WX>W[T&( 
@[ML.8""O/T2H3P U PG%5@+&_.A3IG/H#.5F0 !/<:P 
@*$D^*(DS2L +S-9*8YG(162,Y]J*[W^2*6C@M3=\X*@ 
@@VJBWQ\X A,H]!].M1Z))\I':08)\J_.4[.TO; 1\SP 
@2MN.^Z( _-\&O!1@"3Q7Z#@7-#K++B;58 &C:L!VV+D 
@]?V7NFF029F!UL\:&18+(^%E[!R4KK%(2]U&[,5A+F@ 
@Q.D6N*6.'RR\"<#;DR(/"S6;Q(>')8UMHT)QZG4(_AL 
@W[]=PK78K]7SE<"T<+22X*W]$9FX\LA@Y0(WC!W7$R8 
@=M[1X(&IL"P).#-:S'H>B:N"WJZ^#A_^I%1H*?0+@ET 
@=&_?%XO9Z\!"KX8@S -[:09QR>&#*W_ZUF+ !D;- AP 
@@'R1\*+;UZ"8(E.(>MH$^JL+U,=+!L. QO,D<C&DV>  
@X5#,_<Q";([Z^*:H5;AU'&N?B,1<EZ_\^=Z1#C*' 28 
@YM4V&.AQ [2%$1SUV4XAMY#VD ^+P.#L0/L:9Q03^*$ 
@!IJ3"XENP8)[RKPE*D"/_CCN::LNE0NR#<]<!^H<--\ 
@(R7^T*J'UYDI$G=;@^[E>8PR+DZ%V_D+)B%GL;I8#Y8 
@-LUMCAR^2!/ .'KK,UF@F:QZI5&^HX1PPQO+ES&Y+LL 
@TUL)BL)'-P44+@[1(,J:P+08=V2^:V7>9:R,5L<RU!T 
@V?AJY&SY)>T.?/AUW *499^8"U6*;^RXD9MZW"L^R.L 
@ALR%O';&;GZMN0D^KJ10IW))?#[]'^6^J5 HJC #D=P 
@HLWD'/"463S9V'^%84L=-!9'!;N\BN7+6A_"J[Z+""( 
@T7:%6SH*K88$?>/8:W>T4^ @MSH4O5HT\A^!S7D,\0@ 
@D\&.:CB3$,:JR-C@5!#%AOX_2S%?D-!!HJF0':3#RMP 
@YX[. 1D4@!J/'"*>7)D);G2-CC8E8D(,+@VAG30CHV8 
@((I(F?BQU/)%5Z 2:@JD0.0P7%_-(39I$LS;]\U2&[D 
@!ZBC&]A*I6M8F0WDHG*+BLPC0#EVVD.6LEDK"03D<>  
@'T38S&-_(S,5F!E@67&C_R3G6-0]#.V/GG( .+R>LJ\ 
@3S_EXTCZ]'O:2U+,>;'>FVE90E(9#CSFSPGY  ?2QLX 
@98$7:]L=J9S*6YZY$V,'#^J#Z^=8D5<8 _ML47!J%P4 
@,CYJ6#A2!Q"8'LLGUB,6OBR3/XP>HT]<CI.4H LLVN8 
@\2PSO$DTPD55-9)LO<5MT&JO=16#T4%0(QCC*>KV/0D 
@QP&85^=J8X>6R66S_4$QN:\.%G\P@T"[VVIXA39OE;$ 
@A(7F--F<>.?:C73MBE_J#+*,-E@]H7_LF*"U=J^5MQ4 
@+6$3>NO-$<J>Z=1&<]KGX71H/AF0J"^X499?BTJ,'"\ 
@Q4D44]/9RA0^H2'F4Y5)3!.S;6H&MW-=<&>LS:'+@XX 
@H=<>B#V69_61PZW4DW&Z,DR2UB$^9^G=_5DK)7L]&-  
@\_W:?1P*T\P'37FT%;CGP_^P8#J5% A=D "=6G;B278 
@';1=US6(),LHL9507892N8%(?SE%6"L!F7/.M)DZ"V  
@::Q%Y>?/3V4IJ/%"ZAU0SJZZD&&-VT65<,3O3'7=;V4 
@I#Y];ZP%YI%=F,Z_/@+BBKH>K(JV>"/5!4[97DVC2R@ 
@)+6RT'&8A0W#EFV)5*I&A,K!__GU*)^"H!AB)%KG6TH 
@K67,9A,:;LM+7+CEKA,FS1B_9JG:=!OZ,<!2OQGPU8< 
@>N1#-D%=F=1+-NKKUB7!!DNDJCFV 8AWHYO6\V75RXP 
@Q;W?9JBWDGC)\=FKNW&\<M4F;/)KE&V;)"HX[ZBS /D 
@IM*'.<I:%14J,UW+[MY7"QJEQ;MZK'H*@2,:E0]S9\P 
@,IO[9:! 2NJ$>:X-+M+W-#?]#(\^3]T@Y[W3DK+M1D$ 
@\%95YXR?'^&,'J.>> 08@K]FT]?H-_B=#CD<-1M:(-T 
@-"I]C5OX>NZ#L:YGQ8)?2189@ D0.S*>^5V!76@_L?P 
@,%HI=2&C:)"<W])Y\3G2=?YU_/I_'L)Y<??"3R2;2!@ 
@$BT@/BB ]@8X;)"I_-U!Z'JBZ-\(T![+.75_@[.Z#]8 
@AU>6GX)%>BP1Z6*8#,8$&([=P2Z!1/IP@91,BU=&J3( 
@W06"C8&7_0C1!^7)M)ER"[!^U#V(PD1ICZH&/'@+7Y4 
@K&4^7FYAWU2OI= UT<UN%P**F QC?#'9;7&>493.:T$ 
@#BX5ZEW<%:K_XA%Y&Y?"GIWRI*C$OU8^0BLO)LJWYQH 
@'/WW.#FA>)(+]"'AA,7ZJZ9+"+?VRYYU4,*G%@A?Z=\ 
@IZTU6"\4:^HLX;E,\A#G)T@:2/?EO7;N36?4YA%-;OX 
@UU2@3Y#K<E:4305P>+IUFDMO&'@[F_<"_"P7(JQA9YT 
@#).'<OB"@(TD<0@6,Z,<2=?^WJ8LWYE,59UK6\8Z3 H 
@0?<%//B7WQ'-<<1UA&D7-6APAX:E:YE<6<P=_89X,$0 
@I4,429L?:AF^HK'HY\;QT*J)5R)]WO4#/D7](95]\B\ 
@)^Y<;86[V 1![,\(V",XCZ2;R"ZC*C1BOSH\L+MX4[8 
@<TP@MQ!9'V.:FUVH;>E>=WO0EX@[U<MS^XP=F.FON38 
@?B;VE<';'@N-]/Y/?2&$H527E&&W?'\6,(%K_BX]P2@ 
@X[DS52B-[0X;J!T#NZ"!95= 10TMYK:2^?"ZG8:GC64 
@'WJC(B<1)^V["<6WCI$5BL@ME)XI7+=K[H0/R@1&K+P 
@-$O?4Y[D9V\S,)6@@C@G[84NS>-L/.?TI)WJU0+?K8D 
@!*/'6YF,EX[U/'Z].8L>Z-#D&5*FJ.MY.T5.AC\;,7( 
@" RD1&8"Q0SRKUJV:']&GM&M6H!J'^]X3UJ%'\*TDI\ 
@Z2_12K4,H63A1%I2+:'"UM@RV9((#2"\)\][O(E&XMH 
@Z%(MHA?WO+)<34?6T@0RWD2CDCXN)WVLT% Y]>2O,!  
@Y3_Z5J.?MWF9]BO'FX-H;*!^9G2-O@RU/UQ!M+[[H%H 
@,3L@;B''2M5BB,)_Z,T553."DE\^#O,[UEU)M11;#6T 
@SBOED#'VN-#'*6R'KL@='/LQZ><-Z(U.@X9V7L^M*%< 
@\^B:TEDZQ$%7E!K,DLY'\D!6-BV%T2<%UZ9VMXF!/^4 
@U98N(4FT]%"7H%TZHR+A^Z:UO&/4(^$#34*$3]O!J H 
@CHGZK6AZDQ'28HV7AQ"B[%[O>+3J8"/[M;;B $_C5?, 
@4IBU/3M:(WBQ]FF&"X'OR.W_6N@0V;U^I-4]=8 7S2( 
@_K'?W$I/X^__S1XIS/IK9%1L-3=?OEM]$O/^+YLY9HH 
@(/Z)//1B2.^]=LG4+GETV1*A<)B'K5:N] Y?ZTO6%6T 
@O301T+C#C0^+AXH3Y"F('IT'M6:%81T92K#W+K8HV*, 
@A9^:,/J\ A=I!NF-)X[*78'*>3OS)L"3:7H%MB6*]JP 
@@&V21;O/L"7WR"=E4F>7+O_Z0#G?+:OG@ L#UB4^7<@ 
@^;LI,47X-R$OFX9CI/F>$;%7M=90+9NQ2[T6^*1Z=-4 
@1%BX_]J2J+:$09=4\F$E2+9!T?JCDVAOEPND/<:0=D8 
@-])AADY+2TOO)*))Q1YH)/5P0?<T_@8G7)RN5_FW_H@ 
@IS0NJK&XUDI7F($/VPN8D,<#(',G-_E>[U(_\%PA,?D 
@#4'GO$<X99;+GOUOT.9W#<44NO?IX;7.TF=8DBG"OVT 
@B/I=P4AAQ=#K+$?,[.&.X5R0SC%8-\&A(@BDY#T ^[T 
@IJ8WB!QG,;+(/]3DI^9:M7*\2:2\-0%/3' .>;MQT4@ 
@K=$+F;]"O#H-T3/,&)K_J\BE[J&]<= +$&5UPC@3Y9< 
@8RS!SUSOU*9=!8%E5KSW!:L83)_NEEHVNO0B\6UTF(X 
@$;?_D)'^?/<FH/\3CD9I +"X7VK/K<2$)V3I1AHSA;8 
@1Q5$RK@*L(!%7:$1[^F]96=C"RV/PME CDJ"5P'(V(( 
@UOK1/J_F%DXGMJ&^<P\Y :A:BHN;%!.!=?M1_S(0TJ$ 
@LU_G6X+NK.AUX-6U!&Z$_;T^HD?%4ML$T1E7HD<.?%8 
@U"9HBU0^,=J<J"Y_,#_$PG,8J4DZ>JB=+.ZH!]HM9:0 
@A",U:A^C[9?G!5M4*1XNXY>%';:YUPA.;<Q^4*('IF$ 
@:FO<3#\PJF6>?M1GI^Q1"<MP3Z@LB& GGVRJR$.N;L$ 
@>B_WI]6%">L;@[?(E_'UP]):]5/L-C3YAY-P'#HHEI8 
@^;AX0IFO<\3@SCQV\S\[$3)#14LP(^V-!,S5F--3NF$ 
@]-LX8$J2 G6M,'0/#T(!ZU*)CZM8!'^F6)01/(6"^QX 
@D=;EV5:2=1FL9?4RG$ 54AR6PZJC_/$& A&,$I^XZ(  
@F1;W4OIN"3\M4[7MNF'#MJG&A"Y?#YWIC?Q]:0AR+8\ 
@-!Z%/&D+R;<FVW(,<%("F5K\%NG\FD[LEV^'ZN#FX7  
@_1%F:Y>&.'J>.6L-OL@\85^?=*#7\!"U\)DW0TK(7)4 
@::A>0<)R_VNE$;FA.U';7"^:V5:.Z\#Q-E/ 3I=4XT8 
@ $PN20VW9;<2:C-R'>IOJCEE&28E,)KQ171QV?G_1)0 
@6P '%<LI7T27LPDQVT[\6(;HXN69C&SJ>M,92T0@N64 
@$('G6['R5Q:A3Q$8 Z2+1T/;I;M"B @IUJ8P<W,Q6/  
@H!;KF/V&1[>TQ;[5HL&$[[)0[XO.]A??"NRVB;PIC3X 
@T+A[-.RXIC'5:]5VSC MH-T\H]%-JT] RE"[ZIO=(*0 
@5(R,<:(G5!G+7@3+HJN+&&9[&J "A<O>F2F<%'IE.U@ 
@7)]KI$+BJ-)+#44MA@RMTHN9?ANC%2=GTM%V:!%D$H0 
@^1ICCCY#A<U?;&3%*R.?$NP @5*7*JZJ(0$^"Z1#3@( 
@]"<B.:A:Q87-YS2E<D,SZ^8?\YGW4^:KZ;S6;S&TT=H 
@N(KH/@^ 44*G"C'3N-F#:6[-_L5P]JYUO')'<4P!$^, 
@5Y"H :35N<-26"\T*9%4?AZI3T LC>\0G6[[$]A%I_@ 
@L"@AYAM/1O<E=N#F!IE+0BFQ4_-)&T3P/0#9ZVEEY!< 
@DCZ>7I7)K[L>DJ8R=8EF!SUN SH=3,CO$?V^O!?$7>, 
@'/MHWLPDDX6_<V=V&!H'CU]PC6I4SJF2^XAOE71AA9X 
@/!554W:;XLCAX,XG5O\S_]43:2[\()9GX995//K_ZL8 
@,<6FJ4"FZU.G[93EE?X#@JG$4N<T:*QF>UIQ+Q(M+JT 
@%E7^&F)_7A%'Y"<CWH@\7 )@!+#AB^-5EWX/BCL-#10 
@?0_U(^"_OC!1O<^IL^SAJ26QT7PKS@B<3V^S266_#N8 
@@1 ==71TJQ34MH;P9ONP@P&\ZMWOD/B\P[3-G!GW5Z8 
@$3I[NKLU8W9-7-494,%^$0D^HA>@-0GQ< *.?&!L+SD 
@$WI^LO[>:5O/=$$/Q)E&GG3)7IY*/B"6@5)(G7H3^_X 
@+1>G7C3#NA3Y^]+ /7/$ELS905R;23/39J4$T5K%X80 
@PP>+U^L,A)YF)/VMFCNS5Q$-,GP/A$_YT?,2':;EEL< 
@$NLM*B]0C6%Z^;Y]""F5^N_#*:$7![:=ULGC4R"&<]D 
@"/.@";K_"Q58)UB<!,S<9:(D\?V8$;]\F^-"&A?AFG\ 
@6^J<!R_'I%N^(PDBDTJ=DS"SL*U J+C#[\H?6I7;T60 
@!1UJEJ_6X?OWVXNGT!Q[X[X]1Z9<>^8,+'2>>,'2NQ  
@X?4"O[9:P=I<C>XEP5#@-%+:05T_GF,MG,=GY*]T)!L 
@^)K-FN/_,@_T<L)W<_0#K95S^8@QTZ_F,3(R?D!24TL 
@[D*@WHPC.00,_;?@F632=+Q_Y14"CUU4?$F4$5W#FOL 
@P(L)]I/.:P<T=_\L"0^3B12/,MRL<)ZI#OR]_Y!3$38 
0GKA?^XN3NEX+L7-@%95R<@  
`pragma protect end_protected
