-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Y2QwafDRw7SA/sIv6Vg47fQOhd+lc5O5mIqfkDn1BAH2xZ7SLKPnr+Cv+ig487gU
aQ1re12F/d8IKBwUo8c3WoFayOLfKI+4Sabr0jgkAF05zHJ5D1KmEv3CGElz4m5G
Mzgud2C6D447yGyeqLrLvtlan9QOQ+SEpNAuuZz4PP9iBxovIv6xYg==
--pragma protect end_key_block
--pragma protect digest_block
fPFwi88h0AJDHV4R/s9XV8GvFJQ=
--pragma protect end_digest_block
--pragma protect data_block
YRzv9wQMyBYL5dI3LBqv3CwTej4UeWoqQ2f46vnmEGqJZ5c+XcOYg27kTM29uE5u
EBHT3HiU0jufemi+U5gEBk/VzNc3dvJBCH4OY7YHTGmNN2xWurlwyYAN/OVLshOn
jkcKMgP1ptemXsidFNRASdb3oLkr0vBFlunHPIH3p5AEVK5CMbU1VNC+G4zBVBPD
sT2zP7ib3jETjXC9K1OH2wVYK9BCM7Qa2q0KzhfTETh7apXogAbSZgHP5cCwgdtB
bqs+ahyq3GuUWFrTUAUti5oyd3HgfJOz90MrUukCuaQVqbwY2N+mSY1env1OuZDz
yDv/0M08csVJH/qoXMy+9liYKgyzJSm/4pik1Qz7/8A2jsQkUP4VoE2k/U3u5IoR
m2KD7xPPJxOsezwiMZZ7UzlWZZCgb160TVP3r4A9DlGIQMrmjT8e8MTKC1SCMEN1
PtwsMWdTJ+91E9VT2St40kZYEGkT8BtFjGFZbshMGKKCKzvXYzHYwAp4UqNkIAmK
HpjakIRucHux4o/hvqcaQyFPJ0QCi3LY9/1+BT5r+MC5GH70HbYazWimSvVTxSjT
AQulm/qKiHGenOBRRcWOVyqjP2mzeIz5joHyVtWRITjnL241zSkBVj2YHrQymDgU
A3p7Hy6ghnsrVN/7HowVW5+aCojZsUr3rCcUYkSDl/F0RLCHhV4a2WMwaC2Lu/sH
7Hi/gjBIrLC+M5XkrdtJRZkJrr4ZYxiKbj5wuR6ii1wCJduv/ZTuxwAXznNgQJOy
jgq7KQhU1cLqUN2Rb6PbUMbIp8KlbyUPBy2CmyCbLpsKsQq/+GH2ISHW+eqD1KNc
UIDwrfvLIGUAH8j24ZQkcu1dgQ8jG7w59lEE+SapyyihlUb1InCqR04mhJCysMT8
RVptfBk6gGWA/G/KWio3+/usbB8SL39rAJEtdOEWCnLIR/rBdAsvdtiAatkQsLoc
eh3f5FKfrvd2cBAwsjLyF9WzvXBz2GE15nQFlhd/G7LoOuRzX8B995hBeZxRKDw9
fyHyIycCmG4KDri/207VHY71sN5WdrpJJ6pxD757gj9I3T6Q8V7mj4bjc3NZIN1u
c8VO5qX1kponNailaAxfoC8sNMZ4OV/Ez3F66VAyXW25Y+pdQgeVspxJNqv6S5C3
GUjqcXIsoHFpio4puAnazvSvHETOC2NETdaW7zthny1WE9W6QsbyQTGEGGQC+Ybm
kjj9XbNhRzbzHYGV7Lt34Gwg26/YQUQnAnwjk0icizKQT6q6s9SZD5wzU/k4FcdF
EqWO9aYpPEGr8KPkTry+Z4kKBZURKiog+N9PdSgjRLPMhp8QiLrLSI0BM+d69vTS
XGeCULmdSrhkbn622vOARKePO6gGGeBtE5YkFCKuBC0hCcj6pssfilyMRChU7Igw
irTz1gDisRHQlEP7MkZdbhKEvICNjy6bL9bMTPA/QGV2pnJ3j6Q5EA+KSYHD+TPC
bg8VKm8U0/86ra5l5ZWArdQS+FH+/6bbuqCdZXKTlylHpCUp8tQMJbeuCYVMhck+
QXaK0TNfrvc/ZnwrxmzTONrilfv+sN2yGB0w5iFXoTGPeJsd3HyHoZaslXz9RuVc
n3TE/cHFpMbkhUuqBpUO3ZxuytSU3VYFl7OgGUzbIhUzPibSZk+clEWb7XKWgzF9
e3nnuELpjeLZrJm5sxxtr3GSnHBplDNwL6B1Nrsc7awakyq8x7R84jsrRkqBPDch
kS64wHELtD29Z3M7HMxZbYZpcnpTQsjIA8uTbTQF9AkJEgh9PAruYlB7aU7Q1oCU
m7Ojsr8Gmq4aYzTwyQ7k0xm18GFGIx7KxmxF9E/9ShtKDdt58VmnmDKBz3WRCwTv
KJb0OEE+zPpguked3OxylCpHaYTsXezYvZp82JuR40/coTA5gyAIvDp8M9rpwGGm
TbC/5/0Z3YE+RsFAdFUgPqztgOIZe+P4La2gmiigIYiFkyMdkErOq0baQJ1tljnV
r8Lcd4YyX2zDJP+PU4nHpN3WOzCvNsmjSPpEMe3J90AmHQdGjZ/3uRSoVoe9KGIB
T24lWmbqayBNMvAzJE4uWInaDjqN01CnVTiLTXzg3zJfEa8T2p2fxoi0Doaxa+7p
uTVvI7+UejGLOjbTTrUfo9au2UOFFNGbteBo3ksV+oSOC/oomhry2mhG5iBoxdE5
Rtar/Vy5GEsFFIBm3U8qRQur8CHGkZr2ouanF0XmS4W5M8ds9XT6n4kvvPyAYo43
l4n5nzIzyTiq98xhdpOKifj9q2B5R4+ry5ewUhk8t5+VDerR2KrbKiTa6y+sUwgS
yR+tmaL2rHDiUNvYNR0ecToZ/khEB9ii83OWpdEFW+1MCa7SzIIPOIslwSlXhiv1
5CTqKiz4v+/7nJiDK5VAf3xs67VMJdQXcaBVZvN1Q6Q7xExel/xgLGBBt7+29ORN
hMChLNx1YNJ2uiUTk45XnjyTi2y3keCDV2XIYqts41nL+BWF2Q32Yew+nWDf1i8F
FCbuMdyP+plHvjUsQJDXbURyrnAhNF6LIeYW/6eG609LKDE5ZhkGu9FNIuDRwoG8
LeH3kgrQuJDOI30nBw7ejeIwK39Md099z3o44xpJNVg1h4Eyjx9PJaVbi08aPAEV
Zi2JKymDENkDAzV3RCk8AXz9wTIACgul0qDTUx4j2tPplJwMsMvmybA1kqmfW5f5
UArCjmNcOJwrGzs/EKvEgblX/Tms21ZgLZH8dNaXj8GchBvgkVpahDoCebeZ0Mp6
17ItZEwcgJJj7XcTvh2FoPuBbHF61lvBqaVRPd0r6XlLxp55Q77mfrsloCSfzuTr
2kAzdQfdNN+CcROT89a78MPbVlWITpFk6Jl6QkE8ojv2APc9aezRWd5xpYOFkq2h
sAexJ1MB/D315j5uUN8EHmsj4m9uyOvsDlsV5yYvbgi77r7zTzX6/BHGZ1Zl4d/Z
5Z4PPYBGDZ1q+/bc209Lv1PgmrSUP0B5KEndqftyIo/3uw7EH7Ynj8CLMejr5xfX
2iBSUh43n8q5I7YLkw5SpKOonXObCG8daBH5qKmLu1iyCEJFVNJNZYjp/X63/kEV
aUb5HPB0fdDR31U03Lmq2fjIKXG1/eERrq+oDhVA7fwhIeNKRRSFURh/rHiM32BB
e3EqBiOMcqY0lCUdOqLlQzJH9tn7smYQbmZmB/+/+1rGRxvRyjwc5olaMe4N7t8d
mxxTKbVJhd6Wr9M+qUkZsiJzg2urlSXypWOBN3HNzjkr1JiZ7Ezu4i75MI7FRX/j
GCbrO0P/7eUaG4iAF9GnSizlvM94Dmn8GHuHr1u1fg4g1h2NXeEtBaalMo1PmEFx
ZLNVwCcrjuVCCz96qAzKLkg/7RNWOo4BXZlQVoeBqlNiDHhv6fbsYmNHgihxGTYW
ROkdvQaSBO3nTPXfoxouJs6frZ7goWw/APjg1yfloK+JPdHPxhhN5/1ydFwSWIhm
E8fZ2sJR73EQiIFcMow4tp8on2UOKYV/5r0OJWEhpWf3JyWCg01+AuhXG9MVMbfd
1306SL3lWkQa7IYTaur8FZxH1NlSOMtNwy4QdbVmICW0YeehuF23cry5ctEl30PD
o6V32crnh9ax0/Oob6PCIVqDTDzPY/p6TU2JXRvRv/T6NgU3UuPzBGq8ady0xmql
HdDtEJ8Lb0sKNBBDSBbNDZjMDghrbYq5ZB4uAuQ3JP7hi66s5l4kh+YDW5IEndXi
qhOrtfNRk5XVe3/m571si/szfOK4wZgSWNizWHlHCj8POjnd4HHuRiVze0IuAg7x
CslZQNZIJsZcgXtvdaqmXDCWgbaiS2x1ZcWpOgP+T/F++Dh5mkspTnF2EvVVj7H6
TDWx5ujXaDViPYawo7cXpHIaDUT233rgBPa0ggNr23121dWYCQw58kPTYklqIDEq
04ZKPHaLoMFpJhcGI4lt+n+B4hN2D/k+TU+ldmofwvtiH32fLo6EjTeKf9qnMv8s
KiroiM2t1daSu7RAJfip2zMrY9z8NF2xmApyO6LQtWdmsw/Ao6S73qAD0um6sqCL
QEG28LMhic8C+S02hVAdrH5DJ7/bpXv7Bg20MlY8leDNZd0oMDI2lddu3fhM2BL2
lYLGUmqiF/uHsAkIKPS/lIZ3qWyFq2CuF5O/ctFs+QHxMfO0DighJ4ZEyBPEpOdo
8pAzvuli2FAiS4IfvBX4hm+r9gn7QS7G93LdOONp+BjErEvGMnyobKsYHBQn1UJ5
coJbAuSvvdUIZ6zJ0XKC1Br/0Gt41pVmntCVEjNsJnrNCDBVPxdszGSSLwYglVxo
gCCAnFuGTwaxek4D6FZzqZwYajqqBEd/Dli9N0Psz14Au41/oSw3GeqHsj2AXC+D
rIvbEZZVThyWuXsxDtVPcVDMIwYpacrgKa8N/dHwzeNzrqqNbveCdCqgqe0KaUA0
SN4GTy8ALE/rko3P38m1tlwEhgkJL9lspaiQJ4sYvbV29w9bbKk5tS6Kbn5eJO3i
vFZoeivhmBQCHv8uex9pFMu4HIh8a8KEVB/2jjXFZOfe3Y8aArcjEuYs8UF7hhSd
aPHw7gT0F/3CKd6K8L63OiI7odKZsXbUIWidE/VYFIqmUEmMz9grcifoOD/ltKIY
utNudr9S/XBqt9aJ5Br6uRx0kgv+NAMQjHYuV1qywxtz0pnfIHAqiWkuztTA8BBt
CdzPj7srnmQnmev/DE2mmhVv1ER5kqD5umeT0Qny1zvvzPvzDFVx/ly28oIAqFWf
wJ/aU1kWjLhstxynKjNiiJWeMmNTq2SclT84DOF/nUAOMcufMqWKsYpHDQqWHQ4v
GyFJzxWAkv8MYkSZKXf3YZ7VXY7cyuumDmudEe9lAp3pxUUuYiPXmK9+TYJ8GthF
bHWhG/ZEK3O6+ngfKK/XnmoThsv/CXCCYgcWVTfIK8K20VoJytPAoi1fjfbEtiK8
mGYLeAXStl6lI5VWGsSJy5ZnDuYBw271nOuXlhU3CyawBXuWvFY8XItCCD5BjKia
wEy/QtoAb8iqAJlgZvEtH331eCEexyx26oOPIPUuliTK2qpcVn97nBqT3dZfznIg
tu9jdWY40A/3IGvCB6D3L++X39TeqnGfqHesUkk4s1gm2VtZzXzVygjIAtEbhAfd
9GiWxa9J1aVWPRF4ZSkWM36a5o1oudpAJHMdlVnHSc5l6kw0lgYp3Gyy9vML2JAT
FxXPIagcdtQUT+ztcsFHXrLSVXChrM96aEuZ8bqkxrTajECmmSsnCS+01/mrC3S3
WhOEUb/Qa5bViH0RCPPwI1a3itej+6lsNYwomro/qQF3yj58U98Wf5MLmKq7vh5P
6O50wyYYjJQbm6bpeXo7xlCqQYH1MAW4e5lrbkGKn+1l61VX4GE2cDA+B91gqBJY
WuTk5ZpJdYrAPd2t/XhzKxdaeDOic6hfk5C7WGAxPlP/PeaR0jm8nfC30PMBQJsy
8rNDdgq1D29S6H9k51MdxMgeDyr03zov4qnVfkLv4Geh8heHWbnzy8cFAzhYJDrt
R/aYR4mIoaErl/Q41y5LtV7XgUp/Lf6mlvqW83z/wQlgk0nOkZBEsT4C4ubXIihf
I7DypfxH8TYbHS4wd5G9iZ30ga5MV68CYEkaiWdtd8OK5vQ1Jc2HJZDmCIRzPfal
ljJog+2dRO57OU66u4iVo3OFZXyvMmBZoJWUVM6MNJ5S1f5HfbnVYnr64KPF1lfo
f5KW0sA67bHLTLYTc4B0beKDqY5Sokq6j547AjgJ9KX7kKa2LgHVC/bs4qoHgA8o
5pLXzhknpxZAKCN597W4L/x1yn+Jj2NJPs/l9ddD8ow1LwyAHAgf4mB3myDwWrhD
AII3SHGUyQ1KGW7WsxcPOuaj+GANDrX2Jzb+JZSXobMYexuxNAyULJ35TANFevf5
5tk1uJoHe6TdNmcs6nejZMRsd7u/wxsaAWp6y6iAA7p7cC6PujZ2Txh86hg9lSQb
gcs+bHRL+7A70gesOlc9n4Keqmv5xP2x+KFMpbsCJjQOthzJx69bOqFRBZj9qtfc
ktQwznokm2ZDCuKz40H72YeS8YPw9dK9mRwPaOH+xOLpTPEBDn2/nqmH9qxk6u6w
aN+maOs/V7U5tnQqeJ0MKBZ7PxhE47W3oMO3Ym8S6TF1V/RpXYhW4w8fUZZWpACZ
byQzTLKH7J4d6AGwBU2pTDTA+Sr7IXS3zPvG0LTXoUheV4usaURUb3CziVd+TVNS
2fo4IKQL/nXxZOzqp7jfXaW+zUU8iHg3E4wTPwbOhQLYZqk+/hdrWePv17i3Lc33
ySBGUNMSNIYQJlybdRvqjipDrh6QAyC7n/Vl9RHeaMYgJTbm5wEny3m0OvFNLEJH
3fhyZnYbE//S/k76ych7kbzZV7uxxBZKTVT+YWuz108j09VmpMbirBzOiyigPgia
fBtAzx2PpIz5XbtginCVx9bsYbYeVpFmL4kVh9xKPGqozoRyccuoyz2StRnCgrP6
0mHRQMpD3669m2PqtZ0hduD/2/CvBVYMpRY/T4suo7sM+H3hFNnY4WyMRHY27+tR
/TIMlzzeRteTpKAcdNL9fXXLNzfQ0+jyJqBtV+TzDEKWewmB4/Vsc+xu9mOc/jlZ
uzuMj90gQz1Y03Zptgsxb42x8t801+kyoic95R3uCE3vmT9v8kwXBkRHz8NUsJAU
kP1AFNECEmwr8B0hBR+RH9z5d1dmVOdEBS7jFRSo62xLAz4FZvD/SqrwBMBiKcD2
6LhJHorOWP9DWinj25l221vfYH1HUro/e42WxnH3PtdOCSR1zXRxQIchZjQeodeB
KYqEr/FAziyXgxDHI3c6d0JJlQKcMveQ9UtuzaDoNGBzYoNbDJJCiJQBRNmHK6hq
Huy3dWf5+qCzdXsEZaWIN25lV+IbCkSLJvRQxRJkj9TGyT0eLMGxUP9HdhuSeis7
VvgEm90QRFNnyIz3rAOy0zw6LLafsZoDX29YfccdUnJXEGCjqUwmjcp78opPT1iJ
+iU/FlIAw4TI496iGcXMsMZY+8SKgbM4CGtmoYOLkNv+sdw0pbtCFqDF21KksAvc
lFBuP5JRezaDuxNxGxRFmonyb+F6QA8g342QDxLBvLe3AzWaH4EIt6PUkllSBN3m
lSIESiUJTG/F5Fu7dZ/Q7N5fAp0b6bWVo9eva5dFNrGw+Kcb3GzpaneeZ9qY555b
vhwDb2Rf8Lv2G0Q3PFfLCFhgLjw0V6NqOWxdFt7jG88NW26t9crFhYqF2WGaIgTO
x+UP13z8nB6c33HmiC1s0NXQCz/yoS2SbLAdQIo7gUf7QcSexJlAvage2R0N7VUV
/XHJ7xYzcqX6fB8Cn8ICME0LqiyESH3KTqZrPjuH+SmpxVUEraI9ltB3ZwufvFuL
IyTsevzoU89TUaR/3oMo7GA42RFI6FiEr4LaFTkW7Shr7usVdbUBPlFWkG12fCUL
MBjvHG+MNo8qOyGALnUILFuDc82+jQHGGg56LsZGk4IfISUevnbHZXxjGw2UHy/T
4gub8sWYYicG1/HZYy2baU2mKlVS4AJm2Ck+K1qCztcQFKIReggstand35z0kfOr
5YsNUJvWZxOLk/dKbPD4mhdmwaoHsgL4v9hibKJwy0o7ZBFjWPbqTFMG4k26FoQI
PsJPGY2oszfD/bo0yxb4O0jjAtMzFk08MTNulUPpwRhR192GkqLdiSgL0FAycEH3
xEh1xFSVJX8ADG/he0lR38JKQpJIKCPdeuxAo4D87qH6RLClK6UybIbHBMmc695Q
MqXCIDDTiqKkLjn0uPJRdEPKg0dyGE+rhqJnLBoBEeTUZjiM2Ph76Rc9Kp8dUBUU
sxk9DAdEHaKeT70YJDFf8215TZXn/KYEwSKf8i58xobNFjRGUPrfQAyZ2GeHXhsM
sdQCF4aXJISsjbJ33ePkKpNYda3n+fzV2rh5B/mpbEjBUto77RPHA+SDLWd8Y4ov
Eii72DsqybRPPpUH7EsQfPRLQNPavsM1pi3+tqHzjig7ghn3oi111AKXq1s96Jk8
/7INCA/9kNbPEm51dQz6SXBy+nJaetPYpnBtlt3TQXjCeKlljpm3i4VDKwwJnz+A
EpN8ch0/wf5vMO1BBv/NVEk6zjpyAE+OrnSXGapS09/ihNpD1p1UuUJQfMdQXjYK
iyyP+ZU4YlXaxIzJmBaGoFDLqCFSEv09iOhM4YJZtxZqjE8CBo5V2mTH8nm1P4sB
xkIEP4sw30iM579IkdaLvY2tePmJTjofzfjSFbJ2pZANAknpfqNvGbt+tSxIgD+s
sDIcyC50jPJHhgbJAAo6FYL4Ed6c+hlYYo1xy6uXjsQ+Cwp5BBEcKIVkgq3wRo7h
afgnQAfyWEAlqQRnqGfYtCe+rQ+JheK/VShniDaQ/UkdGcf6+zc34civczfcEere
JTYtZg768XaNytaQ3mIEUCsVqeALj6tez+fKJkq5N+h+syTL/ydBUygqmWs82Gef
DVUPLwZooiLoDrxvrRqDQ5EfnGMmYEelwnIOjcMPbVrfWIAitN9ezsDAubff8KaT
64o61Goq29EnkpSK+pDTxScWF+SiIXO9CQHoRWzpuLXIjYC0KmkukrB7o2U5+UM/
zN6uW8YFLmyKEOeTfhyegt6OJWYUuqOlM3PJpsdW5a2ukeTH8QBRY2j0FinBvZOf
5wI7ztiLDYa9wJwIX1P7nJbUcm4eiTY0zv7bJD8JivUuNsEbAoQcdOFZWW0Nsugh
F5hCUGfYkmjltsT2460CMkJnnuwF76InT5eLV35aMf4OrYSFQ24TygOv0K++62vu
cE1gfiR1BG28nypi/x9jpgiravR5I5wlkO51FMPWmx/3xi/6U2vHdLM5ODH67ojI
e1xh+frfiaxiUe9HNpet2V0hU/IdP/R/GPfJzbNVM//+nI6sUDSGpAjqkmn5j2ur
YiDkeK938mxr2ApvRHCTNYR4/zuxGF9hAKL1f73dE8V+25ezh/eXdzJJc4vjzqhH
JqU8OG+w/3zdx/ZqzbKC2yfQ0O00kZ4WwFkxscanAA05IMJD4w7BJzMhMl1g74oI
vdTp8CZNMyScnWYMjJMc15FgDnKOIDubwofCuYjuqyn9Sr863BjNh4VuEU2pIFXS
Zii3xa4a/Dtl7ozPAHmrNPOXePZFtZN8iwceCeYm/fJ8Ik/1ADgxoTWvYmtqnaCq
tUZFZNmfRf0BVHr7xO1qyx9kFaUBLAVSCaJpeJAjL8T6XHTHeqM/etJYUszCD3VR
/+aIu8osvpGrGJ8yIWyMTI6TKLcU48+RFCHNHC2T6Qp3Gc9FNkWglSa+N6z4UPgq
aE3Vt7ZTeQYW2KKVHzekXBtcayZQbgW8t2DDu0RTC1nEgHxx5+krrnB+bAIG4rka
ic6hpyQcJDhGhnaKL0AIjRmUZuvZTOljuPl3KP9QMnOiDUJLX54KUKsf5KDg7eqN
ZISK4R7uu942EfyDcCVgz9HwMEZ9nKvo1pc5J2cLvxul7VUsHW95zRrCOz4O++1y
v+OZe5GOfjC1Hymp3bQ/R4sF3yFqTmkza/4PsQaX4A+DKyXeWJDw0MCmewAA9Ltv
cm5+EtZkvHpJRzRsqfrQ3L8yrpMd9O9YLwZjudgnQqk6w5DoCOWZf0duf4SKleqh
X2B1KPwq3f6G/fjhfwxRy/ZWmeov5ADCX8jKxP0gjAPCj2z4m6QOw18XVVqQ116/
x+4JersHzLwmImiWGd0WeqKFc+STE6GDTdPhJrro8VechEGQ5QcEsGQdIrktYfHN
oADgX0FoCG6+r0NURCRNCMUil8u+gUlvdzLFQZt8UeNLxybTwjgyNZzYlROczsOE
igvDRm+P4QSe05nJwPRg277DxgYu84G96SVOKGXnYFtuEKfQuQ6b1Cj+B6c+VFfF
DAknYBNQ08fruQkX9GgjDVIPp2eBl6daxYTyseW8/cdTMHwuBDUrFaBck8LQHeaR
PKvFqnnKmKqM6/QdkktGQZeALnd16uxOFVbMKYcjpbgZaHyD5jVZ9vm7QwOlYeHG
Vb1pJLL0JtMuIn99L8qLmmP6k0LErgs0dK/30iYuCSGZQLdNMk8VmpQ5XWVAsZxm
nbEQ5PcZkH07VQUKrkFyDdGBNLjpX8nKn0Ke4OiIad0BwM0mCq/UMjCWFmO2PMW0
4q+mzhatIfM1DJxjZeaOQprcoLbWqdCwhi7pNgcfSMtjYAJqwu88dOEGOFBpAYgL
iwJ1dBL057e1TBUsV9fgR3vPtXsF7+RcrLOkuQ33xiDBBowD4oYIl/8G8EQ/DANg
cXHjn/pBlrd+bftzeWHZGPcQm0wZWiSkW8FSdsqTJcGF3sgNA1tPU6BsasJliBzF
bWIwjOr8EUu8PjORmcQdUK1ppWzSDkKwWT4rFCzGEYZ24yhzB26C+mwnlBpNjhyc
xYeaGiXMSRud6zbZxmS9s2TiHmopi9ShQsZbEuGyN7Ow8AVTvkJZWcb2oJrWdF+n
ITa9hcI+pv42sdH2VholupWNDfhPP/d3MoLTA9893hbSdwa2BFVOK7BbDzKKuGip
F1OCZBuOZStJMlwcW4A0hvyPKISJWP9dsIUYVDuLbOk9K2L34RXin+JIZLY7f1aa
NarbalFGXOpd552e4T7U6JTgEzl1Jur6pwZDr/EcvDzdIf/SKVDi+dXHZTNxqU1z
Pf2U8kTEPfI6Fn9Od4Ow5XMtsST0pvk+hMkQP3pawJroOPfeHS9TJnNClyWxVBrr
QP1igj5n6fz1l0oyx7uys4EudRLVxwdksqEBtvnTL1GlbPRCxt0nXRbi4y8jguai
KSURnXx4NKXmlNnWPOg6lHKUiqfoLN3fA4n4jeDvw93LdxAhQE/9RI6JjwVtmOzv
7LZkOwLrFldHvNRwTceXqvq1wkdrgIXugIc7Bj6Ll5aE1WZRkq7aiFKLTD5jaK9D
Oqv2VoKdo6EUzUlzcMcyYqFZ2l0pabqYCku9qDgVgxVidSuMGQs+skvKQjcfdzwJ
HE6gLhQ5PLek78fE1pKgYhuVhud11vadBIX1g2tQWpWa6wqRHK2nZtQ//+1bivEJ
nB87q37kXVDdhFOLImFU5eEzprfdSaGYoKmUCE4ivdgUvOhHe7+lTayeLl9YZojY
grsu4FEgikm5rlohygV4CqVtgYjiG8UHmPrNQQedmLn7U9PdRSEoxbJa/bKx5BSY
GtS5nhKpf4+ICRIri7vIHeXq66nELu9cZTjm5NhF0UMMB8/9OiwqKwhWn1y0OPmJ
ejFE86vfrW6Yusq1OylyD1P3qgUCk8VrmB1DaCxmSnUYR4akc5oFYnEVqijRF6It
zR5AsEBy613J9ZeyRWydD5S95H6GmEFMzpO60oLzM8vNnO/G+O03WTdHP/GKkxMc
fe/DIz0xnKmDEO5Sygt1v6Iy6ss5Z5qnb6pUQHnDnaF/IAW/DqioVcHMsOnGcp1s
HAFCg7ZGARNudYMO1FyQ1N8Hcoz8yR5q2tWnFlC0/vqXP71SH/iMVdGVl8ijQKPz
d06z/nQ/owjR9R07GHILPEoMy2CBzHYuipGhSFKfDonV/G0zYOseRSPBFhMtXC6R
lD6pEOU4T0QasSlgDQzjmT5HG9G+GLw1/3B9Fzi9lYohUB7Z+1hrVmv5peixNSbs
p6n51dChGgkNtM/3lSGt7psnDxCbkWYaQswVYZdVZ2IkiB3B787a7jqJ0SqQr07F
vc0wueDW98rOtoXGw97GuIDTddqHY3e4s0R2O1jFVkuG5lvWf6LyRaLhl0Vl5YX3
J4nYgTlcwQfJKkArka5I7TlGZ7mrywTAbqaYwknBy2IdfEZpyggEXYm0diNYoygO
FAxtffb1SM0X+VmbDg/OeQ/7uKuXHbe+VYfc29SENslCRymKbBNLm53vHs+Rm+nE
5/9P8Z7H/hZlFkg4HeQK/BVqrG3d1mlOQIojwJ3t8rjojTNjZvcJC8zGhovzzl2V
f0NeVAs4FDneofGXlVBYqVzjOH/qB66f66CfFgiAnCkorF6CPGxCx6iGxXhSCJZ8
JFoaCFs57hIHWmlcPjtWRXF2vHuOtRmlLagf69F6FJG5O3q5PVneUd81O6fnpFRm
hSAgYHXk3nPokGs8oj7Wvke6Abo57N3ZmMtMCKzBS/rlfACz0gHLN3TvHMqiR/UD
TLiNCwl/xxn2anZ8Ad7RMrzK4ENDMv47JTigHROZoXL7vJfC1DyX9dSzkA2m/eZO
f4ypNm2SMhdzAzM8jhv9ZznLP2ksEoy3diSHNvGjYAuEsaFh0X3/eHHnQUlyrHC3
gg4em9NzY0WyB5Cl4pcwREzucxD1zXdXcgX8YvQqoDKoYZC839lw8Hc9mAYGbf1j
Q9JoGfbiPjvk23AD5+Uu7bFPwlAn8ORT781X3GxOVyPRBE7sic9gvQL4K/lQL5C4
m/TMr9VGYrij4uUHjpQOEPR4qAa764MbxH4jpmiEgyfFDKAune14RvSfxB8wKtu1
FPjaZyyv0Aq5ZHam9HJiXoBJPTzcG9oky4oxBNnn5p6Tvg+QPzvSal/ozv2fCl5Y
ZrUQIJuSKK2Jg5VL4Pi680huX3G1Q3mYoYLU6z2mfjxjeDIV9ZGqFyYL2+v+1a9f
AOXIWed2netHYA3XsEu+NQg/g9x82/F16453kk3zkAMhIvqVntZD+hO+Q7pLsa3j
BWKKZgPiUho3H61LXL38Er15wXvMPzi2rlqAJCVISIL2+Fn1bETuOVhxWzTDKDBe
18O6/jSMnNVo0PYi/O7KmT8QY4Rb5e1SEnY5nQkfBJdoSa9u4ByW2nziJrzlnERx
+bKMCz/zvpJ+9wLpnmvLRl3P/zEa/bjNWlb/LCyJ9srjuvxfIAJrqvNY4vZL+NQ3
jgQ/n+ZDr7BiKVJ3yhVi7e3Se9NU0xN6lkkus2Wzo45hI6xeE0bjDEG9b5RT5ZZ4
Q5RMD6PX8MYNOWsj9uWNAmQdURD2jHLk+8uNw43pV6+lLxd+FZe2jL2aNsCPdl0u
xS3pqo/6OYRH8ZLHLXXyTTZ9yZUeZnDw4ZW2r5iEgv3zkC7vV3e2NZVO5+Bd6tvF
YNYufUjAYIJKT0W6Bi+vJiBxfNMtD+NTrv756CudBhn83TTD5jCDD3GA7RsacsCk
JgIiB/wMAtyB3wZdHZOhtIn9kINaabYW8H3oF/njpLCatG7HMDqNzMy7Pg+a9DXm
4l+swRwKXN+tajtuuBv3/hpLNzDVecQeMMld6Zt322rUTTmcJLXIol3lH2vpfk7v
eXq3l3hb3JVvRVsFXzrUP3QdNFztgOyLOqURrL3lwe8H6n6t8c9abHAR/mkywFAc
NI/r8Sx/AUf69FWJMfr3jHdN4iCEz/OQWP27Gnwq+s4ZJLpfQQKuRBloxao1xxoY
mcc6MlUcl1Os1Z8RCuuaXVFAGzd4ErOyTRWdFGapHesok4JdJYxPPR2ChZxVMqCS
/xvuxcuynKcHprhvLHG4g61lf1RpkMmwCApgNljCYwV8l4CuTF6VUicKlG1AML5c
jLbtltUZZZC+WGY2/E6M6SOJGPOzxhsRxlanyVyRUaVj6AfGSHOTRxWnUorM8AvV
QJXNr5V1kqs4uierWwohQTiYJDLm8J7ftt3LMV4w3NybiAbV6+HTMVS9A9cGwOql
3T2VACtbdKCyU/GrGTP8iquK/LnEFM7PJJsTf6U6SwzQAnoAZQtI2bbi/5ewq3gc
wsfB7PVTLJOcPUyax2QisimU6+TyAXvFEnplbGsE9x2F5c6WlKmJLf54TyPaQarm
P+sRFKTX9mHUn/1xh41EEAwIBXCRD8VUqqeKuNqxdwq9xDMTuUt7X3pdQ78KBLy0
yzbaH4R377Ao+PcdZniIsFohhMx3LetuUf+SBf2DHd8JxBP5c9HYJZclDJb4fq3H
8626xUBufAdS8CpLIuy8ozcEDbFijLgYnc/uJAj1LbFcHtOudAPAMsScqjvLwjdL
TovaUjltJsZwtyY/piLHLYvP3vxhZHkgu8EsfqMeUW3AhIPACQc1Kgv3XDzgFErc
WfMtApu9xzq3vm+Vyf2riRVl3sLaf7j+56ry2q3Rdjzf/d/Nry0Lqkpk3t0l6Lj6
35jncsZeBZteBqGxKI/mAMWwmEoNw8J4nxR3RJkdoQp8DDBXMdxMhB8enGMuQEWr
yHBAvWWR5MrREUN3lVyZiijohO/BhgzvODGPLedsFKVrfhKymlhXvyPUAakii06D
96h1S5zMn1a2mdDOWfzsq/w+C4+ZZmtMa+F3q47gJAeDTbJTI0H16grDNF1vS+PH
nB5apE9nnCc/1ZLkmA4iYL8nqfolVoFF9/OoMQFatKoyaQvHQa3g9SzbJ9WDb3qp
LNZkPVJDN2HpRGN3BR9mBT+9kmykfQBIRwoJZUdLEGlK7nFF8fG18dxIxx8DBoz1
qfcFzffEtd81bH8gRX0sTCI3vCpaSQI87cn96z7OXrWs0xv3TKllK7jisIXBdN4Q
U4HcjUgOrjCnklwr+VR1cUcv5EO7CEmVjLz/mKvatgHCoBF02enscq9JV/d1WC0q
ztUybWi5ZjeqlEO/jUzBP8m/IoMRqW01pvfyOYbK1a7IGuoZ/nLkTGbuqQW5zTuW
c2jOw4d2uRCmV8XNB1cxGdD+DQ6Khqfa8nHP4GcuIG12W8aZRbpyReZ78EHGdH+8
saVnXq7UwKWiFmt8lqMQvHdbD9H+X6zcQe+eQ4ugqlEgfIlHXvuFSu9T3ba6B5e4
8ztCvGx6m6gWxjVpKEI87K428w2TPevGl71SweskckQ9bym8mkle47IlEB05ZgUQ
k7K5YDuI64Vddyoc2lQn9635Ddn3BbgVmFFFOwviMiEViXg30+pCFxpT1qdU0ZU3
U2V4r5gZMzGY48crwbAe8HyCTLLvDbTo4dyrQ4uhBBOcHdMXi8c5zv19AH2MbdfX
JZNGsMMutNo5QJL5DyfLr+/yn6c38sAUai353p7H/Zp56Y2p9SQqRsULOF3sEpwl
uLx7BlNWxG2n38QpQVtjrxKMo2/efcWZP06+mTLvE5DvyRv7y6ipbXhVQrAdcRJJ
MpO1WTdEtMq68Pi+bo77QqYbS8tc1Ra7+PEa0iMXQEXueEiFSCnN46VOZ6DmJnIf
torzFB/SmXFAfG2G7oXVwmgyS5GM8UVpNGgHiHJadAmasFwaGwOh7KLMp72ariBR
lCsYJEiqTHERz0vxhihrIu5/yacYJGxdDd5tRqSMBD09b7spsJZZNihgvLeShMMn
TzH92N8+WOnP851SonUpgJUhvBxJF30osuZTLjYXxfU/PpHMz/Zz7WVKcY27T9iD
qAwpGV08LhuVbXGZHNgbslnC5sDRBYnccDW7+SxUjECePDhbIKnAh9CqkBBAF8MP
2f0XqBXyVQaL/yZuCO7upfR5Rz7wFjoBs8eHyODtxLpDqD+weT1q5DOq+jn1gzOU
MkWuAUwbfv71macS5/OUGbLhxFWXPMTZqycMDUBCClByyCxgnACanA9FglaBO4G7
PHAMIzFT1hRSE5jjYU4mQu1T/owIi0XwPfDkbIbi0e0QsTIS12IzUE2C09Z43JeB
sgY2dZPXWrkF2+LNF3Iok4pf8CAC0ipcXZyIC0QbJGv/UHGV20BtgW8pU6PS84M6
PjVKkdUTMo7miaSJzGEQDIRqXV5xIRZcmzuCNCWLrJupiK7/tYJhZmwUIpmNior2
JmLejIJX/oNas8NaN2fGmDHxN9vZmaIxjTj722nnG326TUk/OZncmc7c2poiTgie
jpaBVe9xFdcf3LfmXcmW+dw0ZjX6ZV52iZtdiI4qwdIGGsT9GV60SYNT/tdRHw/k
5/udc1rSdJEGq7TKi1IhAFf6dSDj0N9SG6qDtwbfCtBGpsKHh86S4OdCPk/gms2Z
mUVkqVfCXJYJ7uAIEzpngIozqjNmGCj96D4z+w3VJLq56rGvg/RgOf8NBMBk13a3
QbnDXjAHpACl4MT7HBKJy+ldNGjJXLYkCDRaDHsSlRZk+EN1WN3f8m+RXy9avvMo
WL1s4BMio9HvBxFkt8w/AwiiykYzCWdCKd9VHVe0Y1Tp2S/8iylJ7FyzTOcl1iZr
5+kdVNzJN+JFamsvMxYxH+DGItdZd8MvseSIfWu2TYOwaCyyS43A2onRMux29Um+
EjglJg4Aj5x0wQpXh1pQDlzLKNuFGaq2Z0iWSY2CRYFordMVysYdHwkCZtKiT7bO
msturYK4ZZN14CdnDNB+Je9AIZRAeMNIFC3YpWs50oJ1U+UotMhyuK27qwvGXbSq
zF+Q1IGobPvKrw2DtG/jPzpMu6syRT49eVlSd8s+pltkSwRxaniR1uPji9nFjPLH
0P/2dym7ha73LAkmeN77/OeY8YbEu9p2uYwRM2dKPc/QSiGyRjms0S+NNgE7by5P
W6f+etoby0FUb7p7s9AYrjCuUtjPavuFbyluwLLGi1kuJgoNWcUlqoEJLFa3vohj
UMl/s/Gr2z3Cjty3Fyge4RtwoLOJhJSWYoarBCL39+O08wyJ18WEFBNXQ3Orfkb9
01u+b8CZnMOn4qdse0NPcobloFcFmyHiwH4aLtj+H5ZuySCL6MGy0Qso7lHjaivH
1e4QJv3Tl7noVTSk8QaEzknwIrWgOvKO5XIWyysoVFruLgDykWnRwcDUd6KTdgSJ
rJ9QjPfPUHqKWp/GjJFCLcolD16ROWCdfqQSuaw+ANsB6g8DlsOdcfoV/nUQYOh4
uoFAelimuy8U/HCtvh2xtrhbSletgssDxuRHzD4LEKyrg8YSMgUN+D4lhC+7KqDU
gvU/IG8/EuKT/J0PaoKwRFkATn8c2jM8TY0YWSZng6SNGtboeiL61CHg9o8z08be
BH6lpeXwXT2HJ2u5eKNDe/OEqmd+u8f4fh2HK+2IwaXkoyJtiGNMog1JmST/4Iew
YR4vbG7lney8D3Uo+sUZ989PBPd5P0YxvmIoTzNN8Lvfa4PfPFKEcgP8a8XrhB3h
z5VOsL9zhhjTFOn6UaInE0CmtCN7wQ60sTp6A9qaFZUmvvT0dmMxEokJRETMZXRi
Wwcfkni5lZZX8WMWMFaeOkNA+nVIeYmSgkHLrPkIwoTqMZPECUO8XxEL5eUEzo2g
Fi2DYREZFotOZm/z3/2yscI8LAgHpY0e8GkS00BtyCTYMfGs9+5eodFUXsJTfhb4
RTAtRIaQR5P3T6Z/KlOwo13QsQxjPj9CIfNTa44wFQAhArFfcCGBEx8qcAnFRtEy
aOXc0sJinFQzaYDHIwyJDhumS5KIhYj41N6bXVQ8hCVaWbqkRBh/mQu5whqfk4ob
ebWf4Lo3mvKLnGKj1VjdkaSXX1a6gMHWBrX15zm5dDs0JoS7KjBnd/QsWeKvHUxP
c3el32XoLd1pxuZjROfquCu7+BtcIYUzYNAWsqm8M6ms4cdn2u9ys1oh3Z0KYkmN
mbcbW+Cac6yFmydgY6ec3t/OUprN/rkLM20jTp7bqSNKrxHG8dGX0l4wNij/ReOx
DgAkpnVZz8w1bvxdtmV0q551oNpPMg+3W+GREOOEorJ58XG2rzp21JJKSV3NJa6p
WV4p2JyOwimLKrfPuN/G+8MCi9XAQwzixv+r/f5+ZkdRd367GJg5x+sHUS2Ryi7D
Xcl27eJNaaq3MdDaHhErYUy5lwBvh8j/VcreMB7RGgUKLdThg86ueWTgHlQynoGS
zh/WNM6Rvzv88zws5RKI5b9APaEXHe8m+H8SYondzbMI6AQ5papqaQxajfMMiL4C
2j1GgXYITlPh4n4O1/os97awTGXNcSXs1PsROsCEq3lGBLwPdfHA0xv7YLGRS+ux
aEqkOjCfBW5IVHofoGBX/YFC7yRaCe7z1mGfmPkIriCgdyCJU2cIjlhL4Fxu+2/f
WiQPbk8xz7b4EpE6D/VLg1pYJswQAqpWhNjNUCOjbLRHNkInVzRaBqExl5llMn7u
JvoXqMqHnQ9o44RLG+11MBo5EbvP8kJnUAoEx4C2piqLte0njtx9nDf5OwfhtENg
pIwc4JXhPFunkBkpcsF5kvwGaZyEcwY1tziYHsMzJwlWFk0b9xQ1WlPcT5kWkTTJ
NtZW3rVxkyibTWiS6nrhHTew3GwNPkpS3IOltaVBI/xZkfACVvv6cMZ7UWf3vU+u
pmOSthLCF1bd1oh7KAEl4NKLC7Lf5obFYZjmEvclFxu0B81HBw8oAz9/A5rTdN0+
m1KAuyKCHWExK7+AHKzGSo27PhtQUgKz8CeBIZX3E3/vWfuiKESU2clXHFRr/i9e
sjHk94SMNDvju156bw2pEqFJcu1TbA0n8gQqPgCOnFntMFZQfASUWxn8JoRjNKMX
20SUIeHI7Zo/EgQ+aysolCqQks5pYxdFLcddp80Rx8fOUSrn/t+xcm3a6vgdayRa
/03N4BD15FDsvbfv+8xpsFsDWQDAmFRs5AlOt7rOiPOwsMXmCSH/qXDPnFSXrZiL
Z3/2Qv4tsK23ngY02fcOgthDXRzkKgTSVg3cz+AnDgg465iBrnNSwymHrMyW8npq
6XEvbqjaCeaonuN1cJh0up28pWoApwqr0kYJzN/5pOOIMFQdmkFam1XtVR1y7mI4
MEl9osJ5cz1YtHtdInRRwLDdF38BRo3h4/92A6F1S13ynn/fX5xT3W7CN9Lug8xX
emjQtTHyb4mvhqJjz6C1GHZYySHMrmUIrPVyh3Nwq8xbTwAJT+s7xOEKli1l0mig
k2CkuBVTIq0jBg/e9QmKEDOv2lFQtZGIWgpNK6aotWhFZCf3JOWT7szJnlqqmZ+d
FgdLQyvUkEXur6wRw3Zdkv8aneYc0SAHLSXCVK6zCu14k4uMcWRpf3Cst48dvsXf
fJkThbBq7kD8sAixUOCcl64zNfL+CsPaw+aCNWpe3xjHcG5OzZSMkDLd7GB09oIu
P8RTuZz1GNzKCRGh/7QcmI5IPPIFd3uoOOY0dvW8Y5IJQXTntz8AYdnintyv+nXX
1JDmC+bwkllGgK2waNJot86INBoJASHolimXBqM5oaIrXQN8wCusKJMH9V1kzAoz
1I/e/wHVccc7azjrJLdsT5Mzzc/lr5ZtkN7S6bYPqS2uuAe9f4zdvgCjMGT8xaBH
gbbADQLCiQQF4psnnGE/7sXoHCNZjTKMrPxPYY+xC2ot2b3SUZkJXZG1wJEzTHfq
QL8MvVF8dxUONUdVQ6ZXMHFYN7Ye2K7SoTnPGIr1BI3VlHHIE6V0gfPFejVz0cVN
ixAOZA0e/lIjf9yi0vtBE09dVmySCyGFYN5q2frdcmgZrqUSazGlt0zsN0I4jeA3
h7g89G/A6J7/Po9JjKhygJC0avK66uuNvHvIfkath4Qe7Wrm/nOtFRAZYJr8EVVd
NvWNvormffYUBnxTOeTg9WVCRDcEmNErxwoNdf1R9LP+mn8WuoMv5SPIrWdD3Zot
3+nbzi4cVM1t26N8sfblTT0EuHuKClqNr0tANdH/ri5e7qr4gVGTi0WlrlgwYtyQ
hXE/4dS3PbBVkIp/nT3i5I4LT01K5/UuaClfq3WviSSQifjbDsjZHZ+QfKKUpLYX
f16NlbN+l8MrRyQ/O8w92t2PuvRdLjlVmkeLjEyHDd1PFqhOXZc6kkjBBMJujBB2
WYinTWPgj4wCmWJYTVwmnWiG7d0FPSueRRpyVuYNCH8OsXcIGYErPqUOcq+dpB4W
Dt/rxZufYG7cL+V1307ZTkABnEOpcGC8+l2BYUKbNqoFa6dDPxwV7Mm4nfoCmP1D
fpm+9dc7WWA3WDC7ZM+3DE7DjJ5gUhBzMN3cMeymvxeHdF+Sewigr82aaYrp2Mgi
iS3Cl3opEQJ8r6ZVuGBCCwHMfxSABiZagmwCm+W00xNyjjPGOwQyzAUcmC7IEN2i
tz1XNc6TLMWqVZ9PSSt5EXXMjYSOYBzio8oe/24CghESHmmWLMlKyqsdXy3W2iSe
wogbKen3ZL7WgisQLVOkcuOBnNrJK9G0xwuiCq+BvZqawTBxYB39qOpg78CfeZ+K
VmuqgXDRvPiUvfMWBMte+wiPJA/HvaoURbX6rBQ8eKCd+0WiF2cIx7kUSui9EcAB
sR/zTTTRUxuUajpp90AHlqEuGMAC344J1qQlsVJZvRWAQtFgGAWVYCH7CuV6VC2J
RSdL8G4lo3bcpwqy9Mb9AQzgtrg44UubO++8ahqOSe+R5rAbfMz6ysaDGO0h0JgZ
2xAvHbcS7lE0n6T36D975MMsynQEbrIG02L6Bo3Gq151b6sNcvpT5YEl0dGBxcjc
LKc055tNsZj4+8o3qyM2ug1Ha2rkEd5R8qZWU74iUy9s98Y5MhX5YLTcdjHqsceF
TOOnho+wcD56F6PnyDHf38yQFuMy07xLkdZBzNNJTBEh7RTHeMpffh9tP3zlKbIv
3bxuYntnp/xGYaewHYkhc5Gpc3xmCIJRTnIfBs49cq0ieSwsYTf7Rc/055EOVZPj
VtdteAVqh3nRNoNBgnHypg/uB3j2ZctbWaa5YsRgVzfzftDPaO2/3P5QlplJ/six
xVOEbutHMYHibqzYnvIZzfTI0wVv/Hn3GO3hivzeguUoeYKiHv15B0zPnVW5uytf
/DvwG9WcxaV2WoiiLwIggBAH2XWjbBczymjmfYEfDPGblvJyph9v4PHvPEiimjWx
KY7wRMMfKjJ+cSoHXU351FwxVuo/E0wpNFAZBI8992MB3D/UIYFWGRMFIA2d1E96
d3ZXFI2Mqq57tQEjRpeOiD5cHY2Esa39iOeLk2FaW6WtLECKrWcETIBk9SjCAF13
w2XIkB7JZbjPD9hdATkkEyTvWJR8RyN8vBwzlFpfNQ4uI1m+SlRPNK1jMHgbN7ZQ
/JLtach6OYhRwr8BVgR4kg+EKkIjeZMtF18ARkgFB8+FC5D5vHrON45alFZnStz/
Xc+pbJb8U7wJqt7Tw4vsEzvGoo9TwRSg4s8FHlWnq+arhi72mmu0MafQKwCSCCYh
KqLEqathAsfS1QA5bmfPb8XQNQuvMU+YoN0zpzOuQEQUCu54Pou84uFPiooDo85e
QAPvKqDOXpEumx1Kxse3ivnvgMZmF1CqXYJctTELh346PMWV/h2I4MZY3AtPMMWA
cBqLIUzP5poX1neDhAyWcRHb+nmSCVDqebpeIn2pyNOsaNmV+QpYHCRy49YMD+dL
1eAsgp7mu7jnf1m18jK7vivszPG8uV/8UBU0RlS50BU1kVaKDSUP48pMOD9NrdPG
N0K5OYuegPsBSP9Y24kZSeCzhxGTBGiqrFSsrvN/yAJqoGjQKIVHZptXHQ6Bq/iS
cLvWoN2uTC9nqZoeJxY8GMMq8ERAc2HtWWIcjZiTHUixVewR77yKUrOswmsH8h+p
v43oqG4142iO1Y98AWVrJ2cvzgrQJKT2wg2ALzYa+tHdeoKG6afF/jeIzpuUVZt+
6g7WxewwySsvPrGZ5s2Nu37kxaMCE+lcq/CYwvvKsYUktyA94AwfqW5kpabwIBOH
UD8vESpanh7E+OqWkmf7m7qKUTcIKpu3FLtypzPiDRkdYq3Zh8OLqrG7TrHEjcW4
DNmJv2chFKOL9DElDD0SYcMN8RHJpxe3Y269cg69C6vB0U7lodUchAH1V44l02B2
fMKhkpF/Zo4o23NLl9K+sI64gSPGXBf4XD1DjI9XEqOIDvFxqXNjkTyqAk4IPvsb
FIWfZ7kDo90xapCSKWRoIifea4VE9CQNRDW2ToSHb/tAHaBgi+dl5ZQgW1PgWj74
OPQY9jKg3dlkAxnZ5fNrD3D5+6XRycHOzMd01EcdwIj5pYMN997IM3pfSPCSSxCP
29QWJ+69J4q54+4NRJzP46u0aTXxUhoDMZy2PPgsY2G5pJItZ720XuV4IjOEFxPh
AqQLsrxZsGQGsXWrjUm0fvk1nH8pVfwOPIw+hzj8aw4QJqMVU1bqwU2btbj6tCz7
fy3EZKab2b7Jbu86CPmJoh5cA3K0nMMeAZrhDEUuNo+gEsmMwDAqTTCRawrrWQvs
jYSKd4Vb3d0M46DoIDnR+RyHeIxHWYqDg5voWIFSg8zTBwrtYEzrb9pE/X8TJYX0
U4dXsN/liuLb0gJfPQnfqz5vCSaECvIcmFgvU0KBmasPPcqE+Y6ueg284AVPXWis
zyVVC3u4aTJIemx04TFf8aq6gDkBTHtVJNoXhAXz9gIDz7OkVkPJBwG71iKNTlAm
NWSJMznuiATYCpQZjxuP2IqLiLt+l8TrSqx3SeNe3xbB7yPz2iEDAMu85lJcF9lh
sB10fwgtDnOhuD7FQo+YbZ5zBXXF8Bt2e78rrLZI+l+h/acSiZfW2B/bFGU/S+7N
uYNZhtTCUZ9sjWP/pgYjPmulNf6u0VF8kP17ggoX+gkB0RP4xcpKRjwXbKdJhbEG
wL+Q4RTl4IlVEUjjS7fE4HiIpBosA3NLu+D9XMoyDAvEyZ+Qjo2+gZDNw++Yt/Jh
D5K8nNlOhXrrSJ04SJFIdSr42cS4EpT/CuSY3PYsZY4pqKFApXP611k5KTehdqDL
4o8K4in7vgwQrEM8TT8+3EtVL11xBrtUA0vYAikNNnx8/1D3gHJTrBkHULZtP5bq
Q12FCwsNtkZ7KRrLhmQLvgw1JLm09Lt5XCwxnRex0gQL/vP9S0Woo4XvEVTZ4YgU
jRVNLHydcra146s0wQa6qy7P0CX72U/eUEvndNZ3VPquOhSIX/TxvUxdNZhaXdkd
k1Q+jKir6fNnm3zYEQ6A55GcW07AvMmYV0SBiFYpP11ktZTiBmQzZ2TUS7WzI9bR
w8yYH/EqGTj+vJCtEH63+fKEyj/DrRYgkZzO8/t+ohXziIgpqxkaovdbeVj79AKz
44eVEQVCrXFQXjZAXCVf1VOrZch3cZXJSErrScHBVhIvGKnI/opnZpRh5rcaoFY8
2/htWbGEzEPz7dBEVCSDfRz1OF4uG32go/PrRDBppvaAn3FdTBiaS0er9sXtSqek
EGxiFw1EHwW2pJMgxXvUZ8MUvc+oiIMHPxZQimJWvrNwBcT3dvHaB2UIniVwkUem
2TQEyf1NWddWb0YX9xMgtRNU3Qp3s6rXi1mwecF5jS7zmsvNIg4jLKam28ocyIKg
iktqypzOWske5CkU+x7ZJ6La6JDicCpcmxU2OEwLH4bbkqSldpovpHqqTODbW0pS
5MKzz/09gl2BwaZEqoi5PwzHI9ItQdCxFKyee11TG+0bUyzs4yA3le48MTHSJZCT
2QJ7jxlYbCbIPDSMpWut5Uog0gzV1ZUbI86XuCYvk5NI45K5hH1LuSv8Uk0sHrOT
DpbYaMGTKmBM9vftvyLJQhRlyxdeHYXwyvowRorJMKipZ83TfqDUbXToZ85aKxy3
nvopAT05BWOfbZiVl2FtyOs3vha4ugbMxXIg25CPOhqkzUdFGvbD6TXLepfHcSjo
jesx24DAaw2JnOD0Q7k8SRmWpbKSnAgqkyRa77OzwW9zTf6N361dxCmlVFEQkSzk
4ppcR6fdz264sjuzT+JD/oJD3wB44BUKl1EWzKOcXOs3tazkQ+jmQurzFf0plwMx
9lOp6/0OtT8YzksnmJDolohQDvqT3ZB2KX1FELCBdLbXOVCeji9kTR/zmwZsF5xK
H3N0ATTVxFm07Fgtqg8lmNrzJPJjHaBYvKoPoqCCnI/abetL1wwv7PQRIZWTIwpa
XsQ7IyZJIgQ3CyeEmNlmS5spx3nFHVx4TB6askuKPUSVmvVUe3V6Cin9l4sVBIop
za8z5CTOdSCEmoZDuYt2+zChvqBXRJRwBB7KxkIlx1JzXUP59o/4y+VVAhwRuYpG
3an9Ch5onUxh6Z+VuG6+/6KDDLAx1c8Fqp0+rfiqGtVTc3Dici4OREpH5uun7eNn
RPLJPc16FoLyzFLegbtf6JFGqCdufWVEi4SJstGMJ6tJ9c8hkGJfUfa1ZndBL9Vm
hU01WGYpyqTthVkwyQ3SweEjw4mj0Zk6L+kjnIXRJAS1HsLJGMPJUR3JHakL8i1i
gA3vSH4zqKhM4YUBtj3Nx0My/Bio0Lr+xh/Cy7ybIO30HVT113V94qvXFxrkwYaj
ARMcA5PjihYCesE6/DIigFn5brl59kZLQjHSXVyrJ9ISXo3u4G0jYaa8r1J7HFkj
WC+FQpjDL0xuBdxiwtSvZYjd0w/tZjSYkDu8BZC7uzAD1ckc5lO33etO3hf/qhFd
pAjliX705p0Uo/XEDQEEDogpWj4lXH0U7xkyaYGeCnGFy9xyh89402+WtlnDrBwI
g3Tw/ApgD2SB5xe54erVzmObf4GaddVtfoY+t3/d5AF5BYxzaV0U8ZNtX9PVF2R/
EXIPD6q2LUw/oySk/E+/8D4o5h7cNjhM4+3ENCVt0/apRWyGJ2Gvj2R679UxdmxQ
JOmFlza+irANvors/FSfCeNjVSwBur9JCmM3Dr5ifU1bGLCFJtBXq9XDPWidY3G7
mLexLDgEb+JtcHtbxVy5TBnu8fdyfbwmucC2/MJX2L3aElFqpdEOpoV4Pvw5Vsqn
NZrtPTA/iuLNrHaDbvjOrm8HRW7OVB8w0CpS2khVUJJJP35s+U5eZw+CMPvcUcnq
qeZt4PvFPBrwAAPj+Z0dsPdl75cGELQMFYsA7g7dMkpWLeJsvx7/Qm1r9Cj04UZs
kYe2zZCRpDj706tfxp26g6cqjhOXUyGcb2Lw8Mk1GFQ2NvHXO4wWhxKvH+y8Rhms
yqmpsX/XAA/eKS/Ju6MQ/z++H2GsWngRCXY/N/+wpaD5T+rXPqJvEydKWXRmUTEx
aFIB/khrBRCivQLAh30iLEtW6WJ0aKMQZRP+tE5UUidA10eC5UoYt6PEMhmCy9QF
w//3zTuk2BgksaEGY0BdoiDVNFZl64pP63YsOLRhOTqah8nUCk3h87pSEFQHUZYR
ZyK1qeYAb7nNEFEgpvDt/VlsAS2TSoAlkCV0UGAPIjrddUR4tolqXvVwmZnul9Fm
/NM8h/8QH2CSI0ogNMKDNHI9MkJGJn6h6N2QfP4V9HTT3vlfIqFSmb3pZzo2PQNV
ZHYwF5Ei7pm2zTFgzX06K6Oka9rxA/59M9CBUGaJttA8S0tSftBiRhpRGW9tRp2O
dyJHQsISfkdU6aCSIeXqvBiOnnghX8K7mFDkawhIDVnUBBY1Mnv+Yo+A7i6Rzg5X
//CppwxEMJc68Bn0Aeb6yeqFGuYqkANxM1al8qt3YJS31OVkw4r1m89FoTTxxxN8
8wxl2SFx18ceicbUfAU+dfuHThwm0cN5qjN2MJ9JxnR9hZp8vrtm9QxhjgAA6KJ5
fW2ihO7yi3YsudX/pgHRC39dc79xhHYnn4tdswjgW9T6he4g4UnMyHogmlag2r2g
5oe3r9j0Gwz4XRdROmrP04amh9tW0pS3g5zTRKk3hMc9SEH5SEkVOAjzaswgiArG
IqUaD8yRVcGSzxrvqyXOO824twXpWzeis8pUBtdu8k+vdnIu8JmHPnav3B9Ahpar
mg3OZu9lDNRYRBJea0N33aF4saH3vyauUiBb7gNSYpQm+QNIRrjdlf3Pijl69RXA
bsjjSA2uFWJSkTwzVYbYmfauLKT/YWhnr8bvjnDIIK3ZbImBuoI+MHpJ8U8ifNZg
uIt2U9b3sk9NaeQIsuuQJ04NxsbpQteDr9oBYKE+3bblZ9gg9JIQ/cEkOQsVE1jb
zbi4Ykfn+Januu2PbnC0HsgA7jeTmoJZWdIwhkVKFvvS00Cjx8I+PHPdYtgCHnhy
T2cI/ApvI8e2VbCGZY1ew60qiSM465drIPvTSJuDdDFC0PiIZHJpzfSgoryh5XiK
2fQ43cGIyskjsnIec3J7OQPyPSbXI4rU1lpn9IY9DSF4JlHf9wJS3EvtjCfXEUat
C3p3+JAqceTe2rhE4NfOZSWIvG4wwNgydB82HMl8m1RHo7Cl/jIkUImFjsR6Fwsq
aeaz1ZAr9Yb30A9GC2QjN+vufCpwpT2xctllHb4arUGg2a6Zg9Ye+zyajNvmpZwv
x8IiHwgGfhe0N/HO2A6v0yksXbuSpgs4uVyVriS5EVBxvxFQIExdBqFCbl7k5ZsU
TRToCIsdlOQWBlZ73zA8o4TS6ndGyKWc2JZHvObvmc+BFHoU2rkcaHoEI1XW9ocF
FO0ygnJ8q4Ez3Eutv4bFfLlukKsMoz2raZhs5nPeMCftE6Gn43LNV9+KNJUIj9Yk
WMQMB9FFUP7HLYz+IgU4WZfHHAKbVbD5ivqC29c2nYW/JzcmcClMrsS9Bea5A0fh
r77p9FTI60EUh4+pVFRRpD4pV4epGy8kmWywTliGfGM0lUMPMWpmYoNk1IHV9KCc
/WVmy07aQcGIFlL/K5MuIpc8gwmhZFcm85yLsYqS87LdNbFIA5kjynhgAIZIHZel
kBZdizZhU3OajHUQf5uq1pVvom7Y+PYUDk9JVCexKCUkEavW8MIZxRjzvuHIr66w
YYKukHPIjx7qSeCDF3WMUqpZWBeVPcqEvV1UH9A658UdcKbYBCxYFFnWAB6GG4Ho
Hs5MznVsWDQ89L6mxeiZXf/32Or6I370m6HY1e+gt5NDehzftUgy1AfDxC+T6uV5
RK3d9UDyObG8iKZDNDJPMIVZOpjM0qA1lfbPyIAPop3G4jGhsAwx7tj0RpScAAWG
E78IcLEyedYWthuxmDT/BN2mQZKk+LYbaDGNGxpAb74go4Z5r3j1f8VMFGHpDxPZ
1ZTXUG0tWxkwoqSXL8g+DL6t+iFATsn2EdFxAVivCHQCk77IKWI/x2rwtSdzlGQJ
VBEqs7u0aGHpW3ra/yTMKN+O20BsdG3FBxqZQzBs1mriQ1gaJYCwiqlRwYSQ+T9u
JpI3JO1/eatn6cEIBULX0mSmf63sBGwcyIChZ95VtDBUJ87lEC32GULuBUPv+Tyq
jehSnxjbbl5jRgieukJLwOUeKN7SkjoSTDOtpCwoRpt/6gflCAh9UPrDGR4nqjWO
6Vl+gjI+NebB1oe+kO5R25YJElm/ZzWGySLk9TYs2q1lcTxnMTEnHkYc2G21maFa
q0q3vnCINcRvWMw08qiynkgdKLLpdA+mNy+hTulY7jIPxG75vTrq+p/XUwpqFjCn
zNfUv2Lj2C6QeR820MLpW9kyNWsmAHLUX9MeYG23AmzS7jlGiCJWjoy8CJWDT9RV
Hm478Az9jAn9k7WF710uolbK4eMd0cqNiqdR0EctlXWCB5ScthImYztvWF4bB9l6
xHb5zNCGFBAmsQeUM3mLhf9G3PRPCix9UUhYAPNaiPdVxkfkpP68DuBt3a8hXf9f
/TChAs/0N6aSInLHdUb49x6/FLBcroPskUnFgD+HoxyYsD5nTDLU/lhB5HkfRTWn
JmrxucucUlhJa/WS+nK//zAzpxah53aCQLsThedeLBaEqhSMSvnLSnfNIUH9/Hfr
vu2Sz8frDF78LGtzu6j+5cqfE2KA2ez1du4cTMkQ15z62dfCAwy8mR73/tm1gx/F
GtCh8w2rMHLJx0lGbcpNNwHHWjGUmsXLlqj3esoIfevEOmQ5VhfHiqcvfGscjuAV
cNQWxVv1H3bUolugMebhA0kOAYFaNvscQOy3koY4IJ0vPb1+LkvO1JX6A7iPJM6/
t1RcphcIrM8+ZKFBH7fZuFGBOSEDxp5WvCtRQm+pLTYL+K18gnXXnluhjDdm8EHi
qYAmHf56uLVQ66+CfjuyEDxcwmRY6L28J6PueJ8fEcYYl/HxIJcmwQ+0M3qFjyb1
TmMZ25KBbtC1sfERupO+AAi2EJpAjTSlwmhBYZ6el/Rh5YmAZxi6C3q+fCZZ6jyG
OL5OdGREBQm3/v2Oeg76Z+jnMvJw1YdOfbNz8fEmqJN640/3d/LPPtQTXl7fUt1O
SLwTkIxmk33p7xa95Ildmvrv3xZAf17QRIp7FRTeKW04RJErJodSLjSTUXNsSyWR
CxiYEcUm6bx3EJMEdKXVctJmWdqOCrxVCvWCSaFxddJzF0AKpx8/WAJAGU7biRil
108LGPm8/g7ELPwqXIJGsAQIecECeVmtdwuaGkTQhf63RkYEK8C1FT39i1cXPPpw
GZ1bC/YeHcB5imfPCbL199fyDmOvdQY8WcChDiR5HqkRGXFY48un8vKHGecOZN8E
GDYc8J2WEW1CMoqK/+pRDWeppy6hZLy1sE9CH1mFlbPTK8Cv60y0++vRxpiev3uK
+tJ6FTZcmgoxj9Y4eOVHwO43KAmFGdfrplUG4p46j0UTc/lrimpo3CIAi23kGDRY
uIunDQyeOiU60Q2lPY8H7pVsc6xE5XkzOP40hF1Ob97HxamLDQ8g3UsU2GDV0zDn
N2Qqgr7eTnk1P1UXSG9Ra9xDrJnAw35ZoiLrPSqxPb8Ga9xGGH75w18PAz23J0GU
7SJWYuvisxWTpv0P14vQ8g5lXP8/5Ed6DmcsnhEir6oXHYLFfKyhEDTDokYox5Db
vjDoncs5mg/HSaSj4P65pOjmYyCcutZxS1jXbLJURiDjWX/7HSt0Y3TirFT/P3Se
uLX98hYk7jTmVS+YrfoS53Ib+ruL14AdYDRzwjzBf38PxJ46qYWf3l3nE7z7GyDW
jZ+6xN7CFYxprwYlt2aXreI7Ma9mzVzVvHzlSmiJZxjpPJkQ+GEdeWolJJuO8n1I
4SzIwgsbBqdQqCs6HzndmPABL4TZbPAWrKa1GuoSD7rX2EOmzma3UT6uVGkfgo7i
0ZDRjKBDVeAsWLZXWGmrnGH5PpTBy1KoEfuQxCBvaM3uRM3gxUIKGFzYN2tTNetL
g4me1KAcoGT0kdKo9UVKOhio/sTQ1uN7dsKljMn2cbRv8QN36cQzxoP2Tgsvnya5
LPBQ2eW6NC+q8X91cFS0ggvvPqQJYvXOJqDss5kcwrnPwIb5aQ1oUGELJEW52r91
utFSCnvpBZdXxn6Dkw5yFhf8UICWdnhxU2znntoZSf6B6uCYVE1wp8pbzgOKqqJ5
sF5v4uIOVzUnuXTOvgTX1em5rBwu4J94MFHMifnR2kK3+bvBflZgtQZGIbtVTeOY
meTiip3vZGwhywKZYDhfZTeVOo52rFCdJQ+XmhglLR2beOyDV0f63LJWgxuTAm2a
bnqv/M1pPxwD0Vqiaq+6X5XORin6hrdGgrFJn+lUlpf/SzTe/xYawkqevhrKeJus
jvDpcMQzGez44uH9xd4kdq6msRzFiaOQZKRazjL/okwmZ1q9oSD4Vz7drnLoSDz/
fJKWvyz6pNpZt6S2GuZw3ckJDuUxvYLAG3A04xOp3tAY1mYS6sS6uv/UL5pzeYzv
xRUTaPAsqfKViBOa0MrY5OF1wCXJ5oPTAc6tHDCZyfQS+t4Egrk4f07Wry0lc2nS
Ejh0xii1Yp8/NdoizXUyvctfZ9aofQyABCu9MkKje08C8AdnUrMgDJQ5B838d3VY
TdHozxm3dsPcMe5VdpfhvlFJYswq5BAbGC+j2Y/7wxGxxyia5AcaPept6zF8sMid
LfJ6OtJpzhMHmbHs/lch3XJG0UVI+kj4lSENQFsotGhvOQi19Oh5zVI5J7UzdB3l
MrewLmlJGVOfa1G8N5VzuDCGxKd0iqf/tw3KHiXvwTpLGSdHExAmwGZQdrMclXeY
3UqyJl4TwsC0Ks6ZcvZRMp04J4XLDOHR7edChsTR+tn4P5osaBvr/WNMTgwe2Tym
jHeoGGlua/MvIxFQXQmVA34/5mBG8Moc6W+Qa9XQNTqmQigECc1AjkvzMYKDBLAz
+IsgyeyYPbmJgx5MAOK/QGbUo3Y07GsL+cLPN09FD4D8qvb+eQqjk/bjJLS9/frk
oBLyuSSPXZ9FxkXtGYqrq60zKEw7d5RU6tEPczHbGIUqGPGmXQxORCQ8mQVsJgqM
yAIKNCwTJ+voyIxZ0yzhDjbYA8omaSebSNv5NXa4qFDjTdgU16ktQZIxRvH0UZIs
LLTOFosdHTQxKvrf7un4bnC4VvSDupfkbz2FoGkCNydhJ/BFthGufNjPdfM3/PXb
5NSBLCoprAXpikPyokk2xqVGVzFga7+KL+643mc3JRhx94+tfMPZjrobRVoJ0CaU
JcZYgNSYhIQmdHeaY0ai4LPS7c9qa98+aGGyV5/0YLcDHR6u8irnIiyCe/+kGS25
yAGn5lodL2e77eanmEPPqteqv3JuF4cNEc6XkMLCkqg0WoHXrB0oHoIWWkw9pvVC
07WFILqsggK5HQySzQ6PsGEHh31CEk69D5OJ3ruO4Wnec0nDbGE/fySRrWv31IdE
nfdfi8JvTc8bTJ2EJrhluCxcI8c2cFzoKI1ovHxoLgJwpyxGO6Mj/H8XoR1lFrXI
BKKz/3aa3oFSc50UgbP3+QPoJ8kM2TTrKDRUwPj/NJVVgj2eL2QswAkSBUREU/Qj
+yvrKR6BU6JC+FTdaV91gE66DlDSdLc23803SP5oZisEAJiBBs3MHb6aytfB+xu2
Papo4atUlobGrugOc8P0GwzlccfJlSG16yEERWnjkvivy3IKYnLXa47ku2ufcUH7
hmx4TDCIY4ODimcVl6dKLr8w6+LvOIyRMopTHezhnhLUgE8bRRblnKROUZoCbU+0
vK5ztaVmSsc5KoY7D2STB4zdzMZ/axNNFM/sLFC8LPTcttzCuucXRYMEBofd/AYI
9TaJxEmEHePUVM+Wo31TeTTuOkkuocS3k7rC0RWv302eD1zcVM3anCvEDnu517vZ
9OfAeRx8QjO6yT3iBJ0jJOHvnTQLlrj3X+WF66JA4pvnKoKZSdjGXVezXB82Yfu+
KBlRUIKXhmyKWHrArDcyPi00vAmvjhpiwzHYVfUC0AZcobwIoyVeMaSwAIXufWC0
ssGAHS0TWBb4MyIOt5fawCexh88S7r+Ht1mDc9aIB5ffKjgtnjfnkk9ZZxWNZ2/h
1zfvGDBf1nyYr3YEQyzt607gnMHFW5eQtuo9u2vssMlHQHE12R8OIJTPpgNBzMnY
8FOa7/jgnsuFFB6tuVXH7iONC8LyD2rkTfUop8F1jKv3VZ73qfPfoV0fPIKkxKgU
dCwbz+v60P+KTmHy+j+WqqLARi9RdM9z9/ZIKu6uXczju53yMut7UiN736+SAJcR
PirFNnFtru6kykFgqzWJNjElTHu4ZUd/yxVCG2uMSlgimDAFcVGR+ZT7CeiCVeeD
dP0yoinfza5LrdVbgkxBhKYdmZBeXQ/ln4UsSYfPK3YaEky4+CcMwBgINoGEVNkP
6egmTQuPsZ6XPJNffzMqol0aE0V7n1GfwuLDkU66XyDq8l00e6nAGGh3e1GSV3B6
0jc6vN8LEy63y80LF7oEdWD7nnZM4zzuIzuIizCNTlTl6STzHhIpezBE/ljw2Xnb
oW0g6uoqf+GeWQBiALaiMvnGxTVkd2gX0tLnjbimKAS3mSNRsf2XJiXx3NnxzVhR
/9+V6dSZA89+LfAhhsMD5zJkYOWQgFd2BeXtksvjRXWtHTrOcs74pI0e6mTc0CZx
MFfBmUCwv6cmeS5g3T/NN9WrKZmYbjHlD5gPXGo2wT3VrP0PTf3zxZLDcIMEDcuf
RpuC5vpnUInl4xrC/NOyoL/BO1v7h5+274peRkze5FwHi62+lk/2gwr6lEzWQiWz
9MZdgWRxenwrCKqDxP60gUjByUgovFfjgE6C1d93fW3kZmuLzVudklo2bO3eVj6A
MePdraf7z7wCPUz0SZ8YX51bhmukJri5WoGdN3+HAGdp3cf/fJ6NI3sd+EUQ//9Q
levMgQmaUh0f5Uo0Mxg+67wptGBasNgc9x/XjbJHl0yprziX1+w9jwj6eZJSeQds
HaB6sXWaGtLxmsFB6cv2h6vzkY7hBdhYL49Uy6p5eu43q9p2MJ3ian3EfnnnEils
1Mt4m/8xF4uSOg9NIJScOvF0iqortm1ZBJslpY9OoMwqafdq9bcQAQeN0yUFZznk
xRZpv2oV+CAgBtfUrma5E5HFkGV5FDb9TfyxtjnkqDcdV+ulYnAw1z+n/dL177K6
LJa4KEQdjKq2GIv1CYvxKOKLiLaT8HmmvSryjQiloeW8CRIkScQ4KT3lC8Llkjem
eJBG9wMW1P4S2jE7bqILRpNOnDvg59Cj0Zt5Yw+xsWN0P5kPOaJMlCevB/Ev321p
nPBNlT9jzv34ni4Fzo6GwVzstb2GPnsRCC6dObm6pbP+uSkldi9vkpL212kA9ZIz
7tRlslgYhyhYiJDuXvIBpGTOYtHPSDs2YMkqDHWUQ90XeMKpQKSHzwYWN1neYfzd
TiWUlC9Ey/pxlJjJzpXiRXba92Gd7svAMOWmavlvBtftil2tM/Q2IIV0pM2InZ/3
iKVB54lsA1DwZ59+kZPmRItoY1mbPrJtWYqjsbtDYciWBA2LISXz9Kx1Odbi2gx/
b1WLgbwm/sqWFBJuklAvL4NBkb3VdRyZDH9feklE6MKkscxiJuPpfODdHdJ+lQFT
Nge2i6Fb6GlqglQn39N3XRkURmcdF9xbxNBzJ7wKasbsNey1MPQl6JvEFWwt7NJD
cAORiWLXTgWHsdw08ynDs9pic0hg7TiFn2vYAM0NNzIsJ0EHXCZaS+dLpRUgjWUZ
F9fHbcjZUWoKCuPQRLfP0XMBGhyxqJmwg5S6kzr6KhEd6FCwBKSSM16SBMsE8LHD
fK1voE3UJWS97s/4OwlCW/Ytlr2J4JxqfEZODxiHbkXGH2L9SpbL1a0EcWeh2Cvp
4Qv6lE0+NAfDwrkkzax17HRs7NNcWtKnl311tffj07aYE3J5mVppPGGSqiZ/Bghy
ulrJwkP8YI1xBchT0a1bZVsWwR5UAEpdPN4aR5KreQe+nBl57+G+dFj73xlflCQv
yhNu9Ebp01K7JRwI5uLHdHVvx9wuGzWMMtoQ7sT1wwkkXqeR+b0l6ZYq4OKBrdzT
Qm84IfbyoOhhrpxfoUNegKLXYMhfD7m6Cz3p17EOzv87TXU0hRbKSrZWeKywZqRF
VTJdW9kitG+mR3IfkKXDhrWpEk/IxJoIbH/hXq6KEPtmjxNjuC0XPWG3bSMoMd1D
9QMVgss3iplGTUQHz89OWji/S9UlZksoG1HZJlScpGN9oOEFDiRRY9vLRK4LoZz7
TIKvlaAFZWx1/p+pn5t4hNOXjInngYwvwa/9FQEN4UrgJ49P+43KIgttTljRaOob
r2ojGgaHHk4PcvS/JbI5s5+L7Wv3u9fus4aZf1w8HCX9mFiPU99q03tZSn8qIcK0
yNP8EeJb9LbU4Ng3LXgRZF/2kwLqMzpkHFelm1Jdqm+tmIxM5rs7BTPj975nt5zi
IB/4hPvM04B/CuuLRKONqvN3Fys6wwUarK3QlNSyM4x+xfYPALA/nzpyWS+3gWRa
lgMc8UjWf2eF/rj/Eev/DLaD3Bl3osiVPXuzsjmLPgJrO+RZNklRemF8JNKQoE6O
feopLoekl4cdlwS+hCPTOqdX5yg+RN9F+dAq8vLXdpOozlI0m/eO+hGxzxP5bM2B
KpYQJoQWrlqdb6iLCgtvcQmKsv3pnS4cWwEoG4siDHrV7wlasE5vOF+2jA71nNAA
SsQY9TD40T8zMFFOS/goEqQZA9i96g70NTnmF0VMulAO/qhz1iVj1mf130z3e6cv
ztZeXaGAk3W7nkNANVkeJTvuvhPqa4RGRMfwc6IQpoqAtxxwIcz3Dqk2L0LdHJ7i
RFHRvGnjev+/Hc/srUBeaO/lBCiWUDd3vsDT7omUcQsVBWfru80YBxCkJbk22/HN
L7eVSAenXiMkuOnt5gMsMcbvJwbzO23UQag89oMRXKXSiN02kgzPDcC4x6FKq3OY
6n0pPHt0cx2ltO4lb97r8ELjU03PLU9Uk2tba0b7ZPFn1u1KtQoZcZugruFR5nXn
RMQBDe+Pfb2xqU6JJblUP8p+XlCa2W6MLOo6KRwyTUXS+w6iVaqzhXbpkgBGWB0k
2kE6iGQK+bqXjB/bI58YQWQhqK33IvrH3fQ31Kyf/CqvTwlYLhm1X8exZSFgr+aV
Rx/GDjUGfxLe804d/8EC5vOb4BJZX/APR3uis5HMBKmDxQkyQtu2lLgWov6CWmES
B1nAo7Hc/Ou3AZhIQkP4ktUWBSkR4tx8b3UaNOeTkZWLQizcOI6xBwDithP9iNYi
mT98i5MZ9c04efig3FEU7k/2IsZy4zKl+zoNHa7v4qdSJFCCXC58ZWxJBxfbspPh
zq5z090Dh7bAnBg2E9vRyDhkGV0QA6DFkJNLYYk+og6yLsuFcozxLqrPqsuAGVrA
rYlQ2KCzZ3y/Ma+WVTjhFEcZltBrzzZKcPq+2taAVHeLFw2IHPqzYTIE4gWPF0Mk
ZBxB5jiCUe0RgeJ0ACqeAvTxUQH3c+4nFpSC9lYAORbnzlt2xifWIcWR4XSI1C5L
a5RRSfPUxmGpl+8G72xtArHww2O3ZGc23OcbQBhQKNKdWKxunn3HeXRzjikLfs1X
vJf7uvlUDYjHq/AC3xJq6BT15c2rrl58m28AH/1XSaCTmZ+gMZigssQdgDsTZ11o
bY2AUz4J/7+dLo7uQdQUBep5xW2zLvr/8LixFX6bEu1OurYSIGsxsN3cUCjRqllV
Y5lbtMEUjhK6quMjpsMreWGOr4tGy0to8U4YkArU9bndmvrm1GzxvuS8yXPc3tcU
5iGHPNOKNe7h7dNlpIVjT7IN0i2jmcM/0kx4EiOHvT7FfmRCYCkM0bpfu7x/Y5xH
55dvcNTzj3/8d4lIMf4UJa6eJ3oMn/R63H1+JuNqZnPlnGyJWQvgGw/wgxczVHxm
rbKZxedcTs+0dahA9qhKlxVUsYilJEAklwwoebh6X6zXnAYy5bz7u0RpleZu2dFJ
ze+VnQBBlUgM6JEJ1zg5svffzpGGB4OklN0RAAuJzunjEUnHVcMFBY7UJdnBIgK5
OxJwEsMqCL5X59p6a0WNrMPB8R0bCLRYX5Xdw+ESxPuFXGXbxc1YoUJC/eEm1KUI
29BrCMtqB+/bHHE5wscO8QGDKNCU/oIlnKHQ95uqLGC5UEvF07qaWggmzLpHW/RZ
w2q3hqufvafwpzimJwf9Bx1MoKWu5Ho7z9zG3b5R9DdEF3uoc6gUDikpktyg2B5c
mno/XjrYVfiPU45JTe98KGf7obCHGhTo6MfXGU28DsxgLKItvsI95sgm/lzItLPN
o/zGutmGKaZGKTo8Am8wUnZlvTB8/rBufRulPF2QqHwRFEq5Iv6K2Wm5QSjKPncl
TOCxlphd86MCdewEXQvrdCNR86x53YmSIuZydLENcdSPSZN7OxEPE6HiRPh9E0K/
I2UOLjaaKB3e2L7mzsh8bdmZVZ6KnPeBHDxOXXTN9zSOTlg+ZqfjnCYMymx1UKKM
dq5UPp19NOZ/vjUEqMBGDFcIBGN5VM0C+IoCMGeEoJM9vwEpoByw0b6xSJX3DWkB
qj9edC2GmoFmYj1LJepZc0ibKFpNJi4Nv9VWe42vPUeX7R9wV+qgAn97IZ+ENt6t
L7AXIkD39FxGVhMCkOS28ebbHdb/8A5gh6drLl6LC/TSzHHvl+nWyBrDUtH4qa2N
ZS30qMJitCJSwJ61hrU2Gdb+sEUfWJ0J3SVYXdi8QYNcWHJLs9Hj8NgGgIAgUE3Q
XAQqpRV7dLOTfTo1U+B3zrS2a5SBdI7GlUo5/OQf1SKCcH9rJL1gbTlRh+HM6WjF
HAuyjdIfsCWWtBYGo0ev1F46EJLgNYHabwyjEOQAneGz9oYnDD3qgXbOd2P0LB0B
Ez8OPqGXMwx96IsQ/cfLY7Iip+Jd0QdyiUqGqfcDITilkJLX1RQDtyFJ+YGlAy+O
lqfOa49+TtYbja9qEWJv53gxRiLMEXGra2V1+YrK2tOWxgvY7XxvILmy377GrVdB
lBe9qdjRorTLCmrfA2+iQTJnayozp4Fi67YGVVOjnnhjAhAlWyyYTl/CLockylC0
FFobOvqf5saVdVw/tPS1K/fekr3opG6yiFbhtqx67VcHy+7pmpE4/b8bFWTjINIK
FOD9Puwpg+W3GnVXFi8hLUCe35PgYgvJC8oK1E+c6YfiFK8koo7eZ3tRi/jFAFyr
eDEK/AvE0XHPVHZPMBmoSdvryG8BsYbEKh9j7MrLKmDQZ/vmkdc0/rkL0Qz1SyMx
kZthUO4DgMEZQWUQl5QCzkIXVED+ML0IFdbI35xok8Ka9Q4VXUrKIvdt78C0NYm0
nSwMjEjZGbkqRqLaCf8OpQx2YgYr6t0o20zt/CeoiYV8Nyh7ku4+hf+91Vzn9r6z
vH35JrmrUV8kc/xV+xhG1UvId82s70b4Tlo/H+W7M6JAheDNXnHTBnrX2O80oP90
y7P8t2eKlTuGYfJn89+BozRV4pG45wbLDMC/Ad18sNLMuzBVu6uhLfWknmTIAQZZ
epij+ML8EPteUeKdn1OCEzgDf2fFSPQOjYoPtGLthumSQkHvGE6P+UPrJdjESI9k
YMSez8t5BhG2gW18ijZs3Q+9plUww/RIMfTU8/BnOyDLWUhrrnoXxYUVS6svD7HD
mQHw4YF2DvJdOsmeEER3TJ5nXqJAmOMZcDIcHFfavKZM0U8zg6a8yL44yUvd6I20
JM7OPktv5ys+aDEIdqgkcfbwPxMbJbFcZFXvmyDUEcGjRPhJU4Qm7z/16yARsHxD
3PsyhoxUImYTm/IBiVWFjATEE0E/wFFdbIfKJtTW3ZJ2WTQrFcMXDpJ88knAHJac
9nSzqnRgI9UAfjqEHUNjRe43jQrMa2GG4ieygAAMJXgOdb+zSHiPnqCw3/fU3dm3
NPQgqUGNcnxK4b8Qonc5FyILUQ3FuBCEJG7W+4tVXbiPfvbh8aE4i4jcOZ1h2uWP
vQwCzoEHT7GvpKQEnU5VixOucJVB6N560ZwtjdkkivkcQjktEbuSjz4O/4q2l62/
tsoOGBenWCKup1QQZkq+iyZP1JNEqtTtRUPs0z1d07nXOYmzmkBCTcmEzHJ4Rws/
IDijFveRM5GSXjkEBDuhJAyruoJJD/7Bv5KY7xVqN2FrY/+tLtQE8gxtd13TfksN
cUcsw5d67aMppTxvyH905F4LbdQI4EqCEDdQBfz4/PgCON8dJ2+/SZtRJ1Ia60DP
XtWEjs1//dKkgN+SEI/XZkMagv56wNkuJBI4zghK0o9UAiu9bbQvIfzQecQmKFvo
rENDwqxzoB7Wpo5bmLvldPdtW7QN+HR3lHImqqpHNA85FbQa6rkwi0O2QP5kxNHV
+X0oCrSKvD71WnElY3dMNq1n+Um5RyChmjs7lHKDQ7C6jJT7mfio9CXmT6A8ulXm
MiFxS9lWhqtclA5QFl5NatzsY8JlO8634BVIddC/92NgGsLgVAv/YHIBn6m4YxDm
5F6KkiVab/vDOLlor3sViPjqcFkb+xpvDSxvQZGEcnpUhIRhMZiiH1LLpp0E6OGI
0w/S7vjLFGvQ6MtKr3xZL86D7RgsPybSUX82jNn0/fmQZfufIPaGO/meiZqD6Amn
jrMZXKkmBHuWx3J/db14cOMwRrv3C1q4PLb/zHODkkvQQ17NeMkhTfwKA/F0ICX6
CCeZAjbXn2eEYK/UYNZXocJvUoZiu8w8v/uP+6imJpS9Iphsz2r/5DzpLCIt69Ta
C/uNC9ot2A1x28oybwmnJ/IhmQ1jcCSVlxhhoiy65II/y/h/99sJnRPwv0+Njmt4
cDbg7dFW/BKADw8WZ5+1cvA9UmBeqrHOzPQSzCh+FrGVOl6hA/uvFK2MEo4puQRx
u7hjYmfLS+lSQQK91wf2Uspr4F3jEh+D0DifawXNWV5cAhVqweFgXbO9trXjjdDB
G1qjBj0SZpnI3ykYK78s8Nk0RnCX9duvS3XR7xJ8Cyn0do5ILmS9m7WzXT93i87W
2zUUb+hbBWybwrpNumWBR2IrMEoYZcxF/Eeb3HqS2HITG9eAnoTsibkParosjTym
R9eJ8sOiG5RWa3zoWSu1UrncA4tv1BA5dzI8fbFmJJvzzI3OQ63Vm9M2KVa6Pbch
zTgVdtR4vQz5I6jQdrMQxMkf7gtgQu1cetoCSNiRVs1WJyzpLetE1Q/Rqo4bf4+/
qJZU9CufhW5S/EQubBSlwexfXf0XiLP2K9WlCZbzNlxoGrc5VrTlGMqrtNLBSvjM
Fp5Ajj84HBD1KYMVmaF809tdRE72Tmt64ErC1UFuXqBQ2/6y3Espc9StV8bx7Vgg
Z/2rmaz3LCeJBEOD7wRuylJGgCsfdLFx2Ny2Kfu7VoEybswD071cw6/FZvj6nf5W
mukb1GbyIcYhmr+SRnx4Nflu0zzSYWLILtIxXamT3xFJqB4PiB+AQQ1sxN9SZQWj
sOV6oqW/yvDb5zprdcopVL1Ug1sEi4u2uYiGEhuyusFfuf2NfqkO6zwTVz5JXK/o
zdYeCW28pBK5WSNzG0ESw/gmFy6Ezs+mbFar8QXj3dQ6Uwf5OC2l49JtZMERp0UQ
UAJDVK218kGi5de21D6H+gRngqpOVYOtTBbfg38nSsMTCPMnpWnLBikLExbY7pvu
jUb+UGSgJlAcDXJBgjS0EyMyP33dU8RgWmUJjvpS7GfSOQ8lJIicc7mnUv5fGpbe
gO6lMPIlBAnRBWoRycPrRNWhzGVEDE3iMLcXczeSQuYu9k1Az2wJ7DJvJesMgaXA
QCIc/UtLDqlJBGt1FfX6dvzT0OMAjwfntLxsrIbmTSiNuXkC/uPnQtIxqKV4FpbY
CO8mSnoh3UAmbufTf5AkYxsJuS3lJrBrwLxe9owdQZjMpjFp9y+eWKn7du6uGw4K
UKMKTECfTfaElpMDm0r4zjaO3zxuIUmadHwoorQJw28brqwScU4R9tzsumXrr7Jp
e2AMoT7BkRSiIaK6jDUA90VNd6czPRXmpcxLNEIcj9LMf3RyZ80IRTx1o88HDPzo
+uC/7Swc50ByYe+PwE63ONdUgCxihGxdDRsjmhTiXSbgW03UHVUs3e3jytUrn1jY
U5GxUPCh7FmmMhqWnGeyDOGd82Mrx3pQOzFTbWDEdHs2aDkoMB29ghsvI0wEv3YC
/t0+GzuKfR9SH+Zkl7blGaydamCzHVZPZ0t7+yCaYEtCks8Sfnr2sxBJAkMTe144
fxU7tJQUNIYX/T/L1dkxUY7KKU9fqkBwNxVlLPyTzCLrUw/ooeAxbWwhkID2Kd3U
1sadqkVvbyF4TxOFEhfR3QpKCjdtpsBpkg7qGoYWhk6Sk3Wv/6zKnCumkRZtj/5e
5N2hWYzXUvmoczr/NfMZQdaYJZSzsXhEVcG67OTB9HLWnDtDg2079HqWgPDHqj1Y
TfYI1fIc9v/u7RDcu3rVtqsQnwgxf206VAruJDt/+lFh92ZhM61AsXkU4+5KWDnZ
/1gVE3LWBP1VbGi3MwrljJS7icn71+IyBs5f82rc5kmROfulQrhTOWCSA6Dmj9yJ
pUpbgC8kQpTAxxoMYlKHDlZ5hJbEhQt9Sg37zKeSIRIbnP79lL6sWzZ2qx/4pcVw
euPWSy2bNN0HXYPiFKTWdfvX9nn4wqYER4WOp6tG6TY7vKAo9FOz2UuzNytra6SZ
LBsErKDvCJT6EWiGSDzS+rjuROeoDlnXTy9Nc11J4nN03SuJQnByfypm3LSbBYvd
AapiFAwMs/UhGNptnbaDcSHzZIUXXwqUpApnaotuRx318xfhzukyR+AubbhBzKm1
LvVsIpHdVO+mRxKUvA3Hze+cLROUePxNT9sFmeyX/Ki7UItM1/Mvg8nEr46YJmK9
3IaoX+ykjTKk+ubL4OoeH7Uo/Ltbmo5amQ/a5I7f3BYAdSg28DMyaHUdC49JsVsk
buCSNAbxOx19TwxWREJtujCcXDoy6050I/UTWkvzMMR10t8CIpOFlKc/Wlk5IyZe
vGmCLVFhQeeFXsPcMJapo4wBowtwWg+sJQ8krOOEmgTMik1mxK260ZVrJ+s7GKs0
Jda+LHH/Wmp+yt8c7B3pdo/AHA6CZzB/HNBA75ANBGRnIERfxMll+UKJwR/AFe8W
BXSnj8uW1mwPYs4w8osVLDUxWAPi3ZG9EzqxMbAGpVAgt13US+Ln37Ki9RwIbngp
zNEzbxMCjYhWij+addWvocQYfj+2inZI8dFnsHGQinqUIECPiE/x546qfYwKOPw2
9YgVzPbq1yNY2uApogMkSsZtcZ4a/RgVtfGEqGCz//prnv9Crt9NeSa6JPMv0hIe
0xhYhASl7kKQYftuKUbtcP7Z4/aPSr4i6yCAzUKvV1Ce0cEQe2yuK3A2rzy2wcxm
XOHyS41Ys3pL4COfdo9Ko1AlVTSCsrclCSfn8K7NvEOHCKLMXOHsVS0iTyqbAIBF
krKtFp81hxdUFP0EnF+ZlU6vxGOin5DjvJl5Z/B39IggSDddMIYxb17WsojhyPrC
8MzKaqynH5ma+sMpVPHGEiSkZtbSJDFU7VpbNdc8Wv8nWTTJW0LGphjZDKKzVYeS
RqHK47H09tSn+z/9lcSREd6F7GB3R4xIZ55/CyonEgDm6w71cbcpXP2oOABqxq0d
kO0PPNOFUm3AKzA5qkNKZC70hWL7ZqL/g1FmCX5zsK5AE0TQEy7qc5k8K04wM2dV
uh7HcyT0TYMQFX3yKWOfr4LhNBmOxDWJpsKjTYGzbMAMQAQwC2PEtDfe86MbFNDY
OHfcG1HlkxPZJbMvZWUWYzYkq7BMLvDn5OIYeGy78xg6IvYMggu9kra6aiXJnWEc
ftTskYaIXMrulpccs08Yef9oMA2GdFqmJBhZmQsXmpkkspeDzPUMvSasTDowL566
dUHKZvHXYfH3g9Be101rk/U8cRB7YEonix4lkTuM6t5JiVmecKL0CqjiLAoJJ09D
6d6G4+TCA/wKs29rXo4dnp/R89lEHtdKaaN30Yv1fX0xyWFYGCoU9HV6FcumtVU/
oKSAFrYai/RjZfOAHf4untXOqHNkA1y+NfFIFylbIsGle5mRPtDowGJfd7QEjoER
59SG0Yb2AxKwAkZMrk5Dy9eqyP12lb3O1vSuniEuHg1LO/0JTdrkkb9Ykwz8LxtE
Fe7HPQEw45w45RHOI4AHSB498qJWXCOUEvkkgPT/HJW82Trzn79Xzf4lTY/ZpIhG
c3bG0d2j2ga3lnN3bdP/ErT/QjJ35ZR9vnFDXBebTg/GMtb5bpCG7aDH1NMy6UeB
6Rjdl2Bxqx7X/abfL5rDsqD+vXAeRbf/JJ+Qs2bh4dBI5pHxoFyysIhtr4F+sLJc
DYRqt/YOwRXaT+xbztmsaqA15fWuEsjLjW/A7M9fogSQeBlrCxU4epBUiOIRA8Bp
1PPPnwqzmoYBlXiGIgruyXu4aiZMOq+7kWbE23P9P4a+Kg5dQQqwMEsxdeuPY7SS
RQiqg216Fh3Z6O7rvYKngAaU9OZ+Kvz56xyWL0c1KHlll01EmzzQvWFCZC1EthJE
cuSeIkIjEEshrV6qQoPUj6HJ5+LanCLE0pKwfc0/wr2fFh8UOOsO+mSIECohzVt3
qkisb3+l+Oj6OJLNannyUzcX6hqdBRqESON/papCrWYgGRL+Q6n7/pULPcZ71oFT
OX/qVFWkvcRPUK73Sd4DIBD7H8LHyuHXBZQroAtiDr75txbOtLz9f86L7e2JAbjK
4z5uHDnmJaDizMQurDV1fOHskpqz6mJOkBigF/QYY+ClhxGtH4BN2m+AmFsNkNOc
NFVCilZkqrHyWkRClOaSUmmbw1M+uMIKoi98GtS5oF5VPsG3hrQB1x4qRwkVbNJU
QOWOHhYPzyoH3ch59XCbJnhKSC9kvR2AEAMLBLucbfFwkrMy6eCSStLLpfaPvJk6
0hHV0xCzpx1LCZZ/2JDVNpqpPY5FBP6V7939QFzsl2VSCdj3CZCo3Gu1pKpxTSln
8fT1ommdEzDVyGydfQNz849U1TXTciq49Jsi6Yyo1I6+9ErlfPrwyDyypBfXJ7y2
1AE8RFlJt2UaEE3fJ2SdAJ+KdApYQR5p63AsdGJe5fVmw4J/Fc6Zs8omsV6r40KZ
7ANJtTFXMDLW1Jz6dhE6qXiIV4irJ3xbsl+px+awqlAs6aGUNYNpT+WtPpOR+04R
U4+aViWa7UXUpFOqJV+zagO+2mLBzqK7/4tXv+seBqmP7dVqiQkn/KhOW0/tmsAO
7hjJg9r5LYjZtXlDaNxtk+yrj9ftk0cMCXuFclyggJa2vo3awNrPV78KuiXikj72
GI0Ic4TMriQLh6ndk8XVcWj665ewEAKUyOAUdTjIUaSbGYk5T6cFGbKof6l39iCf
NxCEVL5skB4LAsKEYNE78DiZr2K3xdrFcW0GFppH+ARUFLIGNL+uLqzA/bEJ3+b3
aRekm9W27xX1lPCuaNcpSf0DWZsB8B6Td5aQCtAa1kA7gpGIXK+0ajd2hWlUhrXK
VTKDRH3bc7F+nVFrUFY15P3GXi2IuQqCd/4BQU0e2+ZimxqB2wCVA13g9m9yYUUT
apvo++S/8j66J67yTp+DkG/Hq6FuMtenzGDFk4trGvLYBvyIWCrDubm4AtA6vGWK
kwRgEdIztNUUIgGxrpIFh0E+UMSOdBZHJSfQ7oOFcJ8E8U1XoIiGqst/ZT3uThV1
i6W7s3TMIgeP4lutfJC3xiqndc3d9+DDj2xGEWVlAitOP0SnvLWUi1cTRJKbv88p
+IiOx7TRVoIcNZiWDrbNwEkaoC6Sccy1zA1fv2b3kykYOaqjej4YhR5T11pGp1E6
xrhKEVWKCfN3PgZRxqEJIj09dz3sRGyAZLsN+LHL3RL9UsciD2DulXoeCGjJTZyn
O7jM/ZUfiGpNES/ILsrMJcW+TLoWsJC+BSGuxpPO1V1fffRgNtZbv/wcHUS08IAq
KNCzVYCB3/1iybn5EvfJIZ4RM6YV5i7QbGL321JBIghukcxDFeom1D75/jNZKvDt
oR3N0CtlSSU17ExNcBcW6cG/11IGZ3/pR05wOLxpHUJzRpDhIpwoWU21ZvAD4173
7KueWHfR+L3IHXpDBm9/zIwJbUPAJz1rW6A5mshUMNKU+Ar51/1UPmKCswxraMBf
otvjdrT5BVSO6PgNm+p2OVphPN+BjwbDtUUwWLFRcoP/9ZjwS8QhZpPgERxqP6rP
qE5/E3kIIu6MaoDGByzPKvCg/pyB4KNomwTtlFIDMNiP5UDz7PuODGwNIU2mhpLD
/r2Ofs0w00hI7crpGS4pf+q7a8Q6gHCjIYerSZ9ymbj5J/zl3UmvVRMtK6ChuANE
68FVsK+kqXDmS/KoJtPx3EOgH38vKYvBwZF4b58Ltoh81/VMtOGD6QWZFx3aqDBN
vrXfR2HzTiHsNiSL+v7U6qyJCYzXZ+ESTz5XX6sf2SSrlxOQNeEUa0LbzPUQJBUC
jjR2f8sCs9UiSpZtgSO+MZGpLBgr7bSuwA3Ln6iZJrCTaco8liCctm5TVH53aD9r
YW94E2AfDeJC5r0PQWWoZJF1q0U8k7oQeIi0Oxm0+0XVxc2+k9rcnV/4Wy1Iy2sG
+vA8mPejcNZHH8fC4dntDsOeTgtmddD3SVnbXSW2IwgWvd3sr+HlpZxgJh+l5IvP
sNPuC5qvD1KlrcoE9yKdJQ1ZpAaX3uaTW9VhhWhO1X/U+0sPoo6E5D8N+G8qT/KN
cWijE3tfoERFWH2pXW/hljsYzrLuxlQbVvXyNvv4C3SXfYMmmXWkcvlQCVaSRejo
yupheTu60V/9vowfe5L6vJjrtDb7ab67AH39eVJj13GZb3wI4lfKH6eUinkXDnUg
li9TAdhfJKDv8YQ1hmQNysZb6DWm7MrcMm5QeSX1CymWOY5n0FAsrxLfbJNC5V8k
y4LKJh/1m3237zLeviDU2zobkxtaPlUA1O1/dIN4stPMdXeqg2jV4nDgYHe9oHEk
K0JqQFEHbgS+vEReyhh5CINFtwQzHpQzqSHUW+MlD8i/vFgA1X86pm+RmHHaxd5W
gU3g+7WTLEC3/4JKIuCx6LXs/6vqBb5UefTKfoMmo9AM4DkDHRgIoZVjNoEwJRhW
xYdIM9b0bNXLUQ1RowqZlhw8dk9bQqdFgPFprpzMJsCYE+ksSv20I4h40I04SwUe
B0sALShkwVthKbk7m+ygOA6PUem7iBFd7u4BU6xTlrJw6ko5xdfLNFN25H7gIWLg
kCbrwOAqA5lKlmj6XMrtaaFLPPHPLrfE40U81jGkAesRDn4tSoiH1VbFbTYx4dF7
XrYVcT4C+UFyMFD/icH+gatfrQhwthvMs9El3byPUX86pqAt475lKhdjxe0u3Y7t
db7PULsgTQU0/xyJe4fSUOdE69e+8LLz9S0+xf/GJIGbPBujLnRl3nGznAXfV9D6
fio9gLN+NGox2ILRx1UrWzkGwfrHwsfEnK14AgG4ZLM/YlV/7rBmGyOAMw3u2Aex
OnHKF8XhYEmjop3CROTPxyHmrmSvix4BRNpuddwOZ756Y1jCHoj//yEgWH9c30D8
SY5NaNVEEIEtn07KRrCWPrmQMzxoF2x9gHSx95/iPEUas1ON2DcxNui5VVUGxZwV
nY6+AGaUU1KjAm5skXWT1Q8jHwQvK2Aegx6xCQ0R2DNyPiLwuvP5RbGrGYYyJPYL
LXa/9fes/WV20/9exPB+NBKbir8ly8IOylKnVSZry0jXv6YFfkJTsYxPDHtJcZSe
BfWCiycF9BmmsIa2FAIvpVbmxGyCbeSRx9zAlC45rE8UcuwDQao/UO+yYtbpT0dc
q0DGdGeGHhBD+swm4ZsSYMiXBD0yI7v0urwR3a6UJxuU7PEcGLrPPxDwArDkSzWx
67RuenDwFGldd63DCuwhNO8+jdFMggIrmPncZXwvoAVlLpgpieKnDbkywWCi2KxI
56qMDwi2du1/eYW6Av/BQ42n6QJncQ/T2h5eoikSs2B2tHdYnvCM79wvp1W5onQH
XUXwR43D4brGZEUe+mePxvi7KB/6mD1GArljNHmA3S9XP9pj6u6obg6ec6BvrgIH
8bLriphDKh6MVuBiHOAEQOJl4821iM04oycsfZgSCeQKwfden4fQrvADnGbNFoFo
dF/1gdedRgfrvEDi04lMaN2HtmwyO1lGM+YNnbIKOE0bs8k5Frtvy+Rquls6GFxB
Hjs+wIp4H3rxEOXfpbrvVyKF2YLKonfp4aYAOnh72tj1yH5rdMfOtOEL5ufq7uRl
/Y8PyQsMhVM/piaZPu0lxc5OOtKG2zQWqa2G796T57+QbIdAEaijty9LdROK7jBy
F4HL5RrVJ6xEw8qxR2qYBtekSOGiQZKqZy7PJoUOKQ6lSv44P/57b268VGeqBCA/
w2CcpoSzofo8Zobx6aMhZJWNR1SDxy47ix9G6xZndClOFoJfgDCWpyrxeFRYrQGI
9YJ4MsClsy/buFdA5cr+1vs5VhRodSqgWSE5GcUfK4cD8LHI9ZOQc+SFeezP3/HW
wdJGRFsRvdCnsmob4bucy3wxZod3JYffm/pPIRhUJB9eIrmO182d17K3NW5AqXXu
oNFTMnd8k4g6SO2FKsHYzAAG33jzrnr0ydZ1TsbXo5kNP4KjVqk3NJiuC6qHqhX4
/J8thrTQRtDnuA5xyZD+6SUYa3lYmYnm41zQRMSoj6gKWQf6kCO5Hzddn296uvQR
bg8cE7VxIQfW+23l2UvYWk50zozHSAbJgTNSgLnC0+q6uRssPiRnNbQ2ZcbN2rlo
JBdjFjtKYfnsMSMkSG9d0UuLbzZPXBCG63GskWnTuOBZBlvPb8Dko18CgNrtr49v
cOOZ2Ndfg6y8sHPrU1z6htQAoDKmRYgvetZoKZgYPRp/GLigCWCQw9FiQGt9tjw7
ZkP8aO8KkoYnMhRlwpW5cNVC8ZwU0vJumafLoARfTWYL7fdLYsYd+LTeyvQixqX8
n6CU+VhYea2Phe5bXE1jCD8tiG+NXfrhL3l3uH0JSs7WAQbKsc78Oq9JT9Ke2o8u
1QKkvpvVr88kf9EcYzjSrzu7TyeYE9L2xF4PuZzGSV0IdcIdX4ojCmHAxbDSOOuB
yNwc9UmYgkXvfk5Uqex/9j/PwSR5Nt6l0JVpTloXXAD/8qrZNJviLAISSNszywDn
fjNUINlKS9kRtarcZldwR0PLFHKzyCw37XfETBgW7x2OYRhJ5GPuIkSfPGAxTHtR
rbQ41l9ErUJOJQs68io9SxtfXsEnhzpLtVKt/0uo7tPTUwMoQlII85MtRGYg0Geg
Ojroylh36UG7/J1X59kpGdRhcPIo+MYQBeavc7K7u6DUfMS2rbRGi8ywmKUI+usI
/YhP4Jp4hOnF7sd4wtlYmfyEWM0LH5Mt/mLTKmK5LlssPZSnABr7nb/3eKemiaks
l0h1vgzRh3xCplwqI1VvtOXI0Zw+zaqL6FCGSJKsOuraPMAhjO1jkkxbb2E638uF
p5hH2I6jtK9p7nGrB1Ez3+X+smA4YwuqjPqfCm8ekJk/e7YRTSA/qQt/r62KxVRQ
j1Wj7BvPF7ttxTNprkB6unacidCUl6bs1mEo8PpRbXVMiTXt2eRFbiu4+xhdMST3
comJ6iACo+o5YJDqoH9YvH9metZMH0LztV+KOCIbCausCWeWXbhumcSAfNd3nfy8
TLZk6QrAZnS3bzLDhzOAoWiZBOgjdimbXtxivpOyZvDPhLmIn/kAoUG53v/c17fm
THkiiE6Bp46S9FTnselHu+SmZ4JPWrxAD8E7+a3ed5UNsZEqGs+wplcGq0heh4MJ
xRbnUwiWVNtt0HLz0QvCulk4N3DHVDsaYw6j1kapp4xOFOwgsq404euNkfpULI/U
SKgqr7c7zIMD25fXi1VArRq7rUpXCrIVRAN0fE64ZpP0GGKFFmJk1Gs5r7q79zCT
Z24r4mIh56+hu7WFpRZiywS7uVvm7SGdRbg8y6f1vTf47X31q5vC7WHL8VheQLL9
c8yHXBvAuQWnilf5hgHBa3aCinpvVOImou6q5p+OxN/W6j+ItMtaQqNQ9Zp3eqY4
DPKMKn7DPkU+7HT2B+d10dFS8fhHA8KqSv9wQMKresLL4Go0CqcCvx5K4NXSKp4q
Rbu05iYySDktNwM7ffUjfSSSmGm27utb9l9F/X9Xr+9Z35BsYdqEja3k9dCzoPe+
795rq/HUU7ynJPYmO8tQ6TR6wa0RNu+bbvqcsLqmCetS9qVj1onFx47lTOfLtVh+
98DGxkdgGSM50/vE05OA3NGrKWdBiQawVVtQ9miZB/mE0XMO2IKvp6UXfnT+1owU
CrD5DWtJF5/s1VJEImvr6/BlZADKo2tpwB9uAI7VdcjdC4osxVdFtNNIgFQpsqmU
w+/DK8SJHHUESmy7CMEZtNBptymmIL9dbAriwW8JVUvPzxerfT5y0znyaGETqCmg
Wg160jBCRj1KeLoqeGAqXpvYAtzM9DcijjZJNFN8MlGTVLLQarP/24zN5VxQo6uc
Nul5ACKQ8iEhuhBQc8uiw8sIz10oSQ4gRO2vZH4/fAK4EToBAbI+CASP7oxswumA
E0xCCG+byXunGCaS7o0ztwEzuSi/q4Myl2tItnn8iYk+t4HS/RZjbj1dzoqt7yNN
BTX+sebh/37e1lA33eOYALsRucrH3n2TnewYptTP4ENlzMoKvLK8XhVmz4rhQG0u
oRcU2dmoawcXrR9PxNGlfDu3V8AWsN7zVOP8ajIuwpYYuXY4OcKptY1QgxDHyx17
QB6adS7XcFoWoeb18DF0RmiTpno+idLKufSItr72SEX/IG4E24L4F6tKEHvxORAu
f202XxJ1s5rIe89ZafzVde2tYgLGrx/SiP4zZ5oihgf2ai/kSGvvcOgYV+7L0QOC
+k//84XpqKoln7ouQ5oiwFPfzPZ4ZMDbUPnW2ZmU8sRuvx/VBU7iS/DwLPgM7UkN
Kg47SsLZL6nOCIZv41iM+tSHYH0vdDo1DKh+uyqL8OSsi3pRon9+EAjo9m6hlFhp
t0CsBA5fI4zqn4OV1lblYlpZmvsbGaGR+gyOsNm9k8CNeIX+QRDYJTWht+uKBeOA
WYs0e7S0gvR93ig8XrOATjZmeQOSd684cvMPWo59KhJQ+T6nsaCR+0Fw2CqHcRCX
Vha/ERJN9UCzcWtAsxr5Yee1haEDxLecGVcq9Ku/XAzzRXU5ohbgv7qFZtXeEPn3
nra8Hnf+5F9A/jPvTl/IMS81Uz0yeug8YyrcIdx0awzR+kc+2wv5ceajVyS2lvHj
BmigfN3sZ7v7XGgNcbSnzfryv25JzQN6DT+ACMuW+zPqNw1BNdN5DeX30e2gJuh2
1npGX6x0UCKtzKqwnLhT9m+SrEg+f9ZsuNHOG/8/6yd2Ue/pzqZ8kyZ0ri2RLwv8
Gdc015X0TUb2mcWxxTFybHxFIbBmkCMp15pezKCUg45+IEotZPCM+BamD9QFB0m3
Kq8kY+wtLmw9mJgEzaOXVDnITJOGuOex5UL/bvSgnGH2+WQyP5onWTQ7hyp0Hgif
QTRPJZEWs0lLabafFfG6aegmJgRxJowWF1AyzWKinqMFfRZATlFwRDtx1d1mgM0d
KQvqBgqwbWFArgEEe+yx3b7r6YmABJEhS1EpXWWBBoUVCBLn2G+syW+nk8/fA5Ze
8Nimjh4tZlX79Lij3Rg2GnjBc31Ey9hDptdeAEt2DKn65VOBRDES3TQBrW10wq1h
DyQlBEeHTUyIyh+NqBHhuMRQdo2cg1Fgd72P8PFwaA+6r/fy/I5qbDhbbYwHTXoP
8ARAzsem8wmaT5ac+RXSl6JPgU3pYT1uIXHXE6GW4DLwnMdCatxP7J9PZNxtyUsy
HajHPXZRb/7NCfk61mIlKc+Psym7Hve6eTLBepGxdZjKraUryFs5UIUSue7qfXp9
vFMLB7jd7OTaU+d1ElmbPDBrTsKZkRAiFayNAFzQeW/DkfRWd0Oz2Jj+n7WlbzAp
DRSCQKkl1ddSIk42E8v8AJWpuLqQRycqDAcKol8aCr3ziijn9OmSoHf8hm5KLHkX
0s7vya2N/iLrWWDpK9ZciUxs23zl1lj/0zCp8lnYwhaGOwgPN17a8nPymdtKe9XU
LyDt4sY9qajKW8jxQtMnXcoKA757ZYRNwHdfV6EWKNlCqfn3YxcyCdZbvv1Dw8Ay
PAQ04X0uCHwtUVxrBhEMBDfX25ETnmOVWbRzEq7/MsIPP40GSKs5BcfxuCl8A6Na
anUqOQg+gnbvIZXiH+L88V4Eu1CXZf+yba20Gi5n5lywAjLqhLyZqzDO9xjVY4lZ
ynDcCAkjujtdOev2/G4P5yZvRRSMHNDbed3GHj1s+AKiX1Aiqw2ldBM9+6VswkIQ
xbRMea7OLUlHtBI+2BKwfdgqLW3jWmafHvTMF4IlQGpEYh1XhF/nxDeyz0JJFa52
/XeeoE+xWqLvLZFkHKozlF7QbRfrxqe5Rgxv5vo6wGDr7bDh3IZPGZ0/GoQe5PdM
qqLj2qjKiKMzRG+L9zCIBgiANHpQfGplHLpA/ajvFKF8uuR71AB/0jyjqjUzWagk
Tb6QEIY4v4dDUCqg2bJhzIc1mXfVF4aiZjPEaPZDgwJLM5QZ0W9V4/sVbs8evVR1
UH6+6J2iKeJTYz3MSoegjYjuXQV3cRYaAjmRbcxI6ZvbfTYr8fX3Anj/omPtI64V
cnAtcLKodsOFNb3igUrRjcjqdFqltom/dRzi2yPiMQfS/LKPcgPy2ZzuSRG5Xjcu
KzNw+e05q6LwoNGhWehwiVNwa8YhEMkvoLTDkAkXlZKCgs7fKYLhmWhNzQhAW8u6
LineZKKFTyR9sM3bNwheVdP4fRkbtZv+SRqWmCTRjBtvEpOplYBYTeNUtADOlHO9
v8zbjDpXSXYidr01yfaFHlg5iSKBbP3+7z1JCoWpPctDfc1FuaTR1dkPT6CjXWhC
PFE7na5UKYqHJ0+b8MPl8QRF+7qdMbnRgoNOY5D/G3Z96elx0x/rm6w8ENtekjKp
8XyXKkoMT3baKsNXLNGcziJ1a8teIesqtYxhkWiUJUwACirxtZ55eVv2XwX+5Qco
M3Xvy5mz/AspmVZU90Wx86oPUxBp04PUeI7nMbh8LuhmktbNeKmzJ6Luo+XWwXz5
j30n157Op1nlSwI3OafM0zHgYtj03Tp6lK9HrwHd6sCVcG/Ywa+U1ey/Tm9NGteZ
SHRZd0utlCVyPOl98cbxn96IZFcC37jWfd3/ypBsXCYMJH7Dx8YKo4tb+sklKjwJ
ECqWPlwl3zxtqgel1B8IuwcLUNsa8Jmt3ZctPsXR+PnpHMk3ZQpIGTPERnj5aTUY
OZIt3PyWZzgoL4k1c8WucyBpTO6SckM6AFdxfN+dGqqclvTjJ2A2g2rWQQyTwAEm
tg1zxUReno7uRmT86gyJLuiJMTyYl9Jeqih0pBgA8evLv6vRFIhNKA0vXjW5Q73o
umaMQE1PTydRe9iyk+GLnZ1Am/UsSfcLBik+vJldFUAyX+b7LHASdR0vVWVSuqBC
+lD6/DsNkuZVaqQjIpOkQPJFa4JKMt2TWvxi93tqyxN4NYzExaG6Qfg0WKr5A5jA
Uzu9PW6Ju0VnIXEeT3pvIE+JZtTEbUpxvtuQfyfmZyWyG+P1zjgyPkalA0CSDftv
BqaPNkm3Hy/Yrd6Fif4uf7zwLQmjaPYaa8Tz7kMR+q845xUI2Nz26Oi0enQ+cm9+
kCNBKnb6diqhSDHEsHRZT2vBq3Xg+ixzNtxjv3dvZwH4gURdrMQJsyUzmpmoVzyY
cjO1GnWrwG7sirNwicjq9awnOJjYYA9a4zcO0SEMTF7L3r77eBc2l45fke5q3aqK
QbUJEAUsNZkJVPpOZOyWxlltf43q2enNPsgClG7KEwsCBx8g7AzqDeA1gRAYO/OV
eFF08BlNu8+TLRp3W6B230ZvlSix4fxXiHfi9ThFbxAnSWDvG6EvEAJ/Hzo0GXKH
0ZmmQaqYehM08bvAL1dAbz/wj6VMk3RVNKFuprg2uW5XbqdVJi/+WaUJAgKauBTI
1pgZUslIP1AVWUSl0JVJBfRBvSeyim2lcytXkDUVxCjvjtWSybPW1FROOgIe3GXE
9/0I7swc8/KK9S3vEcxWcgRdUbIji6YAZivu/Ir6DQnBtoDO1Nk6iS54xUCCrFhK
nMatjBt2yAnhMnroIN5kP/bIWnKsX8Km7eOKPjRvjhTcBD4SEZLV03d5mWA/o8eJ
6E36dk/YyP4d0DMOaasUtm9umpRg585axbyiuj8/JAxieNUcBFKk4GAPK+nyDsaO
V0rgtRAQ+KGg9fS4EkRG+gf6X3E9DdFSIP9UPtvc1kG8xt4BJUiqwuyR/exNzSbt
rC+KLR7luDdx5ssqG34UkIoG6cTe97NWotjlaILEzBsPPBpNhzfbljJce2JIYJav
/1hs2Fxqf3wmxA+MvixcmZn5O5gbyowlAQdpzLys5WGOJte7hca6h9kwTs/gaNL9
kg3SqheHXbdRNzyIvtks4+LApeVT/IdrhOq6kkF0ZMgZmDlIAMtjHF0AMAF0GOkw
WrvrqTp0Qu9RxOsJ8mHS7OSBd78hGU5obW5/eT5BKSpmU4l7raBy4whNkhraYxfP
aIn8B/S5OOPGceSs6P/98KV6Z4Vh5JvIk9o0i+XSHKo1BlcKVkXAn80TP5Pq5B6G
PNobOxx5A5PEQpD8gAlsZSYJ2b0eu/9+iOX3MaG5z0riCrJS1UEVI0OjZOEVukdV
7evaDpemW9NUNz4RJxOIAk0QuSmcLq2Zi5tFcmMpu9H8uIhKKCT2MC2X34Bictza
q0hF3sdTFCQp2NSCZyTH+DeQuDjJ71io62jk9pgl66/FEz5p2M3023407hmrSbmZ
xwAlL6D+wakw658p7TMlEXnQzar7kAWcO3iisJfMbbYR5rso7X6QOpgJvvt0r7Mp
AVZE4xQjOzQuJoStnFD3GIUTO5kOzWX4QR/ngfaCsMizFr2JuIXC/mlRpQ2TIByj
wLIE+FIeaDYoXZ2q48YhXQoLNp8VqFJC/2gn8Rbkg05CAk0nH/wXlVlMJCVqGQBr
mayStl+SRwpbgtMyxIisnqppVNs66MA1dfCzfuURjqQSs/K6RrbCQJQ/Um91emAN
Ck8ZyccGOY4rsz6COHCmet8fJcc/LXf7abIAImB5N+56P1dFn6Jv4OsmVCrzTjej
Wihm51/Dm4YLeb6GsURQEaDU7XnE1nM2UjmSWhREknu2e7K4TpYXiqZ48QPUhVju
67mpVTScHCMaEWdrIyrNaCWRun6LoqUaSCZWBd36Q7gT/zDLoIjnQa5JZ8QzMpv4
gJZcT6JM6SmBABbCN5ySMSAtDkop7k9NkpeNtCapk/LrO2v8fw561mq85+bt2H6i
BrrWGRXFFcKFcxcEzeZbt4Ljz7aMEZybuhW7gT3HufJJP0GE44TItvwb2F4hUP1N
HDDcfnR00Z5vPwCQ0JMNFq93lPLmvsevKPcQOLxDu+WjkT/hfn5KjuNc4FB72WnK
errx89xhNoUMj9Yj5pFUKr/4VDkemXn95vr8RAQhoG3L3F0EaFiTh7y+dxYyrdI0
pZMzwH3VkUeX41kmP6J7LkwsWIgSeThrglTinRSU3aQJlo4nGUIT9cRMO1hM/tcw
/q2lSezZIv3z5aNl0ctWUk7R8wBHShU8BnDpJ2/9ptXzB8f9dRQ0y2z36bc5AhOP
rSipUmW5OhiZSp1Zj9+NGN2yO8zZ2TmkIFCLstzzcQUcINanCWXUfp83TktRadi7
sxk8wEVRkLtomYHkq5R95zynSsp2vGW1lDfZIKtG3UsQgerzCShBm1b4WABMwDM4
DqWFrIJMt57ZB+h+r7jLEwRQgWco/QU4gcI39g59mtWXeQOwowvcXSzvWz8pIy7y
1N1d6J8Cf2ryQaiP9egrzD7lPo60UYLisPxKtseWZTG6S34QGNazHpPqOSUoEG5v
JQe9aa8ONOdzHM+t3reu6V/FHfIg6nMXVk2/d8Tmg8CUP/LaHLiRZQRos6nokl/n
CZlsZAe0U0+sZHpcTtZ1/dTy/YEk5DrgEUEvjDWUVBky/4abb2fh8qvuwVrXHG4/
pBek8TAdzANVHPx3SagNlxFLVQrssByTjvl61mQBZ4XQ8jR76Lcwe6U7soMkTwj4
6tu8M0s3Db/EMXYiJKdpLOTk6BtwEBoGEMOBA4ZAVNindHiKkWTnn0sFRjZgWVof
VdO3/C1B2HJHXUQOsJ01X5VREvMqcD3iCrfB704hOYzGT986/NTIIRxJHjq0PNtj
Ldc3fValssQW8aG36/wsK9iBIAGts1Rrsw7L59v6+DzRWI6Qu52nTMhKdTrflxqn
0mO1dP5h8O9n6ypvXysK8nHZXQWOfBxYgaw6u2bpJlm+pAGAX67FJy+LATtOq24L
TEQz/IrkOmazZDfGRThjytdjTNT41Ab4Ky4GOVqOeRmP6gjJ3v4KCKadTE/9t+fN
+kkiX1tXA83lVQfTGBWYQ0Iv8PhAFE0O+fC51/dJhgWY47gZ7iYEWX8/mMkBFzL7
Ut2ZVnaptE0BmhJij2XBTKKEUqDO4eMLPn+qMcqK9g/7SmhzI4QX7sT9SD39S3LA
BOm2+AxoEjQUdnPQl7G7jw58VlVywOemoYTHxPg8pH/c4vrFndZlI0qOSsKCSY2U
0SCoXPHucDpNXD5TJBoVRgIbLnfPzKkeqex07qa+MBSjQDH8E8psVVCpzxzweY+S
K+Uefo4qtgxAvx6gtTc6rm3cPtezVBVTcEpyRk+W6Rd3/PuRmgLMlf+x9oVgNl7k
eXVL/g+zwHtG2PRyVWTxCkUMudBwcD7T4HXoFKxM+Set6ZR+CfEhlTMEg36y/1nF
S0TQgssBF+SIOhj7w+LR7YyhvArTCuL1SE5/GNBLw3EDRUr/RqnlsmmfrNZ/QPcg
0O5atm1d1a0CCj2UoNMvLDohmkRJzf92OWLcJ2cl/8vYMSuRbS9nxv79oVrZuNgL
7GVVoZj3GlGVxbYMNiJXYxr1V1hi664oqaeA+rtzQiYWWxNVKdvkkBdEVJ1qIeEw
OHOSthBKiBlC0py3UOBn8aR98ZKD5GAX6zHhpvS4uLO05z7r3Zx+ysOshHGoFMD4
1TrigDdEpVZ1PaOtN2UgzNB3jvwry40q7LEbq/rhxfBQcxyv5iQh1SPm0koymZvW
1XfLn0/d6fawCj+YegTTlhVxrjbLCJG4pWoUXcsAvhm+B2jLVEcZOsH/E6KYKv2C
9yMxVE9bsjOzeNJA5i70N4j34t2Ia/bdXF9l6pgMrjE/tNXrz9iLDi3nsxNE6t0I
+rVE9RGVhaZ/EXGkHI939sgKeDhyuAMGrt4qFiNUspeG59K25pEbdjFem0Bs5B38
E3sQtbQuprMJho5lGTfKo4VbfrYQ6od5uwvoGq2VlomvV1ZnrGHT1WNLfEDHs82J
4Emz+cjjzAKkMdeC8VopwuyCPtdaSEVcaypDpY7W6MPjcZhuOvxPuqbHGWkfk6a/
dtUvw7f242iUWpIdY+sSku/F6QU7US9laxnU5sq09HZAL7NEb9y6pQMzrXy1vewx
DxjQux0XonQN9oygAlQVhx+C8vjXuboLMN9kmPMgcL35L45Ij6iUHrXgv1uhG4B7
QSNaA+N4rRYTfdA2+CSL8Dcv9vjzLs/wn0+cvB6sb4oKeQvjLF20UOFKFFbcw8tj
R9nbXDnvXMSX2a5ShXe+CiFTr2ItIB6G15Wn2r+zYAPh8ALbp+90D0imvQZoywL/
w4AyMdwf5NHkNioWPYXlHhyYRNkY39mVVEUDrEbSDlajoo+GjRn5z7g0eGbCnm35
5KGwp/78Qa8TAPDCrZl9owU++phlIxg4AylgDFdSsQSmDWqrqmM4cSYcpCtekUPs
RHKenjDW7SbiQmNjVDVxhVY3oEEzmk4qx4sIo09KR5ngicRt6alHgHd0KFTMi3vi
eP5TmcN+k1KrzjsgTBgFiBm2HueXLBLih0nhf2uOF9A0BWtsqOzzcBVX27Kesi4U
0fojBdmpBYL3zyqXIUYbErfbsS/MM29uD8en5jcsU1aamQZQVRAK7FgiJdk6CRDi
VsUUvqErjU0gRmq3bX2BLElNkKNsBaMpxI/SlQif0BaqQi51R0/D1LgzON+Z7rtX
HLGQA95dMdcOHq/aqekN4htEz6a0cRCta/qrQSRHhdxNeDIIPdFqD4ChDTlrxX89
lvflcdExpTjOKwtEUACUGwI2tDgVYRqNjKVt4Kgs4dV03Oj7Hph7YmajDSnF0Tbr
+u3C6l8pHDcX4PGOZcTOfmKSDe+eEq8svj6HLCjKA27KzMOnOaOt5/xVb4qQj2+U
KhWWdWXGue/CzHeWgKVVnItxdF4ch8Ln5pjGo2iJnnVA4NfT8gN4I8jOBygUq4hC
GvmCtlls5DvVgSF/frw9jJuaQD87Y1ZezK6iqmz65v1LVsynAt8XxIwoXnN8YEXe
SJEsCSyGo3F7xpMFTMBryKyHhS3VD6AMuOUVTmyQyhjGc/e7XzswAE3Zdcr30dxO
CuGgctMk3Nepw9D5pzADzBbAFeYkmRntljYJB9FoIwpd6yRCRJv4zc2jR566a/oc
TMTEKCLMq8zZHWtJZfjb3XQrTSHdv7sdkC37Uzi2Sg1cgXZrQQEIhdbLEoZQ0U7Q
cV9mEY2++245xE9Ke67Rx0b2BVvyOL4ZwmuCXSpsz+YkSApUNClj6BAx1NK91k27
QmdYPVyT+nJ+hN7rKLAFF0SZHOLsKAoafwE9LeO0uo9808vrLMPZuTWX0msDxLF3
AJSR1o9RVO8ACggK7FWoG/d+y/iKdwso8twUEo7CoIkjlprzUKvKMSQ1FyQ/E5jx
6LIbDSODiBNYjkW271kjrcKCLIY38nCu4EuK+Qkl7Qkt3gp4BqD2KQARoSMbspgS
0/jm+6loJy5pJASjBVuJevtF5JfKZZmQNjzoFMsRrj10vyD/p6Hxe/OcrzwiPIe2
pbSdtw84OnglRRYwK0f0KRnw0OG8UMrCAxxqhnx2ZyEbv9mkE8CEvLNNrZeoRhRO
V0xzTGIGdufftRX9xtZeIuXH9sa5w5I1H2dtVVib8dfitvNOzvtYGaw7/4OAjoUV
NpzmkTF/de+n414vbYiRNkmJAwyZ1OJQkl2G530u+uDr2kRlkF1wHwsDdT8F5XNq
6J1SieHAjuSyVNE0R7GXjZFYzimZNiOjPh9m+g+dv6FEg97B136cOEdZejVNMWLP
hOks85t7soilWJM5q7qICBMqfPybHTDnXBy59XhX7xQboGtRB+qt9TvPUWJVnsah
RkgWL57SP28npaaSaAJdGtjIbJO44kOvwCF5u0WOLYsonlxHpTZEU83qrSL2CMBx
iXJQ4/DYmTPv9UIY+bAhEe67/9gFeQF/7yIUcAwwzXKlw56b4VTdxMLqgD4QZU6I
kapOavLD40ZKNu/me0nNqga2iT2lTFU64JTxMcfrUraGeXjTAR4bsMQkkE1EEXGb
tfiH7FO5Vec4Eebyi0MtxFVR4y+1OGOu1VL5/gdqx9obmxAJe0gHsLmOJAXWRwbQ
4hm7Ihq5Ul2SZnwLcq5a89Zan6k2qPVONnzUEz6RRx1iEzb4iswv3D5oaTc/XT46
1qUN0xiZ0Ekz1jLPuAs1MjPavQN0u/EKUHS18yX77urf2NsNltwyfay7rNW+caRf
v4E2QKRw8WFP2LAUmKTcTAcAldEGFuB0BswRI6LyFXyVF4jy9nUtXZIZbXgkCdp1
EcPWjZMEEIdYhl0m+6pvL1ulFDk1DaGDjXNm4eaLzD0KrLfXTpM3sZyLg5FEHwb5
lim6CiFQKN2eL3L+BQWu3qU7cbMDHrpWVYYR+dZe6I48PHj8Og+LS7VUG3V5Hmn4
0kzghmuaEbHMG67o/k1aNcf84sDZrgmH3R8FaTe9m1N3xvK3IGxtt5JqcS9WxgO4
OGeK3EKFr7CbpWsaph43fFDRQ08wcjsRBGIg++hv1LSNCl0DNsJ0Up7zgXRGYM9L
nUYScCXU1sUhI3m87EcjlIlhYXUrsJAYHDvWkbc0mDMoangQnO9QKRM/Cr8wZFVI
d/aX0GsXKNB3K9qOQtHTqrw+KDkrRv5YyL/lJEq0swzZALLERAJmO3FlHWBzk9A/
h7f7TB3DiJ9O8izBI2Hn3UXkQ5MN5kh/iu9o/38IrddYFp+HPU14pdi5ByKyGG+R
biutAwU6xI4W/yzRzqx44Wj9jjSou4NfneBGaDUaKP+Pi+cmK8BEuYgYZEC979lh
+dbQrnOW65Ix6/sg6PFZq0YrfxgJdGTaPZCvc57jmztCYZBmAZuW6m4OQvk9BFdN
pen7hGGUAv5Rhvmoi7AcJ9UJoWVrEqBn6XyrT1tO3MQ/xg3TfinQJ66fCje6vPAq
sl4BmtlANinbkw4hKmWhCf2kV5TFymY1cNwVqNLlADzeB+oPbuo48rH56pWRvCdY
E3x4I5fYK3ckUnMmmO41V4tQGEF6utoGW98IzuD1GMrwMYmOofyxd6awzDQuFq5L
GOEjVhbnJ+pIvKhQxORM+scGphALpnIGoj94nSieNek9vq1iZG1X3m+evM5XZbzt
JN07bOxjEKyHPS9PNikzMo+E2tIvS3SeeXw9tAPIZ4nl7TTuchAz3jttSXlBYGSn
S0/+JUrsQs9iuJr9l59OgETAtxesoLaTSbUzx47HVY076xdkzSro/nxD2769Q/eZ
yRf0RdgKoSNKv01bo1LXoiYCripmv331GKzz/OUJ3beztQO/s3yx8rcpQ00U3zgQ
msNlKExElmv2Su3rdOY/8m0WB8OvhpThsSVlTebPY7O17wCOx/CzL06iTt4J+COv
Hvf3p+l4mOX82TRTBpJLik8JYmcOjVLFK2krpOrQsJx9jO9VuMrzQuR04hnuOZw1
iyszSg2Z9M0LAxHVvpoklTxZYzUyT90Vu2FDGzjUpNCFrXzQm9lNKjVeYbsIXC4k
0YS52BdpN1zfPGwh/dxo7U2UJqtdAj1GJwg8B+xG9TCiM5W4SHRTSWPqGm6psR+G
pxXz3SZIGkCuodpqGPjLC+tdE9VRA1JCVLv32on3nVDNdZ2NkBFjo/N/Fo5/ijc/
yclnpoFzBn2lZhywpgxQaK/AKMzfSjrU2hLOrnMIcHJ4+gNeGRbN/KhgRj7mE0lH
npU4gyHu8hEWvV70CuXLSH9FIe2T4sbDVv6D09beTtF8VLqoaHjNhhQuuBiSaG2S
+QOOaK93NzpJzd9O2H1SBS0qs9CTi5s4n36x2AcNhT2FUh4A7rlC5HNXhfYYIMaj
jrTkt6OQFfu/p1d8UuDYY9Zv5EacI6b0pHE3nqOIROyyp+VPLTtXVmZKX9lUXpNk
1czLFCpti4YjKBICUmnyOrXDG1q4T5XdGeVzYGQoJ7924fSfIrOdPf/qGyWuymtQ
aIGXvJ5DDjIek6S4/4JhEzO9r1mnhZRUVW9RoYdXLXPELMCStOMZJAxesdHhI+00
fj72PtOcjsye0I5c00HIqdDeQPh7xAchMlLN/u05RMZXShBVFN3Mvgy+59BzciB0
O54GQuHo0VbQBBFqQkPzDuEStZemTJ9ROzAYub0ypJ3BWIK3QcZUYe/YE3qSoN5I
4YKB5CmImXWw5wLsrboNIYF04vqH7EkgPfklLUZrOc28D9wIKX7CnteEh19xeZvH
uqY50TjhRcMLNp334ZnWbkIlpuW6/fRZrjnOBzm8HmQg+JJjxI0FaNjQ6kWD7u/y
xrlZgFa22L21O6x0uGqUfq7lFdx9E2Z/MAV3IXq9ZEDwyR37Qcc3czBEZy9ZffQf
4j0U4Yd3nGeCQ+ZxZ3iWd9nWHoEeVWwU7qPkxdvDVMd8TvVFvW/+Z5PME4gQ1RGk
x4kR2BORX+iVqtNTG08RLPE6IQlVK0wFuG5AQak33YtcUSbyxfzjKnW+Xv2/zZ/w
h/hTJ547CMNjrEW5INYqHGZ/P+KSP0MYR0QgbnQ46KFC9jGaQK/yLgovuTQWZX/R
gbvQt7AU4Hk6D+yzeWLvq0Q+ZzmZgmKvqCR+ELGnVbcEMINZG6TOz4WftShJD7d1
Qzym9qCqD4t5KMXZMQ3hNqqAKcx3zONkezOEdI9mKxon1FUwNInX+HXvNKLFwlro
6hLQT2xdn3NwJU6LWd0HWpE93QKxb69agXyHmwmv0l9Rf6seQGJY1TgfPf/7kfsY
Bo7oqCZGl+TJ36oxRw1LGr2X5kzkIPYQHLw/0POC6KfWCD/Md+TgwQvWg269jNrc
1Jfgenl//LqWj85SDpJBYqzPwQ6da1h5Teb3Ibf5ffmMcBjWXY5kMbQWBdM3WV1w
0rQGptjgUcQ3agCF1OnhbM6/rAr79f8mnuzRan0gqvGT/pKkmWTXFlqWhR52WIi+
SFq19BYU3xrYTqDViejquQ==
--pragma protect end_data_block
--pragma protect digest_block
zt+5ogxiXiHmKTslf7ek2AWY7jw=
--pragma protect end_digest_block
--pragma protect end_protected
