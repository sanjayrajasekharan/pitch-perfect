-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TG7a1KcNv4UXC7o6qojxswCQ0PNrfWo5a2OhrzHDUvTaLl31IiIH+A1rP6Z0LWoF2j8VXXBE6rvM
mQwiZ0eSGz8wiuevJwuszguuVGpfpsSrmhFob01Itb0AaixVMAx285IhlKwfRWPFUNzYajz9A0KX
RkBQR53TsmGxak03Ncyd+TwXuzxL2cVNsL3mkXBQY+s0SwHve6Eejt/WLMocp56QPkiv/Qglt8hx
/kqWyzJ6pHKv+XzZzqj9NLY0n1vJPBlmmqeAEGQ9RfF9aBmKCVTTivusCzVGX7rzEoDQgO4Rg49A
uwIPkRUwsGTl8Qx1p/ajZadGDy43Hti2hE/h+Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28016)
`protect data_block
rvrs+mmXNGGW+PjHpskRbdiD6Q8N/pFwCQD612RYnxCqaFW5p0eWwEGcE81WLrHiWD+HLttaRYos
rbEYGNt4C5aF9XZHTcaXncMC8Qd9cDk48ojw0mrJPAE5yVOYbpvd/ATFGibIz9kwg5ZNVo/iRYgB
TDZYSlTReZj5IWv6uF7vph9Ut/j0u/36TzHTkEF2yzFRdek3Biq5/mNabrwZu9+tiYXby3FI9Ylp
XG5ig5q3LMCj6JYHueQ23AHXS9zW8sYhMQKfUvURRdhhlFiMPR6Wi6T8oJqRJYgX3h5JxP/74IkH
vlO9VylfolxM5va/yyreHaca/F7g8q6SSX/e51FvTjFi8WoBPNxOJGjppVgprvISygDB8mdzddOp
1sK3ILrIvcUfLwEOqDfVPm/HZwQusnNJLnJPYI5dZq6HnjU0ldvVHyHQXmzdjvLqpmdkRQMbc8bT
GhqkmJiT2LKltGOnbK1OqJ+sRwbgXHhQ6QUxeFyTvkIIiJdCSjtk8GPqdl2+EYTVASWCz+7r7DDa
XjiUtIsG+ZkEgNeryjUW6kjmtQh5Me47Xdne4vqZ9MvWeQnmFv3eZVe0Q3EZIgPU7wp6e7iXnYxf
k/WCziN+FzzuseamAKRBh1dub95Ay2eG6lKzunbTB4r6sdyrB7YXLFprj7p+VSICyIw39aiPoCDv
uVXLOW+jhpjh5SCZtbYblYk5gMtq/Ak6nGIHGK1f8fVKwCTqdHcZssFj/ls2qtEoyQo1r0vyF6j/
kq31I32gt12eHZH2TLh0DvKdM8oRTCGh4hKpvYJDmolMVPbLIgo4+7BuKQffGszhvSzyjhx72Lgq
j73T9wWRJVJRUsIougrXjGFaM24SYwIi6m9nC8IK8Ud4aG/vL5rdC8Hvl9IzsCrFZfmkhujRUvrv
8rF0LCYCOGlOWdOF9YbywZM/or7Sw9Y35Rgj1vZOJuRm01DKZ4LKMlDqMe7usY3rKXlaploWEyDe
wpiKM/kf0XuI7fdWCJRB7bDx/XH1/rgmkjxnr5CpN4rCynfHPn2FMW7TfjfGWaORv+TJmpk5s5Ub
/dpTkcRVAMepbxdbU24gzbjhmqtRR29G5pi74BGPv8aC41V2wlu4wtFKSbTv8DdaMzdi0UWqmY3M
NTshxxEk0Rsyq2bIOXqHd6FJpQsNFx7rqRq+tspx8UZalxpj3befMe2XxQhty2fhTfLr7bRwCS67
xKSJlCEs+bDmFEGqmwZ7d6m/FVCPJ7A+CCKA90U57c0LBeKQrz2RJKvSXX+kWuiO5W7M8cpd8tc1
/m+ztwVYLKxE85DL5Y3T+2gYzmouHwZxjLPY793eXODvyM4Y1y/EKWyJGXCc34wCueTi38VsbuLe
99C9g90YsqFIOMnAvcIL3mTlSlCa2CaUD8MvIb+qw5W1EjNYYKPPj5iE57hOoKmNfV6QVsfkj/o1
JZiHYY1Nr0RZ2EHlx+2lZ5c/HwsIHKvPGK/3G2U2T3PYxL70FG0E3kchXWB+YCewVhZpq0/w0OE1
cwu5UdnNkhqlUx/q6NDh+I/aMp3xSHHQShqUffSGLAmqbBNlij0vTkXuho6OcEtTsq6DZGmI/5D3
7lOih1e3ZSdgifSMKH3d+CdmV3w9C14zge9BI4sb3iu9hElWnpP5byNcvq/DZWTloDABYTH2VVoS
NU3br5uVxJlXENKobbeSC5ZzT9BoluPI7nYOsMRuQVeNoBcrYMwyaHpd4CAYYGrkNEUBISiZ1p5t
5d0UkHxt/s4Jzqpfqufeu+JZnrPG8DSAkfuMTse0+JcJTM/CB790bcZ2mqg7mHZgATRz1WGQF4p+
3Q5ODCrhQke4tt858OrnbVI+7xdSTST+DYkpMF1zlgnGBqlEQ26tGMy1ISLo7sjDvN4Ueq+bPDhE
AotHtU+XY60cuvZsiHMm8oiC3yxy6PzYKW7MF1SaOhzosloKSictJQEOYzUqfAjKpXM9S0vNrSWe
16bPrtVqAICKxLprTz/C/OrQaOd93Godmv6pQSbVmOcjVC+XklP1cQ4l2SEDbqDEebCzFt80KbDm
qsZXl1N/Y6toBQ/xonCABQbVnj/SBNmeoDt6OVFVKAl3xdqJaSYg14X3AJFf6NZ4CLLgHSidzgb0
N3b/MFPGm+mCuWDfYVELzzp7t4RkJgK+TqkAPuX4qAEO5lJHGZ+pC54r7GWWuL1uvI5vWsC4q/vN
FXqMAY9fzg9NWqak3QwjekQu+l2cIXicD/yGLbiyDiwAN7wArRPEb75zH2xgqaXZ0n/UlyFRPSS0
uAn0QceC9hiPWJ035vljJeX5O2HqkZ3RXNnka+bjsYaiHALbdoaSKi6n5GaU8cy4FTPJhguR8maM
FwPkx0lr/PI8mrX1dqW9Ll8Iu6Evlrtz1/4/ite0dZtlDyY2pndipgSWWzK9GaKHxenyv0aEGVBi
1x29W0/NpNGLHPOBaXEzyZ37zIQl98LlRYpbJ6jE3g6fvwgMCoxJL3gav0KmC3Rz4z2rl+5AlKkT
cagjladUtLlcpMS/zDgg0lop1f1VAytb1vZ4SnPKhvl05DAyzmC4jad8xTzziWsUhpzeJT2/tugg
VYvpZmWTFXBhZiqQW98TS1IeS7wCat3V8yKJJTBWMQEIHkjVOqz5clPf67+EzYmVYaIlGjI6D2NR
8vt7V8a8rT/z84Yt8cGnxLFrGjYhFLqPWeNuwCad9CqoTkFvWCl39hxI178xF4LwK/NiKyxzG71I
4LI/LQ3+6Xm2O394zHN5BcZ0BxEzUfvA3xh2X6zIwPTJWrjXbVWPuNOktV2A3zMv9D5+mTCMLTRQ
WooqrEdCHfWrDYSuD6r3k2to95xHA3jsozKK7QJS3AtJPLUqmTN1Rdh+4qKNYQPs3e15SCCHc0bY
ZjYFrYTTzrnVyhOTuhSWpCFcIRMEDobyxaBL2shJjVZkT/nS6Ktevi7ZhrZ2sAFaTMBj+YFAWi47
6K1UkMNcZgPHqQP7wQFpYjYgzdKio7oxElpiDGIx60HNkb19bXnJmgF3h1wooTmVp9Vc8bmK7v4Y
k9WDz0i/+ZMPSpjo3zkEfwpaNgMn5Z2CRQ/ViP4vUxtbEPTFbKyiF/RdQqArhaO6ksJvabgJwdv9
WFybRkQVtVOmbpd/N2nWifFZesxLgmu/80Hmh+p/Sec1GoPsBiBtixP/dGstpgaZe479nfqMvOGx
iszzM3SoRsBtOLtaTvjAE8AvXU9ae1UfyZ1wgHAkWugcAtyPDv2veCkEvtkRpnXInFDFjx4d8oCy
l3FK3qGAUP/q3cvvyvoa7IukyA1OKPTIaVphZUamSd6Am3hK+BaTRhNOuxtp3DVZfSImaLbkyVB5
YSqQX3ESGFs0zSg9X2AQLONMeWTAXVPCzo7k8KAzmVcNi4JoeYzZtzWjCGAOmCVxYUKwFVNsyPHJ
Xcl/zsZQZtoPYV5kyQXMtF6pMxriRrtStjkXb2ft+OIpGSwvAHSah+/EqpxcPSsfKFGc0Dwwt28n
cVdvoGIu7XmVNPhvFJbgh27XAVh/t8n6XqnbgiaFNS+z8FeQi9zlsFb4nAyO7cD9ze1qIFadb/A6
311DTn6cADW1DPECWvI8Sp46uCPaReJoQy816JTCOKRZqwUcmHo6HDgu/LLK4wEVPPoN5Ohe0PKJ
U/aqTuyPQmI5oldnF6/oAW6Ea+8BaJ8czJHj3j6YA+rZTTKP8fqCBvKfJAHHygrDkN2lajGlRf6l
qvM7wVPmoulZeU7TUPK4aIBjpwICUbgaqqwBFLf/83jCiUPlQ2Gf1Cg32Fnr97cZzIbHQW2wITU6
nIyvKLP/kirnXgUsFXNjk4DIkCYOCebfz8IupxRznSUGrGq8LZ93TumL9hA4Fckr64V7id0DZtci
URbzaSC9D3IsG2+WERIFk12nf2+0YP3L+PCFHuctQfLi6AvkAhE6E+RbefJrzqpAMoxAU1xSLqy3
tEjbgyVvMA+Er4lQb/clo9S1mBW+g7zSJrKFIxTOSrt7/7z8YOulYVSg2J8/m1/RV1YI1Hn/xUhR
uloo7UqNoctjxiRoSfUQqwsnQmRRN02mcM76/443rzAGeyXITXBjjTcUUBpF2jLacvB4wx4r5vvI
sosTJ5k7nUDTVa4+SeRmJwUcu4C4nkEozTji0J4CGRCH+SUI3u+zncS875VtdogLaa+Xgzl7dFoZ
dNodS+goE9aMzo/sx1pHQPdVd5HvJlIt80riekYuqBdO0TSG/bBhdZakRIdsHPuwQMvkbnD4U6wD
a8QH+llivCyzNKJ1A0UuANJbXSIq13MtcP1JAtZ63zT7O+kYorswEGvk8A1vvM/ItLNbdejwQamz
ikyh+6pOyRVRga19uWjYB7UVNUCy8xpuEgXF0CpqHsXz7sev0MOFvHgF8hGyakq4MYhqIzRQ/tCs
mCSpvi2nusVxF1Fe7nURWdTujMnCCo1gLHySzVBVchZRQcOxAzCciQafiwQIzl1zE/3lETrPsz4K
3heEQi5NheHeSbMbYw+J4AwS2bDb1jNsl43hpuPd45u8+qoMgHeTGiG8o42tyBcNEsdlcTCnrjs7
7FTeyApQDrDIkhnKO9ZQ7bmuwHS60LYo/mZuG1c+SXrULkvRhVxVIVmoa0E7cZ11Geo6HZYiwss/
mUgREZaE4zYh4mE+26N74ybNw6QvJalgd48lKxC4ET3xv1u7XOf5AJVwqnOW76m15ntFiYQT5BoD
toB7hyP7Jz7ai94Jd+lvVnpd63E5VgrWJ0ObhH/A0ZDETW3XFbqaAK50Xc5TlAebB+rpQh94wvEB
TlpvkZnNoeS0+4/X+KCrDXyIruZ8UB3XV46r7tXKGL4AvSiqCRm8aBWany7gMYnfvICx4PDAsK1n
at5woymrq2HUvrI07tIJKJL8cs9WujxvLe/dLCnUXkuU058H9bYL6V3GRw5IG2FZPM1K179xJaQ1
BWn/MVl0Q8QuccvKfTaMkyokE7pTfTO2TqsrVI//lm0nx8WW4CzS30YxbQvR+6UeOD8+kbnqlqBc
41YmMXKFHsI/AAX3UtanJEo0JAMnKbHSbSYkeVlRr+ie/8bOB+wOXFmflJJ9HvbcshCF7vgEI80d
CGt1bLq8bt+7O51Uk0ImZTJ847ffqtBNn8DC5xuL0b0T+QHPxxpBFUqnN/lol73+8wE8FTGxDeRA
UuDiqOjzAgCfZ0W2E4TlqFDJMLItZcchb4dZbHRdwWYoli9qGwXMrpCjPtWt8hy42jBvVjkNTPeI
nQwH7S00upDgDYXZBOTMNvXL9ZFVYa3jaFSqM/kq0jdkMB1aAN6M5sZlEacZnPAXSfrvoFCgaZHC
e2lssSf/3h7S51sDD7CftzSE0wu4brKzErjP9Ukzc9dLTbl2ZepHgAnOOJRXmMr21OnmyhCr/7yB
+3BOy23WAOrlNMDoP3NebJXWqroer5KuiJ/WPBcjF5DVwPdCXnL/Xh/glU4c81721t3vM5hDXbLs
roeCLRFtAMSiFKGQb2JN5i2HF987FLW5IXvGZ9INNRflfOpZxyfbrBWZhpOwQKniqXgh40TwObdi
DHHE2pW5KrVghK5s5THgod34i5o7WkXDo1bpP39CP0z3MsHyYlTneJLRZWMTiIQhpfPVeetwgtcA
fRU2EBpRpk9OH5OAYXCEvJA/4VOqqb3yvW1R2dI9G4ONf4XjiwFKdTnYdjHmQ3COr0zbBhuFIrHy
sjDUTADXm2hSdAYeUjM+xMfp6WWzto4jPtUCjS7WrgLTbWWlxlA2pACaUlTinS4s/R8P3dVsS5m+
47PkUJp8GnsBFZUga6wiqfNE4x3NC/7iOOMGc32gjLz47zx5lkUY/loAi2wKwkslg6hA7Ieu1lDE
2oppR/JUfXwqyFuqCatOZscnKCyZRBeW1p+OmDn44tszYlaAPBi/hSc7qT8ggINz4at3kOIxQwsp
nNdl45nwZckKy1UtCZNU6pwqSNhIdeBatgUxCoHSDqc8gZ7E5dv+pfT2GmiJDXiSnCFs/o1dLqBB
/8ZtLwNy42UeWni1dXE1Z16sx64FIYbd4am57Y/QLNhjqWn+mskYVBP21WDOVWopNOCzjb7T0715
qxrAf74YOfh0rq6MQgsHyuO7EalNQgJnXnrYgIxVHz+0NKsgPnpiI5g0mwRjLC/Krnh9a9xVxK7l
1jb9euXe57Nt4CQuc+Z8oWyFCFYmOw0Gc/kd70fsg9Cjg4F+LV6IMpgPHH7Q9kv/dUhC1cQMdfhy
Fcy2bRi8+bvyD6qWdi6i9fWKcAQMvvS8jbVYdwytCc5oxGMwdOuKQPLOcj/AvqMuDYYErgTXea9N
6VrZdjJXVkVlwhpPCLLjOyx+taDaGBaDy+7iJqztO9EaZ7+DhbXdRQrL4qpk3Wn/KZGEp7bB6Kty
Yt4f0QO4y64VF/02yyMQf2aI4lc8SEQ/mAuE0WtPW4HN0PZ7/bS5GLI5K3qStud21th3eN+lGeAL
ylRS0W0NrH0qFKKw5Id/aan0poOuv8/KFkDzQ43ltKTJwUmSXEbl9oJDS5WJApHlrnbOxujpjIWO
JDhZviDvS6hUoJ24zXtouvEGGOUF6ssQdYpDeWSC4NajYQIfCtwtxxS8m+0TYy9gwNR9uSi+8vbs
iMRqOsfPmnncuz4K8S8bagQQQYs/tq4iEKwRkzMh/MSsal4GWt9gRzePz49xgFDDBpRxEYtVbZEJ
3Qt0st7WWxMrBNdj7252sM9ldYIVeBk3whShBkXjsmJce1fQk8wZNAXFHWkxC3aqXxRR2ShvECK9
Wi+otYzx3plRfEtsbLm+13E+LwFqltioAd7H4eprF3eAlDzdwae18XLtnCqWMwR3pqcavemCo5Y5
PeHe6neqMO3/grzsJyAZqGhBfk5ZsZqhSkyZaYktBehod1wO75DrwYXaZVOCaT6yx41KFVuP0ZcB
BVc1DaQX/v3qkHDzVmn59tuLzUEmxy/MSEICPtf/S3TaShJi/mqlgFIKimhrd5/3GKIsutRX7oSW
uAhZprMn4GxuyS5Gg/tA2/uccuvNQkUzct6JGc17EeeukozAn1WJ5uyr/apLDDwrm34W3OwvpZl5
kJWfS0IgmPb/P/fJbU28BYWa4kGH52zF/QcJGuNxwXwMjCTgLqRDjspHvNYgUbBze7FUXwe5+LVY
GByEcM0vDlYXeC7xoUYFHvEECS59sJdIUGuhj+F5odMnpSHViR/SU8zkcalCtaoBcW6Uy9OgZifg
BjXr9rHTJJC2Esb3Hxzg+KN5AOAzNx+Hne7J2BxTLppeEbRfy18PCno6e+YUTO2fjjOFHHOgn6ej
DfWMZZFURRPpjI+sBifwroA11SU4L8ewXTs1Z6vktQFkMUDOPEYXVHhO0d1FyXDbgq16S/d1wvqL
hwC1rjj8NsnZMt3eP0l+J2nXJrIi6L+mH73H+OHAFQqgCCb2oyjfzzctedV3+U9LAZcWgXCU3kj7
T4ZqoQM8ntoaCPtO2MABpEA9vQOsJmgwXlAXnMEaxEZ+oHfDSx3KSBe14FP2VbYiZKrYEk2Zh/AN
O8mSw0fYJs1oSf9BY1JkZd+eyFyfSWgik65FRWBBlQ2Ubqv+4w1w7Jr+BRoW90qP+1odHJoitJJM
nBVJCy5yS1n7zsljsp7i5pPck5sjPuKM32CN8TurzrQ9Bmx4uivUrBlRT9Ke+2tT6wiBMLdielX/
6g7qIK8ssHEKze1AMZYoKeWX/jsalWVj3IEVXX/jbd6G3pXf26hfu3hVACxx8H6Pkdr6Mw9uhbkN
Po3uY4bCCGEDiMKEuHw0N/s07ij1ePXrMTwGfoA65SilyhYn7haz3irjY+wiXppGR8NkFQbkChJq
fBj/+OShhlYLs5aDyS+U8DKS1gEXfGjFgxQr6nmx+oUc4yBVoCEooouWBgOygbgoKMNIRTeBr/U2
fz6ANHWRGHb0nXXmM4bHWd0T+voZYxPxApheGpJ2ZFVeSgyex4DTKVuvq2CJl6rIjquC2oiIeOTB
p4goRcXYNgoul2PiAsbQOdIFMcvYVPV37sWYj9EllIytN+TR8Ceufocwy5Zlh/uQDlE8T1oAutuY
wG3U5D87KUNMtyNwY16EgxJXHkbLo/dRvuOo4hRfwntvL+Pr0INJsNSBceIUaSoRTdIDxVgVAYEj
s7tYILgrMNgieUrLgjk3NZgi9v8cqhojr4+rHSzHg4Bne60H9hYGUTQP5bpb/oGnz3yM4NXgNC3y
C4CrqgMuWxOhXyJhuHlh5II8kotLGsW21rAKtyeLrN6PyL4rahwItHX3KBbM7cBPW0kwDGz9Pq84
8eg4zHrGZw1xddCJG1xvV/ZNqV/xIcwNIBYM6bm3p/2/TFzkdepT5ErGJQwNV09EqweqxkN9xbWg
STtyYXaLaeszEhH/P/GTxw1a+qaEQhA0eHzOk1wKh2TxeQyEE7H64TyPv/HnTPtow+vqrQIHE8t6
a+HkF3XF6+KWnOrgj9X+HMRZxvOfmghvxxoNgwFsrNy0e7q0yNFROfN8VBDfu0dkUdS9vW9mKigD
Ww3yIVd6nzxzyHelQbpZ6tYYZjEH+UeoWESqUN31/JZTpW2CfC93BObVzL8yS6ziHcsMKuxv/UUp
gBo4FlIYXnx6LsYOJLdpi7B6mPS+n+g8beO+rjjzALhvnXkg7NLsTp7co7jKgZqy0CMnR2NJBL6r
SdgYpyV4kCEgYPfc8jXUK0ZzDh4S3emlaHAM+J1f0Up2FWNURtmDOeooTHcX4XGweGoENyuhqEh9
CP4w9rKTf+X2Z0I5elVGDq2fchfyEpCRYOU8xzXvGrnngHK0SVu7ZYqL+dLzu2iz2lv3sCqSxhkM
yXxL0iFtICJtB4PrsD9cMAPZPJE5XKzoNnKuT95sGmnF6yUYb3hMaRjyYoklrJruxy1azYNFKAf3
j746vy1erH1dFWge7el/Q8KhUpQjnf1PXOwDnfVW5PF2NUIzplfEf1ZX7YVCs94L7ZGQt7/uGMcq
S/OPfaJM29Oy6OWkl7mmdqstX/AHwZtNBX5K8fWWhJp2ltnxCYgpAtH5O6KQiLvLLmtRCQOFErnf
D5vJ+Xkl8xAJi/CRWVFUSKVYh0KrD5DMIL/dfYnPWAW4M/r67CxdBKw0Rb/naeADTUJtmBkBY1/J
hqt1lY6WzYWqhCMbGyGKbALNNNCw6CK+AXlwuGbR8+/UvpiG7p1y2buAskeBiPT0vMFONnkW3FGi
HxQWANS6PKZsKi3A5i5/UmGSVPK/v1a7NfidntVHuu2+BFD6gu5kmRDGKD1IwM1bX4k4+kuo40zt
IMYAytf3VfeLJpUB1u6l+n3DAOdI0dYc071fcQ9PTdbwR01n73Y+P87UD/ZCaTJ6Tw43v1PVSjVR
uIu1/FIgQh918sve5JujIjA9ZkakUohUTACSQAybyLiqlgzuNEW5r2et9iVNUh7uM5J6UERGJpeo
DNNsrd/Uryd9OvdGkqlOMxfTWMukJB8xaO0r1fvBvy7K6BW+AEhda3+rdXKQCiDpnunqLFCQd92u
90ei/yUIm8Bk2ydeBrb2MJW4pYv5CXADwULwwF9kC8sIxF0UrlWPPCjFVQ5twRAkhQvGsc7iZRY6
LiOdub6/tbjl5hsw8ptvsql+n3dzjREJnOMn59R40F+Oo2yBFVJ2a3ugMmmUMY1Jyf/rpyYD+DbA
QCjHOCunQr3ow4rhHqRVyk7+Pgom1NtQWQFAuKPkM0QDqaYQYwCfZYzELITSIZecXkwf3Wi+uuCy
FHYw6+eDfAo7AP4VoDTnF9CkNyMJlvXydkxThrs6g4lwjBUE5fZJUnGZSOmtqhn1BOI/0rBZNYLF
i4NbAQw04WWC9RWyo3U9WBuQdz/AqRP18QL589iaqKT5ZyoLppZ3wJc3jB1RuHBRZfcJtAqOY4xD
zUUc6tOUOPa1jkfJKVzvb9XNKC6YScrf6ar1TXNUAGHO26hxlJr08nmXIkZjogHmG5dw5mc5BaeM
Uy//kp4nbbzNRi9mx/VWJHr9Sbsmj48doexQmfeR7UEEx41CJcYxd0POi+DXwJr3K60hUcHqnQ4F
PsWgyhlH2Y+6K92APjA9f6Zs5gph5gwtnyNBULddxTw0Q/vrl4gRJJ6BBCf7COU62L7nxAbzdAlw
fMiy3DiM4R5gTKNmHIjdGg1ku18RSuguRSV1pUJs+V6WcU5h5AVHlZ91wq58JFgXKj7x04W6cqlg
dcl8ShbL+xkhkJY8n5saji0BQmTpXL4bWaUG/BXecPI8hCi7UI5obat231NnKDpr8Emtfmkl88fM
NgE/iS/lNpR5uZDifMTPSQovHrOAOf3wjVaMhiPrEz8qRyGwg7r3k2WcSRyi/7sthbT/+G+5PeTA
iIVgbY2q15AGiLUqZCMbTYXDeoV2hhFolWxuyn3XEAIQjV0J12vo0oWAj4qNKEOh3sIAb/bIn53a
1F7fDE0KwQzfuXW/TIzShfpzIL+t3SWBDwSm+H0LjzIH8u0mT8DmGyV+CjvlZN+jVgPhk8LD0N17
iM2O7bQ7MpTXDdAgwhJOE+dxwsBPSB/ErVf797BsGLHBR6k48cjny5AAbjmtPxfbsWxydz+AM7QU
snZDTBt02ZG2kVyz2uYgsXE6FjhhXwxs50x6EiW9NGjpn/fgDOXGRv19Fc1PqC2npnE3UyDnMyNR
zYp1lg75WAVO7ido5Kg7AE99IOj87C1Y5ZmqwLD6L2J+fHgWbhczxNVF0YcyQBkquyNl8Ma1IxSb
+NnOV3ELcQe+hGOY4lZT1SzXJLLYheHbOzteWLjQDZY6MzMMhkH8yP0NkKZ0kKVtqfyjaj1youFn
61w4Brv7SO+Pg6mHbIE09M9Oq+GXylRqWuKWtIeqOQ6hqNjHJtsmFmS/VbC3o5ahR9uZHgUuB7T9
8xyeNRGcBQo55UTQrDgAeiYK2BuUV9JGbvAZS9HmIkYq7KGOqL4434vPc+yQq42euOH/Ml2bPaRs
0hmBud5LdFdzgJdenWfGxkV23LK9xW82BxaXgLOgW4Y4TS1glX2GDJ2q2ell+SweqVBog9P1pHvN
aEEVaBxhPDADZaKkLYBZbCS8JjFnbJWzFoIJ6O/nB868rGLUa8D0qqf2rfo9FaLvULs3Z36w0vVW
UcMqoaTyI2tjCz4WNsNbtO6QeeCP6Mf9d587VuyJzPCE+ubetnpR2nh8LA3PXSC6UKbtpjmJ/aY+
UFBHC5lHU2ObJZ8FN7a3yqezt1JqFXZqnY9MmaUV7sPFvvISI3g5sBYYEk6WN/NCNGUEBzdujexJ
TyjTpFR67iBIcPrFxNwGzbOsyt24SF6UtOk3qM9mfEkcP4DY6lFpuaIMfsy318CrQ3dTcZSLAPZx
+zt50+p1jxKdmYgyvkDXDQh/+0Nrtdb84LBzCdAgTzzn3IyzovBc3bZmGYYY9MlKqRs50KFHeL2+
S1odvfwcUNlx3FJxlYORkKvL+oNShhjKMCqobYjufXkc3l/358dHTMKHt9VfxlmyW1+gTy8BPW8c
1F/zuwZ792U7aRenjVOtbkJJ4u1WKdZZKYFMrY6zoX9m3Ke43MF802qJjM8aFJ/YdeFPoypUj9zA
wF9xMW1AbFYKDiBhKx9GMpoZdGYNbJkxi/hfH4HoT8U+Z4xY5d5RQAS4KBSmtuZLlejPvTYLWb3y
0zHsxhu4b3wPD2DwGhm89W2BeSu8DT3t47RXeHIdwpwSnAReop4zWzimwbA7ZSL9R/SpVKkL3UkY
hPZlwys3/YT3jQWf5fD5JBF1L2lJ2ZMcYm27eAn/5b9AhN0B/bVhGWiYSos47TxHzeQz/7zYxvT5
QXRj3Tr29V8cwRAhdeXSX0cNKl0MU6o2rJquv99lpHbOd0DBd6ZfI5Z880YhfzT1lka7rD8WOt5u
qt1Ti/EDF09SeeYNqMxFfm/uiboe30jV9IDfYZvb9zvQRsmeRPpQucuRcTp00jx2Cf0n5rZOvHLg
cp7RYTWvSEr4qQhROCEUbPz5pslwxw5lnYBI1Pd6u1xcf160l4o7wQOFZ2y1/fdBV/XTJqfJ6eZv
e4bBfTUxXBQxEEQVuYR0imFbKg2uMWZPHGLx33Oh6yLR+KmWGO1ZpdMfKDGqjpUWnrulIwKVB7Js
Rw8WbFEIiuTO2FGtxsjxGoQAYNSUe8QcMgmM/pb4gkQZQf0cRQrrpWz8ijD7nN64GYerPIELWkYF
HI9LQZUwI0zyb0x+33oo4qBLha+DKjSJjWRv33MbYiDdnFZroXR7cp6WU03baeGmwH9SJMYc8dZt
N3AeIvD7Eoo9aUgUSC44rvG60KT/HrlbeBWApHkLkE7zLNzG983B0vJ0WY0YWDiaNAPbt/rQRSv7
O7N9M0IadfJ2x8In0N1pBFue3aUtRSuDQjiKeV6N1T6hjctCHu2YNvIto3j6RMEnHTotoum600zj
r0+VVHJMUriZCp6KnuN3hcap2xZufaxcc4Fw7YN0k+Wso69v+S8a6yojfqdXBkVRvM3oRcY12/tP
9mYRZTsI/MhemmG4KV75p7uy3TwXqunsgXTs7wb4b/ktzSxCKXYlJSp2XxYl76egtk6JB+i+pIoY
ec7sehHOTXMYuTcRMdNpTSukp7fQEWdibuoty5ezLGT6+MRC9kqgs9P7HFPT6jfa2Q66UGsh+h3o
Tub4dee45t2agI6qQBfY1F2NVknL1wXdvG3TEhR9d47WFB+13BTponnNw4UY4uQQjTO5t3pN6CEm
JUacUY91Qk1Za9U8nkehiR49vgCruQDSF4fjg9pPjFunWqYxHl9nl/IzULeQiZ2470+YXQ26A/NR
beIazF9gBcnXd5TeC7RfvVgbu0ksDAFH/JOTcj6sPbD2mTk2VqPV3nvicLPRvo6GhALLWZ/rM7nH
3bHkv02+entRyk+2sGITWC7Z54Ji8WSgUQWD9U4IZsWeVCiENMDAtBIloC/pI3YPshb5J89Up9Sc
QOpEvFvcLknI68pbIW69ZZdzEgcKf1D6xBX09Yh9N/VGhDoLBS4kyeXNNSpEh4DR5znG4h6OxMlr
7o/ku/ImhajL836nKnzMNpYs60khXzZX0+UbqUlZdbT8q6K2HxL921VPTdooRdAOeeCD190rcUsL
uBueY8XOM82rlBxm1PrWAkuvLaQpzncQD8OJhYOGAb5ksAGPvlOt7UggVD1JTAE/+AujXPcrxL+e
eFl4Gl3OiVf+gHxmu4FUobWzxGTszIClGgyUgaKcDM5rUgX8zqBhgaHhNl1QXIulf53XklfcX3vS
GKXT3/5kgM7sFuL4FJV1vm23p74W+X/IrXvtpErIMzEc1nTltCnQ8OmQI62hKwrx/tdx/W5IFMoR
1o3Aib8tKh0PkkkqymbB+aEvE5jZGYGZ6mQj2JWjp/OSm+x4p0vXes01vD77P3ex+R6vNxBk9Ph/
Usaf42+ypGHMb6tNjrN00bGYwdu9a6JVNV42iqAG12wOxO/4ho9E1U0TKRdY0a5jyEIIxS70R2bw
3pjK6XkQ600NLb9VmGWlkMml9X6WE9wcZC2izrEjBqvfgktTVUtxO7v7ctAmgHI6X/ocwAca9XN1
JUtR1e1SWg/vQ9ACg0fLPkYjMWpmFhkEoULvAKIj+tZ2dNKrApDSzP1/Evio56UoZsizrPFDvsWU
l87461nrVik2ra4Y3VQxPgVVsWaiwSQ7uc0/nNruk9hJu9LVjj+/OYay/AWRBUksSzaP4Hwx9gig
/oicjGibHijR0aTku4URJuufCllpFULthL4K5u1UXxQEsuVSOh0ulQ/Z5WICDTiRB1NqNftUFHM2
Q/KGO8JM8/OdzTDEch2Em5teXIjoCAN6NSs42BFBs2V/o4Dvcd7HfULh+TD+fbwBaC7+ELHWP53/
Onw/A4ibPQV95vDoMlDkV2uJV0MD4VdlA9Wgb/4VFiQhTO6rtv10rNrZHcTBlWda4TQCzgTpE0AQ
3IXJd4bY76bMT0rXlvI5ejdGpw0hmcQaho36er0RJHc0nLxpBmOFrk6qU/eShrKZdEtq+3MOgJwB
QkBB02pj1IH0i6espap4BgFMju+Hr8bi6jzUXXhO5UZkIJyCWrinXSurG8bTy64DUErEYhhG4nC2
fphli1TiwjZ4omMqPOgA9X9+w6oFWrCQoesrD8peqiTGHKJSX2T9if5f1f3vV2ZsXOBm6erv8Bu0
aipWR5HjzsAGPAHyLT3PFKUrXSJ2SpHIDqJGUPipvXBHl6rrCiAGtAvhhS/1T3arYCAO4ER53Uoc
z2bOn4EsWSv8W0iuc7/PlMMTv/WOD0KPFDQynxvpwrZR+I/tdH0JjvDW9PJfXQV8E4OWL4mVAxWg
r7sqp/GemuN68Zhs4NthJShmt0/zwQUdg/ZXXRrNxapmzQoApy4h+2Qn6i05YUud7CvrH64dAQrK
22MAWhBFpgAlxYP8y8GfPC5hciQvmoqzbpDXH1+w4u28wFzmfxhYA/2ipOFmhXPiEY7ikT6eKvvs
2iTR0mz2My3LGS+FniIfGrtOrOe4XQv2+Te7b/6rM6NPQgXviiskRDayJTfw4XmqwjKYEtnRoDbF
ixF6pXWR2mGjPJNfn21+1TXbK7jLdEBVIWuYJSZXr+mEnIbI+pSTjSbp78AwvfkszsCP+o1jl4RZ
GaMKiYng7EUKdjR0EWfGC5ouNo7cWBFCoIiGONxZNg3mU+nfxgp647zspvDfVOvLfKPBXfg97FLF
kWMw941H8UlMP6/6KlZ3l9vJNyRNjMc7kiiC8PMXwb2f7WdvUl75e5iq3qeiLwkO2eOVxrb1ij7K
jK2IvT2T/ilyNWTQO7ziwRpBIEZgrf7sFUxTjonGwywPzgi3v0h4F9rV0io8IQbqkBEkyggxO4XG
+FKlcMd5yeQKxt1Oarx6U5c4RZmPIiV4z4ILcQCbJ70UPOHdaJKNtTtgoS77fvNM8jChp+tSKWbK
HIiPwVoR05D6bpa9AgyzojWaT+QitF+cqxBMXmuSABkv9NrMuClVj1gIJIgoM4KiRZCNg8fdwzJF
opBRlvssvEwm6OCQuwWCy1/L8JIQYpHOA3cKDHC7zRzXVuUN3NgnpMDsxMS8soALyXY02FM4MTAA
peUZ4mjHyRmUpeBzLHDTPnS0zxFhlrNNLV6mtot8xPFabd+ztGSjK53rcTwk/a/+D6mugp5YR0yd
n9eY7C2W1539iqBCUI7q/ve61jUrMcoShpk7+gr49hh0mBDMYlNHqRQj+d6rJyx4gAE7riMJQRKv
rcEF07uKfr52qZ++/7VBrbwwGU7I8C0wt8gIUQpqOHWK+7jTvOvQJNyUyV0NlkYTkLMit4/E8Bpw
P0a+wb4vNisgPl1V4yXQ0YeTwvWVFSe03nnR8NlhsOICxP60ksjEuYt55IJkt0oAT/N8stKpE/ZR
wcRuX/BUXTy7umt7XrkK2YPmXoOgX9JD0pucnbbUkCVxtpMlYTUaLe66f8b1L6njN7ZrNUPqzAZ3
rYYiqruXfGdEMg9nGAJ2xbmoBvjphfQbNOFNRs2CAlWl2UTMQhlEW415SbhqJ0PGHnYeCT29UnZ2
+8iBTDlDfIEti/ZsPwCI6j0SDRWjoK/xp1c75KcJeRIhs8B9DaNQPU/OAeNM4lsPSgYdWtLw9p58
hp0mY46PERrxa9ayXBSFJzLetoO0rG2Ed7YOXcy0foZ1fR1ny8y5is5wR2gpvQS5kbLLjt0TwCVE
0U8rXgvMnFLWdDPCujGOfRoTKBkhe6Z+HGPqF++ykHcP1AwPlmlu3DjcvcgS9qNaXGq2hMyhiFK7
E+9ipjYoNlzCsgDeW49n/dfQgDRKj2VGoMyHejeFz/eSP7/fUmMPn9WtVu0pK7Y36LUBTZmcrCrH
hmVIsqWUiwo1gWkvSuCnQkQTmOANPKi3Y4xDyHqT/ia9kl5r2xb5UxBYw9Z2GfnaU+13F3P81+8B
u8RedgZO3XbTBFRcXS7egS/FWAUSdGWq6T7D0GBHaxjC7lhszIjEqFW9JuIkqtFLMqM4pPu6jpc/
uxr0cLuGR1d+Fov42aQ66FPI50YlEsE5/dQN6dE57zI5SmpLdNpv1hbbgEnEmA8769/Jbeo/1tLj
AWhQqpMSJHFNc26LY3Cp2icyBq1RYSQURrra7pUzKHfcXDPGKHWiwG7kVaVZofr+2YGf/OZXLiVJ
kXkN504ZhZgXsFLZHedvZbW5W+DoiMjrHx2jgncy+wq5Cg5bWi9BPedlUnTy+MHMJ4l1JtSliICH
XDKDuOx9zgKuzoe/U+OZQbc7W18+vFQDk+Olcm3C5jL5ouzcXs1lkvtCLe4atV1vEXs9Y17nlhAG
sozRxbXsGcTQtnQrNF49g2upXecKH/NtvnjzyyxT1fOYZvY7rdYZq6FSr0SZjXBhOsSEwhhYdtSf
ikg3yusKISmJx0xiTMiKom0RrYYd/mgZUdqlbbEuJhVjLnf8AieL9PYAg2pmJYn6dVa/cj1/N3JB
5N6ThiVWoQbA7RvEld6D9Z/0EJw4bzbXh1IAcNl4cZ01Z3aw0+F+4aP1S43/GMN3ZKu0YREpg6fI
Lx1zVLcle7XoW60z959VwFrH14h31kPAMke1whVIGdmWUtteY2A+B4cic7imO72oRRd+iQEFOJ84
qkJ+X13D9lz2vXNjKQMQFBsJi4IlL+mF6WEA+5F2ywptpathETg+Dxvav5vfv3BJQ0FdQUuTBJx6
aFdFGozKM93GQD9E19/RzyX0hcjfhUYCYnDzUOXC/XW73Ql000JcKa1A5dBh6LXUbneBBaHVmnNX
8bo5Db8thM1KfY5cShc5S6yU2D+4F8PyAQ1BZiXHLMvLxP2rNkaPiQI0dGnlfOYhcD/C/Z9xgu83
q8jYO25mN2+dz9q73b8nRjk6mTTtQVKLwGJuoA5ftyavHQODYgxuCBPDpZhv6bDO5USJFULG7Zhy
brvGWMkLGkyxtmVr/BwKpDBLhqv0SL/lEQe7eMcGxOFq7L2sRpGYx+XjJtQ8LtW0EDwlN5MqcrfU
C9tg3suNazowQhc6R/G+D7kJXZxFXfjT3LksBQ5YrFbInbhmH+6yTOwfUCLeWvGKAf16XPlKkMxQ
zK3ebQF/CC8g8l7mpffIQvc3ys8WPD2Fcg3Fs0qkbrsp6K9UhxPlm9s0/Kw+qEhQvwHp8DqWZsnN
i1i8Dy4hHJ+lKYqWpzP0BcDTKBoUeHJIDPyyxL25LXulUrAFWbZU0yxdEqm2fPxwB2YVzys0Ur5r
o1b2FZlYsLq8ROibGla5a3PTozaG5kRMgP/w5d24i9KmE/X0tfzXE0P3d0q/bkNZ4+svgoY6TjTN
/3WjrxtIs3KCY+y4mj9/y78R+/PeEZlmUZjIWAoAK63+nA3CS3roa7i8kwyYDGTOlYOLqq/QadfR
ICBP6gvPp/xVgvd4eiz689bKOueZKPOonRntKlT6eg5bz+OILY3pKg+mY3gOllHEnNEqo5jScgtv
ng+4mywyiAAarel2gdeEY7UIpQSOZi+/PxIUBOSIWiUYOgH2ICgGV2tiUdacHj6jR9AkqxqHxUgM
Lk1doeaqc22UBJAAEDV24UcshdnfpJgtM9fnNtD8Cmc8rhWzj/3VMcNXJfpRV7w4xw4ywfnWBeAO
P/sFxYDTQJZeaWFJH3vjFETfEOHvBLk8vo1mRYZ/gVbjuTkvIrYFY2WSFISj0crVzqOneC0ZfRan
iVqfyp1LZLzRjbf+mGonXF1qnGOc8BPecGvRQas8Xh3OuTWrSHOqXvCWksl8k9v3ejsm83T4KSnZ
mcTcNOJmd1284H6cJHtDHOWh+QVRP2oySPw4vcoo8GwmbolG4waf5vth8X2BHKwkt9DauRH4i4Lr
QV3laZaD9jjopX06JR1l514tyAqjjXLO1MMBVI8Q3Q16NaGnTyluxp2HYfF/zKUPJWwI4LceONvI
BFTj1opB5xFJKB9rbSqe4Y7EVhIyAuOoRyOm6aCou4S5QoTTebTX4WbUldHxb8/l5yYIrBJg6WUh
b28U9+VocPdH2QbLwunLlVPOl+dbuZwcnjnRE1wNYvUOPqCBkmy2+qXpHvkDzM4eGgcITYp+VS/9
Fchi5v2nUNQ95Mv4+yKoer3nhzJ+uhAQCOGpXGTPowQoaRQIOL0a6cTzx3+mTrP+p9D0aSmZJOeq
ps4dwgYegqk1jXN7YkAIg4Y6sxuSOIroy6MTgh71w4BVcTXXcmR4qWwnNjuz70CFAaRkpfzb5KSP
rO0AVPHQ/UiFmPl1lEqpbOZknjL8aqeh4dibL/+aj9IUfi3oDR9gPfvh8swRQVipT8TkfZ707Ldq
i6vsaelPr+XsyO03PJjXFHxdfWWsMXOuHjXfsMBDpfUjmw8phV7MVU4yEkB20qJDyucRqsdM5LQV
hrW6gdhkKQDD4ut2QnksCCDakIFQoGhYAtYG9oBwxbs9lbULvo/5Riv5UfM41lKa7n6+EnWi2Tzt
BlvUG6nja/1ULY7b9x7WWyhIVgB/URkLP5nUPMNxw/KcP8i51iyntVwFI6CdBsTgy3ocT7lzoJad
WdspwUx6pAp3tpBD39v0lG9wc83Lkp2J/z5i1oND7RZwAOQ8LKQZPgVYmkhpPbltNHl1RT6gWGsV
EKqNKjl3sH6KozNJ6MIaLsFsLmGwtQpm1Qpe1QczgnOh4k92vzMYZmNeRIrGy7jb9SbquZhOsES7
k8zu7irhEELvkjJCTz7nnEdFrB0xr5slgBrPH1N/h5tQT160eV0oSYzs7Y0qkd7cvvEGhzZqlZ8G
ju7FNeiiIqndAE5wj6VreI5jtDCJ3Zfyq0/AK0a30Uu2G4eSWzsaem2+4fY2reqt3f/UNuqZpV3A
X9KSgGY+IISu0wEGbwVRYRRwyffikxr9aA71QENrKzzdJVyVLyTL6U2vaQFO23fSfhVOeRzw5RTk
5se4LvvWWoAO43tOzJ1Embnetuh2omaggCWkfmh8nf/H+M95fSqqYncZF+REHCc+wgKmGfq0mmEP
+hDAVAAFhDCarvxUAD3fxb6877yz94eBaNv4ltZyLYtxOGEWwcEKll/NNOhW6w2wBulv5WdxRWYR
oZfGGG2LNUf3d0MKElMo6V/30hzwjy/TY0/yCWS7GcgwbROjWkw3nBVH8QPo/ZhLosakaRjIcBBI
zniuSNrAr90qZJv4m0HU88vkiDus5HvpSxFoR9YEdj9VtPGSDWZc53lADI93P0pPSXqyKokypIVC
hoeC3sxp6BeR7CCdPNgY4adL4KTHiHMnIyxkHe7vRWxWzJZuFXUrwT30RhC32DMYhvcFu7GCyd29
UQXnOKR9ymuzzlqvOlEm9pQPjUOY4p1MuivMM8o91WJHtbVbYUZJNhk7ivnJqL7i4gyZghQGbEq1
SXVQvDfVqpwKZjjE9eB5OxDqASSu/SUZF0mSdoSzYzNt503TGl66ijxL2Bp7PNKz4Q9fFiO0fV2q
jhODSpFzGxRObP8pYbbrlwW18O/tuB10y6uSZ0bsdACbsHdCz09SSfqEltMyq7URu5FhVOi8qmeE
ANRRJmMRgSA++K07O+UvvQiFKe9xQpLK49mu88ZPe2JFLSTOWACyqz4AcUUQ/CY+DDS3gYy6u9mK
0ZudI1G0MMeZW8S3PxUfUxlhUzXPwz33bXUflfOMj7Iv8xwESnPR2a/4qXOrYFcIlvLdzjQ2iVjG
CvGbu8WqQmv3iM9yTxeNA2NsnC1SaADrHQGCJ6Ox1uZh1BvZxVGTdN0TcxTiKi5/Mc0Sy7pgEscU
Q2wnkkSq4wSanYU8ZyYETzZH2u7rauqbZu6BBfTH3aXON2/Ss4znkF4BtAPogdbPpvgoj3ewL3no
qZJvC2K1ABWoH0VjTZKZ38YKZ2ci4x4r2Pjcznh7J4kwOsY11S49dZTnwktj8pxVPu4xh40GAP6x
RoBTUzAPFB5Ivw0O/d17As3AxEmKyFJlg5Zm9N1ymxGWI6yZKo3t90rvAGNPAmHs9+kH/i5m3Wfd
QPqQeGcetkk+UwVrugFfo8QJx1MpsoxzfzIjtYshK0fSy65OgdYoa2VNoyPcDWiFVXIKSQ2ItH7p
NJfzWe30PU6cVJU/hHlX1HHREDQy8tNBoSf8sQ03eeEfv+TzI59yMbyHutTR5inpPHJXfshgAFDZ
os/iVdEdnVrOH6s/32YD4pzhJJ/u3WcuGcKsF4MhH1QWm7G+lZGizn+bFjeu2xe1FttYXXn8oznC
5lbPG+/dos5J2v312x3kPSEyiMFDYN+Gbpcbfoytpe80WXTPk4xb4UZXWOlu1jmmkuPgb0Xo9LDh
dCldiKHcLcpWHsI+1h6HC1vHUspN9h01UFoze2WClpR1YuLARFDoXieklReTY7QgC9brAqtFKLh+
pUZQt9wI1sHmJ5lDhzcmxz4BWZEcQfG17a2L0QlPdv8Ro4SBLlvLIk/ijS+RxucbDjJXnqIa6PL3
E1uF0VuTy7nQbpI2AfJ+pRbUxRQ3vQ/qOsLHSV+MpSIBoeBo7ob1eOU8H0vmnXMqh6YzzF818deB
9lOwsk4vv242gMxp/aTanXgKxqzZkZzhddHpKJodE9aIBO/9Km7xA83k2vC35Cu9+/SXfFl8Y8Hf
RYvMeutctt6kpDna7yyL/gLAm4V6WeMTtAjNUohwzUsDxn3mkTjIVF7E/5wpdaneH3u03kX7B2Au
+jpOJ6T31+Sf2FQqC5OKL4A7Ebod3A0Mv297zS3IokkvDb/AqT6X1y7cye0YwvkjOEA+ja738/4j
MT92qaYZWdfeZhXr2JEP5/WL/mf24rBSm6zCuXp/V55PLXOyh5Fh0yIilMCN6QlLOGFjictGcmds
dnntq/O6dRr19V161skGyWzbwWXmLC2MHnhlTQc2SURRXuhUNKB8yukYZmxN/o/Ljv966VhsrdYa
/7tv6L9pJKfRarUtny2pFSKvFNcVf3QloBYkkxo993UzeZpxsyJfzjiFMfVhw2m6pjOysoNNLTX7
ulKNt0tOFrVz61qO4ZPP8vrxWwFTIgjWZXqZFV1Wb/IvaO//3SMVclcgRvbEIfZ7bp/bgj6yxAKD
9BMZ0NgYUd+FlZlfFpXt7QDc2KO9zcUxV3kmY0j8ZruzoEukwBhqdIC30j/8Kw8VTQqZdIK9ddLm
iU3zEi9x7re1sqGOWK6bOxnRStzjGvd2r180EJuCiB3TAoFzWSQ/xNpLLmrjIOj18z6dP4k6HsFl
qJ/8zY5trnVUO/iM5t2qT9mwnLBwRfPL0dTpOY7INaqEMWsucigryvXuy69+Q6AyAsEo5TI2v9Vs
XhSRUtM748rPDHv14BbWpJd/HoyzuqT7IFTSc9p+Cc58vncExssaezGEnCS7/0Ze9pNLudMn8NcJ
DRUJeS7YGh0rv7VHVc2jOl6paT9bDer9NZ0MlrjjNrDi2dhzp3+5zD+5obRvICKlaJ1jUP9pEcA8
PIyWqDawiumn/jYMhhTdXwdrhv2kzsu3dPWpPGh0LUPBK0FgerrZDVlTWvgkJoBU+RaZnjJFMo26
0+WMYY1kbvipC6pHQy0idNvKbb590nxtVs1y6An74ZbzkD814fGdfmqMey6xtZ4RS0SkKpmL04pO
cR7OF9xoyLIyPy6ZvfyPXKNMvi18kEyW3Zspow+puCQsTXX9ozT5QxyepcByTvIjuSNBvgN2+C8r
5JviNZaxuKPH1dGsHPYMjQB68VNINRrTcYY2PhMnMxgKVW9PvOJeB3RVzkc1OBV+68Q8j6Y45HtX
2ppQePd655j4q2pm6/c4uCa9PdiYVMLDZiONTTwMsHHPniyPisoKfSclkWea16wLRqvAdwxc0qcw
qeoGlEAO5v45aSTwvUjh2etS8UoQkQU7BVRB0MezBcKM5vDzcG2gRS0EqINbuoZsqaK230wpbUNZ
xr16utp6cttj10wk0JkYPWG+SRZe8MOQIFVMjzS9t3w32Cif+DHdS3Wn6hVty8ePKPzIZ92c+xIc
VYOUQtclPTjEmHLJFjqpHWpwvgsLaEHeUQnlF52l2jdIZfbZ+2tH3rxhe60FedqjIPIDN7O4JAFl
/80EzyrCC9Hn+F2pt21j4rxXRteuKT6c/WEFX/7Hs8xhpn9P5gsfW1SD/PLWVZrdcG5eybJuLG1+
c8e2XZXSaKaV19As6if3M/dSP+UNioSb/TZFShKOePwqLzxO2S+Y3SyoTpJp/FRgpHLZpM27KCmK
fTKOsbG0FDF5Nv5EIWPHgFvuCWP4xSc18QXdGO0HlNmifRDdo1Is6sk4KzRKOLDy68gYBLVpgit/
Cr2vzjH3cGfyDN2qUc+fD8MT22S5RTblJ62ExNg89KiCCQtX3eoNb+tOup/F3jA/WJejE9JRCXrF
REe3Q8DZqNL26TJciX+FgUqPmAw/ENfgf4emtmKZuR0MHDgCe84qP5YFGN2WWgrhspoFUWgtrR8M
IsHH9GoM5cmmSxKpNLj96zClf63Cnl4KNqkmF1MWP930HK+SE8h2qZM+XSNojhlGD+RwNdXLOSbV
mt9kQ98i6wKMW/rWeVrNojFb8CjmfCf0YRdTszdXJKM8Voy/HUhq0KsPODSXcWUNiykMFmhmFI8Y
yvNCe9IByvRQXNHNTKp4T9s9aRL8dK6BarqdnOavoe90D57IBwl31q/g/cqAGD+659qoltmqgmpg
/M5RTmSGhyWLmeu1ZjlVgLe4btBpS51UVwGvukPEfg1RgdQyzbDYwOUBIBzsTAutOKRSngE11UxN
tfDY1Fhn2tK47eYXWQGcQJgimNTCkDuY11e10MCNMxUHfRK6Xgg7fdBsG3xLKsJYuCeS+rF94PU8
ZoSCvYPz1qV00JvNkHPOXWwOaXGZyn2KTfZTwA13IHxbIlIztH4JwkVAl+udeMh7+wy1xS/F7aNT
BPI07wf6k+vxMNIcvFX8qEaLBwufkik1BHI+udwECDpvd1kC3zkAq1QgOe3LChwrJX0PlYGYGBWg
45jNtSEcBwRb2vPjJfS8DfAVcFSAfNQy8ZuzrlvIFRH6Bfu0ZNsDwaKZKsmLJC/C+BS7/Q5+Kk22
Bt/XorvcFvVUuTly/MeEyIMVqXfPiFL7kISGhuabFgGsK6pISDGh+23QeBJffnJxNXUq3A5Km0jJ
LLDSn02YP30sgtyQKp50tEOPpacJ45ufTBVamJkyD/ffEPcdFQYRET7t/Qw9aPFvAqkjBRSkKcS9
Cy0XawMe6H/od02tQK/Q+XeP2DJ9pFCpj/LC8xIn6fq21z49DgOSzQRjjLogGVj5xiXrqYaKSjam
eS9ijq1LQizSFW2Iux0CSk8BMdHB+2B3cAW/IrYnqB6LHm8G+E37ZxVtrYzriyBBdUtLjrZyS/7X
H0FTH+r/oZtkjA03guwYefFGA8oS5vYtGsBlG4e1mehivE/U1qr7WWaERKVBGMzBfEV6YpaOZYit
bBSeqt075PdNAA6BmDNypWT5p9sZCrHCwBReECWkWW3Mm3Vb6jBH2HdDBX8mc+FIWIiKyIiTAWcV
A4T595A9VcywBxGJy2P/Arth0YwPWOVdvtUnuuPGl1Gn8W2d4V6jhJk3Tw4VKeocW5rZjKQ1Fv5Z
HrD04S0ntK79ldjqN45JRofULJFxhvINePWh6J2Zkx9gnd4AD7g7NCOeSnCf+uBXgoB7C7S1P1LJ
bsFm/ZgzwGr5p9nDPSoqgL3IckRJFPT6Sqd50+/8xP2hOggan9nM+CpkEWh3o+hRs5kQe4IzP5hT
d4aMbIjQ3KE12WXTz6dt8tlRoMkpIUmJphIq+oS1nsFIiBXnV+GL0mlgCnbR7tk37ZkXHlJJBMOh
88Wl3A8PProLQ+xSHV5AKaeRQ/p3PCqmsV75YtDgdKfVx4CCZx9feIVE//4DPNQc8My4iaXE/JYY
vb1p/SCA+rjQMCencP1aWdPlYaSSyuWu5m4Xmtf1AwUwh3338G4W7yZ/WsEnae+ylq8uZp8tx54q
QEKc3mqIAYGPM+p1x45cZkRDE3xQuW+QpGADLQs+GqPDibXyDptlfPd1D1p6izG+vO6HzxZ18cnn
vo/KmFIbPuJmOUABg1RaUhtpGJZgGR4uZ4s8U0xArU+5TQ5XTr8YDOsAIOQtiu8/fQ7Nz5vZBRHi
pv52UlURp8jdfCrfYyMfBUQdYLhjPGsVEZYwNG20aiRbnXX0ywqKykj4RGc7nJcfYnCEwzRuVXyT
dgz8wwDiFkqKfeW4g91U2m4P4H5K2iOG4MccoiMopg7LtBf9B6bBDdyPp3CTc5uZB+BhWOi6dIOu
DdumuCBziLA1rHAGvTdR5o6YA2Jui32gn3jKksUgI4D7IeOLGeOLYa1Kele93YDs1aDtaAvdkvez
txuhhUhIRjOerfq5FzTsPeJjek3uFYL0ILUmTCsk6VB6aFYkl/sja40sAz9VKpNiBu4g4hfNBUj1
ngHuTKR5mrDHRO84KcMet9ixpS+YkCDwOWl2xPaWTiUCErF9CCeB4zq66dswE7iT21+dJlYEzR4/
PmxDd3vhZROr0J38ukPK9X2x8pf7/a/rl54NL8Fde2MLKDnZ3X71adzTg238A1aOObCoa7n62+OE
fXEiH8LGiaeYnEqiD6Uavp3MlMuHMYEzE+fjHkggzZ09qoT30Vgyivg/3lh6deWw18iQh3Zar4RX
PrhBt50xMe2HzYhDw8O11amz+JmimqetcJ3H2CpBPOaiXDk4wLs1mi4hu25TNrnaIQODf6KB5dlv
UR9Y4ceUnoTZT5TaYwk8UnveIPi26UCyoflwXaxlpuB1FEuxVhRNmlPJpnsNcKINKGV/3juaLh58
BAGjK4Lmha/7ILweOzwu0KhVlwIDAAUZJ5JG0Dx2t48qNDmOwCXERIIIT7EchWAwNGBV0B7dnPHX
Jxho/KsKevu6PISyuZBtksS88QNPBoBU3mYGIXOQTlVQT91ogAX/dbGPayVoz6nwyEL1mIZF5BNv
fgAAd6XB6r685Kw96MOdHXrp6lsdtMME5Y5eIPX7VtKq2nCRtPIT4wRTm52uqIYc2Hma9Yslt93J
mAhFYNGS3GiFeXeXFuuKNklhI+dm9IYkmrhgMQd+5WHILNfwRntupdswTdKHzIB/kPhwXQoZ9xnj
UAgNPr9nuAO7WI+mShiARwOmfEOHX6AyImmfnMLJjOVV2qfHjCLJ1ltyYXbvB1YrkffN3EhRHWor
orHJNtzkVWcNLAXW4h0h5i3VjbocBWYw8qzO25HkevqdHnf2fh55+qpXdJf9fWterIPDxU08f40t
6+w2xm1MDEvHJjwPgIlXfETt1T1DOayRpkLxCV0WwUS/pllQtOJvQHpWvejsKeYBX2xg+sRxj0kl
ZHn9O0siEVxtV9q2AZKhsUk22IXAzXTck3CznRX0nhHJsmHgOSQZ7vE96np0vqYNn0WhPverwcx/
M7NK4YzSOH2xha3KNKvW14vSA0uL3IIeEfLrdrczrhqD/3djhyQzEU44FWgAts6Ld9n/UNuOWJeQ
8s4aRCdBZ4PWCgCsQsqCg+OSldywF8pCR7wxkaOmt9nlwUlt1wojqNZJP+5QjOxyk6SNWSVFAX3v
ZZ98MrRuGBzenajDJNQN4+NX/O1h4qZRzTGRmn0nmqQCEeNZI9hEzbeuhIY4jQuQaUVWHxS+mzOL
Ae+OC4QCqG8yxeoCTiokmOEwgLJjSa5HaIS6WTtficM/xLZEIaa3JuP28gXRANBhiVDzc/bzSr2W
13tVJtJo8HnSFIWe2+jak29raSEaJxfM7V4Bx4qqkV/ugULag8JoyJuvsVweQPpjQLpUSizSaZuS
6Gz29IYLbDRkauiEMIYwmxfWBOvHxMguWMYY0hw3MRSLYGCF5ULZxX4R8Pmk54yQgAbpCSPZGDXu
x++zQrXsWFZoITCwFYQcgiNqG2LNeB+QwrtiLSMzw8vtshjJB8rXdeoeRF6AACmiV7a6mJlQ8N0v
vqyJVzb0TjXAkZ4+3hzzAw8yw0/G3G479NuPNrhlkayTuvD15HaE2PcAL0d+rVFErndsbeT6rtrM
ynfvgNIOX6A7t8+4UlY6MhWqSa1wdQOkrzoL94zy619k3PqgbuXYArBwFItomtj+/XOblNHMnZJK
lRqYiqudpw1G369D2UqvULCx1mP3VtWTK3pHWnGwBmWXncqj2W20GHPbYPLSfsiXT8rAX6sOguZL
x6ekOustMmYz91Tp/ELGBI4QyUl71JZRI7q9RnHowUnVYYIjlBfEsgs7a3rCg7mxs7GJvIuRj9b7
2F2HNTQjtkbzbx7zEh/CjmBqJfU/J0N0m3zTW5iKaG6U8SBpvkrCbXExjmzpS2NTP2cIVWlkLzOD
eEpJmHF3Tv49Mbnq+wkwnEcpY1qe4U131/L6CyYkG6zqNXAbpqQVB3MANbZEpgQLqqC3utyD8O5T
vcv+STs1vtKY/tHQDYu3FQU0tMVzfnhXT1wNMlqhefXbqZy2pzPai2gbAZIi5DG2GGkZ7gAL/LJb
kYQ0ZBUED8NnKzMlnmLBlOrZ7JxghoadCXk9bYL878tCfI3zFrZXCgPwQKsVoJ9gnS7vQ9jEPGSQ
QEyxi/mq28E1NpYvjyUAE4oP91GkkVTRfjbzwQbPBJg2g9Z70v1BSF8zZ6wn1dxFjcaMPA9LROI3
RjZu6cFAbOsUGkVCp4Kvqak2tWBlIQWP24nQXscOQ1jxKR66xhylORy+GIOjb9s9gfsrVUV57+Ak
VObuuJrra/lVwy5h+L77G4c/uTIvSrqTHIv5LWThNB9w4hVDbDbZUyexBxvY4mbyGkVa3WkatPiK
J3oOIf29eQghUNvLjRM+RzFBYI3JFm/pnxUj7wRvUJRBh37oYAd7GcMsQB8F1rAwuUBPd5zryMrQ
z8B7egMkouhDRCOuIxk5kKldWz1H5SLoswZxBECe/4yB7Vq82p/isJYnt9v9PILbcf2CfO4lyyZa
p+CXSo1U/EfXWOsIWdwaA4Bgaq9ozfKADzxfvI6TG1kYpD1yn27qRsb0HoeilgsdmjKcJGxC5osr
qV/gIfnRs7Wl9U++fVPaVQJffN2h18H6REmTrCLn7AEgKryAMAnM+8wsbHtaEMqs1675NWtUr9S2
xiK+Y7Wa8gVoqD7ZAWRQwyhvJm5n1bu5lchV/fA3sHSxibcjdPXgrUwcQf5JFGMwEMoG0mfbP4g4
ptXws3Q2BQN1RQxhHFm339KpBLAqvo9fbBs520McsaevZcaJ1d8VlHWRsM0GXhsgdvfdl+OWyuPm
fO5yPTus0RZx119v+6vin3VxiltZ9WFjiE44F8KuNnso8xg8sIyKLTiuZdUcU3Frusba1FjBVwdX
14USFgInpacdtdhdVuC+ed2oddgj4HW3heENWKnQPcBz572xnBAu78LjJU7IYE16kwPDYXwma6D7
oYufVQoWEzv96PmFhCh9g4+j8x4DzUlrZrEOfSPc7u0zVBexj8yChlW+DvP0Cg/j05JyJYxQ/P3j
RuQw29bABG3SgxXoZ1jGnXNk6Jy8R8cYutNDR7pvxcp5hdJ2HgO1sAuWflm8u+ZBPNNe3LiamhAp
vocTJAwvotcI8VcHGBUn+V1x2jFLKZyyxk9B3DfUc9AONtSYzar3NWBXDpkvCjNBgJTghlcwN5VR
Up1ZGWeauxUxt397KG5FesI71d3thr6cd5q6FYKT4AWDnMj56aiXW50yXGobLdjCMnpdvDM2rGwm
d0KWMG+i+1WhLFJ3+gA4tUFJdc3NI8OpU+g26j3ou0Q8xSuJdX+hlcrY4neyTP2YSk6EYH+5UM8Q
OqzB92jRGaIjs5MF5P7lz61jnz6UtN1DMC31sYjyFI3sdrZTCWR1Z1F0I8rEdcWhQmSkIdd1h4Mh
ftOTy5buZPmz4H2p8YRzWFckSSJa9F7c1C/2oll5+nC2+WKGwOO0kBq0so+tmqjZXWp/cTO293ML
udQvWnqh0USQBrGVY5aMTPEMuXxIDZpH0EL7tR1gng/5U1Q5YOvw86v39XcxWzjT1BgRsMxJwsHu
x0W9pof8eUPiRb+t+hbeeNXsVwgXm8HNNiaYubKOii6gUiA5WL16veJfuSlwjnnAI6OuLgWVCWJ2
FgiCUgnRq4iskJMjL7MmdzT5MPo0Ja/+UO1PfmozPT0x8zYEsWFO8ZMUGvI4eH7LkQYCiLqTM2NW
Sw/cCt1BzK4jh/1Vs3DOn3Nbs8Zn4BDJrIG0vYck+WIOkFzXSkFDCXLSrUIKTUJtAMnpmC7/UcBp
SOr8/dQafr0vvZrD0CKr+C1pxmnSUBNjInu/A/kjN/CcSoT+Zmu9C453S6xBHUjvcy7we2+E6PKe
0oLTyerwwiGiiR9opbnkjitleHXoJapkjUYGgyBedyJ+qIQ/9NgNAJ8rHVOgCfmoknIiJV29vRfc
h71hNGF829NZ387dJyk8VajotvEjJO0eu5OcWHBfGNNSNyz2ye/UQz3xe6KXlQFYWO2Y1mZKOOAH
w56xrMS5v5yUBQ8CXRRz26AHTjSl8IXUSyuEJ4qW4QqcpQ5i6IIkNBvxyCQFCPPbUBH9Ymxi5Pgr
iD/l7jqNO74R9mdDYXuCLZdzdiYIVDJm+rCLp/6VOvlC0cbpC5N8gdA2DKSsJPlWr1rwFDMadDe7
JvvDB3sqxuxGrEwM/nNtVQzmwlgVsoY0QmVbkT3KUgoDkK1uGO4tHf1WLtnrXc2zf8GCACySsxR2
a+TsuBhIuXwBSWOYdH/8HjDlEg9AqEAnxmHpTJJglMONyAIUq97oEwfp/Au4q7RF2vjJKo+ZtVvf
EVHhPAdV0k1tJ++DvCg5f0d+2p0Y+kcrBMePLW2WtlMG13QHy3jufAqmtgRA9g/r4+7MzgUGtL2F
WF/65CT6rrCwD2SJXOGnJqgYwLtwtg1SknwCKM75DfHwvaPssnw8aryouW+rPnz0u2B3ywclkBPT
xz0JwyoBitDH4iyXYAGmpjOsFO5p1Fbs+0dXBjGwMhyPTOjdGZtzmH+7q0/60l/sk+tnH2c9z8Kv
4k/Xcx3bjXIHR3eRUFy1+Hu8BuUUX8bz9xDwKE4tWISxHuhz5eVmYS1u/SveKuQP2E6YLJzAANku
8YI9Fge6t7cAvR4TdrOy80FyYzMJUzv41I8xRSqUz4PV7/B1WOO7XXpoEJt7lUqx9LRHAp7h4Khz
13Yqt0ltkEYvHANReDyWF2xHgn1ZnphMEnx1dkUH8U0EXAj3lw69RpdKaJ1xMDPHqYbuPKU6PfFJ
VSWnS0iwzcC1WPyPm9ONaUux2w+3+89sonAaepa2AfOAIXcHtZcaFMH8RiKL67qbyjls9d8QfKki
t1N5ozMR4P/3svOu6hcbX2CN7wyLWF1yUaNpfiNUNwkiG1q0TJSaQbDzqLhc4BiQRLODDjoaT5Hr
+UZgWqJ9haxIiXgxl6XrglkvWaAio5DEgP/v7rwh1g3umk5o76lkxBffMr+pNhdoCLnuZ+nGMLQd
Dush4ZJqJKbNm0PPr7M8oeLUfhVK3CtbFo5mml9nWkglDtVL7OWtXdZzrOk+BMt2HfLixDa4bZI4
C6A5L8NpL0CdknPbZK4gbwWPtCEVLYo04wR6QE3FqFus9NhHhLbNHFZty3uehVphcwkhn0vQSaxW
ga7uIomC9Y0BnJqDPvvSM0jdCogDd1Qw5uAufaG1Xy7F3cDTDdq07F/2ENDDpSWPsPHS8s57yrFY
37w+oyihfZm9CDeL/vmJoIPIz4/4N92lS6eVXLIyJGnIRFXuM4zaYTDKl3qkoFH/egO5U12p/4Ua
USQ3ZDSWFWn+rlwEMG7FoermpV4qCCEAMEF20VyRnVI8n6AVsswB+/8DbilxHuRiq+I0Em3A9tSM
FijjJhkKz0r/L67sf2P5ZyuGBq1iyflhjk0oFLg5B9fc2JuryZEUR25Bn8e8soQBYEUOp8FJaziF
Lo0owgWZHagbT9wcWjnVjnQrsKlfmDlc7jlWz6zkz0kbqUxdZ8IN23Tr5bHI9OInLzlS8PI7LXec
LOBtY2x9fD2v7B1v70sO1eqRKxvknTaZQuZ3900NW9fvQPUSUANRJWDpyEkw0nKsLQZrs0s/a7S2
edJ3Zif8+O1x4eNX12KuTWWChY2PADDuCCu5CyeMgIXZ5aBKFdnoxFtEDoshFQxw1fvYPYNSvF1z
KZtMHWdZZRUBCAG8nElW4y9Zh411PIujmJy/Pvsj9I4wfzf/oXzxbzdYS1uztzMWlFSljeTa585f
opPnNITk8xg7UDVb7KZgRcF7XFCO6UlPfgUP96eOYdZe1j+pT2hKH2DlYw1lDm1m7sOC+VIuE0z8
FLerAOtlZWI7lEEUj9Aqy0kVRQgyyQFGKmJsKu1+sGtX30+eKJAU8EnYWpQRd1/mXWPpNGOAbJ1t
P/7bqOs0U/HwU7hNp5EXZUfXbFKEV7oXGKsNAvXvY/Z1aalQkZgGZ6E5g8MzOXpgz0Ipj2hEj3IQ
5ZsitdjXifzLNyE2dcwhwR0EoPHeuMsdr1ldy40onul8pGxriDnf7HvIV99owWXTuBXizQ8IOS3y
wmqOFM3VN5wHURq7B7FHVtinmQ2G2RhJGKLtrlgMIa/nWPQ9IWJwFOPEh97NCkFfXnJzfwWrvo/X
T5+cn4QQSNbAtJNIdSAmkgqZD16KYWLxGXZqbJYjkbEa+YbRn5MfvSMOzL7yCa8ikrjtpKwAZLfK
ktfjoMH54H0a1qS1qy/XuRM4o/lP0vTb2Dw0hgYGyba2UKYXP+B3TGJnS5q08JWFJUuWOyX0JXP5
YmNZ2MIJBXiUcpcgji9CySfIe+8fcx5lc7xy67qeOpqgLVd+xHEHhKLGiZUfkKjKXbBQU6geD+WX
hDDmqDY7sqCD7PyL6ywzdly5uu9SqFu6R2UYbr6BPFGKWbKhtLTEIIZQKtJ+eRUw2Ko4fchxlCDA
reQiQ0RKV8OiD7MOEqkWQz/ypPV90xa9SWA9zec99P1nf0hGLfnwOZpQxkqIfHgYmR9YDbXKc7oH
JUpWxPWxiHotDoE1/qOhh6abDm1wmk+ua+c/jM/bgy2K8kvoa3RzncoKeK/cMNfdZ4dZuVSV3US4
vyCfm1QvokRZVkfL69cccOGR6HtPpZJk0OWGhLWXMb2btebPJDt4XMTM/g/rC66UWp+r30/hqni2
UMhf8ehK+BlYeWMPajc8s1ew+BDzNewhnkhImXooetpQrD6QJfnAkRvQnuLMqJfAfqpUm16i9tc0
0TtM+TGU/8l6K0Dujr1ztgAMuKIYM4LzIqJRHaNh34yllvCe1tCtH9gaYJ9g8n9ow421Tar6usVJ
NOFr4OEwwlCxS9iMrACDwdkHNgnHJ7dBrPGu3C8k5SQUvVsCF9yBx6tgCi7f8btO+o0mkCExEw+n
J7X+7N3vBx1sqdwV58rL2Bl6VA3icje8aQLrbE7t8RIFgcNISWZ4J6mKb3cAjQAmGts2c3X/bWm2
mU9JBFRvEyf0rsZpsT5rf7rzrSniDEHGwa+aqOLO51VqyRF1hI8z4NIrdnDZbepXiE/dysklPcX6
hKLpW3rK/3s0k47021+H+M+Zm/XCvkrxUR5L967E2UJD6pDMr3hLdnwAH5r+cHro8r38BRK9vRsy
iNdGjUqCLhDLdmKdGx2kyjbr5mD9VsKF1HrGMNW1xU7/trMT3vvfx8w0O8l3mz7Y7NCNX/FMUuIH
JgWZJNMk172jOE0rKVF+gfOXCss9XzDGryUUxec5JU93sH/gga7rrz03lvmBMYN3j+rHSYyqbEpk
eYEL9wgb09IdhePtwDljeotb7EprnuYrXTtw0Q45Z+QGNjzYE1VlXxz7dxuvun0zGmvTfVBBfVPy
r4+8T+945pcuflCq6Nb7maYTPWUwWIbVTcLjYiyPv2EJYg/3OQWOJdyFJD+IxCMZ4oWYqwP0mIRd
kaEkAOCfle5lleihW1I5eY4xnwzF5DN+2+UXQ83IlSn/EwV4rmvEDi8iWRFit/3d5rqJbMoNGmfL
Q9ieVF7TDqa+yvyvIkh8lmoYmFctdKc9da9HwWONA45h9XJxfz4J52gKfkVJHcV5xHWQhkgTbuiZ
0dFPlUiX1hxgrWbmoXj0JCistAYBNsDfSeP1OnQDZ2HJgN8xdxG59op02LipZUtJSFB5vM63oCTY
TyDki9m0Il2GgVRg4M29EyuME/NpM2prR4+uQM14zKXys1+nRadCb2ty+WFXHTQeK/fMUBiJSAxC
mXWpLJVCY4KHLIl+ZMHYTD/h6AB7Z5WeXyuBT8LTdRIJlhu3rGlpfdStWDYuk78rm476Nj/RmZf0
tS2h/ujMmOfV+lTa/8CO4S4EGKERBCBgDdFtw3ytoeNPxSBQNirhPfxFI8/LLRzZd8m0QNY2EYhN
p2nSs6sGD3tMsXattOLEWbj1pKKhQMN+vJaX4hHxQQdgYhU5ukCLCWUnSMA97Mr4BJ1LF5ESyvX4
ibh5AsbbvITus7fu1a0Sro50K2Zvp60azaUelh/H3g0fIaBv72TQ2oofIn+nVk7lCrsOTaJeBxk4
THzBTxDstWAdzZ4UIOObiLGZlsswOx3gwCccD9tWOWhnNv+BGi0o23Ijjtv9gQ1BCYUT3X2dtykV
CzFQ1072bCnqkBE6T5oQQIl+WO8G9NXnNyfJErUEcxkvIaA4WufN5EgeSeBXQ9CEko9uR6uTjAH/
t7ufjzV12t8qz3gCr++lQuciH1G2njAIa0SG7XhsShmDb+osg+Hf+VdhyYN/tpnVEVxcGuh2/F8x
/EdL776c9wW4BsJpeicIO5CEO3QsA6zET/KQ7v6CyhnwNqcZmVzgxxrzSaqj5HWuEjzmOXD/BubR
OxyA5uQMWOx7nDyUQb2mLCRlGXmkBo2YPAdSv4PHWDBLnvLS5aE8jQ8CExNEbNYs5xvc2FV4ZBDS
DDk8xy5IlRkxUDV/O00g1uzYdeJZQfxpEvWmrkM17YbXr5Xb5HxMZwkUA2dUT7ODxMIWaxakUwGG
Hup4ECpO8CiNHodSV7xaitIkCsgBC3Se3bUgw9093zvZuecMAjVqZvbu7t+GS9aGXlLxXHo38qSN
hyiudd4BNcm0CMG3CeuXlMnCtY2hrJrWViAlRmoWd2uzQPx577pbP6Zf8PsllPXjDTz8ID7QjNRt
t+e+kL68Le10Lw/L0+D7yYiMs65bLJ/kpIoZh1OvdUGEeEvf0QXT/HPY33tmNsLtdRWOuDxXKKvG
w15h3swDFZq0eTWiZzgzhJ6a/46AXoZ5EDybKGgW6LYSUQ1H5duKUtalo1ygiJ/5hvll7+dopM8i
B00dJ1RWz98kNt8kQQ36wKy5MgXG+T5j+U+uxw83L1dimcaVV4dPjs1xMuJeT/rzRSyS2N64UrbW
0sBsYLe2yxJCH9RsSIyDDSErqgYRM0SoOnzGDvT65KyY/B/5ayAP1QBRXXs/iMj1OootrpujQQfO
XLjdu0W7ZHcUTs7R44l/5kX74pTfqBuqxvTlCIJocsao5Rjy3ltWTkXby38OvUxHf0LqthVjVE2D
31K/wqj1wjsBl1tFpZm/aHeP2N6O/cl0mfBApD2lOL+IuZob33irOzqMai2JbC16of0cdHnHTcYT
CKYz2wQKCdqGRPqzDH1wgHCtTboOW+Aoael13mWVUua/evU2r+HaKH+xsOhO0kHQGMLorMZAYRmA
mLeDTe0bPOWSfqrI7CjBnoo6wpfjeFzEMVOBDRS//daqoYBzPx2cMDQUj/CBdx56Oo+WNO4kzV3U
rQ+tOoJubPHJJ9kahpLgXXindZgiMoZhiLzoJ8zgR7/XDYAwfMw75XCTW4OpCAJwttvkl4HFbx3z
qrRa/poOx/T4mMvHOquidnQ77lBkqz7eGJsda8V1TsJgSbEG9c4vANOucSVjuwIECN6pt0xvS84F
dZHZWGouxH6f+hk3e0GhjCYs7Au+OS6iC3JMpICHj6JGL5rZ7qxP8op8+KqOpy9e/xuejmd3KykT
PkzgkSm78KhbwuQDNo0/8wxNT7g955DnMkqDgNWCZs0arm1WuriicPH0WPUBSy5vjIUr12UGP4/m
zYFbEEsMLi49CoBeXt2nfVV1EIlqNTD21FPJhcHPqrgJAc0aY4WtmYsnaCmRI1HlhYplUgHlhyQl
ykz59ECv8ta2iJzfA3NPkY55Qqv1SIoqQxXV3zedmzI2lGp6q7v4sx3Wk/gS66ssMj808Nyee9t4
JTr7pIXnr1VjywHm4WpAKirR8UPaGGPF/mT82j9Yx9+u67ejcufECYXnYR5XxMx8VSCVPD+uda33
PlJZcDnmZVO9gDUFZQftHStLUqjl4dhJzXkBU+DHnZZl3ZuHcyhs/ycEODPXMB5Hy0hBWuIY59ue
HAiAyoWMZArTm3Iu7Ds1Tk1LH4OtbnPWtSeWudTG+tbNSr+jiALX64JwN8j/DKXo1JS0YPaDsGZw
pLdetbP0OrwOKN7g2Pa10R/GQhoVLs8Ao4seUdLrkKwCQHe9U2m2gkkZI5nnyKcWwwagVGRoqKsN
I6KBkiK3U+r4SNMt9wcTSxxDAYjmH3Qe1WmrFGp15/TXsfOKq+szMPN+g94dee1NnqSqRvUF4427
W7lVNidYQLAb4w3f0ry40R9S6bsm2a5bzTrsb0e7/13JK3hexfWaE+cLJ/irKHBo1waMYLJ4vPbp
dDhyKhHTp2XSuNm9weXxIwSziuwohOlMpceER2O8obF73l4fAQZh8yMsKpgzVgcf84JEAQiO7Dvw
sjt70IJFWLmnR3hEm48A3mdSDLxeYBPgKv5d5QvE9V6j5M0zHVxVIa7rY7SO/OUk5vgHl2dYm3W6
BxRVm4BEzv80GqLPZJ+qFGCY0jof86RvgzQ5X8ciE/qcC7XLxy2584XGU3FMOl6yW+2C2MiS4SbZ
PFwkJAtGqAQzzS7mAopLGEdKMqDJ/iCwZmJLzIcA6C6me1u2OmlNYAa3gGQFIIfjg5DZXvp4LNzR
M7AaueoyjUBXcHocxRcvOdYPXHMDh1zdY+Ry1OL94J2hNOaXZ7au7LaX4mXweqmegNNXVVeLkvZe
41a/ol9hZaYH4qgOV6sHkNv6budPqu/ctfjkxK0+K7OxfIg4Jd8tK+GIBX/9bf7yXJwpTGnBGaSO
L/FT6hIqF0bceHvX+SZWSSX9AlxJssGD9iInK5gA8flIqjMVMkKQ6g5B9GgGBPHxqeX/8/99c668
8JsJCCukhbWtlJtGndRjEtkWULGj5SiEN5TGq5Pd0YXCS+WG6Ry77UMIRhIcJwo0ziwoa7Wgbnsj
1Ar/TKCMxo54mNcBZxPcF5io7OpDQ/8D+UImpXXcgA4U0uRHC9qEpWAVUHgcGfMcPt95mkg00D6y
aTMKs08uZlAuTsdShbLTyaL4yAhP1S5rcwiBCC3h0oEwqJSM/JtmJ7n/fgAO+9bmweiWjj5JphVT
CnneRTOHxMK/1s172JqTPhpYYd2uJ3twSUCTBrtkPZRtYYioG5QFjr0ZTc7sLgYYSe+ApEFfZ6l8
Mfrw7FVtdoW3o6VLI9MdxkknVoXPINT7jmPfyKNwlqbE6qVM6daQwwHKZsQmfm+RA00h3u8R61jx
x8up1KN0+xpU1QJMLLAuzRUEEkQRJjY6cGPd7NKR7VRgL+ta8aVprVFQ/XOY1AuuH0UXz7VADM8U
bF89LFqL0dZpR4y71+f5yFieufwXT0S1Oidkc8y53xdN9lEwHCvsutn9CYtD0LaknWsuVgjcm7Nd
SbmMguBFrsIDEycBxyNW+/5F7PSOjquMFrV3VXxNycHBqGR9T8w6dasJf/OEbYyUM3KixfHw68gW
yEt53L83SSX7gEubiYFkv/OlUdJ0BwBmNz18ID+gkqWPO+beDjRayEf5whFx0TpQ8EciPtoWYZiL
ZKegOvMKm93G/nBYq1fKM/IT1AEPHCgPLl5jgSrQDkfrzfqKrDdNFVPnsK38KqSiGz0HQj19crsl
b0aErOYP/EbucuQyRaXibVt8ahI6VECsXExrJvB1fbP0ZQ1DkhxDTxkb/Q2dNbp9C4yY1Tl3wpXH
fQR27DAztfCjFjz2TkCiw10AiSQG4lyegam+HMks0yZ/ok6UKj1JQdO6m3GYpbxUa95shonlocZI
KBNhsvYHpSkQU98DSln/xBkJ8k/NfhClKh2OFKnv0e9m3FKusL6orTAaNiw85uHpCWwHPCIIZhpk
qOZWdODEZEqv64dd2RdMEanFxqRBr0Sw9TeweO67CA2E8dRxpN+ZO3rZftnE1Qt1L8YKWnj1mXUu
2lmN8tr9MGiK3+5iYL01/h1nvXab84KaX05UQlmR1eGCQY+I5iOvrksbjTvttVvR3kdjS2X0VB3K
ZRYXu/eZ/6u5VtKsUIdYxzh7mw/UsBkxnRt8K7wdH/exrj57Car/NW4nAZY6e2Zpk70BbU2Wbmc1
HembJbiwYQaf2UWuXrK9kgN7fHSR65RzaK2GNJuuwOUJATyCPl2uCIN3/JrMkLyq4U0gk+q0iuC9
ETN3FxTXkROtlYPE6LLgtpam5cizoNfByEPZnIRai+geMZYbhdeL6pWgdv2vq1MX84eESC2jgNn2
8AZLCSa4FACC8SB1TnB3+14a67ggWkOu5SD+uBmMttOzw5RP5jYJP1cS3a2Z11ajlTL4S5kvLvbC
37gE8Tf25yJb2a6ihfLSKHq1Og4sIesOOGFihZd5to686E61vkkO+QwWbClHPkPf3SoLnQpJbJ/L
80cQHEkn2Xh6MtIMJxYs7flWPVxOd961K0cT7ebcISWdHIiWgH6FBEys43T5/csf+ZlNJQ2/MpGE
GYOztQt66GtH0wEGTWCPVPlzrmixhXKTkdpPw2HX6v6BvtY7rk7wfRoyfkBauF45SBlnrAGCkkjY
+UX1DHD1Qp22LyEoUeH0DzytJf3il+Z1GCllQfrV2KxNzwDqRv4sbaJIxaI9HPeKar4hGD8x596Z
SqOun3wolxWeJvHNf7pPuPgSxnQdOguFvI3zaRWrnhq8AthN4cDnhJwYfLxWdJvnuQFkGhz4w5Nk
tFflD+nfddkHWRJZyH6gHhXrlZKnkyXyR+Vf/zBOWqRI6rTldVy0LWwZDOfz7tNEN4JFdQHVcJpn
2+QkHtShBCF9oxz5o+LpQeiaqcM5/HJO/Gpe9EO48DgJ3OzihXlBw2icrbKcvYBUTsgMPSYcA69n
kq+LrU/7yTSIAyLZkroYdAddjL/twJQq8WxzrmzJ+uBDTLMLot0SrzkTdS0Xp3KlOaaZdWHAwupC
eS/KHvwL6I83B3KsnsQMzlNveKJLiSE+Nu50bEnzRvwfZAJaoFt8w9T1xv5OABTH3q7H+aawmJ52
dZO7d8gSy9q5wmElIVMfmk2XCwDKj2g+l/FItRiqZuHmKMP9ERw4mlzqTKI0dUMxn6XcqWjtrOss
2qEHrxH5DNsUJ/GLe4D6oCd+A/Oy19zoOxHMc7LcCkqrkKCd7ch9DHpJU/iEaO57/EOtpQXeMRGe
yrzR9GXgOSXfrCtPUr7rwRBxp+9lKVuJiUFoyls=
`protect end_protected
