-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
CKmNMWh2yXc3YT2H3upi/2oUdpPdkrABc7mbX1lrt1gqQ3AhbUE3az1/rL5U5ozO
sWJLHtEgvAlEVChy2ASIU5z6DmVHGL4BT3pqiUyCBrfyyvB8M+UFU31M1MBPkKjr
cQoU4v4zZMFhO3KIumotC/1Z+yvHu5aumNcFwzYB3qs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1040)
`protect data_block
i//XozFnFRPTBbfUQj5MUUKd9putJTFak3TWPr8OO7GkBu3cq90gLav5qAbipEDh
hivk+qD5gXpXvui/PR+PMJ40bF4cqMMsDpKACuDAOjBOpIbTEeLLoNTpcSzNyv54
xAC/JofMx5gx4kAlaP7u6CUocOsxx6pPr3VRTuvTLS9v5m5nWT1BFj6tbermYAel
1b7GCM0bLbuXjVaP8MtpZN/fAGOiLfgZ8rlW+JKt7x53oPnLFdILKRjmY0+GuJPh
r4OVRZnDeEmw9+bjFzmybtYX+OEfzeL6A0iYZsH2rU1OZNyZwK9unvRVuOKWUIPR
3MMWUpimc+js/9v7aYa6sxlrlDvQjvDbcyNtEj1zJhI9kGfrPZcCJEHBD1lawqtU
H8T99njAPoiGIXT5dOcLKKK8gSai8CYNk2OwUPuPXuzPQ3Cen1Q045zujzxB8pvu
53cfOApBOL/7iW0udOSBOyu3M1NTn3cqgsBBygGDIomgHu/3mvAQVSg1jAkVJ99T
WC96QWcSRQVTczp4UeH0vmhQ9lFZFHb96aZidix9oMQdQmvJBs1AwS8sH+gt7obG
E7GF4AQ/PTErw7xs0nefAltzLIlMqR+9FaqPSOqauC1ojm+758WVs/GZxN9H0xjA
UL8HA5EOJgC24zNQm7rMbDl25ClWdWs7wZzOyTJBHmj2SsbYckm7MO02judoNb4P
HohxNojyhxBBw0QAQAqKWlfIjgMkZTgE9/Xmn1Rh6ZRfDTZtJZbAFKYJd7B3XDwa
H6J4V2SQV0DzMn/53GkT2am0h9fMp+oqdkOHr7E7wauYdfpif25PhWeKqhINVI5e
PJRnjcBM55sgq/O6o11ELZEifd2QFiTvH14wnJcSFMV/leo4viiMMFnWmg2lFDag
wtMYrPk4o0KFhtMPMWC93wHBT65GdvgLx6umOBJ8aAcFQnoX2U6Q3zsQign8nqB+
BL2mvCJF+Bqsi6oG7vnrN4yKJQacRwkwYXTIZheW2QLfI3LVfZGTds2LD+W2btla
D0Je0mVb1L6oB1ANfqfpETo1ZGArqaKHvRQ875kKAwQ18Sajy0qRw0QK6RAJcpok
7uPX1Cw582xx3SyUuHV+f2E5y1hiOjCdeQiblyyxunl6WZS6yCCm1FluCSiuLYho
qrJkie7wF7ptIQH6K7f0+zlbF4zfEUI8rEoBkLYjwRwvfTRqIfurCuBOV035MXhy
E4OCmZVibkhB4In0kRXIbTOZivr2RNy9q2xAOZtmH/2P7J87IOqsitwQ9oNv3mEa
8VCK/yxZvaQ523sZfNl72ciBQanhnShg1Om9J8A/EQbc5fZpYvex054/NYdNImCd
8Xz3cHaqATghXGryZBFpJLUo2QLFw3z0QNsx7W4uA2A=
`protect end_protected
