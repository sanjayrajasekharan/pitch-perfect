-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
njBMCMx3RIOKf7gyEfs0t93/SYSUwFL9xO6fr+KiYPZ27fO3Sq9MEiQ5NxZ4yYB+
FNjSZgTJPFpUANU7fdebaWoGff1wCx3+4KU7Hi9PxsQtW3USu8NnOyYRWBiNIN+X
VT2ulE8xcGKqAzz/pfBsZ/pxDMTiBc6xex0psw+qaog=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 16507)

`protect DATA_BLOCK
33/5CkKGbpa2GAMwXgLhHCVqgZASXaqlKY00HxM1nlbZJT63/eGSq9kPGSUSerRY
1sZ2eRX2EtHmh2Q5k/Yun7rOtpqnu1alLDfuXCWXr04rR0y/L3OZenKHpRALxdMe
ZgcqT7y8PSTxnWycMdjvS8/NhHiIFQKbFxMIoAbaarUvYN6UAv3D+6rZztcKeNbB
faMrThEnmn6eFLB8ZgxPqstrMZ3RW8stXwdOWxhefCwrjYYF6hwXnUyh/i8Gi8bU
YvO+f57Yl5TtGnkv0SGCeRVrPF7yAzGLd7SYMP4tz3kV1JZ2F3GPlXb239muNfew
ZxqsbPd7fCoRYcKv+uXE+BPei5dWi0a9/duO2OgPVfXYuL7yK77K4Jox1JxI3RXJ
y3qv6XvoguAFAkwzEPRxlmxJQrBykhXsu3Kpk3wOh3fE3qzKtO+UasR3wsa3f99Z
03qg9qA1AQjHMjQVwvX5cZzv/heeBjbwc7FAfJISbwvZMvG77LbqUZBN6wKibczG
tacgz3OfZzK5dIB4hTNufgqSxei2l7gjsx3uMV1tCTFPa5D9J2QNZtFdlTBnNFpE
eHmYHafVT9N0MkN1VIWVSVznYWzU5ktxlgoQzUHL63xZAbqr0vt+OGYacsfNzlWS
+IydsFUeNoN4jVLwP1XX+5qFeKl8/WCdfQ8rvjgNax+N3pbhO/zjQ8RDjGl5lmwL
fRTniLVfCzauDXceBrRlSPHiOXjcW6afUaWf9b/HHfg/5JMvPuyaNkrMQd3rsRyI
KQKgU1x+eRDBfe06OSJ3/FJAVposXbXpokaZbdAKPwQrII+/EBCBgk9z0uKlCNCy
UANYX7RyqrthM6ER16GJPdRv4jTsAIFX0GuODhwyaQml2T0ZPgo5Rk+qdalzZPZw
JP1+Xl5uwHjxljFQIFBOxWz5422cZu5Nl4dCZWpTEQ+gLKdQVAZ43/PRz4yYd7Ya
DsN7VbsXkEmCag1PWxWnxAyNvCUtpEEI8F1Rpa/H0cxsBRbWFD5ZBmUXR8yk9X19
MhIz5iTC3hiOiuDH/hT8gooM6kvB6OG1IhIqU8GMkLIcqT4zkwb3MtklXMZPvnm8
S3D366U3ZuH1AwFY/veObF9FtE1WxzwO23gZt3pjyTJRE5yw9QIYHO5Ack0bmf0y
ZKaWYQNlMOvxNLN2+h3zINzLSkejEZydWt2loHfiSiVbJ7hHiJQ6P/qeV1I97NEq
9K1GZBd2oAFNXfND1d3cZziRYifjrclbEiLyO/rbBU7EA4zzKv15386mk9+X5FzG
6mQw4nrwrAGlH8F4ZI3qYvBg42bipBiMHCmmZ0DDpcXOfp+D5XP8UM5k7F4yD+Gw
CPB9lo6cDLd0uqiLftOuxZhO0bmCW6TEybWxpKoeLHdu0HWC3QCvcjrjZ78eSTw2
gjta44whRwrInj7ucX5JnD+eHzxMCl9lrjRKnSPwXzd5KATjXLWZT8GVUD+Nnllt
RQpiOeb34V8Ee5V8IqiJ2f1fwa+ACShdEpGQPOqblgLtRm5MBs+uCJ1BWO9d44r+
eoCGS0uM3tr7HECOuIex5ZIg8s/BojT8Ufhpy3fTEKMRcl2/fsA54uGiabjSSSXo
G0Oet4G7DCWfiDRLmU3dnTOBxSWMbPNz9DOoDPamP8aojwwHxz+2we+BDvU96D5Z
CRkY12XqN0/vYxNSo3yeUoFMqVQEM8MxmzXc9bIZhU+S6es7bZ4Ql0uEdurHMFwo
enq9psUN4fy1/kx9UPJJEFM02IJpg3SICph5JlHb7TEutqWV9AQB5JxrxlCb1AUD
Oc+/q4VQQBrPbbk6HB7p+mPs+uw3H9fC9niYnu0mQKuu96jHwFWejOz8+cIjZqKL
T4kECPfxV8lALP9QvYd9HN2e9T5ZaJBE7cQdvhxLYrG6UEWWQnD4cDFah4jF80ht
P7T8ttmi+UqgQyLMh2PGJIXZc8XEQF8aeTZYkuZCkIJ39ErPjFeKL62+HBh2wYC8
s9uCF7fhi255k/ZSV+mjKgPQ3MVaNFL2W3Ed4o0xIwmz7D6a3h/jhlxeIiIK1Ao9
feGYYY+prkLLl9kZs9UIZVwTO2uzIHEwSc/7O24HacA8+9wmUIhXD+P85WCyJqXc
OnCJxO5CMin6CR0BOwzS6wvPWcgfxzgXmdL/33bkeQyY0YY5IvMBw4mDHHuNNEyi
dWYuwlqMLWfOEyoMGZCPY0KMYoIGeGtp1nRK9AJyAlvL4QOlTcQgg0ejFyewPnpO
KBdFSBmMffKtPXXD4t6W8WA41E3ups8tRHc2s7WGEPhPjJONP3Zs5bgF38cQP7T1
HpqatgGGQObihtXCoMdUGrxDFlR6VHibfz2LVG7U/z6fYn7CvSSn8W+mAAwg/3HB
Uyxie/k7TAmjNQozUpWKcJU+rxLOP06QmTFncHeYeLP3I4l0NRMhVj5TWyD0N9Kn
sNasOZhMofU80yMdU0U5AI1JayPgX8UrPGpm2MLTT3Frt+fE/2xx4yTZS6JgLgz6
pUmkIVqXWOqO/JbDD7s3JqMjH6G4Woo1b4112/ieWRsEVbjn19L0VDeeZalf7Mow
xLCa1hTPibfJ+1ECXCuiE/obrScJ1nurO5+sHZUvZJ7wgU7POfM6n2h8nsCAzIju
3URi4AjDFCghmRrg2NeSAggebbKZIWzNOVwY2pinh2hOkFOTLlTNylqeYJWbPNke
uhNk9VTtpfspXmo4p1L3AnhHQrC4F00VkosPT/X6iTyfxYknMjNIDIyt1doRQGw8
JK0FsDuNsOHvmKBZ6sA8mo+NA2VFLu7817nnjiDyD4VDSeJ+oYlDvWfSmjX+9teZ
A6O+Y86gIf/BiP7CukCbvCMXf46b4KPGvx3hMkCDuYFHXLSGzl0taOGtO0eeDHtP
aDOyowwiXx9Qwc/C1O0bKiFAVE54KrtTPrYRGl1awo4IdFMTQr/VM+AGw7Dwv4bk
u1b+ezv2+YBFmTYmOwHlnFKXbGUBApjdJmFFeFDTTeCUW/iioXAOo1oR/WooxVb7
64QslQOUSEGL6zS/VIADUk2xodUwIDpsOkQW8wxI/5gD8AkDPQvb6YH7zyMitOoN
zQ/5j69MbNfVhv+Bn7raYSGHkF2Yjd2+wlrAZ44oJ5ppB2qCcT+pQ+85ZWrFK2P2
IKQDKbbDGPWPcbV8g7E5iktNq5QwK3YNhlmFXX7qPyggaDzgetZjVv1gy4byNBU1
yp6cLhWsfyS476woIKHj4EJAjJR14tmvIPTnIUENmLPH9qSY3RX9pttHYvp25fod
Wz+fxuIBP7E1lD4D/jzpvJlBQZKwLZ5VgmBHdmht/LHFZepNJyGSbAQeSbG6G//I
17RqVRTPZqdoSZ7p8GZZQnTsygX0MX7OIr8H4CRPGnmqqoySG1J58wbn3UsHbe6w
9dR2YTOpiqunfpU6mpvcRnMtzOgeebc48ysUFj4kri13ZZ4EohTohWVNzNCEVRyO
tfBWL/qU35vxeKeEcBomKuNcekEfyN3t3dfo10DqK4jpHUkw5KjjHFXsg0kxI+hk
t95ly4SAtjSr8tTmHAkY0ONdLluQXYBXvOn/o5ehonLUmAB+FFNIdR541taY/EUO
ww1AuS0w0ngwk0AUtQm5UKrB1oQYfGSHAKhIbTVmeyyV40P+Edrwc1gqeASlu4V9
Rsu1S+S7WVcb2VxgUtO9hSG3e+DOg9vIkMJsL8iCscJgW7lqJRkRMhEEwMPci6kf
2eK5M5dTcIMaNsiJqiUAqvShkhrPfrscCq/4sc+k9C7JKK5Mqa0PrQaRWzhYf9HV
H9uFawvn8mhGS9RFGVqnZ8EcyF33rbc/3syXk3gKsCmrTyxRYakrZxa3+xatB+8L
/+sMNNr0SXCMrRFjnTR+6DLGJwq9Op4iE0fqduYa4cf9nFUbQycMUuMNKgWl8Iag
gWSRjTBmsAcO+f5Wj/F74PWZPg6/p17+JwBKKCjkE3dVClem8LK4PCc1na/BI2o3
XFjQsUhGUlq8JyC2ZVgj+A6+fXzmvLV5JDWOJorXmNyizT5d1xbdi19HXYTQ2hxE
KG2XBigzakPrv8dJZ05zfjrdTJJfvM/HdbP+o0PFfLWNFk8FZNvwJpSQbc3ZtL5j
GiSsPVgm+q8JgU4FyfWiLr29OpDPn8uGmRWvXRfIj4CZy56WREkgOvNF7mKzfT7+
0bAcjIePX1KNf7PQaFZIPLzDYhvaCv9YqmWckHSO+RES27g5p1e90G7af91If+Pj
RR8oEcquFRGZ0PXCRP1ry/flhcROUb2VlEO/N/nFXgxeKOdDiDed3K7QS39rd0/z
GPNfQ8be4Vkr209sMM2W8NJDO0U1WIJXim2bvw+goh8z7/5/G9FpSQzTqH6Mz/oD
19nqnBi4zmFYwckdBUoF72QvGnorjdpod64ZtEw1KWkNrkpM51HnNYtMVp+OD2Ee
gUI9IcUo1V2FEZUu5SnjT2MHQ0/Og9H6iTsqPMt1e4+jwtwmsq/yKzkkzXaqqyej
z9NTyGtSXuP2qF3ARwxTDdw/MY1yrl7vYKhsJjYmtxm2WTCaTG3Bt0afABWbHSWU
t9Qski5rC3vE4kLKbqA13cX12mHTmpeqk46D66nWHYVoqNlRgMifLOrHBbXNucMv
96/k0BbKX52M5sUfTw26VBm5FkL3N59vQKKuMa63zkEirQJZC8Zv9Z9japnm7ojI
67AypIvqBiTNI6tYU5pvD9KsnT+r+PA0b4gE6HrQQdGm94Bclx9Cfl51lXrOyPdB
YRQRkNje5G6Qd67sx7UOIwOGXZRoW/6F6ch0oYqvsoIloXhbRNixoMj2OtAb3HCQ
D3SVFRMcKoMEI7NGqXIh036OIEdcR1Ny6z2fjRMdgzZL8sb8f8Dkh7+9xuvYRc6W
SNqU6Hr09BJ0WI/mq/imAZ1kJqpEqJVVi6ZLETCaM9q58QN4AIZU4JEgb750gPjB
9L9a/piPw4uCzdIT8d+sYvSkRXF1aRETDncN2jik6zbyCbsUGs5mC/zZR/7u4Tug
NblnFetJz4QdH6Xb2+ivPtg41TrfDm6k2MxT9KVblD7+acqJmssMkCRZ0ipd0XIh
0a3oRVYjrhYcqIiDjJmAbVkUcVEesMw5U30ADsOMM+OdiDOQAUeDQExlW4tMQ7XF
4kuw26QW0H/OtrQWCqhNfJ9a3zAODi76ZzoYt4WFpUpKmA+gdgyio1gmem65E1Xr
vJ+OYh/HjoNV1uihiHO2pcCjBEcbV7doXt2FXuuc9i2smpWwFm0F0uwgd5I4bq/W
Q50zOs1GYV/1YFcbEJ0t3ZoSBay+ABbE5DQuHWUwLrB86HIhwhhq7ICScMK/jurB
ua5N505Dym9nzejnRxDjdMzTPS19JynheBFU/Yb0zRRP0visaflXA6t0nbOi86Ei
Bm20Yj3luty/CBdsEWziMcCHLNjMjPcWYNj0nm08nWNgIOtrc8bAMKD3+4LngwJd
QQyGmL47zO138Kco/9Yu8L6aLUBW72DkRZd8sJQcAlxZDBYqDlSnrjGg1g8CK0JC
dpJjpCRHofdUWJVED8CdQuO7UFxzyw97lzsPsIO+ycFRuMwu1qTFhpqou92QXyDV
FNf5c37hYNoImEjwegJT/4PIpGt+uxEkO9gUbb6vohcqOazPNveTQjo6UqwRmfcB
Grc0B9cgtbXIwECgLGEKf6BT8OjwbX8yttvd/pFK57QJL/lT3mBHO2PAgs257blQ
Z6tCovKemU9hWubjZ26fcagbR7448YhpgAR1wUYGZy89cmy8x77XMUaP0ztGgDcq
50wqsGIFi+S2lIqkJtOeCB21hHKK9U63WYw9bJv9cbCh9XPe9VRjjKjyLhuxpo32
TEDgq9ul97yHLpd/mhElwnaBWF/EQRyvtUAhMwa841naZ/UtRr5Kmxh/BnJoIOrh
p9IR5Rmwkkml1MCLFv7jpMbZNefRuuASOXFr7P0pSBO++JiyAtq6gUozapVsp0r0
1sZN2VB7h2rpfSFQGRNCyvBZmpNQhlfigxrkxPT+lwXVP5ju/ocqjYSI3YCvwvCp
MX/YTqIiRLF6j6r5Hq//Wum2DoImQHjCvYR/yI+m43Q2f2RmoWQePVal5rS9iRMZ
1H2hZhtBAq6EZK/Y6aO197PFJfYq6vNoxk0ML2TLtP09ydt5IrHI0dWkCil8aq1x
fq2PuFi9WGWL/PIZqJF1kWHvyDHL1GtD+yvWcKfopWthsSty2cILRaVWe9GuLW01
jKZkFGoiYxDKlpTchiOl2XmEkjyteMdQaTiJ06x8JMN/4/oVMdPQfX7al9F3v3Y5
UIKvYrd6tMoo9hLCBSZaJPMwkCa0G2xOHSVfYbrm5y1YtnBBo8EYeKkFsBBlOlou
bnobbJx3e1duyHipsP/xIuI9ZXfPNZrFT1bo4d+8nA99E5zMbiE14wjwCpMFUXPK
84OtZltIMZkGM4ZLjtubxKE8NgL7g2wj81XBrBUZyswL0oo27AqWCkCQ2RD0VH1J
TtTgKGVNNukOLlfL7Jt6OGjTXi1qPPqp5aF37Mkbwoc00fFm1jxQ4tJWSNPuzOUh
1WBx3WXy5vWNZZNjZEYBrDFOc89kSje7pHxiNEU1tM010F+2c/9bQEPrtUNNrbrj
gwOAPYZTfexLvrj6+XtRCvfJ6UqWtFGyTpFkEVYxRaAOY/HAyA6NMydv0fFNjcGE
9RsjwZ7MUkmELdNX3IKebVUDwk6lc9C2/NdQ19mGMhJgOrYokg1+BVak55Iqe5oc
oKRuv+pix+huiXYogbeXgoPsAae3hZ60BVr7pgvvO0aNotwETdziYtPIELyRDZle
uth5ACx9lByBPRJJoU0fD2WEF6Aa8mIDGIcSCn4Ei6pD+SO1Oisw0O6KPNHANWaV
Pu5qrQRcUTlE7R0Z/UeYUVCuoGWujr/S9BPHT9ek8TS7m6qqvbykK8RJR2c0B0bX
nxy4Y92eZQSf6WJyQRxLJ9EAECjpcUZGVlYsV7n950quY8QqruAsgV74dlP93Ud0
EegB2nVc5edfCPucrHvDwt41NHo9IB7HI6+JSa3Bb6YGH0e6ldXTzwESKxrUWTql
4xIG758sBVBLs+DC/SS2KZa2E5ZtJJVg5XYPdNetdLt3SWqMxOggLriH1zRi2B4I
vBGKYSGJarBNI6j6AvAOQR1Kkg6RqiU6x0c0zQm4hOcnpPrFsG4uyosO9HEJXtcf
GrC0r48zi4mS+omoSHOtc9PvBQ5P8P58KLkYvvOoPhka9GKr0vHTfzZJyKOEo0l1
VFMX7VP9vevuI/8jgYCqjAjtZ2d5cWlfJ2xAWm272Hd4b6I3W6EDq0IQtpxMipX/
U9cB/iCJkoB/X2BwLkkbXuhRrEZmFUBr971YzpFjRn30LXHFgMLIpwXQ0EknWlgx
YDkS8EEfT2EqH4lzyp5pb7/GblbzFN7dUKj0bAPjM6fxPZmix0kCO3pnH0+WNREt
l8KBBLURsbFX0GXk7OyRK+Gh3a/7JHJMX1TUR/94zbQm+UF5eHpLNZ3oHzFYEh0U
Wev6yXoSFj75PH3rbGYrnj2+KOr4SC2v7RWxcXItVNxW2cjwtwxNgfa6d0O88kOn
Mi0fc65dBs0Ugw8GWdX/rIdW/HnNhIjL1Cmrhb9J69DyJQ33EbVHmuDGQSUYsOzs
RuY2WjjcaL5oznD0Qe8hiU7deb2nxxAHGSWUm+GtuZxILc9fY0fRu8xKzD7sntee
C5Zvx6htIil2D9kQkkUI8wmpwvr8gLTxMMBtWDdY6bfK8ajrj4jhFIcvd4YeNQDs
NkusTcqjCu4oIPekQqt90eKs19Fizt8/YXHRpj2qkmHZMwxqeYzNzdRkrf3WNhtn
tCaQZIGG/HRIrCWnEiCWLrlqOtXKf+HcK1jyt41FU/lWamSqJUR18jsZUuEcsg81
7LWGt1mDgm3NlSgzpqnlGqWBpY1gsFcgDTqPwsgOmLAKh3e1GILnMyXl66TkxwOV
3dzraGk3H3FTOtmkFtr5WwQMjGjKb+QXqMst9o/urW+uUTsmomXMnfN/oRchI/Uo
QRpKVzLSVjnqq5v8MU9pgtrPjJu0wV+VVcjXl4PTzvMVoheB2bNiZ39A8e5dTe6W
lXD1yyzST9wl4mcLXkvGfZKxgez+Xf7PFJ2HWWJ0IoFbemToU0hAMeV/CdItufGL
f+hnNRisgaG2EoxzBhtuNq0dlMr6OlDMtldWbhNSnsjmC4zXuFNkOhnSOS+dUPIM
kHQhc6O9M/u2skzAkzIUmHAlofXaZ3jwvLfuLbzhlR8qmMa5xaWQseaphloKcnai
OjZc2Kbnt7u2A8TFx326nyif6vw5wS8N3rgnbvmD67zUhp8MKkWkA6ehEPRMcArD
IQITnO85gFZi/AbZKGx9yWkLwV/FiU6iSOsQD07vuHdEEprFZKOyTGBghCSDWAf/
HSn44phbuXKF3+ymTysu99cS1uP0MAhwl2iAyH5O9EISWl60TcF7l6rA1iDX2taN
I8Lzuqyl3OXl6B9aPhY9Kss3/THn2Ajkv/FeqrRM6+rYFojZpIQLvFYzyyq50VxL
t5JQGcQL6SiuFM/2VVA/sxHLvtEnmxe1IK4wPN+QqzoXDraX2zQPoTCfLIAet+Zr
moEaK2luHfXqw2YfsTCXjoG3hSb2pkmGukmPjC32R4uVX1bjML1tuWD+4Y1234gk
qf94bJhMT/Qa33vyfJ0mxYJGMrq+p9IukvncuOEm//hThv37slFEtHwLkls8MIw9
8LufmulNe+zTjGG/l1NV5OkVC2cpa+HYdvUjCo2O/uUu4808UXDt0cWQ+OcHkJwu
pFwtbuTBjt7b024cjnJoSXW972y0/HiOrcfzPOHnQEXRZp/G7b7wxJ71bTa2l2em
0m9JMGCvxM4rKK2spMtpZyYX17FmP/REGlKGiPCbyPVGJipI6FWxuevTW4MOC/mZ
xgRpoOBURBTnmj/DRrDK65CCmKAWlEazJqKlE1/6iGGB0Re9z0JewLAwvhbRlLyf
EcNAr+MYvqqVUhCv9revAMbzOGyeUSIx1QGCOUIDIswfEevHZyZLPwLgqiODqjKD
e2W196jORkj9/qUasOCVXRbPRGvHHydD7NkOubDfkM9amYs8tw6lpBTojpd/wUoA
TNlvuET9yGwCu+WCQwraFnxR06GK/9qOIy4waJspoSt1a2qMe7tSBEVS+gXoh5WM
7dlSLKjiHwjkZZMwTZ0mlXgHq18Kjm/jG3n7BduIjoEHHfyniKXBkNpYYrNEN1Ei
NmM5YwrIzypKWek8zrSp2+QMPtJwE7sOzLTIK+fzBHyW9nTjpr9+GgjCRvnffwMK
u05giZVPQC6UYOaxSRy+SisCnDFFxvUTFJ6CYLVqseuM42NyPLfMP4FZ7qg1vXUE
THco7dL05IiiGeitSJTZgrw0sd6NaLpSJ4k0ha6X+aVhq7reH2pz0R3mYUANegk/
mOdFciG3Ps+1L/10qo5WeBXtlTdz81AtMtRBTmRd5k/DHiDd8ThyV19MdpoXDSEO
DigWc8yf5HdlQUQjba13BaxXqMHB6iBrHORyLlHuF7/m9PU4fSyRfUOAy7x/DXLJ
WTBeF8l21QPmlb/nw/B1WZ1ujU5kes4gwCCk3avhpBC1e6pjrhqrSA7RkJtpnYfV
kc0jfmouOB2MswTPKpF441wBQHEzsZyTT0tJTxQRRgen8kD6yaE5Od2mqpQeU31o
FHlXKXhbwuBYQZqMfu66OjfgdVL9cOTMvgC08lDCU+nJFYoBUF1iJvLNY6uGL+Q7
uwrxkZFemIUdC3sWH96qy6tJ0zQ720e/2aEpXFRfNeYz2UsApGRJniKkl7CWF1Ej
AMj61kT5+nnNEFWqbDiQanpttVY3MSUy88XQunVqVCQEnS/1XPagIA/SqFgQ5UVH
6MNEqfnAesy8FSr+9BN/a54yFk4tI5ghu8VJ7nSnz/eLkiiEYYuSsrzgSy17yFUH
VZrhXHO4oreznjSOmb1k/GwmSSRiLwe7D3UiRbi/CnvioMrPQVAi/LBCAKcfTsJO
ku57sVaQlhzDXsjRd9z6LWa8tAbcF+4DeGrrjBY+TmPr74kkIln3WplrQNHAtGPi
QzTRXeq+JF20oBiRF6n7jUykpXlrfP1RFQcMFJRCe9YgXH354kK61bI9a4ZoBLq5
M2GXh0+YnBfY4dOXu0fHOsjRbFD4k0ti4bwgepFUmUxmc5BP3XfV5BozKSFrGiot
8h598GW9KxcY8DPRs0SvR0qn1KOxjH3JPilz33OUly+jw86XcSVl71nVgwgqNzc2
qkI2kpIiSYBIR8TyByWH0wST6f7jNoFtreNn32e+pWgkYiRJDncRRCrkm2JWZ7Mr
whk/FWCdECPG58KkVelyNHZpTLiQt/ENJbOab9CSx2Cq+N9wCBFexb//wKb8Eyct
P6TQCYSSu3diuwUuS6MNQqXC/uZTT+FsVKDrTv/OuUo1LSvLE9EFc60oDzRFiZte
nqBUWcfjtegug5gdoFSqqjWhnVtp/g7CvMrPGvIS6KGTDsyNXiSiI7A1z0c3A2i7
B8BA5DVAL8vNOTUNQCZtfwkn3RzN47WIQ0G+Nw2IstnBlPzthTybR6J5L7IOwfLu
vdbC/0xT2y7Nrj10MXkKI5KXy0KEx6qj4wdldcgPrg/QtIzcEnJ2c8Av708wOC/2
x8uhGNVQt4RDBP9FVahJBMMD/h/Ybj8qi9wRmHAbXXpTkbzxFCm0rddhGcRsU03i
tnq3+FSNzVbn3smSkvdd8Ld8qj+da1GCmSug+BYeDtYE4isWAvbeV3FxHLrlJQu3
MO42+xYwK+nciB35P/idyoJ2POQFGBhxQ0P+TzMEZ/Xi2miT/+AyNXxnAkJHYde1
BijbcnMY54YMVP4T9ksh/80Thvtm4tWHtCPinfnwFMdT/9vUhKYm+5+yUwX3DE5A
8Q14lJayJTG207qvvQO2zqtYKAjqMU0r80AXETqa9qUD9AdWLoNyG8NYGgBAddov
AAxWFN6FxGRGWZbg4BOsYlKf5UVQe7ITfP/o1A9+e//MqrYCxCu2/zaJHL/VCBV3
G1ESFG+iXqsugCDLxlX/ni8U+Y/dnfoOB3+V43tI6QIWfAz4TLLE9/e2SuH8CVBf
PRLP0L/DRuzAzHK6zPxhWrCkXJZV7YJ38YQAXBKuKwAR7n7k5JgsWn7606Ev1FUa
svXqo72DuE/F0HwnIvfV1pyuVGqH09lK11sFoXRNN706scMfPhqxRGzUZ1ng4fEO
QEVnBucyiv1pJU1a6R9dNDIFst30tCdEsQ3xHEh2uUXC6SPV8kIO9P5XCi5nUDZa
2wav4I+rVDTDaYn1jBhlRx/XlfYpSn/3RHpoMzIqLzI8UgfVEhIzC1Nh4VZkiTLN
/l+9eJ58Yd2Yl2IAxb1S+Dbjv3qhPBLh+4AclX/9dBttABJUNxjXfzE73Sk3fS4V
Re6Ln1JSVc/n3IzHAro/h7o0KIR5+dhtP/R6sbDDJjITJc5zFwkPbPro54XwbR6t
l/bzNh0vDBkzCAca0/2WuvoigyrsaAItLFZRmJOuXklvFUNoLb6Fp7DbyixGHaBA
SZrwCVFJcEA75vk/p83uVgYttISziS2YnXQCXl1Scd6jJT6KEuWLRDK4ZnTC4/iH
exoOEg8HTqqK+zHjn8GlVcjfIs+5hCu8VMEdpjZz3PFliWK5qvxivRI+LeRhSH9H
bAFHKj2QqFRbo7A4FVGuhPQ3rfi8Pl/9hebTXU4M7wNe/328kw5I0wIuiCeUQifd
GjNGTUjYiQ7CnV3dS6Q5vc8PjpHcJC52MvWU6S3yaLhFhBKMaUC0NAFVSn+rrFzz
zk/eA5wHv5gQcnv7jifwsPuZU9zBiyuM1WIPVmsN9I27DojpzogIlczQsg+xYiHJ
SGIkdYSWGt/6OFHqJIhKlTIhze5/q8X5IGG1yjXHxIDO1CXo4pRf1hy+4VmNVY/F
kGNEvjDSPhAWEMfmrv9mu6vOeQE9DU35ZdmBCv/44ivusLzta8dSJ6vh9aco7aCo
22BCdrY4+XntMXLhtFdSGmxfPepGWvJTwZ9VOLccLeXYXFNQshoaXPWVptupTisH
5QpAyZ2sX88ZHeVcJXNuRdkQw+qABoO4zcOXWpcsBlkKI5wQ/FgJLWXeKeK53osR
raN5InNcb0ZrIKKBxcqwghIJKXWWEGsQ/b8ykmwPbnTYi4UbpVT/hZRBzvnsTFC7
wmfd1/SQ3S63dNqH4OucPr0qFOqknZD/5chUxZtj0vW+SOO2EiZi/8zzj0UrqA6H
U2m+0z0ovasjqtDyxDFnI3VuUxOjb+X0RTyE2Wx9I2GlTcC1WSfiui8LTHyipxsl
5jqOEOZ8/eHrHFd2sbH784Gt78o5OdV45gEXq8QD4CTfHL12N/5ZZP3U8XcHMrHj
oadmfhiVH3OmjCmg6kOBFKvpsW/7FFg3dSmxLECB6tQmwQMGNzY4iSaNfyuylfLP
CD7oQ+5BLIyTuG2riOQvoKdOmR8N7ZkF+KYnnr5FuaVu+fCND10Z2KIi7pJGAKmg
XVrMz9plLZ8PXpi1wdH+noeWM0NUsh4BUGDcqzItA42l5OJDpbiBcNU1SlcUzhEQ
hXOaIAu3oOYusgF0OAs2c9cV5S0C5BrdzhtoyVqS4lGQN/R96PSuTF59kptJ+RIT
lE5Eb5iId3ET+qUcYUEyMPzcXvQCOueSN03+4XSaIAmP2xqNBVmuJSRk6SbUkJge
9VlTZ6jKFdp6kqsmASJzm6D/wPH0H0cWnWXIx+UoIzIEnFomekdrpnHmk6qDhSPE
AH5Pi2izADl7XOFXcfexrlCRdN8Clk9cUJRadK8XcEYpqf6Oe+37MlLD1x0Q2YKM
w2idQNjTOkR09n6PRhnzue+bFF1M5eMY2k6o27MJ3Ow1xAPXae+Y+KCIYyowbrGW
57iCPIw4xi5Ow4mnp3ArdmtjCKbnODyRwiK/lr6c/3TYLO7jzu1vVNUC+x3cjFsb
NSn3d61MGWUkRatAG/Jz8MLsaEL/NxGQWZG/Ypg4NeDSF0ihJV/pAzKCXzvetbHK
vepd0Ar5cUTEQhVdT1umwjxBnGMiEyo1tjzwIFRqnx0ja860uOqMHegid/do/N12
8zu+ZiVEE2euBJ/7Fo9qnn2p3dGyY1tMLXy/o4F+exBuhNobYKF0+JYv/8h5G71G
2f9xWMFMcjQI0gAk22VgL0Shkk09FdHq/VYUxfZF1L3y0PnPzdfcxNkrp7Y5X6OK
WhbmF4V+szr6c5yN8JiGQ7l1m2SaMCRjx5rnt71o3QDvUXTrMekyALI65SMfQZhm
oLQeZI/S6YzcV4AxsT3jDWo5Im/MaXcYIxAXjf/34nRun8kf6cU3q8q598t5+L9J
AORV2BdNlbZIPSSYRBqJ5189TpsE49zMi291R5s0MzoCGA5JjB+Xc0NL0Rxa4u2r
0HCbjwBpAKyysNQZCO33v5kOrKCOyk8hC+zU/wDvhQptDLJOqCosmppfim/tVmU3
Xyp4oR3wKI6JSotvFndbLZbPKjYbg57LMUwzjcI4Cp5dW10acK2jzVwgTChNeJDY
NbQ/0RAk+cu1TWEhDDyW3fNlx2/huR6/EHa+CyVOFHdXYpvOdpLrXtrQhIUrETxv
zdq5YHqckU//c+Fy0o0m8Y3lTi7rRe5PQhFD4Df+ruJjfB4OIOzCaJKMVEEerAZh
LmZqDApLJCr6EE9TIVbPN9WQlmqYp2/ssK5NUl2tpSi4EK/0fxPGyXSCULWyLDro
Gp03B50q3Fzb+v0mzZq41gd/oXFeK1JahWSfflOLWWI4t495J8PHDsjOGz7di1kY
yjw68aU72QxdyACyv3AgC05sgdmGXxi8e83EpIJkClKZT9Xx+XEp75/EjcHTzRY2
byKNJM2MjWAOysZCspsFKW/xJorswCg8sXi1WPgcI6iW8EP8OOYP6Ox5usiRDJX/
7rixtj4I9Zz7y/zb1llBH2Lmp5ZINh3etEQTFR6PixzBaWKG1wnFhgppogNjZhY4
F8owfk0A1Zt+ne5zZfuBotFit2X9fwW7FFJtYiXOHWaG5u4AUnDThIq+IoT4vTfO
1nGh8rIRiyR0qbx1iKp7yP0KEUWDis5kOgOO7dB3OBwtkEPyYG1ANoOWxSgf+xHz
tgtWwvaKt+re9TYnA6pKeplg2KxaU5GAjRBopynuVEhhDzxzKvSlL9WEUztPY/Oi
7E+grxvARnmll+jWE25r/MuKc5JvLrSOqb8rHZq9itEF9SW45XLBSXyNkw9IOb/O
cN9IFFLBxhabuR/JrpKfZF31HwKTII+rKdVNeU84n8u1RxAr2VRxCjCnazWgComt
lMaV8s+O+xtWaDiemszb2gXzRXEpHY5SCT+9un5SM0unmepoKUVj5t04REveXUeH
FjF4sWJTKbXfKUT/GHhZ1LkOQD9qwe8rJz5TBfoATVJzOhqKdq+46SzjYg/YIa4M
3GKIMG3ZmLtA/yOlW7FUE3fpeh6NSIXY8WCgEIpG+BNYU+7g1tyrxnA9LSdPw5lg
nZplG6EEczfA4fG7hDEa3eAymiZcxVrHlu1T6yVqEl0iMLK6qqg6DLNrnAqRKsN+
Ss1+bTeHUf6DuRscsvqWG/mkB0YsilemPO9Ab1efdJ4ky/7ebi0ou4xnH2eEygcr
3IdH/7UL8pv8fA3gj/vNaTECEiN/SIfk6OLOlU+i6976FNDbrd93zkzchTLeesLM
0TLy2kFNfRlYWnpeDypK9EgQ37gHR/FVyc/Q0HgE8Umwl9LQE7W+MyUIne4deiCK
M4/U2MC25WjnPiJvK5If6L2i6BfTIadRqbGYaLcaVEGsva9y863JO+/GguBkw5f+
5lrLflzlW8At1FJ3OENcq0golNonMrBzFUWWIoqeeTLBPvHnE0Yw8PRahnnz6kTs
z3nlzv6V5PzRhc3DlBNkDjw/742iY/6e6Pxwdhs42DDT38RCTtqC7tHlMVhG0DGQ
Tl2AZsyQyPniC9+dx3/Vd0wzwP4p8Z0yYCiL19SrI3MwuxK9eDVTd1XTz/Axptwo
IJaQXkr17MbKrFViNsPZ3ko3ztAgJem32s3c5P4GE1SeudOAA/Xe/KYXyAPJvRwt
wQM9aWsIVwyA0dy4YvAIWJBAmq66YeK4RsgnQjEnLXCrOWC6hMLXvBWXJJev6xUL
tajrd//3OQbIN/humYosEgqrMeEoi5dukkqC7k2bAFYHjj0PzGjYi8oOtI8ndhZe
El9M0zn8b0WBVK28YX1Lwm+D1TQFYa1j19a9NpjwQ4mhnWL5OK23hYjmf3VXi+un
KCt011Qg59sojy/1DeDSR/Sr+UQ0Sb9y+tTIlKO8MhUJFlO/fjgTHfKF7fheSk9B
W0axCTkGwnwmHcMYYXHDC2/BaXLv+y8DcwAZyYF8QGmPDf2WJ0LFyqGME8RrfLIF
RdtzXuPE7qaP3CDpTXgKBowQ6ZyTyRQ7/Qbn18tKMjmduPYr79CaLIdAl9OqAH2Z
ER0nF0uViupLHYQhki06wXXAg9RJJPeJv1ZjFjuWMROhkZxz8BQ17yvSv+d3VOvb
pxuz30VqcYLpnQWE5r53G6PC9jahSor4TEVVy583wVMcI7tpXL2kvIdk086eo20W
dLrJr2r+lSxxGFvadJ+pRb0fZbpcC6K9IkdidWSuM8RguyLEAdlbK4nPvQvJYUmw
rldcbWG90q3zcTNdAYlTwDJmM4SrZh5JsYKomNtfvWT4ny9xLFet82NVQ8+ymxuD
0v27FF5Ie9CX6DaLlEzkGrBTeVdn/OLnfgk9MMoPoB39yojXxDtGfZHcFq+9RiBv
aTmQrrTYnrTyZ7nsUE5a4eVWmlkYbZnYh1Ijy0asvNzLwD64EafFwnXmdhHA6Q/J
jW7SxAnIFHckN4MTFEiAwxM9KdqDLIZGTmbMtlG5Y/kOLamTAiBNgsYTSfa9Qab9
4AwiiPLtaIlBKUkdUkyH7VGmQuAxGeXLRfPZUCfFUPRHh2rptEBp7at0WAvmoeZr
lQ3rOBz+eKTACR2p91k15hscSVYKWMrr6RmY54zhf8gSwDWW/Fd7wMMkYYGQbKX+
yFkYt/Zyua1qLjgOeJHp9o5N4LRfGtMryWKvTEOOhtYKP+wfx/tiwIn3osYTpFix
SnnI/i5mHNX68A5Gy1XMJW1pkZhyVwHPRtXQFX9qWnhcGaRXKUWTCMz/zOWyUvgN
mT/F7xt/gskANcfKehHnDKIQTqzHnIuwEMjEsLF7QCSCyhovdeK9sJ/OHZlbLHXe
nsZ/oYAXScVpUEBbbceyco2iiyUiPQRMjeyCXSfYjCQLEtpErteNozz53avrvqKP
CRWB47zIOnpAGVe7eHWlN8wtPNtYx2hVPmBAV/yNOOW/H9suNrs2dAQbAmZ4Db0p
pAU5NzThLeWFwB1lhFEIB5e4VdcvVHhT6gnxRGFLQHOatUxEskTNwhx8IJxa9dlq
GCXVnA/O/u6hM5wnV8iW/E/djjQim6FhYZTcK0pntfwhsCm7zMkxN4MigDcvMSR8
GfbqMoA7EJ8zn8IwdkCz9v57e7DT9Ut3xtZPm/Th75TmRqFajCYHND2qpwybeg9q
c5Tj1humVCv/afIWV+47gUeYBNwYA1ZpDeHUoT45lkFisQRs0CrFjHuaJUMQI/2H
Xp7jXxockVfOrA7PasX2eQq4p5mRqNj4Ik0l1+ae7FR4Dp86z8nRjzYMTH/HTeED
W+qv6QtGWQymCQ2GBE+Ui3fcfm+8I0zKHWyqhdKEZxlt29HwuIdk+OMZyvrcdTJj
2pjqVGdjmVS9lVR0YTkRHPRkfWU3jH1xc9g11ghHInVuGDXGUYFfWDwpgNGIy1hj
yN6asQmpbUDInMsoz9Fce0NwFbsaDMR/qfu0UKee0/o71Y+O3urW5X9mSu6cQnIo
ASwjql2DwxrBu9slEOoVE+JQVMogBzVxBJW39K/Lu5VhiVzXXj6iRahKqUxhWJ5e
B73MXHF0iaYfxyWK+4No+tcQyF8u9BDbrU52R/+OlhrMAeEUE+1f+vGzHv5RQVR7
IAupkF2eqfsKf0lbKJmQjsaWhKgryCJQxmnsu/UuE9mIbCPP1TAukPPHzjYEMFZj
aAJB+zqHt816jeCpot6w5ygDHVCHkSGD8jUAqlZmmCVRjljLR9tCraME0l/lLY9T
LOJTaDwRmBdVzyEwPN6oHsDhH1L0CzNjyhsyjPH+xSxvJ85Ko1v3Qc5bIpiiMfVf
6On/Z3K9UYzHCDvtO06rUey+f+HO8OpSbNtlzJO7attxAVSQBTItVnTrKEFnZ9GW
MhI1RDjJl9QYASipjkQLzWaC0HtlXMgSfj4j26mYXvqb+hH4fr3b1sezzUrb7Mk3
eyjCil+os5AbWJxp/FqVn7+KyU4nkVoQVwROznmdf+25Rh7Q/WROIc5OxSi9uXQR
6VaUxL4aJVtAyR20GX4dkSX6aY56aphmLvSnnJwfrgaKoh8MI9ZDYYQsFtOGYlPY
PIDXHHQITtlAt6MGPbtr3XamefUFDzMUxmVrHE4S3hGFlaUdazwtLI+/4L9iD7kA
/xYmDA1Au9O0qrrDvCazp13OvhqQgyuBTnwQCwHxqH9B1Qmi85xKtw0bOhZwwC+W
UlsAhQ0PtMBMSMU2/gQMkEhnVbNs1YaAFw7KqIyi0jrLsFVr+N6jOh1tBc7Xwh9v
CIReE8/5aMsnYsOdQZNTWUFfV1yRwjLYRd6Zg3pdYzMC4Jw5kGNo2zcKHrszMymV
Qto50SadJ9dGRxXnD2K0Y/BLIG0IhXLmzTmO/WHHZrqlEDKqObl/UhoerGHjGCqd
FtHsO6phNCCg9B/MRNsLsta2iW1kM5e4JCjnxIcSDH649LACuupBFdqQ06gO0RzL
+JDw2ClHvNIyOXnPqHXofUl58ZE32ej19xUXve9ncQDItDoy5Bf8jczA3NB8LtH4
cxInwH7J+9CUuZ1I2L/ltd72kpfkQ2VVlVxlTeDepQg6JcOBceQ+8ewOse/6gz1v
o9or21+vhvukSKZYaB3+NqPhfzjXGqvYnrsyIr83KP563J6tpa2KZaKDXgcdINa8
fCheXM2v8EkjXZwOgkSpvbQhuWvLxHZ/uircxzf2xcKVEhHXy1Lc0xmHb5cygdE9
T5VyTxRBSQXNsC6dooBAcbCFte/CyigccEgZyYNRXvUqJTUFqDyCXuIgIGnAc5P1
KLkKMLnxFjv68VNXcl9gt20kBAv2CdO2hK3ttA2l6YNymsYrDw7RxiFhX+pb3Y1X
hkdX/wPgql1lX5u7wuowPM46Uo6DVnshg51zfsQq7djr84w7hL5MKKsNF7IpPSBQ
XSms2AYJqzN+LAaAZBthCEbYv1TpXryz3nseugpn7zWNn5UvzH9oZn7Qtb0X1tHm
JuvvgXGXwqG3T9vJ81Tdkj2HgYTgs16e+4WZ/SeZvwfGVn5xvbPWXpe5bAW0q2Y0
TgAXTgr3H5lEob5EuJWM+7KPcGLHrTn+Eundqj0R8mBqDPj0pYLEVG9f3zHj9JCY
wRG5dETUI2EP95zV+Hs6HjlguQrUWNr2mRYjovUXIcy2BgMjOIT9/AMyAq2eNF9e
NzSe7pc3U7Bbk6c9ee5/YXnG75V6t1AKGSTYacR3krgybrRJhmecSqohneyUn4BB
qbcBM/8ZjV02inDhe4m4Ihhfcu6RRiUsh+QMxdEK8FWS0ipYUudNCv9rPcqjqAoD
CsbLx9mT3Slem5UPiWjSRS7M0epFnKh2QaT4ocPTeoY4cEsnvgMleA0biRo8+6qp
0a+eOL4KSCCfabTeEdxU95FYMMF7SOQeAkBiGDAXo82cPPSSuWZGkjREDOoa6r3x
h0cBeQkaiooWOnW8mBzl7yM9891u3AL/dda0FST/ajqRwbvTXZW1kYms2EJftfci
pi+upx14YxHKxBRRboClwZ90YUdWW560Z/NV4zf3ZrKjXk70BJ1ACCkpCy+x5+pX
8iHLxx9ngSLh2lIwtI374PZcur1vrWwjMN3volckNb49CqO1x8EpO8pwzYLorIn/
6cZJ0jFZrjw/CvrVxDr3Ghg85A+MaeM4hrpj9c4DXayoU7KT84FLS1cCzmO0bJYk
oQU5hfGxoOu5NyT2o1kEDp9iKN9xf/ePLza5+D0fjfoxd+chT8sKwIv8cwkhSMAs
SgIn+rJNX9ZXCf4w17qlJC5OsvM64/HKOkoMbdWC6atIjDRzV6xJW77m+R6EvBdr
GAZz9UBWiNlTJ3vd+e05O0XR2q56yNins0tIzgBK1ktImHMjwDu7DHm+eooXhnLH
+L0kZd7ZXwbda3hKD5o2fBUg1mipPK7Fsw6Vfq3QcmnJh1KZ/ahA7s+dCNNl8ZTQ
gyoTx8ZMeaK/U22haB00L7bMLEtKndqmbKmNB/13AFPq8NCMFN7+WKO/IlNQ57TY
whCunpM+AyhUhuiVEU3Aye+uCZOSvtmEaCcJFG+4tQfjLrdk3zx0aDNx9CDP9B4o
I6pDFA/JD6CA/tKvDFdS7FMVeuR6/ISddcsAqu7uCt5MYNym6vd2Q8yNh9xOVdSC
5+W63OD5c5LAi6LgY3Q/sVqU/1ZdTQxJgxm3dX8G3kAteVLsLWCqVzJ9xbwHLf0Y
FF1S2rTHfycoclcqOfKZ8VkiSRDUNa3ZKwi4Q6Cqwflde+tktQ0uUBiAjWIfeJc5
08Ml31vj0ZDbzjpUmxyjzF2uA4+38Won0SIiCkU/Cj9hMLHbSE97MtEBKwc9RtsP
NYMzwyjX/g/2HAplrSCSeoVgUXX6e9Tg7srkot/PJSXIRN4PTnC28kP9hdXdPRPm
d/YBls8OdtMQ3N4fXClSUSZBcexyzwI1EtToDcl2FUGVdP5nviLtozv0I65ZkcFV
L0VzyjdIA8pVvmX2olga6t7Qxqjpj+3TVHuFYWpqGloU/6jqdx5EnSEldF3qYan0
CnV1GM7e6HM/Xu9prYSDQ+N3CIrc/01Q/ZfazQJYrf4y5Yc1SotZwVT5MFWyWPSX
vOD1yZboH+OL162q+yczf/gBihjMpttRCG2AM6s3+AH2DOPzRAs0bS9c6tmTZjjI
x+Fqca17EDexhwB6kjNVq4xCI1O4P50n61Q1bHkokdttNM7mBD2f5U43FpPzpc3g
bE7Yms1apoTJW3bUtaITkOwR0WLASQOLWRCUFxO1oP6RvRulyYuJGFgZbq+TJ9QL
aSccXdH2lRilQ5w9i0m3j9RoDgrjTzxeRZjfgNX0AvV1+jvCo+uSvfD6CSilRleQ
9XYxreMe9z7D0fKb61BFheY0wpLEZyzKmoDzV7irECy5yz/3PRqJQGfQsAwy1DD/
uvQ2l4WUipEqDj46y4/oBtqtpa1ZU1w+/zWNnkNdzRuDfaiEJ/gXgMOOwFqIM2uf
xwvEbEvusPJ0XexVCWx9H0yZSPorMdeFmBgQxUEKqk7676YqKI7875Iz/8vZUJgD
APODEMrlXU1uswpgbtVqa9rrShLtosfQM71Zkzg3AgSYNLr0kZfwOlK7qdQ+k47d
vJK68AvAkYIZ2ygl4MDqa9LD40bmQObtrnUgk31E9/iBKC/Bf7O+24v7DmEGb2Rx
ZY2MJe3tsRgUCEKk7aBTSa7uv+gDMXEf3XpY71QQQg+Gco+WZw6xBsr78l0yo96p
3sWNXqy4fMj6Dxk/O8FPpcXx8fhYGH97n2P6o9d/wRy+fvEoq36jnvxSR0DQozHF
Buv0x+NPp9G+tTjOdDB9qcYX4Iqg1+JFQ3ijKMLEE5PcqKd1282fn7Zjer0Gazuo
gxrC+R+i8whiEtrWWlJvgwHepojkus8TuIaefnK5hlfc1M19hNZ0e6BwMp/g85Yr
3OI+Gp+qTBQbjGcDQf6B3Ttzv881Cih4qq8tutn58s9d/5FDlezNZxjyu9xxdDz5
FdOZ5Vqs3hQTsWTfmH11v8Wb4EHfT+nCjvMUzCnPLqN7aIJWCDb5ghKgSzyGqgWQ
xq/ZzcgGynYNhnwh+8vvFQyP6vFUjOTebhZ+qEvEPXExn82HtTJKTjmDY8fKqgNU
S9/HAySaL/i+RhO1DvkLgLYnhDJt5kxrLuozeGkgqLE+suWFclA8qlK8mbcTrbos
5M6soW+3N9UKBSQ/DvpUVAwYGuXg8XJ8NPf7vYGe5S9mIimwM5Hbj8A4oIrEBuqG
bfz5yQmPtFzJN3Lqq0W2siEi2IUAHDWiWbcTles0gs2Zfq5Uru7MHwVax0lIywXl
2Kq0tELAkz3kWaRNyfUhtp1ubPHIABnItnj5tHt9l2K2f5DXHlwKKcuW2Wh7OCDm
vxszg8e5UOHSp/LAT9VwKOxRhE0aCmkZ4W1R5MfK9Yuqk0mq4zvDFD551C5Xtq3m
QKBkuqk+1yF/KP2shW7Yuo+/v1KICapHI0RFENfIH40gPf5E4QTbTWGlBSzlw++s
Oys4I8AHEI4PAHpkmQKZhL1azNf0ZB76WEkRltbnZa/eypeCSeWRSGt39aw+Bro0
AsM6vXtZpCPZWH+hWH+QW3EG972J7yn8hKb0lTCKOYCDGdvFPsMxjlxws+sJ6L/R
e1WS6a3/ywTMnaDCe/+F8TqhpfH/8TyKs+OMqgp9lwkFdstcYWEHhrADTApU9M20
XaNDjOW374dJuIgv2ic0OQZYT9VabvPH4kB3MJ6nlt2RQa/Pc48ttFOhkKvKCCJU
8xSGEpAtb+80BJMaFAZKAn8FG7ZioijzfSfM+LvBOzTi8OCEFqeV86nkGW1nXVJA
YcDIx2nUhH161z6imd7G/XkeWDvONKz7p0yGTghRnp/LvCxEa8SWRRobLqZAPMZ9
ZQ9dupGuqdxdz2IgEfCem1eyBR6U+WeKWUedvM5rJ893d6MjrrJecQd8ZF+Kkum0
oKYtKhIMODSihA8pWkieaEmC6aKVi2f8xjZ5E+d75VRb6E7QonFrOTAxU67QmAxj
bqgD6sQjzeLgVtiisYXoDT/jnkriffWj6RAGGUZHxZp9o/0hO12ZYceuf60UAn96
cL4hxEjhMjgR0UmbW5LqfoRCBj30wR4MK3ldkQCqHsokKjDOnO5HgsaFwcoq79m3
x1/mLgN+dajuvnn8UqKwyEq93fi5ZlFzudxYnWsMcsZh3iqyjpl3whPOLAJukMHZ
lC1ht4L1maQJ7nu5wCo/KA==
`protect END_PROTECTED