-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Bv2COXC1zf/uVM0NXMdRhK9dilmkRY2p/7lDmTGa19K/iGlnVVu3Ldn3CbMhTzPX
LV9I8pg6ytNb2K4m1ftBDF4ytnq31RtCZbcoE2tSV70Lj1LT9CT+Kg3/dauYKw+V
dVYiDQGCYShbf1QMAMlRs+1Tcu91QAmImO2sENE8mU4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5560)

`protect DATA_BLOCK
DiTusFJcpUfwTROz9c9WVhpXcK7bA23A8MjOZBUIabqxKj3keR5dSORm7MWWc4BZ
6ZA93ehXD0HNZgVlIZDN9IAIkyj0YYeH8Mk1sKRM5WfYJVNDbuNpgr6jJD/thmtj
mwiQhE3GrDTaf4OCpmIGKj1LqA7hsXQdCY0JD7ox13L2yTphruBuHnVLumE1w7A2
Ob5Y4jKGCmNX7FcyzTtAlOkdsWU3ah/Un8y3gdrymVhv+IrvxTEQjueWqvi7vB4u
9Shk+PnLLfVe8oI3LI+06ZmJFUzM0oWagtagBj6RYy0AnYfrlraAoDObXzQ0z4+J
aO5/iKNkuB6xLFG7K4VANlmdSyoMylycVBzlGvhLcuU/XtzoDZv3bmlO9LJei+s3
x8WcUV+yikcsa7AbZRKvKCNhBuLwCXXTy61XmDh7QNVyJf8GpX79wmRj4qI6HkzU
1xYazrmXhAmQlg+p1uYWaD4Tk0/o12rGSnWWy4OgdifQG8Octog/ld06uVGY9vjw
35XvPMX5g+dh8G8s1P54BkVtrQ7E93ED4S7iaB43GLDRgldpwmsnV+gCmK6IT8sz
v7L4gfRTCokkkqk+rMFi5LTWM7LmvEZitfwJjT27Qk+Oy9rODlfXsVgvB0uIStn1
1JVbTpqBvFySeCwmrEJsEB+L0Zg1caEbb1zgFyK88SAZWvGfHMyzh7129G4pMI4Z
eL9BCy3heynvbB6OiCs3L5ZgeTDOb7K/emxs7fEKUR3kBx0+Uk/5lxH5vxEYgR2A
qg0dcTVWVJ42TH5jKhPafXEnTnMTXtaQOxX3puTCrfz6kkKj1O7dYhcR85txo0vU
5n5AQWwFyd0c5du+o27G8DntP622Pdur/eSvmRPYQyE+B3n4gkha04SG61djSiJt
U6cQT15bBUyk2lmVr60Lj/duuHGz0D2DqLAwTM8s5oWVJRkCvO8P/yoPbzzvBgus
5a94HFLBmgteNBx8jOIOqI4NKwYeWZ965vc3xwY+PTfktX+zjDumI86t2gN0c2cB
o/hDgDjf5hrxpvsyaPKdE+cQxrOTaTOcIBDdLslhnKiOD/VhqiVxOq8Iqw7tfyc/
wmfjc1hTReo0bqyDgx9Xt5VF9CiJma4i/ughR7tHBpN47/FErZfFdoZd51k9qPNN
zkbXXcm8cxk+4x5vEDdn9VbI1nS8k5URO02MgDheVcQHLkwz7ZQGA2Sb56LOGEO5
DgoSzmVHwUpQajtgUw0blWT0qvggrw2SxgAywEwCMqiulbRV7nejqZSiY6Xey8hS
uJy0xsQ+Y37boB0VDEcrrwdmM9KV2rThIGDayAk6x33uxqDw7rmWbluUMjuVLWWY
nIAPux5czQbcPyXv/zlMVqSYC8zh7Ml3CJGLYOE89kGSF3PzNELpy4vHk8VLUODm
9G7H2yd5YA+Wd5Ky1QmIixuTEYmC35y2uxWTb/ZhQM6ruDCzkpjIOJXTb3t3toBB
bbz9sNfhjRWRTyu4yprnsrfGGxwfQQpL3AqD103VLaFIg4JHmnDopCtGoIrAhvpO
SKjlEmuULowBtJbzBzx//vC5qJn4zw5qMHeLLyNas5xQeOebSVwwm95rSwWcWwzI
zsSdNsZUlw9jPYjTugomuL9ed7b05LWuJKbJiIbi56NnZQh+Oqgyn5PiXoNRgSjX
XRZQfCRGL6Vlr5GgI5BA7bn2GIL3L4o5jpkCG4aVWmzA7ULF+TB2us8F/b24WNWv
HvrZSGdjOjVgzl6Bzo6ZFR579Iagwcqng8JMwxPE/jKT4M7NHh/L1QPVrtdslFP2
pd/HIUjqai6tC9fJ9BuiwoqogLG3ykaCE3eUAV3vKoUWEf1vvz1ZK/B3k2ZHuccJ
Xb6LPKKtmB/vIPtAuOLtHdFOwrNTLhtFWIb8KRbjgRWw4So31eI/zcltEWuNOYgM
iRbmk7o9AgcDrtncG1kGHqfgyVWDCI43Dzt6zE5x0DBTvSupc26nSg0W7PY+5IMW
99Cdd3xnWsUAqM+FclaExsiD9hUhhcN6i6Swwoa8cluiY5VZsJgT5gIFIsevylMl
XNR+xTPB+3rZ727AfBpMQbxHyV0ARvqaguiVcqEy9H+hiweIf2y3/wNgn92nQsMQ
VBRH38SeT/LIpbMD7gJQ93ycrZ9weB6DP2hEno64EQ8h6HDK/+t6+n874X21704K
rlSEalriCn2ceVMN9YSRxwI6SPH90/73MrZuPaGNw4GpizMv4xT6Na4DOjRwzeDB
drHmU1cjbesUyjF+sWfDCYrg7OR12rpc41mpWYLWojrlkThXw9q3evk5J+ai+LQb
82zDG2BP7q6lOcmR4j/XmShdM2CTCtzydOjhL8c+HHkNIA7ePnl6Z9oPeN/UXipS
3rG8V8B055jOwku2Jclw4yiRKSEbHzZPlQo0CuT8h/9cXPwCojo2uYx/upz9G2Nv
jdKPdPQLR09CnOyw5vm4acfztQBKh9zaPiZqfESTm7rcjTjR6f2qksn4gEmOr+T3
8QDGPzk5QKeb20os4JfoSFNLVCE1BUY3wUM61aKx73I231eFK66yekDyjDHRKdCJ
DKSGxMcijrnWzPmeHNEUThf5DOA32qZJyLSF5HO/Q5IwXKAD071v7oCmYssa/20l
y45qyAK+TIYFNEtCmuEav8dX0zcXUTc0owYG5BtMF/5VDaOH5nTyJ/hziapEhr3m
X8qyhPb+7ejLbsRFZQrKFI0yZb6o1Qzp/lZ1S5cO6q+5tT/DPZ+AWeFc9qQhdEB0
X/W9sTN7Il4Htm3AzY39MhHi6I3bP6xQehAIS+jlMsIYiyuoCCMnDQhr9a/pazyS
srCC+247/Vz/0DMfI1kplODaqFFfPxQg5deIAoh7SSBZKADmX0fNH1c4IZerEc5x
YOmwDBnHXFyhwQ59/NjwmzPfwVQJs7QuUE/QRtvvlKIVn/bFeCjBa/tJZ/Dh+Adm
l4rZN1urswmYyQPlc1attya4bwr6e5d5F12FmEeUXgnxZaZyYzLaVVKPM4Ar8qxq
B7uouNgE5/lWB948IgcDqS4FtoRIPCZMBJMzJyUchnxlNWnwAgH7sRYlrRkka0qs
PEhUoyux8sodn4UQg3NdaURND+O5BYYjHLPEtXGmq6IQ7Ac1u4wj6CdI5KJmyZDH
qA1pq9dmXNkmUOkAaByKgNIuptOIlKU/sWk/XuzXuFmpO/i6BIj3KwbphT86Fn7z
jO/KGfbf4qL1TqJZTLS26b74q2Kmb4w5VODeFR9V14BkjmsJFRfT7r6xTtNTGzR6
NdaNdunRtOyIyDujnE4plxrEf3bmGbdAFSSeApQYm5A2Cf09poosHevlNfTRZpej
ajELA3tiaELY7xXgvHOMFa/qDrd3PAlvvMPPEYWdvVxIA9FPtCM0w3SE74ysJACF
hJuXBxzP/3DOFRhsTMqvA1g8dczHZJ3ISZjQ1QxTuTP7uOmyZG/WU+ALczsRopMH
miIshGWA9B2MAM4TOJjfyY71Z3SOk3JgtdIp/190dzMHzKWwWACbjfgGJ5mZxczd
VQFtcfYtldEiEzdKuetrhEUYdYgGpOR6FIBrr1cKIs5XU/Zx39fMwq6EYvzGKcbc
D2B14SZQtKdRHeFk9/QVR0vNWWtKM1bA7cXNCrsQdBha4vHFa62KqOL9SW3oFtAi
zIX2u/0GNprrdT7VPz6IeN8/sgHV9zNdMmQ1kYHBfQPQ+eJXM9ZDpIhlJ1eY0k0z
2PzKFmMq+OBaYUfYLj82xIqLCziV3vXvi+j43RThxPNxqhz8GuL4IF4z4Iype8Lx
rEwREHL9FLhVR1lD3vuhsyJ5+xRYHU7G9und6/YRnp1SGZRu4c+vLyqFCE6XF2bJ
hlgJFnVw7j2cZuct9NaCgzXZ5d7BBWnkwPiG1osv+x0j0lpiGhU54Sw5Cu1J6Jj1
Yi52EBv9r5N/hJriWocXNHMTw7KBoE++kePGRNwsq2sQPVpM4+KMTf+Oy4ngUaL3
vGAwA29DFlAw2Dl/TiaJMQSUNjKJFXEanwoOWH27zlqKcznuSNQXZFfHUnifafjd
6PuG6pESK6L4vv2yphe37mNulGSnl0PNQNA8I7gveP4x2eyxrEtF4JjytYs9FdPd
7y8bjlplgHqKLzL1SGUFpW859m7936Mhdql4wabxdVYNi9u7KJ92iORe/Q8Q9ccr
oPMiuQUJ2kaQhy0U5X9bFiFrVRW2rEA3gxPwxCNIPjgmgxpE89AH5jST6pgDn9Fv
JH6wXknJHSZYoXzqaLQN4q8oa5sS30uI3+Raa5MLDnOxL3ZtZ5E7qIR4NTAVyMC9
s5ycBA9uo7Hwir6qfnwf2nAtvzjdizGAP9oOFL3D6obsxTCWuStjID9ETYxhFyCq
DPKQJBf2CZvnBxyio3yEl4gT2H9gq69V2CAIlpEWgbSac/X2OMrmUqwxITpjv/tC
8q9HRlZjn6BXUz160VBaJIDAAQo0BFB0Tx1tDpGJBSUYqDwdlzNwRU5OR8x/zlbA
01u++meTjM+DzR3vEDIcB4lhW6XNleMUxXukVm0mUORHwxyuD70iiliGaWbtwatT
E4Lhp91fyB4W+gdahV9JT8eYH/Iml+U+ow+Of8MBTMkjytuGtcR7J3u5CV5QPl5k
h2uWl8hxqwwr0U7B7EOQWskCjLPsKtrc0kNSjIPUOcS3ebE/UnJs3KZJXq9fvtRM
gDs1ZE2QS8A406Yb/gRuzSrXul937SRNF8e2R705PVjU8sPhEwiJYacqiQW5Bd11
452G5XvRRY3u9FeyXS09QJ2rS+Zivgf8I8P1W2CJQnjKv8v84PljJQ5Ira5tNHKV
Tw5PET0Z+JmkY3LWH778qnBng/FGqEc+vib2mpeb0wSb9HcWjd96qP6mdK+5ub3t
nIkNcxUjhG9pY/F6sk5f4M13pjIVIlkQnAzmGmntWBxk1Dz+bx4CXqDbT7zJfRxE
jZppr8twui70SwzzpJUgkLHKJUN2YEh2320iw7yOpMinCAXJnxTDM3f+fAXLEHw2
mm+ufqhGxy/DGNV7xcAUO3snUTl9JPMhkGYMTRNp7/sjdEl3Glo4jJhlBRfvbiHU
YZ5ENJ5NpEalcvp7h0Ff6Cidq7wrXyFR3MmPTwNsB+CcQn7flSUhXq+sHO3U+FNZ
f8dobV2IlLZKLjP0GunNMN6ifW/AtJA59WD4OgOB9IHMr/g9C71vqD9WKVOL20Sp
xXLCyVWIMLHhos2s04cDg7V9HgzdEhtVp9+YAGQ0aPHd+eHFh0TWBGUAn7O5XDOC
I6137vuLMfXvlECvWR+kb9rRGoYsjK8qEe6s1vcHFQsnBFn3DL+LERP947+/NtSB
YaCyZuAYuDvPBJUsATCoiX/bm/rlpk7C6jK8JDFgHIiy7hDU9PDT1aX0kiBnMRto
mjjtXmMnfyJCDZXIqxofvvwMUuWx8WtSuGbjVWLvq84TJMom1zGAyOED2HX+WEBd
tQ0UCZHLlxinLtLXsm17YhP8ZDbZpz7RYW9wxCoNTY0OqR7zH8l22u6/dNPD2FsZ
Z9KVA3O7NnucOMLuE9AHyHOGfffaDkANoxD7vdpChwn2MQPyF6fiKkQkIv6UYYET
+e2sFFhkxkFQH26dFUXp6LO5sTLccY1KImiBtn6dNiNufkXIQxqvWBpWqvrK6jrc
KDyUuoLdrI13lY62iW+iEY9Frys0TV/RJz8NEHokFxAOGeiSl8PTDwi7KLvGMKy0
cU7LPBzTg6aZAhKBvFk/8QcS2pXMAFlf+C1elPYYkoYh2bMBy3u24tY/JcJwCavo
lZ/uylemoWWPdvFJnfT3QlVuQc3icIo3yq3jV7MgMbs4N7W4hg0lQ6Gevsoirpdc
OhyBU2tRq/1EwZ2cxNREQSTM2Vw4oX/UTO9Ccvev4KAI15lGvJT3VY8BwhyKszQd
aPX2vc4vM5VzWS2LY/gXCbYdYSpycAC/e3t6lOyTpX9vKVZmGC0H7YjVvEf+3uAO
+B3OkJ/oG1j5V4pLAmQ51zzsyqUqHcsNfen9HjOUIgl0jC/5/g8zLN6V0tErQNwA
nuevlYBpvrkTk3LKvUVIqzmH6KKVBEIWIw5hL6rqJ6W27ADj4Ugybl0Ne42/ikKg
gyXS5PRnT6qFXcD0v/RqNR+VQF/JdA/owjluUlRu2ZKgLgzw4gW2LDsgDXdySzO/
RU4LD86JODYoZp3LrIguaGi2JO/ZEjYYxqjBMKfFVxAb9/ciEcBnsmzH5Vmedp/1
2/wGViKHTKZaJy6WXwvxhyWwxS6irdtKyOeuvkSUHQqRk8Kz3Zl1SRYQ2jZU8lfy
yiiavVebMalRP0EOfO2dp3mAkc69COAPeh38i4oSZQHTpIZUvM2RR7LYKs7Ge5zw
cdGF7GV5+h93bnxTf6BY7Qgd6QsNjlx+AD2ZQBLfwE9M2sgbyt8URjojzZvidcEr
TcciXaaQfCM4v7WoDhRtI0xEoCSjU9Oi52NddQuDOCT2qk5Xxc1kmlqz6MEMqtLK
wVQ59egd/5MU2W2eMhV7rlebJDaPuOJ10YqvAsZF6znMBOnJTQpEta6vUMydtakW
/Z1T7S+dzU5nGTKRKoLvPI9+KTy0aO7luxzgpI7pHS5LzFdjNq1/ERSLvqVA1l9C
slh1KAFKyy3/WqQZxsMXuKIyZJJjjUF1QUlwPVd3rzapnA6JV8pyX5UO2KbpCG0M
EpVjLBAL2M1ihmMI6e9LHqW2Zy3zPi0If68Qat/2em/B27tKAusT0YAnj33r3POm
LCa4b86xhc8GIDCgCnjNryRjIREV3xx/Pwna1VeInBGDQ98auUF6k2UDXbjjkJOj
sxogmwU3Fusp+0+DIwjTuCo9PdDnhYhDHgFJ5fNRfDIMJE5kpbYRIXFU6aAG6lDS
7dKec8Dvp/iDc58hMbPZ7oCyBy0kFm5BhXafwr5kGj0hYZn0WqWWCOTsU+pgRvQW
Lh0jY34zkJh7/A4wdnnPt6FrWiEmA9gvro8mkY2Jun+RmZhd4nKFW6BmtXgx+nja
EAPtHXZ52G9KFzgOGRAva8llCGDspgFvtl8EgFnggYZRulena9nXpx+QZmPz/Rf3
KXA5yd8zl5z1ys1ifFkny2kwCkQ8MNeXfckNwuKmaVIlwOkfUvFekuzXYcbFNyww
s4TZnRy07Ku+Gaw+BRxQiOIOOeViyEdFplb57AlgBWoCE71yDlv3Fod9c2I3oZEl
UkFSLFKGKNdVQz36ckbzdz0nI0f6Q6Pl0AeoqFW5ZRU0C9kCezLrmVwYR/qiFU6s
8xaECamFmLOsoFnGOCTcgcECr4Q7D6lZsNQqBp2fRKQl3i93hLRElG1LZlcoTZ60
2bYhqlIhbRq/1NBaKe6kh1jFdiKd78kHxkHwVKI4vGxSuif/OQJ90pfTKgCXHuGt
sVx2sIaVBsTF12qlxpRnNspsixHsNlbZu9S2qeayz27Ii20hICc4cU1eCqHTYt9N
DW9i+CptPmquDzZ+OFpmSQ==
`protect END_PROTECTED