-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
11BVBzCjm51ZlEqFqrvYOTt9XIMsjoWIsjy0rCoc1KoXI2nNf231qiQqZbA44k5d
LDba+Y9rObhLgOLzqNJoSEBrSDJrVvAj3rhoe7sKVJCluqYc72ujB+KFXtFBM+7d
KWMxVg7hRP2dbZ3phgqXsVO0Dbab/Iic40aSqx3rOqY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13056)
`protect data_block
CdMEnKgwgee6eUHcBYg8r9yLR5ksdSKqHxzUgD1z4fPflUI7vDYqrbQIvJ3vfGfu
AfIZZ+icHhmAEVcnjwn853MPIoU3ep/ZJ0zpbnfWFV5a7t5EPr0677qSIqHkPa1m
4MPsb639cP/62AgCnQyLTg4Ei4COcXXbJtvUFPTepu0xsS306a2wRJCt2ea/WjdQ
0LjrTHbpCiQUu2ec975MEmDxRNP+CEGq4HNSgNtRJ5+3O1xTK3Cm7cMNAz7lwCMO
dqd75MdsUhkRw+xRYjf8NZf6Q6ro0ExOEP9sMyxHV53MQy5rysOPl1tvCwSduNlm
HmxJEdY5P5QtNftrnMF4KpOwRnYfO/s1q33G0rAuLkNcQ845zlr2bXAZRCJJA44r
nsm9MIG1D9wKeZkb4XGp8hN6HNGJJR+6ukV8N2K7yPO4OPwJUVltCb6Uh2DDVv1e
8X15pc79A3axZVblMFPRPbnhvWimPHWllyeNXoXoq3nQHo02uIjNKAEbTgTgCt5r
TrmX0VMFHVksAMmgKWe7koSEosJRBqfqeJZvBZ9rIZns84f7+aPKvDA4zv+vKsZC
ZS7rFRWtXCOw7PkSYKSnS6rwqgSk4BsKvQH8w2lV2s6rs2uyq5eOcKWxqYryoWa/
z1rdrDk0A3xfBrlV4xTrK6RXKjjJQ0GADIu92MFRW7SZaG9YgkA8X++pp4Nn2gWT
+vtEd8FM9Cd9CeokRbCi2McBIokOPNUor+j563S4P2DnFQuQSmL/r+Q+XTYNqt7n
HtcHJz1e7LcPuqZg/n8q/xDbGClAaxg1wdBeDWsGQbJgkg6pGlsnBghAfJd06uHW
WYzSoK9Nw9qE+YIHd1FZRkpJk+nYi5Z685sCbA2DnIDB1lvXgL8PF5BVDWIF8lSf
qL4NUfldqd4++2cGCKc4qsY22Crnmz0hmRfNTyqIbhQPb0g2LNm9mdYehvUaZBnf
aPDosMsu45FuSU/c0bEDm1qIn9vGssjB14XnWHamW8aaSwTSPPbVpK9pJCPC+/k5
hUsxPJPa1H0DXbA5f/i+mYct+FzbNrL8k5OKg47FCLHLsy24vHUFgqdTpciLPIT3
IKpYKFjyqFEzgB+TeivD2rAcM1+mc+k/VIB5x2gbaKXJwL2JFHtnQwbHjaZGLrZ9
IYzLEssB78qrBMbMib3MweE0q+PZiPy4Z/3KJIJn9Ps9WXmkAI33YoaS9ogFckem
bOtKXKwwcsO+cinXVC3cyKpRSk8jdyd/UsQ+2g4a5BJdX/nvaseCYXS3JipOAoof
9xEYp95FM4we3XRNduaL24okI358ciyC1Ty2mOPpAJjDa/huyDAWlgmSJsNPqPTH
PVu3b2L8LHKWctgCP7edWKaHJ07qZpR8RVgGm7r6JxKlJt/Gvn+PE8b8kQIXABv1
Q77dolVQ7QYpQTJszbni/7PScOrhVXYGwSdGF5AmLu+oB9rnZyFDfKtgNtGnASR+
dByKRls23NNkIrYB3vmmuhs/PsVJ4M/sj3bPfLWWZ/lCFHEjGG1yLLysldna8fxy
tyIVj4ldIH0xRm5dc6pzr3sgD9CAdmcCfoJJdUjYvuhi7CdGSqZVQ/bzhyWfftzj
uL+paq6ZWu+Woxq6SpGoS7T8hNMyYnJO+Y2j1ok48q1JK2AsKWOldbe/h3LMvmJT
/q0gEJuZUcKX/jZYQq/X0OLEGn9QdhLEJmt1WsG+V/BSR1kh1ts1jNcdRTCaWVx7
x6Gu+B05OhJuIMD0F666Od4hIBET7U5yRtcvvhmVgewp9CI+kE/Bw29524NsB4Y7
epLBJy/cTsJ/FPQoFAa/LjS3hIQEYkjTTYfcFPkTp4Y4/zB7bke1/VwHSj4ldV88
6xFMmSLAdFnWqrfZOChCmQFv2A1HzY9WWkQITEQcA7ti+2JEj4L08woyCLbfnD7+
zJlN+DLXhizBg7zjoHEjVDb/ZvXc3gj7teM9o77Znua93yX4dg/3A2cqCTkJq4tc
f+l5CHcPjE9COVoMSKw3G7WRExI0FAkSGSs/24jlc2M3wyY2je+6Q4oMSAc0nbPW
3O7UQVZc0qQ0B4BfDVJlbVcZ0m9ddeFcs32IoXjVkoou5y4zmLj5xdqrrCkJBxLD
YedQoaC1sfq4D9aqnPLVR2UMuzkH2JFj+80fG3ejWnta62WcKfTsFRnr2DWO64xp
Tog5gHM8WRuXVccrV3eV0VnBuGQ6KPqV+KGvK6FlkDTDmDCKwLGUpljIVfLACKpZ
1wTef2q7rOzzpst5bhltDCIp/FSTghBQ5QFK9/2X8otov8+H7ig5JMIL/gt6sxse
wabG7NoujLy9BwROVHlYHowj42E5YrWcI9qOO8hdCfDbWSmpZ/rXCpdOg+Vm/yxl
FRbIGYdBPzPC2EO2v9eVNi7AcXJtOUOls9El3TbyEWuGib1iUuxvnxVBKUPo1p9A
vdzUtiHYkPS724M7hMyhYvZjOHRGUnPAnnexmrXegwgqXmpp3gpaoaKI8+E5qQVs
sAL4VKaw5q4rU9Rl/0zviCr+tjnNfKj/OkK5glp4k9pTGnViFQieKxBK0IbOxx6+
sr8sMjFpKeuVoTmw3U6+ILttSno7fkEfIS418oD5j3dpKDIcPw/yRIGgU+uswZ6C
uLgCjZaLOf/Lt1jWh/6YYgEAXynqAwiwWCcbjXMFfa5XlnNunk9K+qQqf8nr/JHS
JSOBS+EsEb0kw2jqEEglYBE+zusQ9gT1D6vfO2edq5gXADmfUgGfrzqR3C8NPV9c
UiSI09tx4OyV8rBhMWC5931aQHcbPNGMIGbArq29du/1kQp7DUHUPDK2Cap4aJPx
jsSiUkKdf2xr95HYWP89Lt9c4Lj8xdPuLAwAoJ23XRngJzqPfi5UZNmXkbMScPZS
kfAoDZsHF3s2bIwykiYQ9WMvkU+h1qBj0BGGz6DcNxS9M6oz1MpDYGk4ZpqrMFxK
wfFmCcSmtYHe1Ik1Mmji9fWaEQXQ4+gLEAvfpcdU5CkqXyZoF6a8Ldkk+46cUEe4
U5n+Gf4VPW1SjRDxkE96+lovcxqx9L9P+kKUUDCQ1/tzlL8/XrpfluVC9CtvRgCM
8aJPtQkCaQjOS9GpE2M9daLQ+kRXWhDtzYbCdBeGdeeTBkuBh5sq2u+g2hEJ+R1T
o6Yd4S82KWxiIhXWK3ZSZAQasmaa0SKLaHrCjiBvniZnJnvJx/SyvVUog0GpYd2v
dXJNDzN6BSgkZn+1Qw5QI6SHM5iZx0B9/cazuuiPWckkxNh6n+Vw5e2sPloM/nhp
GcgI71kQq+NBrVXGvt6ncom45hWYrqF0L/Fe7qBiH35otJK96JbN6pccjRHbN7di
Txhxj8+MV0GaLRwMpHCEts5rNIdM4aSGOGOq5yUlDO+tbtfdznUIXnzthdc8sc7K
LBVV9A3NE9UT1JZLjGrGbwAvDvl3KneFmvo0iBOjJx93hGfi7v2DfMBdFf1+gKrS
OCBWGSzxFFuF36+4D6mBzkakK9qTXIX07nn1f292vlHPiLVPl6xybf7AaajB8851
K5s8NuvSLhbqas9mW1jsKznCipPUUxV12h+bJ3Od3swH/+MIyxxblZirsIj7x9nF
Et4s+UMlFNzuN3bDPuwrg/8uX+XUK6xKxBYk761KU88xZR5YSuUeINZQcIU1VQZH
xZ7R/rs9DgC9NTPPlTARcW8eIOavrqwY5fQJ9tVDYUpJgSVVk0SyEtKNG8l0b/wK
QS/1Pgb9ZiEgLHfYG8bHKSPrDB/JweqaFNKz9uSJ6RqR0aUtu8kFSPSJ7M1zJJud
m+SDV3rfkry/PPOgETuSmPB1s9V0ByST7dIsLoVLFY9ZAevsAwaoTBGM9D/j1PSU
26S6T422T575HG9IyvhpgiOTvjCqkQbcr6fglFAvRm7OA0jcFzGQkfnkqVKH4r23
4hQC3tFWcvzyEKc32dwcrprWXU4r7lY8Bvy9rf7mCfM4bvizc53A9c2QCR5PgWR0
itzBBsqu3GsRAQFsyLz/WAmcMgHju0ZAk9fRyqxmiBNWAQu/tkg2VdTr5NE0QMQA
mSMvWOQiQ1Tuxk4aLRy5Ppdl5vO8+60mQhoMWfZ8sI1ppMUmbLHhHX3aMVIqINFM
5mtXkc6nWuVQeFFX4WUgm2fO4G+xQPTHFZ+FblQLPsGQRJFExDvN20FIllpEKMKD
t7+KzL4AQplU4PyQx5iG+pUvGjnArqzJCahvnGG0Aa8kcorGVh+540+6y118MpOl
I9HH5u1GqF+WSO/IwscrQA6Zny1bpRVQpPTw7XkwKR923DyBRQzQ6OKnLEYDoN82
pMa72cuqxCo7uei7Lq73GGXJtJ2sErmkfuZ6rV6UbwFoyG2eqKwGxHONgZhMJyEW
Ty5WTcH/GsgAgIdGKYBM4LFly7id869nhUXMj7LAjwyh8LZ8a6Ppu0nLvFsQcR2b
WqU7UafmdVK3iWhYhOH3UzoWB3j5yLkSRqaQdreFEOX7CDl8NI0B6l+oi5nZAFCj
1vrjTRoNi8SGIs/XCJ25qJBxHoLc8OKovfNYOuJXE8+AyvYVD0nRyLBCJnBzaGUG
Q3GL6pXDM6pwPbz3g4mg9gJwXZ8rhzD4vhyDP6j8NFRubp7SiaCYvrNVSxCVQfGA
dpY4/6oAWmm/4Mtp3l+6mZFIXbuRODU51oJXhLkps4vlFWCZm/FGPB/1rgZTkuV/
H6YQWUdwoMViBgouPc8OpCJdoKYMdDiCGVsHMgI7jk0Efgl/ioQFwm+yT07n0egV
iRpxsWnOLlQeXXGptNgHsDZcWXDMZpTHI7agoyWfGfweiF4ZYvI+KHbNiPvJvykl
mRk7GpnwWKBXfN/xSMsyTN/le7JgnThPQX3exdG9auuK58uA0LC8QWfeMaCErbpJ
O38CeX7kkSIytfH2aeqoguuZ7fk6QKGd+uTKbIyFlef/m/cusHcwh6KhLEFKhLBL
qdUOMConGN58OvrROdLi7IFghldt6faklT8tLDY9eqxiQrxro/+2pZAlkpSCHp6t
Sphgi/34vjnLbmX5GlipeNrRbunXbohIg/BwX8nUWyrlvsmgMVMSvgi9P9BiG98E
/z+gNL0PtKHVEeFM+fOysJ2WavJnvhbhoxliPuRluYa7k1Q5S1x/D2ZlyhcIwkMM
hiYfnsLD4fErickWQ1lOQVhZbYa9keeizpa3x9ZNkfDaeEWHfKSALTc4jSSGRaHW
gaUoqgyDa63Ae+f9JcFRJee3cDpd9jPi2Wm6s1P1oOazAVxY3a6xp5kMRAB2NEyb
Ndf1E9EMXtd/4PTmwOK1Ja6SAiXLAWqjEkmwWlE0Jctl1TIL3DbweTUK4X0Qfq32
MpFGbm0S004gSAinT0CUs0gUrYVi2TsGgh7cpDzk7GYeBYl9hp7YzcWWV5PtpMCS
LkZElyB2k//X8KlFQcawsVWkrwkZ2QtRLBRkMbt3CFSyAXn5FSy9X1xY0CIiPyil
nWypC3TEbEZN+aJ15MK+WxX0L8SYrt65Sw8Ldqk7tUn9xVXhnMywtuU0tDPm0a60
k78UL3CzxXmhR9rqIjYy7SFpMBQeNtaUM8s0NWSOUud43i34K07dW4VDBZX/q6lh
YLX7/md2xtyvNoq5lpQB23WQ4UF9EEUY13fYhnaQn/sBtFNt5HI273GnPQKT63ps
KW+i66fNlO+1vup9XVkPYfWyIrqyljFzYt/GwrcELmOMrRkljROyGJhWz+FPHfxX
Hzt/T3hUZACy3Vk0LhsYfugZq2X0nG9NoZuJ12fDsi3Sk0nP8w375o+JBg8AzCuw
+zubB8tXN6AxCL9LOEnPxjdCl+C7pwdOaj7BLwzo41YGByPMR2mKsdQx38tH4uAV
3vE2epAV05H5g6Q7gvq/pHwXPtTsK5JSrsy2ih4QjpK89o9yDDeR2NCmFqGsUMMF
HVz4izaHArm1hEOX8e0Itxql/xSvryIEjcxzQPyomylD6lMW9Eh2Us2txl815Qaw
WY0NKoRbYNLvhuQ6owDxI3XvUL7lo/kw9I8/aKY/VqG8f9uIC+Nk43RsXashljbf
SDqc8veqAHIC9TXkX4tkkJyGL/TIF4sMBFLRYRp6mP/UY6PrfpqGkyUMaBobp74B
03gDjDE8TJf8HJ4WiwgjOg3pMpFLrVw2OJaj9usQgAVrFFExFX530IEhBj4EC05D
G/Ks91iB+6TjvvnlvMly/+EpIefIdDAweY15lMA7rx6F88K//KK4tOJ0efIOSIc1
8+Hz6OY5M9L17SSZtOESqTl00nQiF/7U2QCuR6gdL5dgR6DYuWcfvaChQMXSNIJi
zjPZzYu9++7DSCUaG2XJT9MK61AY1djsZgn3o8d5Q0Jeoa8GpaWy8yCyMi/+9hu4
qrNHN7xN08s6rchYiJgUnWNe/yeDzpn7chAM62QLNugt1VD/ewLsXGDnMupo5EdT
fseukGIm8pooSzLT3Cb4o15mYhaGnbKwGKLDe7Ox3QVC2/SFNk9gS6J3+8QYIIFG
4nBMgiAydpp8HC+3ghTh9uNjJvolMSocx5kVlIr12ndWGb47doRY5cxsfaXeYJeO
3mqlZC0X3wIHyKUYxdE0O5vXMKq3bussfzSxX9XY6YgtRZVwxPNRC3E71yyc/lq6
/uEZLDXlWhwHYybQt4oJX4Yv8bwynJFy/mcmLYos1IBsCrHOSJ0L8MIKT0MK8OiS
zuGNNOjILFIJDNy5QczwmK9yGkfraDwHskzA1Srs8nkU1AmJ/smu4x1I0+gjG1vu
GYIjslu+qhTYdvyzQhyloRs/7hfwEnW6raWroMQeScoxoedlsf+BR/mPPEzEL2P6
enMLHglcTPG5J27SUmSmWMMFWhSCvTu90X9ltloTs6/BFy2fggxgV69/s7F9nmD7
6GBnX4tqdJoEWZZKyMScHgTRUycWiiFzsdjap4QKc6XDP6g24cApdafz6740w3/Y
K5sKEX9/X1NxrSl5jds67CrAnLkF7Q3Wl0YAmxS5YYId4se2dVVrZpFZPz6/8sKC
nKLC0iVpuNHGjoaA4CcXjf9a7fgGRx48pkpi0kT+yVcngzeKdKz15KljsuMM0y2J
JfbM7g4JZtLUio6di425K6eDKrVmcwSTDlRfWid97l8JfU/nT5ilUdMQ+Ip4dyxw
2Y6HSguA6GJU0gSRjv7kyzIDLIwoSb63TF66A8+PE6u42dEDUq4rM/1zrxplEgpu
gKnL4HpqvQjhfWRUE8UeOdxsgxeqr/+8TFztVH78hjqcYWJhI830fsQ/Q7FtzLZC
ZLW/5/mdpQsHxguZeRBTT8bcW872oK2rC/7mX1qcoOYgwxA1ruriMbVrTwHHGCji
ZLbgHv9X69jBOp+IoT0Ead32lLQLEB3DguxqTQ1uhhCHpg0goGPsxxrtgdojxdxv
Gtqjj27T7U1OAqZDB2gOc2XDF+8HA99D6E7HbKNFgWwxcK8KLo798V6xawNHWz5Y
3zuT+ac8rFy1p3/1Bp3gsod6qEtJv9fb5+8NCMG+dK/lwdyqmspYf1nnSxrrOEII
CqJZPcEwqHbUjqxO/+xDWSDB4cq+986wGWZ0EwAPapr7tYeoDFr2qXyXjWsNoTGz
IN4Q4o3Z1PD5c9jajpUMvHVUF8siJ8RRQTfvW33loJYgMIuBDYn0g+Q26SXLdDk4
GTuqKkR1io6G4pEmx7ap+w5duLrOgrkOPzzy4pF7B1ofHvrY+0A9BOIZHJYsnm8e
O76B0c1ikZApWonM5OGIS2QloBSoZe/DXsrzZ1Mnt3a5d3OMALxhs30RsXjTkenc
9lw4YBjdl1nvJwcCsjuw0RxAmydd47GCXgs1IBmcMjkrqbHXJq1RbwVsjeKODZPL
LRBvVHloJ+DPsAWVykyxueWP2mXM/e7r4zu1Py/cMcX67qGzlgy/AWE/RwKnqDpR
Cdb52jlQJke4jdmVWVEm6019qGSsdjP1zAHvdeagwypmZLqJ8Rk2wGIaRu8Fqf4s
ELjIfGfwVQIQPI0KUsO9bZLw592xq1hAr9vsgdxMFszhnV6vHedZEAP7YetH0ONP
Uva0L0QPZdd3c11h1nD7kdy0709rH+N+04DsEN2MuGe5h1PfTrHNTLAHWEnaKM4U
QMSHonBm3nx86aqtJhdNhkcjnyOXPUrpDcVkD8CxbiG27UlHV7avJpNzLTUPwfNt
aIYoT5nWX08/Zz2sdAne/g/YyP3FESaZnUBeLa0+kqCtqunbHAkQiINdMqKC/REb
NBAI9QI06KMNuty9cq2UKazk3IOXqMvmgocyn6319OJ5DOreqyt/C+BkHeGLqmRe
MgAiZlCttd0CY9aa65vCPxmJ1Re15NnCKrGHI5htFzcno5K0PBGYrtUOl9qvjW/P
8q2trZcVlLqzSHVtwlqEas0MNUgxtfm0qlhEckaAacZpDxz8bDFDjZYLUqy09Xu+
IbdN0AdTS74pm4HO/16toNVonZSqBtVDv59Mefxq3dfKWTGJSzEf69f4zEgXZGKb
HhNIbi10vENdBiz1Kbp4KkSR8552gm4aQOWJ7xpqQFWdIZZpFdhxmXKzOPJc1gDC
/g5+leH9Gb4RoP62hGjfgaJz+AFleI7BJfsdMj61VgnxGuTlSSHy+PLjXME8AOGf
S11fENd4r8lEQETAvmSAokwCh3oZozwQFZm7irmdBuUQhqilPcu/P59ySArwz0Uv
vXDu20J50QOFzBEMtffJLhago74TlNC029e3HFTPTDX1wr9XQpzktwhOIDvIwzKs
Ftxn5kE9IWCE0d7GwZchPVLU9dS/JA531cADVGHCrpM3wyQqgPWNLueCgBH4mgL0
24M7Ejbeu7S4Sb7ak3xedEPx8lWIGp8NwEL16myQesTEAlQZx0bav1vtwfwc7yBu
95EBalkAaGjYF4HFcfB71k8f3cUaQUjiXK6/18UBNvfXXm1m41KQlKFe/JJK0iY9
935pgI6CIizjLfiTeVglQg2YafzWb74lL2/5WD1864VJvcXzvSqbwa2pP/OPPBVf
GXh+ANSuV/zsO2KEpRMQBN6b6pi3129N+hV92o4AnyTCWD/4nMHoMu5u2RPdEerT
Va5ABsKaTL0e6WE5zug4zJGLCKQhBoQKyOo8mz6wV0izpnKoyA2CqYAujhSU9ZHk
31wOjex5nMRrXU6+QtF0um1K1abrjISRpxG3V6Ox5v+z+BNfvs/fWH3hnkidH7Uc
GSU1Ni6TcIFEzozHBx4FDftOI3DQOV1oMVR10WFVZcntyT1/4gj81TATVNF6A4Im
GLxjOItBIZ5pe7qVOcNuMYLDi8pqZSe7Z3j6Beqo8yocFuucCKxm0MdVM9taa1ww
rIcE0TgyNQRSqVTk8QUK0bt59L87+nZ8VIV2zNVtFtdlNy3jNSUILnapnEaMvan0
+B76IOOciQC1HZwYlkk7W+s5lzIZRnAiVoZXMLQBxAdzRrM0ufyBujAM1/BJPsr3
MJQ0lIqleOEWbq8Txn1zo3OSrDPSMqaVknzbctzvWHdvQJTuxiQEm8Q3aBoriW2h
XPsR9RM5kNgXXJtkcENBfet25vPdqrIItIKWpJ82tzqhUCvD3gk4/xGF26YzZcUZ
c5IlCttMaOzdLcRGOaphkubybYeuatmhnKvQtJEof4PhgXYsQFNhRhP0PrHiQRj4
2FbCtkxHauOhTM5lhFRSMVVWm9MzH1mMePSxPLkXQHNe0aT6+uURBs3LV6GJutaP
8KEKu8NmRcQJ1ahKnyrW3y9ogVlXD8oWuQ2Fzs/DrQCB2pOEJh0uEhc78hbYZ20H
tP28++SC93Zp0N98SL3GDxQNase8aabij8mQpzqSUdkA9bkKRnSsWdjnnxWawfpS
qO0lBY2wd9ey883Z0XApTG/ky6Q2/VVPksVz9oLVn5CTlVAoB7mkSodfHHyYF5/E
+0R+Q90aHCj2HERRh9xsWO9TY4t1a85IsNdHdHeKE7CDt4pOptST8EX1i0ZcwUAT
382A+XUlvETQbiaiSKkZ23ZKS0jOCzJyqBNZ4vIs/WMj17x6W4ipJf0bD5fOkX53
wTmEwLUAqJLpKpaHc6OxIiS+Aaq4re1PHAMGej/Dltl4agUIMHDjqyLAuajL2Pee
f3vnzYoLZu1RV1r6kbTOxb2XhYHN4SsqfclswDXenw+XbRg4bmARnYOJnQWW0Rik
aiciiM9jm/ocRGyL+drbQ16OOxYNbUaGvSvH0mDkNip7+QTKuHJGjOzPXelqYWrv
I+iMj9XzkBM6kOGg/+LOczTSaJKUNk9svtrOrco85PVm9WlvJDQfmzkZZqwZ0mIN
64ZPQWdWZoURcE7RTAnhkxnBxDZkxx1wu4rq8WX7ekcowFVQUM7GGYkfesu4USn5
JCSxI+ZOD+/XKLOLzQJGi+Womf/XifVzL+ojkd74e6MtUXmMnw9zyOaxEWJlXRc+
tIw7tbdf8sCP0ujc5qKp0yeLgYg9fSgM2rmWy5tCcUKDiOiW5CLxLQt8+KSgiWTe
MfFwqLmGA6Ec9kmyvol8XzrzAh6ado17fhEeGzatDrzkNIxtnoOy5c9dHC6UT4oR
c87FJ8k2mM3f9ibxGWHuTSk42frG8cDR1Mn9qGFijaJJHemQQddtb5aw8IHXOMt0
xMivoQBY0y0xeces68j0tr0T3pj3uAyxAAW5fpTCe0VdXjwxMty+KKn23aBLgqgH
Dx2k1DubKEITCZJejreCLpwGyouAfjqoZb64wRqMcRvV+sAHJFi8O6+YjEVxoMhD
Iywf+IHcQ3YynWUJxImpeCfsJhd2dIF+vU+X0abjQ11SZfMIYfEH+TyuphnB8bob
yLBN7MbygJKIjWgs1japyeLGH0SQkRwI19e7R1qW5seQQJsg0aVRAiAGnXAAoOks
Kegkk974YH+0moiWzPD9Xu8u2uqDx2zR3O9h5f2Y6y1+EcBWQ/8c8pQ1mRRrKejr
d/Ta7c0ZcUYCmngmAw+of8BULqiQa5PuC3cnXhp8ik1jj2TmuDrioozjknph//Vm
t9PKKW/LfWIZ7ZMJ96XABVRwcQ0/wi2SMn/NWVbA5g54tdKeKiWark0i7q4OmPts
hsP5MlFf9hrwte1PyiLqdnN5VvATFRTp+xQTvCieeFlAWwL1NJ1GxxCYK5D4Udeq
ix7nA4aEH5gErbzQD3onVRT6pYf27Hvha7mnsrVz/8vrIvhUgLYTWazpiC+4IFl1
AdQKpcHtpX2jQtV60+n81yFqJAgfsI+wyyJ9Cph/0VLlez4b0OVhVPo2W94ICuHs
LKSk+qK8HF8aY2ClXq7LY/3NFM36HXEoonDV1+ml8Y/7UdVwvcQk99WyM1cbyXF7
pm5YRisYsp4jDyXvV9qFvUIflolBGUq/jyW6coaQLWH+kZl+bHCG8kZD42x6ktb5
iOyd9cLahu3PvffKkqfmmq7RgJ52qJ6/hMLd1RyNO0GpSsoP1PFSoalQQURnia82
17++p0X/M6qWaabNr34JN4JA94Wv6hW4gSiyOtwHAvkKsHlIMxkkq3pwRamWy8hd
6/zIE99nd4Fum8XCmiJxhGBNFLtjlh2CV+m7HzZCEg3ANDglB+bet8rcL4zgw+lW
0hCT/UzyUAhWQ3YK1ZebVaRvhx1qyblmAVVKMbZPRJc2eT0VBZO+rinYrGISBCjZ
s9oSda9kKjQvDGKMR4CQZIky51cPOg/ah3DPfwv+L2c2mO+MkPDE3v3e0DOz7tsN
p0UyNF+mYI9gbSJOOO1v6SfPraYNrw6lf8mh9ZwxiSC4COMkzqxwjKPXfr2ZwbPD
z/OIVBq2BZwIavPjnArLEbeDc6IYLz2eTpmmA2rKMGdp9iuLiiYgjz2biu+3T8Me
LLMicL+JPwa1Lvzk56tpHccQJi2oyR55sAuwtIIBEZpncXTmZyMYRotBvbH43r3Q
hhvYsOGmlNggMSh/ovhU2muzWOucQnuZKtdoBI5xBmH6PYDhX/yCzy4u5KaEiJSB
r20E5+OBeeBLnGgfOB7X9kTXGp3Y6HSk+k93nzUmJVPH591UrZV076xszlJoY1Jk
9ypWAFl7Ft2vN4yGQVbktcatbRtGmpzYMod2w7WYpnweQfZlgUtn4weeBpK9x03n
7W8qkTY77uBM+f+hI/TujVgrO6P1j0Dkfug1DtW5QqN7CpgcrpF2ADYaBZZCVT3+
LVa5diN/kPaNvvsXPyOs8BRlGsVW4QuOxT+/MBHBJq6v3Dft+/vitqe7x0R5pjN8
DTK0/ipBsvC3jF2TuGNLp8JASJE61RCtJTDzvYLqoyCJEXoePLygPckSLIijHV7/
BfcBzGY/ZSiXygji61MawBc/zUHOqkdcQi47uXlFsCNKxHPJHDzeDzZEh3OvG8NU
OaFF+0kp0PQ7/xccQBel5vTdieu3U6jp7wpIG38JtK7ih8EEvWNlVsiN6EBkmGhJ
12KH0TLyG0OcbY4BN11g3pB1B18dYUNP6oBf6fk7mP8slzceMAZ9kiA399c/DBkN
vsG018+1xDZS0r1h0ScpO9hf5x9OTokuKZo076mfsz2yiTHvgMvNY6bMmAkdlvi3
0IwdCRKitngfGQhVUKJo+z8qP6ysQcKqrGXF/NaUXdp3vODn6NbvJh/xZx2O/R6l
qto60p0fskcTKw8dpyUKtBrifXiS+08QzUCZVciBzUuYbh8iI0ryNC/8jUgeI9Nv
mANJej0sOeNLFVvAPztCcyh3/zm0zHcJeOCiBJyNX++zf/PijhPfuCRK6554ZnLe
4Ku7Ei/0eLVEaKpjjS1mcRxD6dEFJN/sQ7LoZAZLiDYER6ubL/iQk3SPjbnWTUhB
lA+G12aP0sYgxDyRFIiQ5eHn/tHFm7ufnnGsQ/2yzuy1Xj7MobIlub1kzlCcntCz
na0ZBmsC4N/HoYsW+l7NtN0+JKmWs1b4jhw9rm6pMizOmRtEBYjLmj68RSLPL8br
aNAjFxWjga0jJlO5GH6Df18iYltrgh3oerie7VxVMP7tjtiBuInAZTp+FFPIH/Kd
/sDnHJt0aHLFayadg65xvb0val2oo5Q+h1YKnQYCED/vs3Tram93WAb5Bbt8PoTI
l9mVYaN5WF8MtYWnNYuBtxoIZ+f1VbsQ7KK3fbfhyKhf0xVhU7sPmQDbXXru6hbm
u3L5mRiPKUbe/nzRQ5QQ1t0VOOs9PeSyBuWfr50gbOCtqnFWzSFiruuo/uc+mRMX
Heg7Gy+npvBxFFD/2hU5DidIwXvRCuHMAJ0CpB8JR+foKd2fdQyE+GpvAfRB/U/j
e96rra+R8hiVBD837JJd0cHwviMawLNNceSA9oqJ1zfuGGk2Wn4iyUqFfc6t7qOJ
o0nME4EnTdkMeWwwIOpdMcxWOY1PxfFHidW3p4WAWyCFWmw64sTv2xfKOORiBx06
lKIvqGK2L9H4DFWemEeUOZ0laYKH/56Gu6i/G4BDpK7XqY/UUJdasruDx6c9HIY9
i+4yc3IpOVY80R8/IxGad3wIYxfz/gtLBeil6yyPDFLH/9O2D10/Pz/c6DBYwnKm
u3hp/JvARxVyuAcwEvq8DRnjYY0Q74RmT2niWb1OBtyS6Cs5ACwqBbTki8v+hPNA
b3JG7PVeopqT4UOu1d5N609+UPYdB7S7WbAnnfYCn3HMCp6znNizdjT+x9aiQzuW
HQg1QoNHvOysZmYr9fbRwpuKaWs7kJzCKv3A8yIiqZGBFY1q9AhtYQcdKZU1DcLH
YYcgnLieSCQmhOOtvVsZ8AmgJpmP04H0bufEhhaW3N7OFlZt5GAfTdrPnAupy0nw
NFfg+6syUJTRIYEz7OrhOL0LOjcDeBFQy8PlXZI+rmCePhrcZgpmfbgPaz0S2Sv6
GW4H96JJyEJSOKda2Cjce7ad4/aoZMnXKeE/SOhYEtqOgXVMUToMsIFgntdSjbNi
FEFULBssoAV7/MfUIru12C87/XkrofOhCKCqXZLMJhYqNm1B0k7b2wTxCzufxM24
OqzAY60oBnLXR3RMv73yxAVFHPTG3GIFu060lNJe/3obECKzm22toR+NJr3rcx6I
bvGn+PM7F8h8LAKSfbKVt8SOIwBAjT4WdU7JZ4v6cixoWsbsCys5RL/Zh1YD2qF5
tCHrDxEnJcf/olTaDpmG765bIwS66D0pCxVfCEboJhh7Y//wtOkRzmg+o+7cxxPG
vFkv/XbY6RqtQAqPKgZbS4QR4fUa5NEu3N6xHEWIxxVouP278kLI6eMPwBSF5AS8
jDifSWPrmna6eHbNfXdImeMyCkif6HMSgLbr9vcZA+Zcr5mZ3bl0U6UFm+ClYiTC
nsQDKhteNLLQkBDPWRXVJSTHIn4HwJnLYe00DMSzLhTYRljIF+oEkrVKsvB0XfqI
yqdA9RHI7A+/8WYZQrvkrJQQ56eSkkLz2UQq4Yp9K6jHtmExwP9djjE4prv5Okzy
zh4pyeyZjE8Fyo55jsnfMUrnk8GhU6btX5NwlpIIJfT8RECg+54sIRCfXo1woHpN
ZwpSK9XeS7xxIymTgta2UBVsJAHj8yMoOX3AKZlKf6CGt2OVoW7vvA8xVssLAJmb
qifYE7dsc7JyJls2COSJ2/kRmGFq9eMozbaCTzh8T637Ad1Vc1HFZXwn/cZIhYAQ
oBpERPX5AJMn0AlPZjDhKreKRytKNIafedYXR+d8XWAs4l62ktI7Fq8Sbvpe8Njo
CQUI8Aoqr+ZXeS1Pyq3q0Q6FsfVqUF8Zup3ldMeuUD1KUjpgy+V52SeBibCOunLM
WFg7DlPNtjQm/WmsWI5sWtfEML17evfxJBpXMxh3TJkMRnU8J7r33Iuj3u0gSWsA
b/TpcGWcekiCONlXuY9r6R7FPC+j9YPRIredwr3mSo3Rdzhvkg4Kvm0/FIgxxir4
hsRSFvQcyzs0j90k0TjUajNkw1qnffVDHH+4QRHVKFjw4wcEjDYNZkWhouDhST2c
lPeJzrQdev/iJa5ZgwN1ctrB8kUXsRfKuQVu5FQ5F/rhPwg0YGQsXJMOxffwmPM9
qNoAK/6WkwPXB/k66u4fJ2jptWE093PGfl3bkoh6CKoAEjZDEbn6EKExfEmQQmPc
rVFjm6sytnCYUvN2Uo4ek4OJcB52S/cGVQEmA4j3ST0TNOYRP5BcW9kd5Waedy8X
tcYysiTjrO7Zgw7XrduoXwrJHmE6jmeVr6sGQHqOoEYcPb/Qr3GrAp+55sm987It
1GEa+Q0KekDO7yZpzDRao1BI6LuQ/dJ1K/1llSoP71YBevBIASVA3E/WCbYHwpUS
i0b2LB4KD+8d+9dVbzmA/uMkbirg3qUGloL7JnbkM7bXbAGdhja5cJUW07Tq4r+1
2tYQfTxv8LAZJd5S1J38KLsclvVAUPu2peuRmla6p2atAHrBticgki8v4LVzcics
1m0bpYeEEPmWTsRGfrmlmIuMTGmqsJDRSaxtfV0o/ypag7Plfq6ZUHOXBJk3YzNM
HHjUns17ApJ3agR7EntJ30TDn2LHfGTn/ovnOIcllSsVulugTh93rq+ECRGUDD+K
1j1tzEy4uw9PyaRX8V1sJBGOeW2W4zhJdy8/2PVy1nFVJpgAc9I/xOj58F7KlFOO
Ldkx6FaZm4hD6f0T6srofya0Qlvr0szwQhmvDMUAlQRJsJV0ouZekyIN24pMbwV+
NBdiyr4ipJYESfaaERMXEg/aoTLeRn2NScgtumM62ZVWmnl6f0Gt+KRRO7UuDByL
yQjzQwNAubysR5oteidoejK1BmpbFaahomjiyfdtX0GgEwSH0FPYhtu9o5cil6wm
jlIjH9TCh4y696p/Lw+p0EzxMCNyYuiZvQ4WvpgiZ9Hq1GDNiF2uY8S35hdp0JC9
yKlwpobh+FetRE6PyOB1U8HTmhCZ6DBeW2+ZcfpmBHpPUlsmvpyG9G6ZIdiYDb5J
JeUbJ2n6EgLxwYJ+cCLun1JXK4tyWttDeSfe0TvpL6wIw4U3PbC6u9uFdf4nDR96
9EpJ7CiWdZC8FryHq+LV7l9S8tWhGiW09mi7m8Q5ad7Rrd2t4JpfPM7cxFqHNcFj
ZvG6Ob5NTCCW7ZBY1C/idz8+unBcf+dsinwG+a4NKqi7HsU7x0+UkpRBqlwphXYc
JY8t9sWamdecT1kg4/WHmi3v7p0rEZkXLGDwkOXOAKyns1PS41ZZcN0BtslyQ1b6
2PtEt+en/gYec1JnEjGBrZQpbrhLGzQtBy+WckExVzjz+nmtck+hYn60a/FHXScd
8J2HwbGa/8A9AhktRbQmofq1wI0bVvPCibQsoip8f9CnGPh8OWbMnkhTY39KcxhI
Varv2D6DII6P1KwpesBlambkF0Wl+yzf5RkyicpGBZE+Fh3BJ+gW9Xq0EWz5AgpT
fxW1jkbPB3O1fnEEIHhv2UMKkQTCom+ChB8ZvMqw0RB2f0qOzRx67xSCjGHKYkv4
YRIEXriByYhf2K3+8k4rbuCOtGiIfZlgF3k++ICiaf/WDNWdinlQ1lQK8mkDzgfX
sA+ToOuH+pxyQeujAOx5o/EXCKgBVUnd1+oET692Ab+5lQaewcFiJFL8bm98oPVR
S8K7cB7QVD8GC9Rl6IfejQcZinmEgb8WeY4PMwoJbIn6wpqmVZ54BkQph8e5hXR8
lZ+RaJoowgjaqc+f4nAgdhsaB3PGcNEKaz32WtDI1GOqF+PqglvVZzbGJjj4HsbG
4LrJjrcKBP0+kUl7DCvjBcLWwPD1bEAl0Lki8SlVrgApkVlXOFj2DT4KEsMz8AXc
bnJJSdY1tSoD2926UfhRPfzxlZ34NAeK5UFaSS7Q6JGWCTh9CPfwMtCbmotFVdfo
U9CRlVgHcf0Z1MVnfTnfBPa6TOtMkl6fZxprkkvMS+xLLpXPAi9pQOdQJTJluCfm
0r5izYzQWOgPLgUG8dOTt8eHp7QauNGTS6OEeH2XQs7ANtqdOSOOtGtuUQazaFys
fUxc43F3b26qBGm5T5RKMW/vIkSp2t1oEY5yGmVtKGSt8jLEiunN6aoLU71TY2LZ
96X2bHLVAhgb4hKzMCW54ui01M5lgHFZ2OrMgU09YNsOMzeMhk9ofU8k5mJDGPpm
JP7PWxhYLDweN1Ujbyw5RkHpOZ7qXqITATywrGZpa4oip95GA9fCxz5BNKuQxUsi
XREECcQZcgeo2u8DvQtzhdI3Grc7jRtyti6pnIhfqy00reArtCkJFgeO3sPSeZyL
4JCbQnRR8gLtGWZ3A4XwSq/ov704oUzg/yqvjLQDZpIYMpk/QpNLiz2+YP5mml4y
cyKs0ZHJo9LI9qT10b/kBHK0wXPYBXBYk/Ywd5JC67S4q0MtL94NJkIl8dMzYN8V
UWLjDtRengWRYjgNNsN400C06Qa4Xaz6PdOdIZ5Eqzi8sj/YrurvrJAati2ewExY
RoZBl+JV5tzMwZNWPl9jOUNXjNDrhshO8y2HCyvwq+2CFh4A1X5QqtipYaJCdu4F
Ed7gl/9HwYFQkS8pPbDgVgaqhxXumDzcoIQFi9NX8gdqkI/Hu2pWUe1i/d6t8Sc0
`protect end_protected
