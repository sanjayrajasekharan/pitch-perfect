-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TLsdEhtMiNDDp2tF5VW7WOu8k76gABKHzd0FicLS5AYJxP313rcZPDzaL8L52QknxvG66f8B/Jrd
VmLfhhEXE5l70xuVDF9srMAX5dRLzlz3mwB6asIG5ajUsX0NbAKucOUDGIQDJdoy4QK1c5ByjeyB
Zo4BryuzkHpMebwwpZ3IBALlRmOhduw4YY8Am+uU0TNd5oy9DgfAUSeuduIkWd0WWgJMFwS8cJ6e
Q/j9FVeKewRXdT6c609tX69toO8xW0+/Mx+/KUfEX2Y73zpsuc/iYKdLZBUD5E3ibJF+ggZJsTmE
QWAinf6bOT5txxQsx/7yW1qUtnjWJajOq4OkmQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18320)
`protect data_block
cPdVp3t1Am9epxp9kVf4YKYg+YRaJh2FfgmFykU96PRWO97ikp6yuuiNn150qgNY1U2IGA4bbVOt
wAkHTdyX36N6H6uZ3HFBAoNBTPhbd+Dd+QSqGtheo9lgzD/gmlyNFn4xOdniP5i0PtjzUR9me1R1
x5BzBEWpEcFL0kRiRZ/v0ZtOYnVwR7dJettBI0DVRfiSKggIBMSCVatjk+3GrPjYZZxZRMgK3xST
XwR+p98PAsO5WDCuVjByuKuzQFauXHt0Fyr7DlY62+Kv2Kl3vpCHjHNmebNIB1Vb/hMnRngWdYVc
irX+DnZy0Fv/C/o+vdhWdxOWgguK5a82NaeLQy9Hhl71IvaobqTrzwsxDhK9r0vmk6ImD9Y5qdEY
X86VjMmcV63hTsiu/hlJaPtF4tSTmjNPrJsYJDlIxWVdHE1urjE3+05Taec4R2EJj+xGlaNHmUx7
YTr/lgkl2y6Un6QcqrWFL6R6mkYga7ydyFIjx5pIXCedqjketzQXHaaslXum9WNrl4ZneJmZNvOU
Tdj2F3Q3nDxPT9uWNTi3mOUmBTeT3mv/68D2ELagmLnAkY+9poCWsBYz16Mk7NccjKUmCjjgr180
nHeRrGzDkFWf0F5Bn89bKqMb2gcL9hlKdqmhf6nlNdcrgGSXQhrEMXvqMZTnkBK6a7pQlA4MIOLc
/cwi3SiHJgeByx6RjcfhI5Io1/ZROWgOsD7UI/ONQgSWEqe9gTeLeL4DVMIg64a6deZEz26ZK9U3
jZz6w1IK4m7xpsSAtAQ2Qsv4ovHDN/ZApAJhkff4vbrGjkLoQ1/OLdv0yFQ7L6/urrBbzsjmA9gT
e1CYocpW7PjU8MDv3FwRT0XW0qQdFFbCJ4AkNvhQYEnhqBcErIi83gB/3mxsCBACmQuS83uVjYPU
Tk10VxUyDsC4XfWQ2yYuxdRCTG/z9BpfCz6tgX8YNmWHB8M4NkTCYH2lUN0oE9bUfoELQvxPU4qR
9ehtIniu4nK2TMvCgEozll+TY/YOmMZv/PW8TB6oUDwf6dhQ9R+89d8GZviQeKcXfUjgIOzcA3yb
qb6xJJTxBKo3xkI97NtaHgG6cI/UXEjcT2LQ16RKuCCs0/fA1RamkxLY0M6rI/XaI4ZVn+psc5wa
y9SkQn/nz1nWpLLsU7qjOFozJDGiUWkndgA1FQPavBES6IOjHKsOUYLcIv5jjLz4JJmXszSpmPyr
dlw9kiTHZ1wQzuoU8A0nmivEdUfBOG4YIvNohZFPPeerCBk7BHry1Kb0YH/6DrjEeK9v4Q8Vdbds
OjaVp7fyFx9FRzXcAROU7UBJ+7CQFFnd2Rodz2IiiG2ZU8uZbS9Nsjf9wztEpOKc0hizMEbTYeW6
gb80nEFJ7rqRbGZ9sX/TFimvXc4mqkIWY1fHHdfUTRQwx5KFto6YEfMfAbGGjN/GME8Jv1AjIDJa
jlYd0CgyvXZfVpMrzidjaBS9IWGefu27FhzPwsBIgB/fmJUzhAiSr346Kt8WeJ3eJUi/H/qc4pzY
h9V23YF2edP/6w8BHZnK5ocI5712QpGT2d1rmlvfrL0a0uu4LTmSC1GY+VZZJIObOccLu3ZC4ozO
e1Fm7cTf6vesqpMPU9SEuT3kdXmb7TDQMKQT0tjmfJpSl66yjhlO307L+DHpxOdwLhSj1LhMzy7Y
fi/zfU7eSaa3sGeY6H5StEhqaa0a+xEhxyB0l00BEOezbFnbxaRcYQZDA/lVvJy7X04GsXp+6fAj
2gWXRvk0akVEQnfYU1L7yJVqIhgV2YLc+KaCYlzoJAJjOa01eLQwzA09J3juiOZZyYtx4ge61pdA
mVIuU1gxnrYgfYYlCWY5Jd3qMTm4kpcJOvWbJ5a6EfCP0GehbO4a0ugdF0wGaA9FS9QiaCklAruO
HxLMjdJIL7oRuMddeKvrYt8d9ttHppsQdTls+MwuUdGA3rr26okQpnz35VK23aE3Wqrr0LXbZoqH
SoOJOW5KxD/rOB9fCUD+xEsYqsdwy8aNEEvELsBJdpadCy709QZTQbgXjWUMgfCuOeG85VO25frM
GpSBMg4LVw6fwbJFgvejqUMu9EjPKHHgWqquUP2Wxlm+nIuqdWXksPY+YdCPunahd/ala4Q2B0B9
8eE5FJcvklKvgszAcAEYwHzlMo9xM2IMC1+NAU5hgBOnOgn0X7Zs1jUFyTlOfrYigyzufQjWZYaJ
7WZlp7LJpEcn8VjgbJQCGONXxcIhU9P1XuYxvzYw5Q97I8JbNi2xKbe9ZRQV5Wog7j0fckS2snx1
bAEBuuyfMvmxHsP2ohACyHELGl2fX0A3HtApMwd4cpdY+uYWdnbX1+z8hN0QUG907Wl6/fs23b+X
GOMvY5qLc8yZJ7Xyu7aEQDT09klQYFUMxOKa3BFA4/tAVf+WElpR78h02k//Jc3IO5/px1iLZvDH
4KLgvQJhhR8+BxC6Sw+zG+YzpwZm4Nf184w0OUmK7jr5NwfYQjocQ2rEWutEAZQM8Sc35h22mMPW
sj7Mb78qTSqYCy3K4ge3GrMeA2PbvI2MI7jYNybw8bzquy9fLmqBwAJhd13/91+s1XgCSauVygTI
wSPDCZIFTQ++b1QQbokxnOQR+da30ee0zBUttyK8oZdD++8VHJ8UCgLqZb0MZUKUaXs6VBfp29sE
lya+Kc+ZrzGqOApzBIANCm0+pUXWjsi7NFPhQY9LePfj5iqUo6T2lznfMxh7mupQPuKPWZhaq0+5
tgMss2lUeHtkoIQ3AmGH/tSFFNcg5Xx+FhT4UxoDekLckc6yP/wyb58WZrH0lhrR/G/TR4FD+L8G
r7S5Gt0PWZUpmov3JMCsg/VMdeUCayKW0xrX2lwkKhWsQ/IpCM0ffjtD5HRRVKmMT4nVq6qHpNg3
R3Lrp8ECutzN/Pnu1kx8l1d1w2MEGbLRME1MJYtqgGD77JieimNSCtJLCnxrlxS++NtGVcJxhgap
xr1rSgxT+jgDi9ohqR1aOyXY4KwVitC5i1nQeQ+mLcwWy2QQn2p0AN2gMUFJdK47IrQVs19pGcP/
ukor9D0Ij7GQhAvM+Du2e753pVVYJCMAEOkKcdfXbCT9X+UJnOEQMXC78MAjZprR2PgcHgnPZqt3
72J80yVrvzUu3Jd04Z7kWTV/2aNvPRIfKUDDV0xD3TnZlloySkaUJ1/PIBDj/WhhkOcbHNjMiT6v
4hU8URuVIEN9IrUjYJbWH6HZSeJbyYcQeyPMp5BoNxxuqQwRuupshQ2fmXWcgRQm7OP08WnQCEip
B0n91d+dEfcjrnct8TGJHJaH2KY2Zptb/sXUe2Zmd2EBDOxhzUhBlAEEtFdZQvbe6UUfFFDFM/IN
AkSAPnQ26MEuu9pUBRwkaaRS4tsT1VhJ+2estd6Wqk1ZSh1ASt7i9y547meHoD5biflkywa7QAME
9vhlFcRHrGSVhIh/9CM6dYHx8cOuaLYGHwdhhxbPARhNhdzGyDS8X57OsbqR4V5FuRrNrzNcZMnL
m48ynkKUBJJslVNFJb6Q7+QBlSLzEhtD3Gy6cD7dpOLhlS7SAH6RNqgNrzR1dOQoZffx12ma9BGg
4txyoYte8BARCdjDamQtrqmQxyyZ598zUiTt/wDmJW/Dx1/DLYy6QywCoazSt8cZQjb34Fu7t5v4
v1DgQs6WTl573kdq0E3SSXbwPpJ+benxlmndbSoqUL5QYVMtI/RRPfxZrii8PilRyiruj/pAanaq
r54RNSOn8WlCic2NZwL0/1vWzxdIYVh0o1GE3znriH22ZZ7GI4sa4sS4Y5jIlNKlSfj8rM1ove5u
8xvL2dQMPRmKRfMCvZ21kDZJZF2DvXb8pomIpG4c8ChMia3wM0BF0bpCrJi+9edXq/L9jBoQ+6u0
4XTqZiSimwbVK2tGfd7CgTAkvBmjfwUU06VpaY5GhKqUyXFHFWNlF8xrqz+SR5FzjzXzDOhCQzvv
U7EYBSX9NpRzI232x8s+D7+FNho+SB018Ukb9aTrkmOOSNwuWGohsv0n5S2kFYK9Wv4RrdWKVUxU
Flh+t7OI23y/H3xM7Vw0DnxLBPTz+uaG7uALraykRKs/XWOfLlWy1RZX3IfKHlOGLsHM7esdZRoe
sikJKUeno2VoYTV1FcQcH1O35jdXyxf6lcZx2DndvZzc8W9lTwlmzlhjrIC6SQ0543L5HadUkTmg
TvnRxT13xLBItT0btyemu/knsuKT3Od97YFDl4GvTasfelXzAq06dK+oJNxRa6sD5GhAdakBOmYt
p1xtteabNRkjIeJLaQbtn2Uff+8Ldmh6irYYaAwd2YAnRMwZaWFDJkH4fVgps/80FkLUr9AoECF0
xiPsxeYhfwoRNi1YOwC9GKPlmjuwnepI0VXNPnjLuU6pCspjL4+UgwQhnSgXl1wlzkdHft/BUnIH
etqiMyAoDGXkRRbBpe4yIHLRXmgIA3mXbC/Qbr0saKM2Big3Bpr9e8aXJvwu89BQxU/2+UXnxkXg
sGLAk54RtDMeJA5+iwdgaM/2CbZIhCCDPyOA6psCn9a9uXIECSZ2Q/+ehWQDBkLsSCHW/U0kuMyD
wptafe4mhUKQBSDRTYl7iofrMynHREIDJUlBofCX0LZ6YWsUCFgSZeWZO4j9K9N4pSS5jtNAJlDU
JZck/5PvP7IEkq9vSSx3tD6mgBuzKd/kxXhiu/oMHBqKllhpxJgu74M1xwW3AiUzh1ppisAiAX8a
AZ5iF7ysp5Xa9mTp7u6Ozx7dSObr5VH5GVsdNKbeIAGHbd27DboqIn5wG9hAYj6ZnT/NaE7n5yn6
XhUw6L7R2tyPaFtf4C9qoJuDg5iwo8gdiJwl3khnwTlsKR8AyUgdw3eL9nuoh2FejmjQfoUahToR
8L9dz3LDv3tYlnBjrxfzvP64DvxxbW0kg3CElqSSeOzEFl5FP0x82UPztcnX5L2h1j1Iik9lJu7U
Z6pc2wIjhJhO+t5vwsaipqF/FkIKdvLBYHKDRuIIHxsstakwHk8kxBa2DGZNeYLeuodjl1W7Bupa
idCK3vlUsRX/IwWgxtNZdstn0tPkm3NBxLMKfUMfuhiCTzgEyScvdRhjf6cq3wMhNol6nNHs7hBc
aeJklFVSpd7k71OQjzvAQv4MM80LZPZOGCzmfuJxjMYw477IRrmfKGZOQZAVUB9Rc/qi7Dzm3MX6
pJukc/nKBbTbaW93hYA6pL7B1GFDVFbWlqGFk/xiPanknBUP2jz7q82uJfzS1ALkWa5NlNTttmRr
3KxW/iOKI269pKuDG4QL8qhx4bjVkATkVlkzZ8ym6970nXvr3rIdKqF9eEYpD70ywIUJAZPEUvW0
BrXIVsRFL7SeVZZB2vAQy+Wmchi2x6KnMiQHxpT9GltAaI8StpkJRtEOwLKW2ARIuPzQ1nCJk21f
3xLxOQY/j+EanJPyO9vK86OjOtXP156MPLvQ1AvkiFFQ+xf1cwKC86pP4vdPhcfv9az9nwLoKsuq
9F6FKS0YX4nNXsgPAlRv23Y4iBlg2/T72/qHcxyljjf0J4pKtG2zFZq2VERHONPC2dfHjus25XXU
tPVYm/p0rZ9wXFstsLHK+LoEavvu1HhjU9z8y4eIM/8Zl9m+Zz+y4PFctNX74bX11aCJKWtmqLUB
645KdU5fZs4bLv78tkro18SngUP6NY12u+qvBDlhTQBQFmKXzYdk/pTPpyT9zroOFMyWQOGOSJl/
YBbCtieJ6LLPMorWlIaxk5Gdc977kvGwa/7ZPaL6GHO4MZkeV00VZYVVsJ8J1YzySxQdatCY774l
x9nQGHyYm9J2xLrdy5GxJ7r5SpMW9a22mYzg9atZh+YQ0OlgKZ8x5qeiQj+VuukrtfKHa+e4uxxK
CYS09fPnnE18DEV2h0G2sVxy4EJL5aDziNtr88ZpP2qzOT4GbUGbcSxXYCoij7cBPspOJhFizeuf
AjU6/nsix7gXdGzubrrBSadLLJ2P+mchOCZFEfCtlgoqKROIO6q5WcrdmzYR0+/TVq9ofIwNIkBu
lwywRprLxILocooq/0TSVa1gc+h64HJ9+UJ+rPhRS3o9keaVe7+7daZsr1waR4wRrB/Biz0BAyvE
dCStZTcfA3eBIWWA6Hkp90HEVLdY5YDxDwClFGdvK9NpAl2Pxb4x/LSDqxdp7VqlYVe0gwBQ0zeb
l1rrfVvI32gcx9aHsbhjLYuVxIOeOx/qmFHveiovg97HgwR45916sbz3QkMe5ir5WuumGUIvkvad
MpzU5tOYv/tIyMnVpnnCx1P200BBAKMR7v6NvwvMZDlMg9zkAi4LYX1zWIKp/XdDF+a03ethdCfB
AcfsTPWC7Vew5SDidiK34ncRoizHzH1A+ohxCVWtRnfDKZU6U2Ddp6lR3Ir24MkxGzgnaIjBwQzO
1GCGunZ8pNBM9JZojHbLE/u/OCQC63UHkFpj+sqhOaVS1rYp33Yyr9THMd0TzT4n9eMCDnRptQy6
/oD4lAfIoZTqr6ufo41FBP6G1dVxZXuGxZl8N4405peUZXJD9ih0SM7Ry7qI3W03u9a2fpgjAPAf
STyTEgy8z4mJz3yGNn17mzayplEZrgbqhr4qxAdWv2ue/6G0jYjQJzCzVqiLKSyYmsv3d92bFSVU
VsO69QzfUHDTArNtzEel5clfbXl/PR2IBY+8ZeUC9xSmlOADbL200v2vEEhvaQ5wOmSNmHlz2fUD
ZDLyZnjIlCE1WLGcKJLyCltMipIG76tmcs+0cM/UTsfTllaZnHRlnRU7ldJkZDYdbi0xvuoFOGsk
B6Y3IwxiNkAGdq6juRVY0CwJek+6O+W+4FUVeZtydwHBq/bwlMJVRAlSAq/YfOXAFscyjVcZH61V
bmKKxYSmoyAVjKEQ/K5hnxCiL3m2Bx+cbi8IzOBQ01Iry9P2TXL7f3bzMtAwdIB7z3eNR6AUBrF8
PqCIE1wjmR8RmdTQT/LHL9LlNtFEKxET1raKodNxxFOWFpOeSCcuARj6RBQ0aHhQ3Rn0+13dK/ma
CbfLfd9I0xeXIg5qQ7FxKEUV5N3lePYAl4anA2XqUvZ5JPRYSGHDPxgoLLbSCvDECqag1QIAznGE
+drtBleL4KiyJFRbeq7TsDagz5uRopqm6V2WGZJtc3Nepsc3i8Ny14A83XOKfqC0HzgrhKoFvjBM
01QvFTklRyo8anmmeVNsDdmv4PgxmwBwP76mWLrI5tKR9SveI8ayzrQk3bMLnXmi7ZgHqa5nUbM2
4rHSaEFYv4L6ppm20T82Wn8GPnVAPkq2zsM+UHvwr1LsOaZuQlVgs1erNJvfiBspi+1w8H/b6y/l
2b3B9WhMhpmqAv/ea4UNtu7tWfVG0FfAVkn5yUjt6VdlrIinallFzFm0Y+32cNeOkWAG91+WxXBF
qEuzafUoKFUsT0BvULjOPskMV8EbvXHg15Je5iW9y+WA/XBTF3FveYamg+vh75/FbJ7lc0Kk8YoI
gb+gKBOWDYOdNRsuUIhpF3AVFpH6VyjXdQujhW1ip00b/f2Ou+EXSmVF6wIh5LyLnHfac5pEwzhG
WfS7/5YuK4ielhdBD+EblMivJP/MxdINiZIKFyIhbpPNJnteHeyCIQcbwaknb2oLZgE9nlmLMBkr
d8St+jk7JP7YeAc1hk2Xr9N07OoMbSLThk6Sao81ppBV85w0JNwVtrnIBx27gi7G18yuSk5rDQRd
4+Zu3hCdHPJYQRtuea7OCT4bfJnKVb2bO6cjgq2m3tQWOC95o3qDhec1mF4UQqWVVi64R5UrYiJ2
6B6FDLVKfGnyr9wrO18XX4MO+rn+btzxe2Xd9sh/XujKAOybQ/7Xz/XIeyNACpGGgPF2zURWHB0A
dDVXBmQ+XbKjzJmRn5Kz0mqVAVeLAUd0I2z/LE7aDnxCUYpMhsQvj5JOgJ+iOQdi8UGTf/Tk4iRJ
U+QhUk+zPSukev4VAHm3l8NonIF0aijR7GBJbheu0gd48sIBTIHKv74jn2nQyN4WmOLzQa7yaOU8
M/hcp/rfTWySCohR5FmF94D0TNQ/oInfyZuYaxZ+zAe1WHlY0NKdVVicthPckVvUyoahxLcYca/1
n4vP89onpL81dUJjrnBIzK0VTrBlEsPFucx6V65lHT02YwADS4UKglPOX0HGJrfuwm2fepGwdE2T
/rFJha8ZJ0BtKe6ZRgUnUxlw9NGK+SrGlXilDb2wjvj6ghANFBcKp0t4rfDhtTmmdn6n1AP4OlgO
AV2FhhAm9g+18EepISuINOiy/xTNvvsalUpolYucrVHnhLg65rHufQVOWvClLl3xbxjKHTHSMALs
IiL0qduy8uzq87EVxrQxGoM7OE8xR8os8FkyXVNRMD4JlqhcNeYAJJsOi+FoCKDabUWrNtYDjONn
lTNFK/uDAKa/L2Gatr3z0Z+z/NGVSUFl124OQTbOtoTBRaArDQ+CMTSynTsujQx6RYcgs0h/5g9F
ZJD90IggNJhZbqYgwJafwPknLm33fi5AYqap/Xs9JD9b3g1bMg2IGbCL8qYRE0HuqyZq9dW4X5tN
vtEBCp/xQVlgoqNookIZOw+NOaBnMQYmMA5/VEc3dJAj65ZdnW1AefMalyD2Gdk2zPRkbc7tC+XF
zuEJTsn8WFqMUazzCdKH8xTspvZt9WfeABlTXP8Zu8Z3a75+nh4kqxevVXfb7FH0n7vkJyZdQCUf
XzrogAOuiiCYEvwkKMmcaF8qCzhnq99nYujQb2fL3qnmm69V3UpSLystayjISjCxuGza3WBWLFRE
Ii4iFTg9TIHkU2gRE/+J6ZMFGXweipKl3qS4rOk/Wgudcwmh+gRH+HTV++nSfp9QvbAlJSgDW8vK
c5Azk0+QyCEXg9WV1qHBMp4TOopk4lI2CI58xYdtQWQIZNpGtpCswUgShuTWP/LWOHpUAIAuM6Cy
jkQzi5zuPA9IE3t5kBdPEeItOWVk+LcXzTSdQT9EBhRcWu0Ak6Dp6vWZIBiSzNGEfWgJPOi74TH9
00ktt5Ln7RN7AxTBPrMSi5+u0jUuP4KRAQBnO1A3vfJFeiRfa2iaclMG/sOrM80r3rjbSurVqptp
2ujX6ZHtiqqPrQhdadBk5XxAtDo9yNTGtjPdNG6nbjNf6Haq4LPmRP5yE9+JQFgDGKZHM6PI+yZK
c9AZqSfO8+LqeNEVV2WZ2HmIw+aaRrwXxZbVtp6MhIS15FQ/GEggPVlXyghE/ZGqd65G8iC3Lttc
1N6gQ/I6Xgj+Aaqw41CDlsEGLcBZZofh+mlKLM1HuM0Tq+AXP0sZUZ9D14iG9tq72n5KJToBqSiF
vNacKx+CUsbAzhcHc45QyuTMqtj/nl9AKEfi3r4E3JtsTDpJqFczNuAqNux6XBXyWZGW7U++kJT8
Umn07Koc5au0KGu/7dJE2fF7aZFsybGFdwSUmyuNraj4t2yCm68HYuLbg3mJ28auLKcNSrDfHI0l
NlcutIRt0hM+itzoKPbVXWSfaKQOygu1/c5jFQn+4jvlUEXhwViNem4lVPHx3UZcdGk1cN+86uay
sLQfm/934XCaiqK7R3BoY+keifGgLXqTqtU4ik4DOszF/U0rzq6PrtYuH+Yj9HpaGpUa5I7fLT6m
E2/UkKf3rtVxltE1eo4fl2x02uVFsHcYKNBfs6jwOrqtf5g57K6RvjkeK+KP2HWTPvRfEM8rsbUp
Sk8jwOgVkl6euUG3KIFBzSPh68orE6lvEIR8oFQP7tbchpX4sSfwm0P9EdrYHlwQD+yUExtUR3pK
Sa/s1gfZlfUR67l7LYafWTXmgY110McwBSumfwAD0PXS8nDQOZzJNI/Uify2YxlWjzISmOeGEdtQ
DaTx29BLpbMEJaTOcD4a2CFxp66ULTGZe9eJfz0/QPTP8tig5RRcAoE3Ls9O5bq0jk2HZs2dNOTk
5hDOR6283LLNMDSP53J/yhJ89XWyq2cG8/ntI+4RhWDTPXtrd9WlUFdX2S/NPZHFh+OpbgmEB1xN
Fy+FDFmsKPvR4kfau0Ggk8A2R/dsBTCowd2VLqhfbLMo8EhMJ5ruvTXuBtmXlOBkY2Qi42LRCZfn
nFjQbcHatX+7sccuMkcNYp/PMtIpQGzqk8K/Ij6AeZBIvjO2aSaNN8TOWiQoXsc/xHCdmpeSVRNx
8PIZYmbwHKZrRrV7hzHO8aO0N9dRYU7sO5UTqpNm6gSakREsbd36cC21uWYVO9pEUu6utt44QyI3
tI5MZUs+VNPg6ux5a7Tn9pB+0X1SqMGujML0iYWm/3YBkrExnJYFUFfgTNEiRyb2G03XHoGN0FCU
NO9Ejhlru3LYYZ2lfJF68jHp8a7LURpwTxbo1O4O6PnWCRahCedOPid8vpTbaKqKZO5KVCj+Vpf8
5yNJLUuahY4CPsPUDhiiizHXKTpLx5Z27XW4fcB/le6njr+bkM0N0d/5wGAaN8srHrGgwicO7ap+
+z3ZibomS3QHGtMiJdqCLCUEeZ4SmocwLKxKydYj+Xq1+scIklA+/tzEVUPvqMIs5VwiLnmYn+6w
29LzMwvu7QLwEOcGT4LCN73b9e7cQfWD3czqYz0nF5sVlvoi3Bwu+zj/zzR0Va8M4J1vzSvAtFOa
YEu9ub/wu8Dd0vr423KZw8EmiFSsYjm9KHaOZZ5YvxoY00Ucdl8mUehOJQTu00RGwnEushOVoqJH
RMMKb6UaoZVMHOWhxLq+wSBouPThwQfOdWGb2wuJupeGv+n9eHeUCNZBjEmTfVdEDROk7aChRi6B
ot0ez0QbQNtPjrod5Hik9MfaeDV8/GvWWechoGrajTdZHEW4upoK2tPLigDmlHphVi840iR6rI/K
fQVnb7elqoLFbdiVg4GEsmf/QJQLWGxTWkK9XmuAlhTYXzwJ5OYShbaK8uHx9itpR3NTqCWiAYRl
T9RhQQOVlAJCnCgjDVMr0umSONCkdnTPzW/OBmdTWrRbOQCTQNtJAYzvgZgiEHTtr//MtKoa53mp
jeORiSpOoEZiDLrM5c3cNboitAa2gHg1QLpq+px4T9Sfr8gWon1W7k5WWLfULQdDQfzuA6IbJKCx
bc3KawveR0pLTAocpx2ur7wzb7o4e5qEVYFJ06jgoRadU7WJ6cC2vDpq3VU1bEln7P0v4+w3DTto
aJH9pFVSyf28PczdoyWTIjMbtyWHMn/NmXaCOyK+mpcQMK0ollOT2bouN5JU5Qv+m+igS4JMuvn6
f893O7EP+i4wd2UyjVJwIPVU+fnnYilAqcHLsK5h6BGTCPirs8vI/hPGDHhcB2IkDYI4Ysm3hRxD
bB/Ow2Vpa3b6+VIFq2BLAovQZXfJ/SK4/eN4AEAaaGWnF4c74Of8WDnLyuML8gc9EuT/kHUJHsro
PvQZ6ppE6R3l1zLa0udHIN/7PxozQoC+zHklf2hbh8cp4smPuIAcyBOvT94ZG+ZAHMwLcsNZZ5TF
tavIZccAUHz9HbIolLFF7Kb838gzZ81ogOAKsCjUlzWj/ZrssSeNHwHrTq+B86YLXV9KhJLNwr76
U70P9lKFnSC1X+0kRn8rBPO37Hu6EYYTBqE9MvFmDqCAQNVS5K4m6pnS3PO0tnHViWr/yqKviMEC
XTADzgnbfAYuzk6mTo16MD46DLGh8lpvyO9vJ17lXrSXOPsta2JXmmiOG4enHdTsEtevAgUO0Wu8
FgoN/VzK2xt0elEFLYVGNhBW39sh7MDt4x2/K268PKtN2Gdnyb9nqYo5YgTaO8wX+xqsMlcREoZC
WGVbpDv4nCdgjgWibXHrXLowBZgki4jeZpHqlaE2NdEE8uL7mc9wBbTSWLN1C+J/dfGlYCK0ywVE
MGIPpK8RT2X0CDO1XSKHLOlgeDPDnV3/dRK2pUnSzlXw6efxsPhV/rcQqRuGJJ2GDczKhkyXnZBO
Wiw8/hHS5Yji22MWnkb3hkGukrWb134siDMBQB01xA71qLt7xaaCp/3D86lgPsMlgvn0xOy4pOwd
ZVM2n953ygebR2/TQ9bK3oJKBftum7KQv2bPExmPThchs1FpsTMBknQkr4TOXrvjQV/0TchPbenF
MKnEmApkINJPVqQEg59Q3MvaQZMaGZHMRdXfKnijVt06VqE1kojRLcWcko24jOoh3PHcQq40w0ce
tLVwAsGafOeP0/pZzk2tM2NOh6uCk10iOSpk1XthDBDiUQuAsOp4lwNATyHxKyoXHIDcOwwiVkqR
1e37zzaVIEs/714YgNwF9AaJR2tKfNNNzXHVwUikd+NafeE7gnKSqJbxD2ERC0xnbP6rVCHv8urR
mL3dMXsf+zWD1ofpBTrkFwKeWrZCto4JHl4CexjjPrBgjCGcJXZO7MqRtSfptvM9G/Vr2PaPpv4X
wWmnyYhYhNqsBrUr3xXNokOELi93xW7OHMutnVHps/M14UoWR+Fy9IJHfjROeXMSgUeSsmWLMWuK
vbqCQHSMz6/AfaAklMv27m8ws1SM3nEquakOwDO9VpAaiohcLS68jnzAOstIPvN1qlQ1O7pR3Pyp
fhDow7xDyAARW79mowAMzjdk/psXJDjzXU/OK1c+OzaSZEWoiJw2JIvakb4z5x7agr+uWklpFp5Q
vTOoPe319U/0LRQUNHlgowmlAmZeW5EwPNS6dmB5uyNjnaFGrY/yK71mg/7xaWWk6Q23i3HY2Ydp
N7MrlZ0kFWa67EtgR6foGYf6xge6h4mL2dad9NX59MiLQvo4fCtCRsGJL3+oYzXasl6c45aSu5eV
rmXEEmhef5WzlZMOAQ/oa31LYhryR1L8Byl4GSdso1WfbUZbYMbb8diVqe+CPTppDBrWlJnkHvgJ
F9K+Rorszqx9mEPP+OX9KQ8RiI6mlOjLGXqp3dtmXVANTAPDe9mnAX+ld5pjOJCVaTl1LBeDg1pk
emOT0ZHBPZcov+bJKPlM5aS+sMo5IpBhtEl3Tkk0nhhOuHVrIPgAadkNzMwkPxYP4epcmWDqHiUj
ZEtDsbOb5Sp5uQxw0P/4So3kayCkDBk+QmaLHSu1nrBs4XeCDncEkvhwsRFDjx8CaNnU0DQIhPIl
VHIJSGqLdq4v3p51jBX3zEERhr/nH4DZKUGal3WD2VSm35kzqgakF7To6mgCROssenSJb1HNpuVZ
A2fosbP4ICDh18QuHWo8lRC8pvY82H8NoYV98l4K2mTM2mPHbbPunzuYRaoFCo36qKEKnmO8fpuk
XhTu03zin2WFqjbVI3iZE5UaDCZxdMB0yMjCG9Bg4kHTd/O4PZrcUMvU1K+aU3h9kQJQXk8jVHu4
Uxvnkw+y4m9BdhUq5bpKk3SY1P/gEm5igC0Cd8tCjZQYr1md4NrjLroxm8RfRkKRjJbDZjWpUUR4
7YA3VsJNWcP4J+xXq7MppjM2p339lz9Nl4r7Bp6WvUyYaOtSQJVLwImHAXaWttGsNZqIjsx3QxTU
+6K8dlJbUcIALVP1YVdnXwXhjjpdiWNKyddhpzFrU2ag4NLXpVdUncElbbbMYzUSkqnkSsSiXjtj
NlIyr2N7EL2oIitdlUz6I9DTB41dSR/3vmzdwpo+mFLabihx/y6J/Ko+YLBhGHewm9iRujzxwlOT
/fAXNSq/5TceS0FLqNSY7ZGmdY1mGfBOlatY+9DFjmZWw0yjjQn+HKrTtJeTrnU8oivyblEWKfZU
o6nlgOU4Hcj1JqADMPuecOSXWigxtRTsdpFZGs9W9EG5HYoOYkvxtEukJO43BrlI2dF1lM/kBaG4
1n1PEaGhUSTyBwmMpCtGcCyBN4tDfFQAuwuHg5V6GYncL5r2S5BgZ47D2bd6F+4FMhVNhblyUX1n
6bWJPCZXUa9/892dyBsUPBFhz1izpy9zKsCw3hp/PBzBs9+qjl4D1o/61ThtKDp8Z7ScTh7c49lG
EW1II9X4N8mJG8uSseFTY9XiAKCzdksbnIxRr+sCGUDyxPzKhfkFWSuIXoWO4rl0v+Bs322nFQam
ejzsBxd7hCJYGBVF3aODrF9OAtA2451FZuMLfOqfzTbP30/IaVo0Mq0BjBCGHUwxSBhOtHM0Us5y
FcCdsZgJsat7leajW666lLeQVkwWStrxJwHXjigluHxT4Et4AnJuxYNLwPWTVwdZ8dxO2+yKoi4+
xm+MYUW2zqd4/GqK6LLDpMWFclYYObOqEKUeJNzOk96qKiO52EGkUA5m8jcsWp5/b2XoywS95i4X
q6AxQLxPAksCw0ozpSCZLd9CZGy3t0BQZfmWCIy9dcry4WO62cZULYLVq2io5RD2jlh50BvLga25
GAuPUWkqlVLQ1j7e/YnEUo/LWCz993/2FQIoMA18gPepkxQbJZ3TY6+ZZ60xQXgPdfNgMi0tDHyC
sGy9Ui8pzurauzfIi492tB6h9Q+fOom2gcHak1Ftt5IU5ie1OxASPaT+BC9XgmHgjf5UHl9kr9R2
lgpbrPMHciyDKSBuzi4cMs0mJKWW2T9IXvtSvYDObWr1SicLP51xxAt2qFAVPQ6QQOhn/aqbVNX/
6BIjIxb/+FvYst8+KDshO8i4GJIkcM+fLkX/S+LJUU7aQYq5weTsAySPsyWGbYFqNZPqgRNK81jU
O4r4zrb+bXR3jLCRVnmx7l9Bu7MOtIz3Gy80BjvTFEtyUoYgac4QAv4OMdjpjHCxLEw9th+M4xIZ
EkSqoy5odOY3QfMcOjKfyfZhFDO6A4RcG0gIcECcakTUiXqCVSdsrAwP13BNGhUuT78shPGhVzhN
JQAGHRv2+/zKCmNj4n9fG/v9f4KtZU+VbkJ52Ak5ci2fKn4e8WvWv11unkUYBnv4gw20SIDfRvWI
8+4t1upZZoBdn8H3gsO+ctc1hyGsELRboJSP/rkFK/hPplJgTUikVw4W5BUZjfCOEgZ2geq/INMK
a8Du2A9js26MG6ReTc/8Wny+ViA2qYidpdEXbz1ivi5EetgZtTCFr/Z/RluqwP+DJ3Tp5ORHzPtf
Ptb7h9hLax5FgBBejgRK8nM/NkgzMpfIQ/tKULfDPcy7OlOhH944i8dmX+0cY9C4W32x5zIFO0wo
abnccOOk8ooJJR2iHw2jOxQsMLaXJEVQTOF6/DGxMLnA6CSxYEJxo8igD709BDh8mlucSpHCS0EI
nkKV1WLiJJYB2OpDdcgKAJvfl5ZhWPul/xNb43AX11uo/P4Rx0zxlgBElR4gWfdBlnvF5RMzvd70
vlcQRLCcaiD6kFfYqlOIxZfUF9umiezR1Sp43Z2303qqpnIVw9pYIOGC7ZOPIZnzsimGmLkObWSi
/gU6f3l3w5fLfI80vbi3vzYJX2NiXyh1Egv+UVHqhCiwrLbfDARi4xWlf/hQZtYvtYyvtiJ4WErP
BOxm1iZURknidUQCyGNsNUo031CPG/H7QYEnY8XdiHKMDs/zygI55xYutUIAuYpLYBhm4YPd4aKA
2UqSXymJGEbDy82HSorkncsfWusqFIHlG8jiqNv8kkjK/eDN4zYILSlvQWMZcj2tgwaofpVWMrsj
FSjH3RHD4ugoVL1I/tdi9dtczETSfBEh+PywIn5VCfMc61lkRYLIg+nvZTK6T54EPGZj3RpQppIH
lv2YRw7RTY8timrJr7co6iWUtsNW+KR7pZmAD+0dDRVmrofRxDxnmUQo/fDUByZ3IuLX5+nXsepj
BN1KlHA7L8pqtLtrbSJHjz8VgWDHSZtWnncpHDU8KMYgMS1P39Z+6Xx6AZ/otcn13OLwcglk6Wqb
vBSbPAQV3DI7exaD0qCrztIm8LWnZ+o+aB2J9DaDeqXh2B+prEdTbASFz12SwwAQy7oXX3hm+xYP
fY5qlZDI8NLU9rnuRlbcakY6WLJK9DY+T53Mi2b5EWxcXkiEnyOWBaB0B0iV//s0h/9u4S8stRXL
MI+1k2EOSeAwWYPQcj0CE5luT7Zcd3P0tAyz9E6sn93zri/RwjwkwWOA7JMk3zhx9r3CX0FaWdIC
Evj9HR6SZ5G6ZmeuXfu2Zx1wKQECIpyf6OqCCNcSNKr1YYuHih3Bk/mdG2Qvej4QiNK3xOWqGb4I
fnsJdSgxWxBa3boPgFry58hwGKnu8V5QoVaT1vR2B7PJHmeDgewIfTTVoq3hORLHz0SCRZu3EmYx
8D+eTc0RqTOnosgUuvUhtCks+LVLLdT50wxq/q9WMl7diMel234li8bkRFwvhsHF638tWUX3TpD7
kczsBNoUWO5Z2H3pswXDl4zVGU0k+4dHjTN3r6liSyCafS+gxxzLMiRrvtp04Ad99gexEn9A1nBf
8zjTwOXaJQpHEm3HdZ0yZTTxp7Ku0UoEyZmAe4pvhT4jOhxAPLUvnqtFkZC2hacqzfaIOVO25U0w
ADSUQBamYnJ599Ngp2Ayo+urKeoMwGZ/89g87EF8HamkYEL8EpfL8m/6OJcCp5l0aQspGuo/Gnf5
hYkee+GpbaSrK6ALL8bu3LWjOajRaWdWFFr18kDjc9XQwN6EPT1UgYR4KSYWhG9ttFp5DHZV/T7b
T+1Um1wJvDHSYSEpO2fSxA5cmGYtL1Bp8KTirWs28VXf42iepVjaNHKfbusjIekie8x3m9Rtol3R
qZdNGO3bJw0mOIeaZbY2ttkQ3lh2JavNcG42qxgpUxAO+UNvk7wnX8zrgTIIES1rpdmd1KztY8c5
E3h+vTXp902Duz2o/eczmZAzD5nAK7EIbyeXwuA/5dO72xUaOWdNgU6qsgaHvgRjlyZMN4e9S2LM
CoARmby9K+MCOpW9XNwp7MixEF/R/llDj21r9rNeoS7D91KlPVcWVx9NMpWTWpm9BQJL5H5vGV7X
yjmUM0fRgHPpDzTuImYt9d40kfqASFjbQLLnS7j43qk62jfeL7E7ygfA4XvpLJ7hms//9DuNh7Ad
0HGn7nMHfy3qiSBmAvLjT9nRIJj5mL9W31vWc3NZTDR6xWTvwGIpx7Fd8HF54aq0Z5gSW+8e17qO
rDkDH6RAwV3UhBbWhkL5lynaz6SXFeTwXvkmNCCTJLQjLl0wXcKtGB4Xym12Y+nMUoHXeQGCtcN4
ofVLRFrHdVMxjOImJPeMPhsbh1BLTJR8JANiHE9wBYpbrN2gid6jZvgD2jZMQmqlWlSdvc+lg/oz
z87JgsdKYrcceuWHgJBecVAyoccExuSZYKTFZozs7ed9+SZCDTr3PZ/TyPj9oxvUADWJ3CX/tbkk
Ev6Dw0/kZp65JBzVddcORcsYRsAZSqBKWqx3tF/NRxc43blf5fhtf3PLhJkIB2fvYMJ2uv1VTEIk
VsVKO2G4HhfL7LsiOSRvBo2tltQKEgORVFGZymKMFKDcZaHfYXQ/RWqB/lG3ZxT/fKyuJZbhV4Lj
g2xgnUhRftQnTAizGgnd0YKo55IQoFiXkuC5y7TrK5Y3cvBvDZP3si8IHp8alPl5vTOj9iFhT+U+
Ggr81vS6ddNuzEfQdCoknROxqvglIiK7AMR4fnujEnFJaHVc1+nUG7asg30UiMUOXpA1T/E4c3bo
lQ8iu7/peMq+JkmGMzT1XaZnX52CE5shve8lsJyb4du/UCd9PjM1/oA0KpKI3JvlPTJI1uJK0yyU
ibP18nSJNkhKK/ryLFPHcOf0lmfjgjMBI5a1MPuimVI8ivD6ADFgsMmeP2m5udw9aCMlnZB72bnN
8zdnCmBoeZl5ApJSn6+LeteusGjGN9XMHpMlmcisXKjvFOgnI8AERxEptz0WVU+feiCJ/S3E6t+J
UkfHYBc0o4RwRNyhDDe8CebgR+fDrv901Qn4UPvch+XB7pCrN+HIy1Jy/JKGEk9iD1tmrFU254XG
BGY193xp0weOsu9keEvS3Z1CT5cyx0pr+TQaRZaXZhU2LR449//LL+guir7t2xLr61W+WBX9a9Vz
GeXR/8FCwDzZTZE5Onpu3lmyE9rDbPa2qPe/htlRTEdGM9y7bUXHXVBqgc+5gQRrjNPt4fslnmmX
F6Bpep5umaxtgs2GxVyucsciePujRWvx7pGmbzV52xziPmvcoDLDCAbm0WH15LQ3XrdDZ9jJtU9g
z9k1kXoghJCp5FqLnHLilMNED6ASgedIHt5PPPdu+V4Hy+dj9mUQ2qOteQ4xLS6cCeq4LqeBzGZZ
SEOOPXgWolF7KwEsLuKsw6gupTc+DuB9+1YJI3oRCAx/yhyKTJKPCkcV437pMP+SWkxCEoed80Wv
0LLGtfogC8Fsiho9ahcBOc+0K1mfIyf66gDDsKE29u3uWa34LWX+301MAYPGgizuJk9vbVl44mpi
vAq+f/a8OF7xGRQ+zD/OkpAwM3328jqM5GKZpO8NN1yqDB7T3IhSWT8mFcqLVBFr8Jqlxg8kDMu1
9aZidPVUpaAppm+hvLl/pPcgXHH1qEQE4wj2BqQmnYEtUrk+G6sfltYkAn8bkxHEPO74rj1nf8Pm
osMBY8uCZi0ijV5PXCtUrr7T8+ML+ehQwW7a5Lqq4yi8jRjPidtwNB/lH0r+egY0V1CxWnyuarD0
uvnIYRauA3KCWyQR3ml+y4lQJHV3ElEuyJEZn521oJ90TQFNglbm23N/EqF+4ZF/dU77LmPLy3KM
UM1VwRlc4fWUsZowaigkYA6NisQf/9T5mg35kOHfSao9th4LqeK96/dZGEwUPrOJadcNbUoYndvR
1b0ff2OlClgyFq9i3h4bUmb0XI3wX+sdEpR7P8dKb4FllgvH63MfWL5gwFWDoNRNZ66SZj3olmwZ
6tD47GbjosjAc++hSfne65jXq2bgG75w+6Uml6Zkw3MwhUwduGPNG2HoIkOAq/mPeO/6jFS4hDtS
ocOVT1dErm92/9wrzg7nxPo8Vmh0RyRlxgBIJ4Jv4CXgWn2HylCWzfrACwoLcV4y6E8iZqIXbzQ9
U2Xdee9tytDedu+VBVIa1z+JeHwHZEenGoesOTE/y0Rx3gvABJcqxQ/tCAVFT47o9/TnjiOWt3ZL
QWzdYic9q0F8iqxvWsl6VqsEI8iTCBG64412aaPLNLjFH7odad5iTFX2isEgS/RYiKc7/gApeXcI
SqY00oKj4FynMSgLXoO47Kc1SPww50gMh7wDU+PQWan+R3aKuT3lfjvN+p+nvdTvfXEC68nce3Sf
VX1E0w3P3MN51RTR2dYAqNPWm6wBryZlBwXyPKTQIxrJgqWyPfANdf/bstKCk7uo3wn9RKlEQp50
5VswpC+sw+CNHB0UOH6TfTRPcuE5UOzERRyDWfIlfgLJARUMqHhNAr1Xp0FE7UcayfVedxj+zpk8
Kq9A/kPrM7ByhlA0iVwIC/+7Vh34RVnNwbSTtyg4AUwvDgIXRYvEGJdV8wkPUR6PoUBmQDwgqmKG
2s4pa7NJzJvprHN0e4gdAuDfrKDpeBDvvksNH8MozQhZQ4kKK9ZmMSG40sihcGkA+ks1pSDMxwTc
oklvuCCxWMPMDmlGoTD3GS4U2GdZB8wmC4EM/l5Ku1c0s3wOD6phCIhSGlC1ALr6ou196QkVR1da
wMZDvSUm+6dg+pNHFUt15Uo/rhLs+d3rkOx5xfegKeX6DRl/3VF5uAaNFgN1CXxY1WiO49CjSW67
YlYxt9wJJNJEZ5YDG/ifuQWeLfMm2qWt9czybyz++5jPPPmgnUbA998Zkeo3ZTfJIIILEOsWuM1C
gaxQRkmUjlmnwG39hrmJmOGmX/p510lZYEOUot/Goj1LqQIoEdUjkn5DRMIrLYdrAZ+KwpeOb0OS
PpAHIsqytgoPdh4MngHXXsNsOtGJFc5Mu4q6gGuPEN4JgumUaUt2Hw/CzKw6i2JgR9Mqtyef1qzp
Y0J+yVkdFzH+CDuBg403NZ1VN/bqoSJwnUr+8Rn/Z4aO/4FEjTgd5n3AFSjjzii0Cnlfu6oEmEG7
MwxuZUdXJxsXUYdzYqo97BZ+qZF4sr8Lno4rVad7iE+Xj29BFJa/PTtVKKHXnsydnN0b0bvsfR7K
jItBvxBTimNYKgHgvMPbOUL5IJeeyiRYWTdH0j2X62KQUNiM0wqAmEjvWrLEirpPDYMHPOH76Q/F
2nTo78B0OhcqIIm4eM9uIPIjLGsllZ+94aY3sq6aEFWSybAqC/rXq09uv4O1kq/n3wuQ7KvdZOZK
k3ckWsk6Knu2k5fHfKB9Woa7xbwZVToFNnjiCnGV+RrNFHxAsHx6M4qI/tS9I0SEUedQ9jAp3vzI
yyymGiGLp/BafQrdrkO9fyqh3toRmQwAXzBw9294dL4mzc4Yd7dxSTXsr45MoiTdg1Bkfxm3CwAi
1Ntq1ChuXiUjUi58ep5vJgWTLL6b0NUc6XG8OezVv1tl6YfamBnPiy6hulvHD+Es9YcGDftrq93f
+bFPXbssxoiBhLF2/vn5my29gF1+fx1FKPnIFP6RtWELdnwNX/vUbcESJhh6JEsPyOsFtsri0WCv
/Ox/3Pl53/g84GRwscuuBElEVMFJEF5z9jDPdXfR2uSHIF63XJE8gicHGUONW7SzqrP8twLpG09O
PUrx4GpdVRpQhL0JcKiKTE+GLPj7BkWZ0J7V9XjHl+P4HVZsIe9LzcIRxbGr7hShoV2JPqGYWTKo
41rn9J6kh+gPUxD03pHvMU1NQH2RBF9u7hrwT/E45rnYYtyZ/Ujc2E0HEnzEjaVfVWOE2o4f6w+f
5nUbSFwtImImTuMe8Karbf1crpkXPyL7P+2A9c/PtZqlPpOo9NxsJZATTNKhDbl1jO+0Z7Mm/trk
xuiHgTN7BSH2ygNY3dmg9WAY0ZfkN85Iut6cqJqbQx16tAGoOb/NLdOTjO0/okghNJ6He85g7+Bm
IcLVzaXdeiPTbuFdGcE+JBgiqccAgOF0beG0cbnhnDJBUnukGNnDWs4xBlWVhagccDwfEDx2XToW
uDTQJJev99XlY2PytkXBWWOtND083yYdV06ImoEC9vqj4MuxVp3v9QmO5aQJNERKi/SiiRwTa1/R
kCwvUje9OAbYBuIO7P6QfhCjmBzUIYiNw+3RTZBsfuhyDsk36e395QKdmYymMofcep51S1WNJnno
knv877nX8AB8SGphZIgG+5/fhb3LkGE4EzE1S6xhWUl1Z4fwYHI+rWUL2hfzkrkeePPl7M5iweCq
oJ6AQlhZaOlJ3ebilpVCehfDXwtaeZdNNW1WtqLqZPkDC0rKL2jD6hhkgvz1D495mUHKfnw6RuSC
+xDrYI2jPeU3OGP/FPEAf00JIPdS5UmSyOqvN/3pher3PLyGchdvuxHpTDH4Bmk4yzB1nhs4OEgP
QmL0SZwgf8yuzPSGW1+wuesudDI/NTitZtWd3qLVB2K8mzy1tdiTLaA22j9aVCd4gfs3r8AffrSp
z3b4CFQiQ96b8YpVmowhT7n/I+HJdYqLkO3W/zL6eR7F/hylRnGWs4ZbvWQH9x6QkAMkBxi1FYR7
hKkAn3FqnNl+09eJrMWZXfGmHXkGER9RBeA7N3Q3hSc93zcGi0EU7mx8+/FEdRlbmjtwTvpqIFGV
1G4Hf0Ekhe0YhrmV+aNOxyBr6PxOQd7olVAE+s8khq0RdZCmJ51lXRrm2Tr63tOXiWPGak7T5MI8
mDE2w4glu/2bC9+HOhrBHwbO6xUXKXJ1SAzg3DR/+8RO2YSuht+Ec50AdZbnpWzuodAhoEz15+a0
CeDgEVKqg7Cg0w62XIwh1EvVTSCAIptv+mjdVu9L8taOd4UQvM80w/sBUj5FupTdnxKUTc17tCrH
FYu7EXx2LgYtQlySMQzag0cVHl8Us5WjGznfmtayzDLA0tcY9Vt4VVZkUm2Z45mb0D25nffcYcJt
GS7EGSnKzRpHtjA9OeNW4dC8Q89ryGzwYLQhnodpsczz7EXDka4RTnhaGORoHzcD/jRzFzriZ68O
tGDqgdV7RpMqQn1OtQD01RZxk1Df0sQXUkAM+tOd0ZRAPr/iDkv4IU5o/tWMaKXYxgl1lhXh9Qoa
2dE51ED1UyfAsmTmYlnhFPcZ2k/cFwbNJ9Qt9Xq1YOFA1b2lWP5byyB//VMPbLx/LQ6bGwQWz/sD
+SUdx1CcJB7wnqsqmbkwxRedsx9SmbeQBoPdbWzmymlhpus6/57LlfdlULrxpSzaO/Jr5KkGFPqk
jYb+eqibObHP8rJ7Rs3hUccfst0pwZJm+OD4Gc+T+u97SwcOAbF1zLtZip4frTxGPldkqC/Bg5q5
m83S842ZYyV7UKPTPbprbuBandzomI6Tn+bQjsssaQ70EulphGRqZgJbQzWcET6o0jCA9DijPC4Q
JGmWggOqN0LXcR8ZwUX3DgWXQxWQgRFh6amvU9b4l9PjYLbmcmIs00OYnDX1hCFvU1jKUiCCoB5/
C57vFbG2BA17Pj2Q+x9DyGahqeLrRveTWJvhV5iPkrCBhwDo4tRwtNFcDBvB2gcotr+xBmXLc1tG
s97Vlwho0twELk3U9zhDCQ8WILJ8ND4DYDCtjG3Hm/LgPRjXSRh7kPDOwKLeQlSgorpI1TS4oIza
cdPrLrzw2ThhgVT3MEp9VkVOPymkH99uKKm1v+/fxHXNZOtQgiIf7cZBreg+pOXWgX1Y8N/+fLaa
8THEaLmk97PAPwAzoO7LG5jEeDWr8Gahube0ovbD6M5p+3pYdC4JZx3JUixfiWXoZzXzBEwqE3aD
IAxXez9yz/62bzKHzMX9vctRsjFO2Ek0IX5ZCUpHIqvcDBAnBaOPjBxsQF4ilBMWW67bFiLzTOMi
R0QDBU39FsbAhPN9D0HtMdk2IqbAaDsie6mO7uYk9uUS8yAk7SnU8/LVN+4aoDJUbUb5wD/5ASdf
wh0L3mAcV55nN8OJFEBaDhqZE9uLhta6UwUW/NNoqWgJLK2bDoHqpzIDBNa23eaQcL+E/EoLfmWB
S7xnodQ62Z6YhPJ7K363hRvwiO9LRaYuKiAngfJi/fVmLVV03ERlpgVUqzwx+ON7quQiHv78BEwS
O3J0Urbq/3H1a075X+mcSdeygo1nNGHfX1UVVwYmYAO7Gn7kT+B+IY2MzSBucUdkBEg+v0OvvQPI
C8aEI2FE30+1ZaykESGbJQ+mLiL+kGQhF6af3S14H1Pep9OzIv276B/VL4hcNez3yqxfRlM3+Wbs
AC/+K7RaSCtKaO9Dnkm6Frn47d25cDDnTEo6v4vhhCgpaGTxScXJjd66tpMU+XXTWVIT2woByfoR
5HDTEgA7ClZsvSFEg4hm2zyxt08jYFfxp+wMQHexjq/YMN9pmzGuD2f+pYercLAgNQYIcejSkVJF
2oqA4i+e/UpXXj6Vw5M+/wF5QFR2F4XGMCyEZYjPWt1P/tbQRifn46h2uKMHZguTsg5CKvPCMpxU
3Az+b6S6UVko7jXLVzda2AL22GGzFFaONR9/IwT2Smx5Bwwdh8zm9vfdw9+9TC9V+TVOn8q/Lxp8
hJGScPmQYmSOiBw9Arw6WFAjJu1N3t6nFUeTi2CFuAbbBDBBJZsx8OH3rgkgjWoxzCVq1w1l038O
zs2Bwnynf50FYnEbHM27KBrzWw9wjSPNR7gINmRZo6HSJnY0A1KZteq7OvKR0vfmOHyAwthdimKa
4P+/4Gl4b5+pkTmTBb8VYtxxB5jnGWZZRwwImoadLP0DXuPLc8h8vNesm4IUnnsiWsJx4IvOwuhJ
o3TRZc277wsafMmn822z2n7fFrexp7o7PFBFfql7o1yqRec1WMdBanrKrwClGxFzQGYNQUa8rTPu
KaZ5D+hEvbofisVPS23EMNzmLKL7zfkbxZql2odgVx5pDHL//wUu+VyBuJTwZHQoG5XakkCMydPO
1LZwBPSf5CVbCSH4HeQiQlUGamPJ7nvsNivpRYcBf5E/XCwEWaEUL9tBNMVFRaruUQ5cWT6MWliL
BkLX20JWcwGZYuYsPdPGIJcEnvdAYg6RMWjOvxLb83DtjN6xpYiKd4NGZaOzwH0bUohmAWldVeCK
BXb4HX4otpeUJETh1+0PvWuWR2QvBaDmfwXIj3OoiskrRQpntAGEnMT33rJpu5BTNjb5ekqMguOz
TAcbGA9vkp9Hk13xrG2HHbWei/t2qb0XBLxeNAg9TggNzK53PbB5eDUm49Bobq7ZhQCukRcIbxJP
TfBuLHq2QVKQAu7aSYV8mden1psa7dU8Tig1k1cfiChZGaP5d2ZFO/TyBePW9gfKMHk5cW59dDtP
x0ulYZbxeGshozLqsMklAnthGJdKzo+ueaQAuWfP9gcgjYyeVpGmNUTsBNfLoIInex0Uk8wTlyjG
gm8DLRF0AVVGmhfSuZVPKv4xusbySYYQMtgjx0DKWq6IynSAaDbZ3EVh2+ipT6St+Z915ftvfWQm
TCCuKFKgHY8KJuV1FrroOXYMCSbwoV7DthA9sgGNw5hfU+dYUBvc82EwIqjgAYeFOdNr0H3PBbxr
4ph9e3as1y8SlrGDWendjGK9sMM71D8QzUMgGvQplsm0mTkhpNnGha+WAgMofsMPD1J8SZw87ExM
blVSkC+CZxIiv/VKshb8FADmerXDjANVf92UtDjL26crIhxuPhCRk9PwQQ79xd45x4TW/u75MtF3
+gVX/LTQ81p+yB6cRROSmW2uDZU2Ql8=
`protect end_protected
