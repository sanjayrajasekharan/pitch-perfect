// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
MXhf6xtC/ZC8UE2fEB9Oqw+dMZyTuszM30QpGn2ziD9W8LPArzWDLUi70LkwDJeodsUug2gMgGHF
aJhpsk5IR4/bCbU/WFuD80UaK2XIPhtKgRRRX04wRexuWVb4EA4GmPUgdjpci6FzlXXkiYsgv0oR
NVVXx+HsW42m3i3GVZAYlZC2G60Thx+LbbvjnngjF428RkFiTsLV7pT0Mec+fsx0HjLDFjHt2Ssk
SGNzPraAkGbyTejhUJD2G3sEgsC+vDz+f4zYS7c2gYTPkSFD90XQpJY/waXkE/G4RdkWC22tjMtQ
MUtGsx0e9k3rPkqufxxGB6J2/JslGkApBqr87A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10864)
L6MtNACBeOMX8oG3MDpCTY2IHskWQYqwdVyDrICccyKmOQyd1R3czHlOzD5g1iTO1MYNzK4+i1cc
F9VcQKeLCaT79ASjNkpEvyq7nsSZhWpvDfHmfFFqx1u+iVsFKYCDVdQ7WubEoHamHYPUyqu41CML
lFX38zZXBnv5gEmspPP5//zSoA3Qdbsgfasc5aMnVQwaZrtcmxVHNI3ghXcqVfmrh1ws7RbU4oQM
2fm4/ZbtfAdfiLUZaKsmGyxlqZeSarKBGcub7quvFFJS2F9GL93ScJEVJiNtTKFNu2mlDKM0DM7Y
KnhIbYQ0Ir3oIaiyiasKdiabzu6ZlRduVKDFsxhcAlawhOeeiHZ8wyqteOAwafTEmbcyHarvNhZR
oduixMAfhRIWh+6jIhUFk5JatzRdQ5JWeBfllr5/+//2PRuMKpf8yRnXlWMENQdUbVqhYJ/lEYhY
kQGgT0ZZMIKIY+86achyV0Sx5ap9sDFyuL2RlBPY+y/hzDQTttjagJT9Eb2B5aw4Id+47vd7ZyGZ
LzoQDBMVwrNt1Jt/bqFcm2Gv1sOhb8U4RGU2jI+BAu+rqJpAS54VXPVTHoguEmHy18koOzhzADYt
COzxPG65/keEudD0bn9YsmmTHNk9RaHAXpAcIqiDi1oqINb18PUyq392z2zyULypBkxrVC5vYu0c
VlqDxFGVH/RbognBaj2IylryrdmFfgCi4VIRd9zraLC59YPTMztyc92yuscjUAH4echz/6kTGXMl
UafL/UQXwirMHNcyAAEKtnbIBYvo3Kt2V9+aA2Cz1YlxBcqVNZnpiYlMM6MYctVuvbQGS6xljdP1
D8nTIKTiIvM7LBEctrxjyWP0rij3bhzjiduX/06pArGS4pkYU/RdRi0zBH+85zU0HJzZYpk1RNb2
4Ut1/A4lCgOk5Rfiug0YMdwa62zg/QjIyOoY0MixYXeX+3Y9alqQEUDmidEtbvtag4tWrW3TameZ
HPwZRThGlJpEO+gpwoT3mBIZ4YOTZ9tq6pZdaZ/OMFSnomqCDKQtBw9k1CuR0/Tt6bkgE2i09+nr
sRJTVGfeTxAWCw6ZayQYNiqBdozCczOv5vEzPc8ZhK2oYUYjjEMFqUfrN6KLzUlvkHbbnDeh4/du
1xP8wgkNM6prNOVLKkEAQcagguU7goDBETQSdE6ueKQOtN3s+Z0jC7nPVJnfkkNmiA14At9XEyN4
aGFR4uZm2GOXbQL3DyxXikJyjXraAGNZACf0J1w7k6AvS4KDFZOi6p6igWpZow6aJv22BGG8f+0q
ePR1BWKt1wgq/dIqmk12gm99jQkJTVHUjNl6sbp6WbFMHZmAPBQHJk+oJmK0I1bh7o+XyoqgWeTv
U/ZbPumwmbsveJ/Vp48wmVYgGSHVRcj7BPSRiQjZwL2AA/hSeSpx5pl9V+empSxBrALPdqtb93gB
yJR4J1xa83COgrlm/4iFZDQva+BiZezII/DDmxSz4XdQRGrWhLh7waOQjHfjdZDtaliZYrpF7dJx
7tjkfv7+P8zA7WjJblkkhhhSRezMkmi4PB2fyZafcCww6pT3AoUzX80nvMM7Rce0c4OuXzIynm2V
XR8sIScXKQRi3C3JhpDURsaspMo2Nzh+m6V6Tt+cMII3TkM+FDVVauHqxVSZl6uiXuesHfTEthai
c/7SDJDgqrMw6AySVYjnT5EYT7/h06bhzDL7cn7R4214LfDyPI1KxVl3uwrXmJmGL7BuHo2/Hhsc
8K7E+TdwDe8z7I7YksMfgbkS6MQir0Fw7/SSu5ArOTAzNtUCT0zmmfV73P2wWRePAeTcoGIBEEAr
hgusb5H0i9LUZlyzZJA84l5nhsIc+HxMqoN0DcUiPo8wI9l0ivu2w9pzMq/3882zVaAQaXjxpv7t
+GYY4WFt8w8zJSBBNR11ecXMn1djdEH8qZKO3UI98HDB37uOP7G84xs+SXamLiDJp4yp+m9yrmdA
nAa5I/skOAPuciqvG11GtPF2Ge9ywiMB1euPyDpqnPvqx1TecL11gWWqs06OiCvuEJonFRtANMpO
PtoAln8hkB7HGkemGPREikZhAIBwX6I+pGYyOez1x7zWFyLrFsR+SaEgOY4xyI1Ii3vOwA+UdN4z
RiRfTP48hDP6hPEUQqLGOlf3u2g5R+S9TLdlsbRswUTKDQsOChcKBwwMIM15EhJQ9O7pfLLc5ITL
JIbWslFF23MT9/rHnmTW1YAbHMtw5K3ki9M+32C+oJeyc4MzSSW3s1msm7TZNbiHV5KgS1N1M1TA
po3r+BvNGbT9Rlq83fV3Y9Cb8INJM54+MqvudWL56dESIaXaD0HhQ4f2e89MgmNRCLFtYPyJLR/G
6CbPhE7vAObAxCdLx9prJCkNsGcmkJob566BcLJaWvPoOMuMrNxJnpHfwnf1tYh/nI7CcsnOiukf
/7EciIWX1WxUihhsFomgnt6mobAtRwKU9gA7q+ocgwEJeWbzOJGzB4KT9VwaafiRnbGTU/bqh3le
06xmgXwReN/mZebbg3mKv9wTaE6FfU4YV4xxAtww5kWTpLi/C8+Mi5lCKQ2IOFpNBYa71GCnZBJI
LGzvT6e32nLXawCd4w4QLs4BXLuDj7mcGr1k7xYFCdW6z/fgEjGLD6+CZmsS693SHhXAQxGLXUSD
+1NArRWFNf3zeC4SZxzGZ+KplVNkVtoppY/1yZsUFIdWCRMZ9tcoeBNArsoUSD1LHgaoUdVgkhsi
yotruT39ikW94W5kFue5OjVk9DJ9qmyIMYt+fVZZjLgCgBVECwAL+O2w+L8uy+EMuMUej343/mcn
vQ+ozrBD9vAZvVfH8VJ2EetIQpPDTK/H4e2mHtK8Z29VgFyCHNC0y38ebY2Bn5lCQIqz3rpmBToD
t55Bew0ATrbd8RbPAS9JRPWDUlQ+7bvixRS/qWoWl3bIqfveVRy2T2e5pHK/dxYy2ldnuREsSRSI
ZDYCrjfnzZftxmZw69gyraqGsSguwQa8Bnf87sY06Y9Na9lmcb/5ygKDIGb8LzFgfYg4lDuY1fJX
My1bppKfqeGrOqikZjUzBH0lnmVd8B8bAtSfYPyouE5sFsSfdsuIF2VPjGXLlZRlUIGEQDp6bFkn
NlZLmG5cXQXyv9QEe8Y8uQqTq1pT2NE3zonIyBtey3b0J3NPCinX+h8Fc7YFu8cSlqEL6wNZDtHf
aUaCIcWXDlg+D0huUSsxffzSou0bWvQKR4hYuN7mFIIzfs1Z2gNdS2ncuHkqnu7Jt7Iiuroeikab
mSIupYuhmGnNT45XQ/BgAOCmqpvGkPhNgIHgmunU7qIqO18t77hqz4IG9LZw5IWB0DWaxboII9kN
7oSKnQYjSRIj3wZHpGXME+KYojoJ/Lc/K5aF/6hjflsAKBeyGh5hXSUHz75gb+paxnDQO/oMzScm
7Be76y7r6yz9X++0hhqIflYUnz8H6AM9JdP2W3ClmwqD3mQBtREdXlpX8PXVj8rZWOeuRVLVAAc/
ZcYGd2XmbVS7ME00YkoQN3nqn2v4xU9niUq/VM4udjsWtjXd6J11hjNmzmBtW5PdDTm136sgvj+V
j9TKLwFKVa6YrlVACM7WdXvVWSV/ihN4zBaF2FzpyPg5Q0fAtDhdOkw4GZaZrPJ3PWBhY84IRGkn
PDt+/3tPZaOR3Yccy2nA8cCEI/+4/wonZueYCAhSEzgoRxrnqtrCscv8eTfplN2dliSovwYDKX8k
aib5365pAIJfut+Y8N/mtrm6/dZau7J1Ppf9K3N4/ma7IVBCO4sRZxxFd5lEdyMN5/Zva9te/yjm
v2Qo7pOEUWh7WfiaWZpbL+4orn8lLtWoUf/PecDYKflXrlJaSE3KuPrgO/58PT5i1JcFZNN8M6L+
pVI0sxqHTCXU6spHD1bbPEg+JnD0rMJxHJ/LRiX95uaMRXGUy07sFOU3hJPk2ibKczwiu+LHXODR
2GGgO3RnR8G1U5V16CQ0ExI8dVnqUQuMwXZpEByQeYtngnmkx3+uqnqQLxL9scBoD4MyIpu4k5KH
PlN/1UcFeoEkRjpvqbgjYd0jtXYbPROYHrJELVa5uFnGfSOmEhqYOKxYsYxuUKyEsvBUw1olDz+o
SOfI5vQq5e4xgGpdzEfgE2WFJPvWiKICFRDawOkR4c91uJHNT0g8cU2O4Fbnyxket8Lkrk+6rPS8
iZr46S3l+BavT+lUAQCPFBjplv7XMuldZENQBHPQMuM9fIUNxHzFTAit3y6kIRdtWnGGypsjfqHE
WgY2L4GYQIPEFHuZSKsx1eZU6YFmbDNs3smMkAV70xBGOlb/B3K/ypmFmUfIRvz1AYKPmGU1LJGl
lwhdn7ZOvmvhVqYE0YdwvYfWxFkAqte1oQuiQY5Rl+PVywNinog7yJjQ+2OKII1WC2MO40VAsiXR
vUUriDldtL2CoiW7RbB+scvymD694bU/vnnHQkB4cRyrre2ni3LKY8vVUW/dk0TWRbs5r6s0L5Ff
vcq0g8pvUHNaVQIA77L0AT8+sUhcnndJebEwp7Ia9h/eqAA6rHR+b00XNOhVIk8wOs+bhLsf0kJZ
TiwEZSketRUJo4ob0tx0ZGxQo4ouJ9XGQVZjszn08YUb/P7kiAtn+6YxUursp0mh0qrbKPrPkFqf
CIF4VOdUYFVxd2BxB3fJAQ7rhbi3sgYznpKVcv2fScP8+JbsiLT8j+/5MPVfuco8GOw7SZUPfmp2
aH/pSquxo829/06rLkOjKyup2xMdz5XKfxWvpaOj3JUjWOMRnh2OIdj6UwkT4yO8avvAfbWuZRKu
NVag3MiO2VgQvb7/W4BXELtfiwrUH5GEn2MZYjaFikChr+4Gol050yVyspI7iQxoJF+ZI1BAORWR
GCwybD7O1j0og0wPv0P2+EMU6AzCV+KUimZQlu8SMhrZefO/5AnQ5VN/UEucoM/8UqNTA7YAzrod
JAMtuzkSa5jhz4KB2FfI370NbRM4/9oGWfIrUsddgnpwwl/OPiKHOGodzfT1D1ud2j8Tzy8JkTbZ
Q6KfPcOdxv05iIFd0t4PVMzT3nQNm8KKm1jxikW0ALRwsiDmL4m9BFpuR5hFVJYzUDcLKC92FvTn
sSjK9n8F3gz3bTmtOGEz5CyUmWqFR4jcL4LFe6bl2CT4kUHimfDKtVP2Na6t0D6fK/2r/izuIAUk
SwbZaxmTcRTUDwDOQNYL/rM31j3fMZTcyA1Bm3FA5y7AeSepFtyUd0DhH7O8Sy72Rsy018e2T/V3
H/1RNdOhHu3T4zGvZlBrfCxTyitDGIgXifJh+Po9wDYMBSxNNq/AQowxAOLGZ0U8lZNpue46Sqve
O1DDJ9rOjuog/euBtHamVPVklxMzj0azyiSAYJq8iCUtkomSDGJWhLnmzNT3SYlchO9rsL18pBUA
DMdQlw1BMdNxcmbQCjr6Kp7ORlN+dE5tO4/kx3ktnu6aHHq9jHpgekcJuqeOVufwR5rWFctPbNg3
SJiNOh7K/fl1GZe8toKZUCnZ461u+nJhQ+Mjj0Db+c7RM3pahIajTtu/163aaYElbYpkrZACvxNd
bpvWrUCKE9QWLIKy9+NI5AHyctAiISyuVNqEaIh8v31oGN6OISSWx3Lp6KAgfmJuhxsFrafZe4uZ
TnKwFMuIbG7P+6GWUMMyydNx5T1fM5yJ6F3qWMfEXzY8uKvRYrmEeJot9x4g7UDqQ+agaqFUgymo
qSMcdTjvWHyO1VXstGDYmZRiKuRkSoxFnt32zPxMz/6/MHfFZbPaKsNSPdZxuE7vnTxuCzTaUJd6
HnQlQfIJBHEMuME9N4/p+8j4RtCE3zO2EoEStHp/q8/nQIxjkFXGmWBu38ExAYxwoisf4MRc67Tp
cTLNinxqFCX9jbUbVTRVCbytBBD9n4iOXP1JyMjUvZ5qwwrasW7QqibIgbfrp4nHBQe4qDl16Bme
wbLDZbco6trf4YXLn9ZBZ/RyrV2wDaGcJ6ZRbVLkA4XDWLPKVCaaY0zKPfIp0YHedLoISx0sY68w
fQfELlSe1QfN+/MKiTE31hBJKSxsqXokl5wZkD2agMfhHnSb1g/0uUYwrZGqMOadJUh90PVJEPQy
UKITlef1cIxIFz001N+5cdMCp4SN2/y2sF7wyrza0/VixxpdYUVm8nfPz8FhNvrm/0LHRWePtQXg
G0Fu55CsKlo8y1GcK7GPvfviMYwLKTsZ1nVR+/NO4B7f7B2LSuQMFSF75IR2382RCAkuY30lzc10
Rnz04iemirlSsuTgSaqErGsZ1bYert8WWjUuvhtgNxW5fSK2eld+ANtkiQyqjKSVSp+2vxkkJyU6
J3JENhBzMrRaSNkZE0GDSysDAQ/1rgI8ctcGJKCZ12L/B3qozWnc2UakV2ralEHvJJmdD+KP/tIZ
byqc6Z+CiyQzg5SiIL721VupE5jz2bQ3l/yF5ApJbDTp4EwgGXd+K1Ms9cT4oPRVqjRPq8JOGRLV
Z6wfZfVfvq2uAJMPbbzCz98bwlpaZgNbkYBLlkhjQdbBQL57u4zY3z4IR2jAPjwTTbE9WVBKJU01
nQ+xu3UBmEPl6LTbjXQAOMTKnH52aiHKv5DwCM0au8OGBw8P+qymHBuxHYe6F59GBM55IE2NU98g
fxGTr4So94BiR8tTBJp/Ex7PbQFlMbEctGWtQo8M/okDupWNqoMBT7CI23MLPLwfNv2ug0pqLRnR
3tR8FctOdS35ebAUFFAxNo3tfzwqyoILoinA7itqrdc/88CkqOrSoUHIzXlL3D7cVFwk3T9XdOWG
Uy4GPhZrJxHYJxwNIzvuKdnJ1dQ92AoAmWNLLrz/iGp8W1g281W5kjTf24iZAcwYa8hRySwS6JAz
DcE0iupkii+r5BFk7dEeOyAtg2lsUR900vjL6HPKhoCYhDd+Amf1ykeXRExmpl0AG5iKIyPf4VT2
SKsUkPxtPVyeK0Q//hdttUQ/L2PZA0edSBp4hl7XcnuhWBt32xRUpSTElbiAIpBNQU2f4BuAaPcu
FHagqy4kMPyJ5nX8jI56XjGL5/fhixpd7WB1iwJOm4YqSBBNwZfJk2vu4QwjQMxOjFFjjhXQyt8w
t7cTDOXXmVIg5bQqkA+qxSt9DU5C57DOiS3X0PoXKwxGqaqt81jNp4qYQ/zLo8YQwqwZmbRhw2qC
GyU1yP4PY3UoQLGXVQmgfdZpf0QtEpTOQIJFbi6Qr0DXAOS7GUTeFVoLYb7wvAMz8HirZS8SJq9t
PelttP/C33j5QTbrGvqTMUv4Ik80QPuzTTx/tBLnuZ4rPYYLE6CQGpuChE5ArN4Lwio95bcMLD88
t+DsYHmne0GwZUJIPurVFHArO0zl468oFhOWOERTmTXeXxLdIYX3kkR/rc17ghsBWXWfrjajLB0o
uIc45zz+URYAfq9BoZD0WNCoWlQFsjua3N0jXNDgA2chED5EZqDag4Ydai6Ua3rz+GhuMmswYcxE
zvlKPPlnggWp29Xqbtbpx/tPF3I0FPpzzp8+eIRyQlc+CC/uttj01QfvXVCkc71FUiKV75ENPBBd
lOPUBG3RJYmbBbgEYpDJG+b0aKyPh0w+YefPCnsrRqWLocKvuPht1n0gC/IE+bwi9bv+8kH8K3T2
4Aw9zVwHYSXlFazXF5y/toSID3YD8Sn64jKOerrdwF2rc5i7kI2AhFNscYry0kgReDgF8W0++YiX
aHeoCbsJQn+aOWYeRiXINO27pgWrzENlFbt3WLIwzrixTZ9cgbaCZYixP51cTZF3o0dkgam32HxF
yQ5BzuOy8MAytXQfCP8I8hcx5c/PRBIV9Qr3eM70Le3rM8/Pp8JO6Qihwz2TfgfmWaSY9R7wHf0Z
L1g24QHc8JaxNwl/RuAds68Tj55BIwJH3QVStLFQuZYRgXp8PR8XFI6xFTVrVYwEPKmhDUSTt6o6
WZImZCCgcYwB2RYTNoQE1BHLeG6igA/XOf4zXgJqXwnsS/iutcCkWQa6AUloyZK4H2TUPnKlcrf6
dA/SisBuSfrZTLQt1DbfLQEWFe+PYbmCLG3+Ak48zsXdO0NlAis2d4Rg5ZbgVMuoslUwi7BWge7E
9ZRDEcAHTMZaoJEZQ+aR0z7sTxUOCpXBCOzzXpUzAisktHHCUpbE1AAysa4GnXKAiiWePcmlEdcj
X7eH5ZEik+07dd2H61Qi48tQnOGQKU0wIWAwqL5O5MfgCqn8W8+SpQNZ4lw99cX0wBW9GvI5Bt4Z
W92vtsyyD+d4dV0BM3cKUBzGqRjrqtwHVgRpZE3ZjkO4iBibU9eJoSHpe3/oRmoL+D8sit5nMskt
Oh6jhFYvQuoEEAdEPViSsj1t+xzCpWP4cgfBOBcB9pbBB3Be0LpYpjB+omgRvlgJtuLSmmwGK0Cb
n4bdUb5RX7hLLELOKrEdrVsGqstRREBxknhQCZXeuCXwOV1SOKzKVjefUdLAwBMA/p6uqqFIkSvq
Abl86PCdn3LNMzODfA4lhFQUZUjl+4v7cDFwI8xWrwiWb8jkLiPwywBhnKiOTJWmoBWtz5FhHGnf
YwKic4Q804ohjOGtn6iMEqFewF3de/GlDiJJzNE8qyg7QJjmhdxX7qjJ7dfK0jecHVzsoY2hp8YX
kCF8ySS+cJzcCL7mV9Rqv5Pq7jkm+iTjDCFXYw7/Vku2/LvCxNSsXYaXkzLEBe42LFflUbw8FowT
mifVTECVHFPhYQr8EJ9Vbd97bNPwKrL4sMya982fK8ECiTrBy/u4mn9+fy/B+6DP1MJgL/AZmp/U
TVFfrPdaN2NmU4egx6L/CehdOmZxnIzaYwmfx5BOnDSLFbY/R9CB88WLGWSwMtcXchgfiWAFABrd
UBq6fJoEkgqxoamcW4j5WRULUrLkalmdacrWLoPiigtqTwRIpQ9wkOmIqGWpoG2PDrS7qufiN2Fw
pOapxuXv6yy6DTp/94aE+hyNiX1/EB07MVB9gwOB9AFhyATEHXBOTs3KP4GDwAgsDmp+2rFKxQy6
HdMyDkso+Ez9/0NG1GIguzLEkqO8o0oqPFbb9IHNAf1T+AttOodF1zde1eMcYpUvzrIOXKEz9lRn
n0RK/G2Mq21Qcc2W+LwazlIZjFaFKH/X9HcHt1ZBV/CqC3haV0lYIIA3hisd+TSwHOdPCRrPwkhe
d7472/KMQ2AdgjR2pcDUu5eDEGKptQRYUghUDTee0y6upmUlSzxMGxeSZWkcvqN3ak7YcN/lQJaZ
RLHi/sXDem6tF11lKh9vCoymUnRFugq9Agw8mv2Ud7ysP8aMbFnaKD7svoq8s1woLK5o0e4lZjc9
FPY/Hdzm8v+yU9DKdzLB40RhXFvNflv8d3h8O49oF+JBMBHKm7CKYDcxFr2XM2OUO+pHrF84Gdsw
BJfBuA7ysbo2y9tXqLVbFThtQOV1TovPhu9cAXtGajhE4O2GZqEkp45jMlm8vViH5MXUsjubTxPx
me0eNGEpDgY6UM1PHoEoVylKDPbYXQwBDg+4he02GgxcaFD2BYqLu76hSVPZgqXgCXNPpm4JkjGR
RPQGgd3UwYEqpvp0uIpU7/v41KRd3k8DA7I6k+UJKiXYWBCCn55b1XydUX/JzsdY8BzTP0fVrYTj
ZcpL8v1m+4W6ZEwe2hK0jv9xVMOa8tLdFjVIUE/p2OWsfk7+h0BqS48V8KL6iIeKmgUsIApYwqBc
b0XPgsWCuNvehrWuoYxlVEljX6l3QQqJg8srAENj9TF+yBr6bEZCbVr2KEDIOmNmJnj8ZMbL3JOX
H/gCVEbI2CMI/h3Wj0m9DX3FJnSTTnp6+naxHH8no9rouX1Tc7KImjb8glLQIvkmyGY31rkzl3IG
V1voxELiusGM0QwLW5Qd1xHDCmYndMBQbm6xqGWPSeSf70PNAzvoU3+hN5bLrVYrKNwXeyLWuJ/h
Rvv0KzSKezgFBdlRNPzZ3Kv2kNRxKX9IemMTqdw/kx5ITwzmYONQD6SA+aWuE4tznk9MXeHfqSxE
NlxgRZvxdlQCHr3ZBXGJ8fN65Fo02ToVZ/arLFopv6BGrs2MhYGUTmVuDCVFW+/HxW9+135C1gQr
ZT+VGGn2lMeT3HMDNwRl9kD3rJNRAWCvyWL7vmWBf2DeRo7ojlh7KLb+siFa1xkFecrt/b3ptZfu
rCNUeYSIZ9gfTE8In5tbx6+jnC2ejv95w7ziRE2pd4CGboTMBtaX5v+ArlKa7bAxd8y0OjIlUUnU
1QMYDHdZ2RPeWE9d+nfkZOfuqTIOxwyKC4Rlxu4N6HNCNi+O029WQT9Gw4NkUJB0ClnB8mY+pmzI
u0cxAQuu410hDenWi2n8pY9hZEoZkygSbZgvsUN/kC8PdQ348QKSpF5z98tj7s8RVEV5NGNoPK59
a4f2rd/Rsfvze3YqvMlhcVaoCgQAgimBXL3VYYHD0XyHTDgDCgV7maNMkLyb0X5LHlLpfwecGhGr
7HzcRp3dHCR9zfYoC5h5TZGShhltGtOFKrad92NcWHjO3Fwq0gjN6u2Z9Ggh9tnhUh6bJZHQfqKe
Ego/6kKBnvsn5XHmj9TYOR6c1QnYxCMZfXBr/DSIKUuJ3YvpF6Z8H2d78D1ccXYmqD1SUGh6AxZN
7vvGlcfw4TcgRsuW6d5BtQfn0fZF+A5SyM7DEkHzZoOkNrHjlS3cS1eG64jvKzUbG1zYB9X+H+mc
cjEKEx+yuT9BRs+wFaQUWo/vMYq8d97s8Iw2x8G7TLFTKp2rV0eCjPhwht8+i2BU+3Q9v9zzRB1w
8DTwxhW1J7I1AOiQ4wGw4xMyFYaoVRovY+8tIbx+4CHDgLHNoJcWgo8KfaGWHXyR3e2FtavUtsDb
hky1XW6UKuvyKbcFjIM/urB/t+eYFRv6ayQR+Cy/o+/BEgJd4xxkayDPVS+dtstaqFY+rI/FIULj
2acdN76x5chayThiomPyprh3tXfdhUP8JLpVN1zkK1OlABarxZCPuwJlYyUu0YvR/9o2l3kNReyV
8wZ+l2c4hEoKWHKCS7YSNIes9YqgcXVwwX9A3XeN8D2CwN6ilSK3x4ItPM5cXaOpFPZAZWwd9W3T
UFDbZa8ryJc8l6AJtSNpMJwx6fp/rGdl3Lk1hJSLGaiOiynOZ4trp99KA5kXBR9EynpeqF3jbufj
p9DhKTfC3xIAwPIg2fWFmCWueFUd5IphrzHedSg7XTwCl3Ov39THAqJlL5BdkDcVeY9WbldkbUxa
D5XpngADgl+YXXhNYjmfEaMMUFwMJksw+2n45WBGr4fcE7CNvMtMMCcKbQErSGIifwfvJzaB/x+1
EoTLrn2fplRwiKMIloTW+3rko/ehtj/pr7xRstPWV5UK+cTvolW+IFy7cQ1nyU8/kwvPfOk7Jz4U
XWU6ypilcfOHXWI2QIq5jgTMSLghkgHDxPTCRcqoxSuCHSp6DFwjEjhzqSMrqzeUmnPXP1fT2k8V
IDaXbHshB13qgL4DqG5jfk0jDBmfVWQu2zLV7YgT5a/sw5M6FmTaaED7IVVy9fCXQsrVHRb70Cgy
iM0f9Ytpn2nYQ3oE+Cthy7YQ4Zh5w3mMXrZ7Grn32NsU1D8QipGukklFfkKG/pIurp9lV649TKDO
yUYTvEPcQ1qL8kX/5rITKkn/6egyvfuzMngpijFZ4jP7k4v3+fUXFGN9GvTZd0TD8IBaF7GzmXHT
n8RtM3sEwWkkQ4v7bxIwi8w2DHcb2D+8jD4uQR4gQjriHm/Ul6BlBnx+J/4zLT0nNvOcZK5XLEaK
nZZuNPiXLJUKFJ75mXPwjrCoPkQB1+iqRNF3KQ5iquKGD1ffiBLpwIX67aQJKrjER2FQJgm5IvgC
9KLvOgP2TFAwbclGolkelHB5gloYTZOqyMaEbi+wU1kbc5q2fTDMG35kJUx8c+RYaBSI3zPojBs8
yifZd7NqqxTRl2UOF9gtMt2gYx5yDUuPykFUWWVNzSwbjwZr5MGzQp9+txzFUtkeXHCmCMSikS79
aSGGAVb1LjNXebp50i2vs5vETwVkcobioDWn3a7LNkaigyCQ+t+A/QR7b9hbqCz9aD+jhH+zdeZF
K+oLgwV+OPhHJaTTKSrsZadrAOkR9g5M+h1gf39R/PrWCdM0EqqU3Dbigjm58yDR9QHYC+WraDfz
1tDeVmYoKohYN4FsHCX6VQlqijPmDLU7NRmfA+f7lo4lN+0NyW/wPwwfqegRoIKYYxt8764byB4p
MEe+th6xptr/IjIMWtPqLokmH9W2ukkakIiSZuFrA9st1xJ72IICtb321ovgNck5XIThVktApsj7
Ve3Xg9Q+kWwYy8Kk6hEKasIXFcEAQ/8/EmrJR/3oDpr6Q/UyBlsRq+/I3Srjoa/fA+C4uXz7HJdN
fUvi20TDM1lh2HQzm+AoYYL8n72JQ1EcqHI+TnhB1HnjeL4ecV220rH8qMzRrlrwUteSGOKA+VSY
Bt1lG+BjqV1FjcoPYFxqzduIrAehiZOUOmz4XfIbcMsSEIM6TlMz089VM58W0fFGILRVPsGo1TNM
QPQX8wr6riy2qvvSVROmWv+4tW2yxJiRSvzVVa2l8qoloisgxH9xI1tkWFMhwVgFK57ahW3EjQmW
eC7hVUTQ7wL4qdW7AtRbKplgsXYso5eKmBwm+le5EcacggQq5TLxFTY2P1LBoPdQCbSUrx7EY2zn
Pa3/gJ6ZGonyLuZ6zQXEoDBzLs3fwf8FvfVgKUyISgSM9y3tYZrgA0s7IT7chLRbYUv3Q9TJCIEm
W//mmIxTKlxSOrt+K2AfncqUznOUG/WPeRamJsx83ViACaFmfUHtu1AXT/vhlsV2bN2i5+BUpHcA
wt4FE1g7VfyILD8qWOJkL2VzC71m9Ym9n7CH0bVP9hT21xFBaLEOXJ2gFnKgk9SSoyHhRNQjwSPf
t8z78l4eX+3sZdZUnYx1nX8fz7+MeFDga0W3SF4oEPqaQuRX5UwJW/66bTnZYGK0ClT+biwwepQ+
DOx5dfqezxKB6T/14MWHghRdC558ol3ueRSr3jPUt/kghOUX+V7YJ0cVrM7ywM24bwXEceQHJdfY
cYWiVXdBudzPBAY9GXCpn55xsyOi/nhPWFJYZL4XCh/krQsp1NYInVuJhPTFL9tVbRylerkZ3nqE
TCvyNigZJvFe8wXzeVpuuPZIWfs+mc+4rvRt419yTdz8Oyx9s3dlr0qf1tZmtnVFrqIRToR/pDDY
h+ACXP6QrbRcOzKqqrE8BNlUxD+h3kP1zDeduMRbbvlgcEKXCbHmwoOFd/23Yx/AMiG1Fx0X7Muh
O4mdGBQQeDkogYECcdMUU86bSmoJ3rvbbyNVSSm4OexjQsx28b6/EebqgxUpAguzxyQdbWLnN0II
1QW6ENdg7lAC9AA+8C9Ujb+odYHTnywOib/O5ZK2DDOrkWKxdk0sc5Z0WyoG+crHu401GmqGHkvn
Z+gnABgEKq3b/42Kv7Nu9yEByeWPW5MDHf7dnb5Lf3J0d+HNTfsiVs5cCgg+PKnNQigHE56LaY2j
snpVaOb+F1NevJE+l7aRDptHz/3ZSFnfzyNJLrvb6RwuCMyZY3KfgoQYCkAaW7qioMWUBPgGAPe6
yAtviOF2mugcQCSroRcB8zql1dNZTTdsZor2ZOURNS0CTrBLTNJLPr2oh3iP0biTiVkjK4B/HnSK
a8Uj8ZNXJvzoRVNxtHsOjXnvH8Ahqv2sweAYLTWhehDaeQAZvi675VaISYPDz4j0efZTnqbhc8or
8oX7Gg5yMCAhYw/i5qMzb/mLkuFVR0JLK8ARdc4VpTQRiePQZWBWdCZSiPOrlLm84tjULQgNhcwS
ZK9JTkRuS4LvS2tFmb3rw4E6MkA/JIRHBAWJVQdVwD+N9EiaQWqud9qvoMuOz67yOTxkZEw/q7aA
+dTsJlnNMiBiptXw2eWdnhp2Gq5NrGMA2zwPPLwqMAWd/bnXgXr8IpPK7eNY382W5h9jdwEdGWdS
bu55XX1sJvMp3tsAUzXz77TiDFCsblmtcgdct6KBYkCUL9FzhmYOnRU7s9CHRC3s6n60VNnxyrND
/iKV0wPr/7a6UfV1C/+sFjCqPXdm0VaF2yI1K+IGN/IvhivgFI4cvAmkNT07NHhqBlhF2NBnMwWA
iw5KvcvpAczOKdGODec6L+Qs+tWLHxmaGEUcL8IchBqpzmV20DQLcC0JEeV3cg35qNBFFeCsnI5y
ClBoZHhKeK7ZK61pt9b1wJHEDDUu0cg7J+8BbBWYHrYsJEkTrt660m4DmMsL+glVvQWbCJclyV/f
QlF6tdJA03KQfdYao7tuTQKaWf4UatXnt+yFbAelzmvWjsr0Tr2vCHr9jeHphFrj6cU3iXN1I0gU
/VAz3UScePDPpafBUsDmB63PHahzg/S4uuPlJWtUMgrE56LrmZEPA6Nbe0rroetn+ODM/lf6BwsH
IiwLwNEf/Z0xzncWG+UupI7+YkKEMVcwdufLTOwmopwtWReM4A76W1e9VXBswFMhoP4df9Hlmwgj
6q6u39NPMQniQe0PG5Ty31QWcy5BIDzSufVr/tIi5iZvOg==
`pragma protect end_protected
