��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�Eʾ)?f�6e��>jH�x��Ɠ}�����$/�o>��x���,��yC��m��U��;S��}���j}כ��#"O���քq_i��c�WVcr2}6[�4/Q���牴;���x':r�c	�K������Xݢ��J*3g*���X�IVQ[H.\�b�@u��]��I��e3D�똂N��g��6�O���z5E��\Jy������rlj`"�8&(+˶Z�KԘ�!���>���+��X�N��	�PgZw;ғj\�7�Ź?;q]���b�
�d�6��7��G�@����#p�)u�:��'�R���(�Y�ɿ'J��gN2@i��eI��H���w�W�V��}����ED�1G�@+I��U~ro(�eM2�E�y�S�7w��!!����$�az��f���~���/���ݽH^��f�E�`!q�O����b =14� +-��>�pic�� U�cfg"Tď��7]�[��(�n���ԏ����T�W�
MW=�����@HK�df�C�k��79�CY-,�RO�������D�7y��(M�Ut��($RU'}+��rc�N^_T1�y�K�����Ză����o�)G�22�)�J�=c��cjZ�`��&՞�-�0fQ���%�Bh�A���]m+�w��v�,H�%��YК�����%>V�Y�Y.�jEX�s�;Ò��_o%nX*��ݐ�$�E[	4s��`��(p�o
E��\��P�ņ�g sA��P�vS�
/�V형��9��6]a-�v)a��j�$;"ȩ�T-����w�̞�}>"e������zVQ��^/H2싪+�� �5�YHۇTCwH��O>4>3M��-�[jl��B��,
N:�q��\<�����(y��c��Lm�����ב�p#�6	hu���3
�Oxd|�ܔS�@����'�U�U����/Xݔ�I+ 3�F��\�9;,O�bx�)���8Mtd@���<�,r\e�Cy��8G!�Z_�s���D���)�onzL��v�g�Hg���v�"�]h��Ǟ,DuM�JZ�[�}���i�@!iF3�g�6�@$w��JgL����^+$�i_V�6T��
�Q�<r��	����`��V��[�+.n�(��.*͍�~�<<��B�{É1Հ�ߘ]�ܒx �ä`�gO������7�dX��$4Jm���O�!��Ɏ��'��cw�J$��f]���es�_*��+9�Lrx�-����T�k�/�Ͽ����{8t�۶�n��a���}/�.sbϟg�\� �ɏ��p�d���mR"��p�%0�B��=������K�V0�DJ��g
vFÂ}��:A%m��<��4؛c�P��I��l�Ш/l!�J1�~���F�=��әg0ݴ�V��cg����ޫ����U�����ӧ�����cr�H�F�ߚ
�]����d�dM�b>�]����͖�i����$�$����d��%��ӕ!�����6*����D=0�ԁ� �<ݵ�XO�:��r�rc3��ĝ�$hD ln�sR!}8[ <EC�q���.�ĬǺ��.XA�8a��q
E�#��]2�T[��T�4j�r�W�/�X��?��v�4�'��O������堍 �� �:���T|��+W�2�Oɯjf朅=��wXV�\�3��4Ԛ�����&}k�BV>[0х��e]\���6�����/�@`D��|I<�+ �V[Q��ΑVG, r�b !�z������,��7C��P�lN�pM����o�H6D�zI�WhO�M���q���jȏ��!Oъ��W5_nu��FpL����}r���R�Jʪ�?J�O��h<E��ĺ^iE"�I��q���!^��f�sH��?0���BPH,����c��es��'�NJ�V!�@nT#��s����J"��>�q�T��ԟr��׏&��~У�}V�X%�d��{�CY[�EY���̃��M�xFC����#S������0��Ls�X���曵�r�O�ij�*D]S�-'X&8�Ӆ)��d�P��%
P5i8RԔ爘������=:s�S����4 �эP+n�9����;=7;Y���av��
�D�זC��Jxe�m����,��&*QV;��|�)���OEۄ{��u����O�.݇���i�~�
?�&����%gp������m
�naR��L�i���S�t�Q