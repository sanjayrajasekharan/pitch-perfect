-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2t2nae5HBl0m0JbmeH8kr6N7ansGR/5QxZdLMj28m6tGTl3G72gy/+GmLRZiCARn
E5YI4q7jwaCQYuFw0PlILPpwsmThkppnJwMl4izZYjlKtj4o8BPT10GijvxTUdx+
i78RaV2eLYWoBjCKB+dxRrnzhE6ggbmWXTrfkVlfphI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 111872)
`protect data_block
S+I+FO9IdRO+ZyNkj2GxO9FfnxrXZWvDJvJv0Czk9ukfmPVPcxQgTp5tZkcqzpeZ
UOV6vZCwHmVgsbzy8Kt/0iiI3J3T65qqv+mKuKGO9BcmfOGBp2YKOyRpBU7u/+1u
xMW9M5Q/yY+JSofhVRLruSuHucFfbAsXutR+8z9jbAk9tt5NnA69/VHqbRqF/rDy
lPj0AvDNFuiO1uOsalObIV7cNlRZRjT7pZuYXOGv37ZLi34/srm5C8C91DS0tKZI
lvgndUsOcWIvAoG8a43tsBZ3TQZ6xayK1nEPlinrb0vAp5D6RxEJHd/uhJp3A9fy
58HbIl2Pk/4qiaEj6Jt3u/4SQAS3KUu/Klb2UJYkSR1lsTIN6sD0OfbEGqg4yB9T
i5iFVBls1EFerBoR7a8y0P7WYb1CboZnaezjxvwMNLJ5H1ZrpogHetO2gV/MyjFX
f7vqdXUkQix3xIQysFPr6fRoi1C6Hcs7GFJHEy9kVWHkJqMFJXd3HjVfEiDA2aaV
BJ/8VdjIKfah4H281Gb+gkqEvoNK/UDla+I7lmM37/9HLBB1cFyaw442w++ePB3n
SO0O7gC+JZ+xIbgaC5Ty4t3T7v0TTRkbI4CnXzNJIpOXAc8n2yc0HPk+Ga2You+O
hr7oPXLVg7JtYJRclZxYarB/xjNf1ZcUH3p7QLDgTotE7OKAovFZe2fihNM40UZH
sUgSAo3vUk1HdKyt20KFv4g3fJtYOeDwus2QyD1acgFR1I7vaZpMV7cry0ZQ9ow2
9RGJdJi3c6Jgh2RVsYM8wzeGvDR4oGRtHgCb0uYhRqNlv9Zt19sHPyiJmLbSqt/e
hGvd3mXPuEUyV08h4OV/zV3ypU2xyWIhVNySzChU0Yot/aekNfDEjRXhJCqk9Sa3
1JyEuLDU4J0a0l7z68MjaWf1O7QYSV5iWhrm3nYYkQY9/XRM4dgarcgCSet0rcHv
2jEbarsjnvchnsZeEZPE3+114jIvHoVClNDsPn2vkZAB8fKw/decL/3RZ9wA9S2I
/VKia7YJYNWafkntFCQJgKSve6t4Q9zIVr9Nl/dyH9Y2qh0ys+A17qimCAD4lI/l
prenUgJDpi4TQFDmOS6ArSMffLWglzcW/LOF2jB6xLBeaSsAzfKEaQNTw1sj9zY1
lvSMDF1t5mZ9xa8WCPO/04bi8kVIoMEU3+QokxCZp0+F953mwJNGPEd5XQbXokEK
6Pzj8qrbE7i5bT8Qw+jicZ4F1MdcDPeOAZh9LDS/4A7GqCiof58amvR/AKpyoGxQ
ztHaC4ksCaOSE1ULnWo6ZtotIyQNS3Ms0IttmfD4P/wLGpW5Hgc+xy/tSsKhYm1x
7d1LqmuqCkVT0W1U/QwEyRLElzTdAOrhzmRTv3ZS3rvYYoRUDXKmq8XMUjHp1+/o
EImd1N7niGv/TN9m+7SCZeyxLL+ULmIfZF2amcs2JYVbKVoNkf6MNRCEn0hnly8j
JqYkIIpEh2uEUipBjeWF5EYdKJHTY4IS46xrQgp9+ROUtHJEpBP9xkF22i8qj+sv
33V1ERXRPM+iYUQC5odQixvw62+P4iedPEvfZn40N61dvVhTr/Tfuig2u7dyBjyg
4TfFYnXDv9sAy7FIlYnvlh762PLOIIju87rqo4F0ypX+3WMrJCkNhlZHPGlfY9x7
SO9n56jB/fuyJgkhQZQE0RRweIrMBXxEKbRpchhsVsRZSKcdVlKK9vGTrHqmYk3Y
KwWKcLatI+WIjw7n4ZpnFUsybwdcuYx12OOvILT1lzjxriZJSzxEdXZVGOyylkJi
VeaS19noc7Vhit4jxPEy+LLc3sMrX/hplPojs+3si5r5lEJT5Xb037qeqkc8v6mo
COReZlKUvpfAVCwxAEpXTrq3xxiOnIefA8YOZlJMQCFx1JfZjXFiF7UzAjHvrR2e
odSrezxVXJs9Sje/MwC1L8lSJVri4K8azbHHJIo/w67+zCVUMARSpe/CDxXelOxm
kL6iZ1JoH7kK9+heCMvsl2JWDoqWC3dOZZ380pW22sj0xiO9QziK/mJ3M4fJsxN1
V8fbl5e/Q9OOO2LUpgQGzWPlDNoS/aWi3XvEGZ8lqujdnDHkc5yM/H1keSSnDIQP
V+6A0/wBF4rcbeslEb8spzzLAx2yGxpFokpP0NzrbhgASHxmHaaNVZSRCD4WRCLG
mnFo5zZDnGMnprcxuDDkjxuFPgdLvhlXpz6jT8TGDhXzn2M/9BuLb1jwLdp3D3Gd
Pjbo9u4HCqQQZprfyeh9JPbiAX4S/9SFiwisvxn+0RXHUUxWAsQFk2spZMvgdQHn
TQZCY4iDxIcnELR/BW3YL8T0tXJZd5THS34Tbi3O17bhTKKfengwqYufdjDeRnID
Bnjb9I32z/OB1E7hlQzRDuS/WWNbcovsZuPmnX4AE8ghox2Y6E4z2eETJnIr1RL4
E1nGD/XC3hNInmd9YPm7kt5myt6jdZzmS3l8chgC9Uh+umXXvDCnP0eHt4TAU49Z
Eup5AOSkD7HBsjkBNZmKA1yWMM2JN9R+fO8l63EjIDVi74yiydu1dXi6ACcDcyTh
e/WR4gSq4N//msia9SB8XOjFBILLeL1YNmVbQumupJb4K9rZHysVj6kKpIwpbJMO
ROrJqCW7TC0+0+sBmVB2u4ZbhZYexOp+eMEiogHkn4Oeygf+zgQXQzVaTKDeAbDf
QC5F7LISq2p7qhv365kghgfNyhaXmz2VMC6eYjuyKNRtaf+QXTJBzXkREgiggqdK
ZVXr6YN3GYdD+J95xf1nWPXJ/dlHzRp0sk4NoFOjBcTfanDEtTiXRH3mHv9O35pm
KgVIr8HJ2SSINDnvCX7qfhCWzY+FYaTF3nsT0KAA4Ex61R1nMII2dJKnTbEVB2vi
tSfxIqaffDfajnnQMWsXPcu+WP425CDBnvVxKFT5yzGxCVQ3uTAI99NbwZW4juNk
mgMcvgCZVZxW4nQyLSc89hn0ggX9PGLF4RWA6Q8tGCd0psNCUBetH8psz/wDGYZP
j9Sn33M8gGXodAvhXfes5kxnj9DXjfnaMMk68ln0qKFLHS2KxGXF8PJNvJ0g++zZ
DmDbvU6nEbR50I24z63gtYtAAslK1hyxTAtDVkb98JM0xl4+goyHPU1SDjIs75NQ
UYEL9+c9cCJytCDrX94lflJaLYsaSXIeB4X4cMmP2taPrLAMqlwVEo1CckP+xZGO
NGibCBRf9KU4ApxUHQV4fFB/PwBOAgqL2UGSTH0sMFtTwGaEtcZ2U8HQUnoHTnZ6
gs+WSXYmTVSCqyhyCNP+hvQRMRpV159xT9SeMtPYsd+eIftaWfsrsgI114wMhMuj
pREPs9i+PHio4rZgK+bXDyhZpyZUmlciFTlO3BaGFQgKe3TiyJCgHE4GR/luVKw3
tRuCHMTzZa88D7eJHfI0HJhNsz57wdVs9mtE37h8ngDVBQN7azBUoA52HLbE4rB0
eQf5J9sCx1IWgv7fXfPjlSHks+FXSskfgVq0vRQBdWG7wxsc2vSqnwmEpJSwzOCx
5oZuY1s4Hv25CqG1v0vv3UUBd/OeWGKkcFX6wHWqNwb7VLP46ofakwrnKy4Y0TYX
23FfIgEmCV3tes4bOEWGJ3dYhTyB3iE06w3SmOtwBRQyujCRVfIl0joENPkxqnNL
XmoOmg9FNohY0K+ITeD2tuxMbhi/1B9b5kXomA6zrfl4o/GkGkSbWCcArVoPt5bI
M7X8UQmUYv5Yzw5NY3sWLNGXGPDE+pCU7NVGIItw88C22BpE9l6f7unZyPrwADH3
ozggT7NLELm4UQJUDSuqjSrFHU536+2TavUzTk4UcbToCnTSSOs1Ogxq5p7oTocm
Ov7hO0Y11zpixuiLU0MkzMrrvLdtaGfSKo+FVHW9A3IDbTT0dQFRTykAYVanPpwb
VjMR585pTzM7NQC8WihEW37ZHxhpj1fWSq0bpwuGJFKEj3Iih2nlnchkaEs7keA1
sWuHnsmfdojzJyyXgfPiJQrQhVNECEkqtyQkjg/1FdqKW2OuMuR6okeUSSspOmvG
4U+a3tuaaBnYewech3FwZm3GwGT1XvDOXcHSVWnjd+MtmQCGFWIscgvEJB9Gtj3p
VasG7yuaBIIq0a9KjGaX3Ntcg8CmLwX8it3DKVS7tT2OC4JUlpH3b6DJy6ViNluE
gVcOZjbN257k3zfkOWAoHCy0Mds437iBpN14VxJJF+6zbdVEX7Nqml7nY+3TK7IT
5DHX1dlSp3QasA2R8ekRdRTLQatj+u0iRQJd79W0ITp+NxhHyByNDcyg0d8KQzwy
tADn1YenE2o5RoYASOZX7Rs8FGeBEzaxO6BfditQfXxV3T54OlrFwVemice109+W
BBnyBNNR+FkXHKfIhkvOawjZaDoD6YoKdy6w7TtxhS2r8Be98nUQAH8+yxvp6ly4
eG4pBWUppA5CZbdjvBtXPRhhco0Y2L2lSoET7OgdNBUiRo+hR6ato1GiqiirefMe
/J7v6KTtMI8TG1lZPEVHqaaeVoPk0McTYw8AJLINFi5aZLrC9RHFx10JehN7a9nw
w2tfhBRARzJS8Qra7Oiox5lJgvWWj0qdiLUigZflFaVKGTHcHRhfXu4+6hR/okYP
vrmKDZ7BuhHB8SZ5vZbleugALWK12WjV9xuunSX6PtMdluRC/4k3+WH7IdH3Bvtu
gF4WAjI68F+stucTGwNY+3nsiXG/uGuyUZVypMiJYYXwJsucE2/fOwE0NcMEpLvs
J/zjTrMbcPgyktdVX3JH2VlTW1ruB2T0/nLIdFxwM/MdHPZv8tLjRV6LqYMvugZt
xQMT2bVJCq/kJkY5B2KIvswuY9Uh3twwcB4ddadm1chWKoNAuZ6LCkdpaFXo+xQy
zdil/u0mGAvS+8pIAVp09mSGwujGzHSZIrSbVRtVtTUlssdBfvIieesYx6nAhQX+
Fz/k5TFenUv9wHbDNKTydgwHktH4tIh7yncGjE/CxreNIqyP9iFmHGXa/wQLsKZO
eL4VGOqKjGEwceicUL+Bwx+uZsw3DazpaBIXxRHWhjIEKJeDw+EQBgAC6GAeVzWH
qmxzzXWNdekN4TrchbYveqBdn02G12NVcQ5RcroVVzTkakqo+LrQZ/w8+XZjTsti
r6U/c+A4zHuEmReC2sET7mdhsBvA4un5rZkTnErCllhuaJox2iM2BtEOX1SnimmM
k5xIJf4g0VWRitvLTiROOh32nfCn27ZNnFPKLjRyPNsTRYE92HEZzMuTJR4eVd6K
yJJPVNu5P+tUvyhF0fpksAsxdiepydpS+ayiEgw2Fm5XZtWhHx6LyRth3TzIgkek
3JvvLKyo6YtKSywo2JBrp6vIOp82DwujEmAga2o2VpodH864A/Au9vRkP4A2HdUt
hOQLQX/5NumFfFdPAqcEtFf585KD9nNX018rWXNyzgnRfmEFZU7Dh/jS8aQD0Otl
F01zgFLnJ/cyy8jmV/Cq49qXGjK5kodeFZ3cGWJI/IAAW/Q0E5zeGYt0gJL+X9tA
8mPWeW+ZHANVdz7jZzgOSC5xRRhTT29UySAeTWN71UGTRW1nUSCr1Q7xHM+Ew1f6
yLCycD3I7GG6vaVBM/BkKmrPEkOh7MH3/9dZldnAvs50pNLI32Sy6uuFJFzw1Z6H
x26QjqQF//B68VT9lAmAURSQhak+FPSdfGSRAx6ct8boQzre+Vo4XPTW0SwexjXW
CcaiAIPuMh5X8qlUNntgF8s3oVeWZdephGs30giH5GKVeMMF7nATP+S6oUd9D1k/
yMGFS3YHdgfrPKHzkq03C6ExdY+7PEYN3UuQJJpvszrgUZ4aIqk6SGqDmFInpAhM
zy9PUWgwgt1T/EHjF2AR71lqFCsNmXLwjtmvTXBnub0ofKuIsfU1wIyEenGMk72N
aFjKokSd1Hxulv73fQhbzBOa3LqNjR508343KEOXvraNG0rbGOZ4XkJJnol8EWJ3
Bu9bjsOgD1oMZYjbasEJL0ZjruGcZHM/gcZdOoXWsq+zCTxAUeI2fcJwfcBelHz6
Hsy9Ahg/iOnbexnGN1TWukQtUVGzsszVYChxuwuErc49xN7ASyLiP246ECWDXhMV
+tNaGsVC+rY7/QwgJW/IG8MQ6ZW7Wf8DZpgoVCi/B+A+8ZRQyixtmqDoRtXhPw6c
kcn8F9IhiPyPokmGylDHOElinW9ZjWrvR7kqstrI+gxTSJrIHFx2LL+c3w56jXOv
Ij++s5OLWz7ywv70qI6F27fJPg4UOlc/8NYPRC5N99bpkIUfB4y1pOtjEgI0Kcu6
pGhEvo9vSIN4Y6i4kAQajLR3nHdziNJMwerTosFbn/F3fiMFq00p9FmekQzyWxYG
7t0jZ5SnZNJRgFLwnjZ0j+BdQ2XLk6NW9W9srdkNk0P/1/+KPtgsHLX+0CU9RHlT
1Jd4EPz3sN/UR0NrbSuWmr5JD2J//sTpI1dUJLRQIVekbqdUXM82nIRyW28cazaW
nKKTZsyW1uO78CYjrVNs18Qo8iAyO45Eq3RQCJJIlY+0n99UeeyBwBi2oKY2FJpx
IMoofEinK0lNFme8XfnfYUP9rE5rVvB+qln1idLOU6jtB1q/ObS7MP8BjrGk46ls
kmGAQXmYulBjFI9R+FTHBx2g/0P3Iks8zyphRGEv5UxD8WkF9e79cq1DiFfL9jRz
joQBki029D3N1xbZIbztrr6dFeM9IweOdJKO6ngMbctaajnDC/FTRzte8sLCUBBz
EbjYsiuPn8oGlvODuOvpW6C8mUq8gXKsIpG15NSJB2m3ClJjl3hdOjoTvmom49Mg
uM4rhu3tE/cx4ddCX+RLgqYMpcXBkkmpfotGXrG22RHYFsMruDRwVK8rroNT8aXg
p9wzmaL0Tv8vpWwdPTJE+lO0iWZwEsMtK2umKWfgOpAyzQhmIBrzdD1OjtTUC3u8
1D3F27gOBj/ub7+eARrbhSgGfAX1rsXCP5yu+VMQ9qfO4GIaWe1DU6NglWWyLH5k
OsyMorVMVkB3vZykBaP0mfrygx+rVjpUJB2RFqKp3sBdl6snBsZzIG20SULbK/Hr
SiXBLtQ5w3ChV0hYvD8NVqnOkZPyR7+J+yIA/okgzIfmDiJZFdkrR0fJtPOmwgP2
MaItuNk8Yk5t452GZkqWveEXz8th1qOkoN3Itcy1k1DjpcR/JAms7o4PSqjrpGpg
jYb077yuODhb8prQ4RJOUtOVMjhPyWE7EBAq7aMH4uMQqjxlazWBbcAdR9E9aVXK
Le7yUzS68sCGysMMvPl1qDDhw4HnHTqi9CyumoxPBNU3gHr4Wh+nvssvjzSbgsCU
CZemia4HqbTDECykxrTSpeFiLS4znXyPRkjBCCg01QPL1KDm7kFBDbqzjQD8KtAq
GgxXpDN8WLTSMmIfMznWV+WDmKK49vVMwyg2Nu/FfBVUQcLYQ58PIwPRBEMrooei
tNSwdwQMbPpf18tGk21YJolOFhFK4nte2f6ZrMIv3dFTRQ4fiUJvKq1GTvpwBT7P
KGQnziIolgLhse/Hju6BhtzbIHDp8phHU7rmdIvTtSK8a8q9BhMKSQ4MVYjz5usK
GKW2lRcyDwdg8QSu+d0XBXGHOo2lZpbbCOxjLabyOCy9uVU+aD28H4euDAvXR5BB
fTxrDxumqvlT7HIvS6YDZZ+HVBhp1eXnZCF2t5Av/7C9SUgqHKF51PFt57Fu5cVm
YG7LB+hTOkEh/wP+1pPsMKujTfbkmG2ZjPFI9Vpi5OgINrwV6v7l4cQ9pL+3cVsq
NmLeo9ala6UK/Tq2pQGUeeBMqmckq+zfY+XXnx5d7j7A6kahkACYMvnRNL2Jh90S
yKC/oUIkiH0d2/YoSUunhyxtMxVdRLB4PfgOwio89TEeZJWuZqwRixGNjlsOdJ6z
3M8k9EKjthw4xyIac9ulxQiNJCgAOehK6hhcKiKsAWqUAqu0CtHwNGRX88Kuzm+J
LqRC5GHMxfC0QfQJjib82Ex/5WmU1c7Ny+HGNCv1/o8oLd/6npDlKILFYjJg3vv+
+zxO5mTMR6b4QxUAwFWoflyO42VwurwC0exvAhwWjl0XYhJFBuuiDqRpB6hSFzqV
o5XszzIPmsQ/gm7YNzWX5qMIsn3t9uUzBMT/+GzxoJY0bwjKoLTHpZC3cUdHF4QS
aKZC7H6L+/5RWLjdkoAhqewykIbnvS2Y56mWrpnAyvhGCursKwUcaL6z+S1P7/1a
4Zg+WWtX0C53WSljQasAf7vFDyZzNB2DL6Gx4mAbMGQNHzdrGZVL0Ku0irblNWqC
XM66SAXOU0XY726z8nW+GAKSyVKoPfsMfSaIXs4KjrUNZGh7Mit7KO9MB5O/76Eh
Ia192ZdPSoB7IXLnZGtYl9VlE7E3KM8sVoAKJBzu0nuabjMghLSQCQakPAX/09IE
KQG2AT/aSvcqx8hzj+DHugTYarYmI3auRlyYBbbEAiG89OBK0WVZqD+DN56EYWIu
DnOXM3dzhUKvEqVgqi3LUQZmpreufdWiIKlvMYt48E1Jk3ZJha1hxa0duaIFIrQr
fk8+/yfrkKSpA+ox3ipfPPUEd4uFbeGcqxKzCQ3omK1rN/xvm2/BK3dKQgYIpd18
bc2mKgnJHy1Jh3qYdlyMIioJTMSS+VEpkf6gvVzXNVxIJPl9sRjDZ/ZouQURGKdx
WNiCQ9mGZpuc9eBSk2L57dkyw4iYz+zUAW2kXaebMrJj+f2v0loIzjiG86c1PjnP
LJ3n1w8R3ZSQa563sDM87pJja0lt3kCYhnamFuJGl8Y8XFPhyHxeB5ueSXugvGmQ
UFDRyB/qCut0NSn6H5wqBR7i5uOF1vS0sZJdmn34lT1MAde+hPF2rf/YmON0iOPX
tgLICl2TN1pPOUFKc3j6vEw2M01nM4jDeeuh2SVNNNdTxBbGsCwEg5lTIS8e/4s6
2Qn5Bv6rLDtOHTURtr74voEYc/+1IjSajlAspUL4yNApKBB8UOX9iU7LXZJk68Kr
lq8akoJ0UUFY7u7QGaI1QU1RS1ELurVJqz8svItpEOrLn0bjzajp8EiUwhMbHyz9
nEd+78sRQvLwADi+Q0oAHVEQ7AWM6wm5LTy5U6YkaZqUpLubmtYh6LDKBZHIjOEH
hMAGc5lyZCN+FxIKR2Oot+pKELoRB+pWXr7Ix8hK6EV8lvy5a/kOCz0vi85QcpXv
r9ICZt80siFi6ufhPvQgs/S/TbJp6ujq/ssoynGC/QZmlSOTGGFqfyO3D7iIgzg6
Nv+wurXFC91DpH2zkt0/1+rBbszcQr6WvKcB/F5ghKSuekuxFy+8ji5LR4f4P6N4
5AC7Yf58CMPM1QuaZeGGIAiOb1X/qBfjvKn+C8rjMp1wiPLQL5KYuqw0MW5ALv3+
oU0jLOzDQpS5LMZh+1xE0q54GuHLkYFk1IPbqf2pA+iXF1h6FreKjsDNkDdUv/ex
GM5/ydNCSHIBcI4jseyEZC6IqbqBowjqJj8gVFdLdNgDJ2DRYzeGHVfLMZMVQmNX
8Mr9dAeWhBfW9E8L8lgFkAfVYEG9RHcBdAaFHd2YACkmsniKsclMDmOpFCyN6fcS
usHhZxW0N7ViZP5oZPnthPFYYxsmaYGMq1jEUdooR0tDPELiWou69ZeNqCigp55B
DCSx6dokzVKWX/YhWOvvL7ogdlW8ASYyghZ3fbNsNRrMeDhBLPwi5y30nxSkp13w
aCT2ezcAEnNfjIRmA3takfWDW7FUbh52DEGiSUnMjWrRnxFB+ik5RRakz4XYFxta
4ZIyvntZw+uwt1+U6V+pNLmJAc2/aqX+F1Ln1qzgq0WlZh9omMpRuu9s+wd4LF5M
gdmdVJPlJiBpyUaSwC9kX7cHcoiUYQBu3dhDNFHjJDDlRpKpuzmrrVtOeRT18Grp
uJrjh9qBKTqrrLOH/iNJvpcekAqZfsu+LAhDXr0Z0vFz3nZzX2r1oy4OIO8Moun3
MrlCA0vQt+JNK9ydnffdrYX+u6FYgethVidTNwCglREuDkl2DcmedsEPS4lr3RBS
l7zO18jCRBlWNMt+XCkvRj94xhSWTX6vEGDbjq098XwvU6jzbuiWFMSRl/rpkjcQ
YfMXD8VA/7Nm0EVKgnjcTPsl6cYi+7qj0yOEDXtz77w6mRsaxPeOQWBLLD97T1fR
NuiMviohLDM9ytZp0HngVNXv1/3Uqw+tPl46ThpvoCIjMykrisG7NKkXqvn1jGix
xgiR6b8Tpd6gvo8y4pirPFBrQAUKeBb2xYcrTw4JWCUzPA9yazNrDiqmoC+OhtHb
Ylk7xC+b16HeO0uYe6R/L2xTvyiA+MHNC/ZZBQ1Oc5NC1kFUr2oH4MLupgHWmFLq
f+mHzJTd/hu8X2bJ/NEwvP3Ag79w1hmZq4AYuNcv+eGD2aehrm0G6mXtlCfPyMNA
B67O+r3fLWoCONElHsliqh7IVEC+Zoj67+lop3DuIMfiLAh6CEUAHOqJ9M1pFr8G
AATU8dK7Kl+aiRr/KWGA8FYnsB4+WtVJ80PZR1LqfC2hdIZQMQsncH/DIVfWmREc
A1i2zlJ+GK25h3xkLAaIrJ7VlRDNlWNjjc6f1IKtXwkTmMfgJYYPcXiZ/NgusMoV
KEQ/pU4gTUJHgnIIJ1nS0ykrp5YbOW5dye+rTSaq46BNoF2RrKC49JTLPMlGixVq
3U+abwsrAzOAcj2gX2t7tFxmNO4ZJea7FCyUVCnzAJzm7JceN5ZKUrTWf22FWAFj
WOvwoThiXPXFixLiMz5rzMS3w4gPFeGSyoAHueGVUqC8j9I4KbWPosN+8AdPZMxM
/FEmm+w6AsxXEPcmpmLZ/5w+KrB0XULtTwlIGui4AyeO3lRRQlFdUTlES9gg1g3J
ux/pAm3M44qzIeeBPDbVHfRxnIXz3wI9s9p2bGZdag8WsxeLmX+VXD7I1GHlTUfG
D4a4gP/AO3zWFbIzThai+iM2n5k0R22x1/pH6W3Pn6C7V14uodp4QUHsW6vJC7cZ
TWJ3FtG5XulsteWzcvfqF+XYbusEjHRMo3kDwWHWF0C6Ro4NIb7XlQ8B2g1yEbxf
T/bn4mgFlkkwPguNDgVO95xHFO3b7lgAzXamwQ3FKvsesf0kfOW/qzX9fyF45ZOC
U9GOIfN1JlEcQ2LtVOr30K2tQgeW+Q2I/pCg5dXGtZGOIXO0zeszd7y26YHjqyAv
SYwNQbZhdCMx4bxh9Vch5RGTAYMoAjkZ7fmS6GH5TwJg9CzveYb489jRSKXv2xy/
KhavuowbCKwZOnov3PDG2lp6z+Dt9/PZ8Rb4GlN+5f5EPN9QM2/7JqwuSu9asxqI
+fSmkYYe5M2d/i04io47R91B+GBexwuH87D2e2z7hBR/Hc1R7sHXu9sDIcqgYbX5
Bu/dL/8NLnW6hNXZ3SvFqEy0NANmdl1x0wg9YleJzIKCF0LZG6GSTPMVMc0MC4t8
hhYp3thPVjWel+K6hbOmA7Y5VV53IDLloA6ZeX0RoolPDmEQfsr7og5jevmoLVyl
KHR8OYwzck0hFZ2boFhvXzH0t3YyyLrlDXXSC4uoHtQgrT/jT5OY4WDWxCZew9qy
12j4P2/K34Wjl2cnK6h8YggAs2l+TDgyuIwWdsUqRkcovLhrKemRCtRsvYu6rZR1
sRNgusS73QiCc+M4yP6vsiiyqWWXZR0I0BtN+PbJHKERTv1f+2f5TYe/9spwj3GO
sK69+2dc7NI3fu6nUdu/0P8VrSownaFfGu5qIZ0MgQo/HKbYRcRZLRACrU6p+ldG
3ibvhUmoJ7ujb2RKKsrfjv/b5FLwOWa3LmNw5jHbr+6lyQV/L8RwvbUTeStz9RuO
1lgj2bcDmy8mn8nM07G3eceYeSudICQhDstLIxHUvpX0fwCc3GYF7c17y37Bqunq
yn4SaE3pwdcKNDr9lD6KD87oSISSu1kD65y5DQmvPfbHIGNpvlQTsS12woke4X0e
r5WBUdjbHSVqIBfCkEZB0QS6Y7a6QivEXSjdSUl/J/KBhZhgy1ZJm1yGAMI5Po9v
ee5MC4ANZnmEDMMKGlJMtA78yZI++lc0NLqgn6VXx8Vx72VAE4eML3nfzA130zh0
TxiJHWvd84TmPwwvZXcskA9gC0FNP8U+7RXJefMvEc7MdxH8jRvmBAXnHPE9PEab
EeyBRYfVLQA7G8xMu/CThZ2OafoDc9Qn9auo1A6G95eUoyofhwfU7lyLgq/gXvB5
zBg8eWdWzooXQCXoVVHZWrEnNoWavYpjzPE1MAvRme3c9KOehyJUU+nR/vJn3Uc1
AjzSqkCHSfRftNhqzydsQfP0leSVrwT5WPiN4HRwRZm7kCHJFk6zr6e9TsP5exgo
xDy6Fxmuf0AGLAOTXrlQ4cZZhcCB87w31sXZjcxv71KqbciBiAXiEtyyRmSDUZNC
0L31qsHJCFzict4EQ9CB8JKyfOU07qNRFLeX7s8e8QQ7zqD6Dry0603REP0cUy64
Bc/pnqn5Xd3d/PVn7qOmmAPlQpjMFUwznZb9N8Tg2Ic2Qonw0zqDqmOGC+NyVZGc
b2J1h7mMugU0owxWquy+B1lVYh7G/2tXiJWjkFzQCesBnsh2ZmeqR8AGnrYGEOBd
/pmoJB+hlOB65m0AuhU8q+jMevJJQ5GdIGeKWv80RjMb7+gAPm/26wJCfuEmZHxY
zi9T5PzQzFmedaicHF5cItfsMXmbfKI6xwbVsLPTg0puHpSRxTunAPzqku2HWBpv
19RG+ArkhSv6dMXl+ix3+Je6bd4U980o4vPIjGlOStQh+M/uAqGfN9I06u0NiEUv
ymLUBQckpeJO73c06yE+srsLR9ZAgcteNhoaHFClSxU/IKQ/O+Bv/kY5T+KcehbS
7fk0p7ku+6SvlMVmCJRoutBdoeLY6qYooNbU5CUrYNivOcPHe6YvZePcmQB4SiIO
gSvLjhXfhMW5NaSLHZTxOueV4NU9i9WXcuLHtn3WFLzdUrb6U0lKty/mIe4J8YsM
+4ta8jKf4gs52okNgKUZavHP4zwwckHkHUhsAwo+LXEl5yEP+P1gZqSQQYec0W9q
88uqHx+TkhmNxnyr4ICre40NbOdiYdB+rBTR6kVKto7V8w7h+I+DZOxC8s+EMVqY
SVmn4r/gqcOeOovsseVim9SK643uqsqAbbJS6XKpPldsEzQoqcI4/EKQmYwRnpvq
vBMnqCzXP6zJ4iBslchNfNZiP6S9JSKAA44WCGQK9T+2VMeKUGUEUv1MDkL56iSf
5k/8efIAuWuJGOQNuWQEAOj0+9kT4B6AwxR/eBHsaaG8VrO8j5orkA3b4w4AI8Aw
782WOj4mJh4AYgHTkv3npoKCGNyPUT8QrwVAwOyT7CaTLKXRk9UcILk/z80r5zd9
Ca6DxxpVeQdJUbs9fpslBoEgJsgeOguVLqH2BzZPmHEdmJfpRX+C5K55mJqSJSOM
Xg89wyPjATVeWH3l91ZjxrweR+QUC0gFm6QgMJwKfWAzcN43c47PpOAru9TWW8SR
4zi21JRZrLWSb+PCyQorCd2Aw0r1t58JDjo7Xs8hGqbFCmzENA/dGVtZRLXzNHHl
0tiNS5/5ZiqHbCLkbWI0zo4IPgmPz2ag8rn7NltOfHou8QtbzOOk/x3w1lArBKiD
VAIfzoDYuv+WqmpEewmBXeMFfEe2RZZJfGU5qQ/iu/iLU2JKJ7NZAYv06/kVTRIi
21vTLqLX3h+vZvEepTNMIUOMUbrr5u/c8as4q/lt7yv4dW6Aj276sSjsNN+IzD8n
2pelUiSb4b+/XOc2Re6vuQcPI7WjgvsKfPg7J25AvZuZbd0YOltYQO0nPUvnW+Fa
urMUnF3TbonhvxZaHv/J5uPtEzNXphe6h/tGAkq23oK91u3s9r0vH4uJrBhTgGtD
Nk0kHNl8uo5gVuqvJv8C7RHi4gxS8pZ8uRcoVjRA8pS/XixamGLI47ppD3la/iMs
mgamqsyPIAKm9eTlDgWTUGgb0xGg/N80ObYgWMoytia8G/jrswQLvxxoI8BzuTLI
UjsMpwUSatdeOcJrLzmi/QZgqa3c7S9QTQ0jmgOeZ6UN7fGSBy0Jt6ohjQJWAqUo
7mdPtM1A1PmVN1xzLZUUn8jqembq0yDsRly+/3hD5gKzdKlKxj2L44k9v+BTVMC6
lKecJRTQMySUG/0popD2otgzBdP79qRP7XMv0C5n1kCNxqY5608dITNEDmmtCgkp
/vatfI1iZa0bOSdx4jFEmw2GM5O7MLbhsKeYMqj/XYUs58YPG4CEY3C+DEDS9rIG
QhHp8sciCq0N6WNXwwwEsKV9GDtY9AFi7wBp0rXAhXTYr7DNZVKnldWDPKdcbZHM
AKiSr+StFXD87+X12UTIRiayQ4sDdJ1y6UqcxMxlJSE++4Iy0rcJKstlCxxvYqrH
Z3hAf/v48lY2TWhNrCvxxpiSZ2kPmlvfQzdHStDF5L/NA1utLcA00YBYgN65OhUi
IVIRCvV7t8lFMzijp/e2WzwbEmKwWgnUhXOzHshSpmz8T5olHiq2cOccRyE11RaK
QMshkpBEbGo70WYFMn0ICWlbnvq8SiCVNGwgw80yn/ji/cS8teJwf48KyQfX6tST
tn7WgiJX2A16wWsaG5PYGzUXPwgE+Rgpnf1JIJa1XtDjJKbWMZ+rUf7T/YmcbFE7
GwxauWMiktiJJ14zTo3mNJtvP5NUtcnFhOG3l0ya4hw0Gc+5KY/T8bhSNPXUulTS
Nj+jJPJZvD61n0etWN3e8ewwqHfvl+IUJXSsZcQYG17rTxI8VNHU1vsVXgxqRxRp
x3Igyd04OaHQWODqYWJzVl2zaCp4Wz2HLFJAFjcZhmYQkd52XXY9aSCN57ZNpE7S
cdbKOG3MKUDa+lhCXSc5Ht3xRo5EA0uDWPfKNYlXUBCIPVWXpklO9IHp3nAU0MVz
1I/6DSG9PMAe79VWaQbgE3B6YM647mWkiuxwwofIMQBoglwjWuVNbPCYWmjikCqB
AKnfY3pD6HL7yTVQ2ynHQzTSJmDgZ0KuZJd+OE7FeMf3opFYq5dsprjQqLUdf2qg
2SaJURh+Jytn+Fa9Rsd6FdCMvmJ7a8lOMsA1O+8r7PaN3Yu0uGHJRRKyrhVbN2Ug
abVgGHmp2vvu93OYh5xo6Mlof26orSUHrJ7chZg6hkHGSAulODKY4ClVqd3Y5nG2
oPNX2XvUg0SZJdOVLGLyhxLZKT1gppIhBVzBG8Qs8TgU9qT7NAc9o1gJvVOS1OVz
XwOj8mQIrYZmuqC6E21OxC+RAHkJ8HHhHxIHwqwmzk2M8Te9SgYn/St7/KZ1F3K2
u51g5PxUTWssHhwnWEM71lPyN0IYIo1tRJEMHreHu6bqJO8w1grL1JJudL5C6rYS
3Aak5dcUYzMwAzOgcooet0BByDX7hXJNzLiYU27aGFPTogut/DK5ZNiJMH9SYB7a
GbFMGX3pKsHaseFDmu4527+kW1TSpR/iquIwrvHsasZ6kmmUL45Loa50M4qtlX8l
Se+TGt/xPOszhqNWkdqOJTVbEPEXbh1/iIq9We7b51XcW2vsowKY3NB7hEZTVV4d
C/jk0Qos0WWXEacmV27daIfW32UW3Rm/219rciMG+FCMd/d6Zo2vVS3l6gbCGnyR
N3fbu3rlBzMOxAbGA1KbQsBAgRtX7+dgFlvjDxCntouhoN0UJJsXPZWsJceao4Rn
VEck2RYiptYlEGrlEWJ44DSY2FhLHKSt6bmksZRtsLewSTb5NimN1COXHYR/A/Ng
gJioHFQ8g/pt5xCK1zrDlUMqZkIB54xJVE58uFHVL80yXp0U8gLtmZPEg7p20L81
UtWknxyjdQCkux5ZmYc5Ul5Qg/wJsYVV6DwA9KvwYid6asBQSR3LRWV5pWZrAKHl
Uj60nqvf2POV/CXtLu28AO/e1bKRxzk+bBbPX0YzRWGccPqHQE89BX/H83S52Pu+
/X1jCRvkDxzyAhwtnEo/yZyepIeCAoRsDcv3mYe9aqbSo5vQt58haIBAsPSDceW7
qHncWMUHitCwzOrSEmVIXyvGZ2Swt4awiHV7IRBaBek11VL8UV1MIFBxkQGeV9Oj
T4pHVrZRHo4o+lJ7eutZvrIJOPAxCDWS3kInZvd5cM18lHng+VbZUsMR7UcKr5dg
q2al8t8oKEmaQ/I2rwgowO4iMXbpTxYv/e8HReoX+p54Vd8e0FBL5mDyOuqPqHqb
MUJ/OdvBqc1ftoIb85tndLHmiyu+1lUCST5fMI+2EYtSCKbHJUnsl4JmyHoOsAAH
ZsNk2y3VEywLm59M+RuaOkD9gE1/v79DeUCb9mz6IyyNFS9Q/yx5+P2gpZgxBru4
Ei7lY2VEPThMogU21+X6cnIDECj5pBoE/kDjluUSxqNa45iAZAOs1WsrV3rkrk4T
9xsHx0hhc86ytJzASOS/+LchSdxqarjNJXPyx4NLyMiNjXeJBUsqEorfA/l3op0t
XYm3hqonC8h/fpxJTkmFC+UqQ8lbb6rrCWug96De1JsylLbND39h1E0K9ZuJdKe2
peJksMuE8Pqkgs674lL8VvsHm2JoxXP+SG9Qhl9IicmBZe+Ro9dvQ3yd+Wd9Ar7v
c2OAoPQbm6SWmMI0VQv56QC5aSlhGCiJNKIBbGM1EtsxApd5f4i03KmV7kl3/FQo
b2thCDV2uwopOWKBXDeSFwnEdSkLnfpswDiRxugRwTff8ATVmhHA+FLQzzICvFfg
7iNVMQ202bgYA38oZtP1wMcULakRyicSecyYHbrro6vcbcQKM43l1KsfMb4v3XoX
LgP8lmrZdm8vX9ywhKItrZtS5POOmJJCW6Xfi9VFPDEglFQNDEiSpbMZb6nCWc5N
42EEVeTztZrHsTryMs7l6zGOO3TOwtnD+/61sO0p85iFuLxFZHSia1H5sHHWExS/
yGUvTtJWOIKuDIZuEu8dxwidqKNTXhDm6DPerHq59NCoFlgYaqaOVlQpss8uQpOx
AF5XApiyWHrC5NQIn8C4pxqYGvDkVa26yDpuqxvdH4YPgUL37sKowvgiIUge2opx
W1v8HIQq2iPr//LFqXwa3fgXIGPjqbYuXTLA0HQn2dh4AjSPRdeG8AGj9h64I7ww
wPwecZw+AqVlqNLVtrfHnftm/PTn3OcmcWnzWZV+Srg25sGyX49KDfHw9VTFaGzZ
9kgB8RlDi1m3i+Yf0Ary8WZrNqzxrgJYMRDwNY3jbKn9KW/r4izEjybWGtrMO101
B+buB1mdQeQ08f2OesE1zy5EOgUbpGTY6TFecR9Hm6a0TCsvkZiDR7UkXoVtQ83c
bwuRapUcvUHTd9H0uA+QnOD9YUd10QG6BlL52XpHPzh2FSyd1d5Die870vx+NCcg
MD/ygWrAweK8L6TXXSkJACUg1MKDeDvNE7Ta1rHPZB5iEIFR/Rq6SrZN9AMmSMCF
hdoVRKKL3FCMVskK0vnUhj6W7GeCeVsxKi4J6ZjVMJQmseMnynF1AkTt0kxROgC4
FumwoFvWIO1HA8TpLqA6LCCm3o4AaSPxUPQ+/4U8c4DkivYqOS7Y2AZ5L2t1nptP
DFskm8h63MOSLe38SWVgNXC1+9sCHs+73T8e1P+mCCiPApNxbfFvWhbnudp40G/O
OLI0aB/sZx2fSry2oYA0mL8/2SIhLYskfJGm8JwTIB6i/vn1s8xHDxFrMVT85bO2
JfaEARm7T441yhF7/yXb5bNCueEuSL9Ichwh9eKCc2Xk7dcawkl0hkusVDK47Lg0
Uv5b11BIfq6hEidHgsjB7u1VqYLmXhNtxhm7+PYHEmRiCsQ3Akg6T27QgUD7Z6LB
8OW+P9VH5OXAC4MUMMjShJ2yD9YI2OSovI9II4UO+VH+qXSxr9Lmbs9hDC/daABp
QDo+Pl1Lddju20IaYKR8jbRgsAtg6cd2tfNEtfYzKpcSSCEnZL0BcZINI/QjuLbg
cKdanSTt6Zbpli1tyKWJdAW+3OusnEK3pTyI/qqpD34npCf8RVfgyxpFp0/J//Jx
RCo3m9/k0ohYvKjQ8XOQBgxXh3Y4WkcnIbGbE9ik9/lX1fJV1SzbD8i0Ri3/KoRl
VaABP4uaMkDIpMCptziDwEbMbzxjhdEs1qYcIwxnLcC+ydp7v32Fol6GU4AWenyT
LiEsAqPMQsmpsg83/2NXTt03q0zh27m87Jx4GVShhLJfWvUq9je3Jm6H0WJokxsO
OMaHuwh9a4s+GW9mzfQWGh6G5QzNtqf/CfAWRTkJv27N3p106zITW4N8bkagQnyP
TXjukJxJLZ6OwYkX1ZI+FIiK/BzlIM0wpPSssxEbOGALlTV974ivbDfzZBNI3IHG
i01VeZAJajtIF3cxtz/ZTtRBAju7cw/8dGcD2tQWbsJN1vaO9iqTt60BHK1V1u6i
swKGc+tM08ZwPfpLFGuJPcsFwDIvY7qtF4HHfymMvwZdduhyIJ800+GuGxYJBLsq
CK4WcVcya9g/3nzL9wm6lz+sk4+5iV+04a6VUzum4zRf084PGWdth4WKSFLDqyJn
/ZMlQ0Jsh9/lcIvGDINQ6JvTesgk9ss5UxMIEAQuHKJjTjPjCXru2HSHETBGkTss
O/+5Bn+M9Vpgqmx5Em3NqsIk/NLSUqsGT8ikGiVXJURjXIxDc/JI8HcnkQL6Pd5h
aquEzjwYteeTZnSGFQSX+QdL1E74eFPCXZ6LwoETKVLCD2+JqS2wcnUoZ9ViPYTm
cbaItBJorRYqdXZpCtOTZikFelONF3FFfgDkT1YmVZqh7aBGvOqtpz/PHMVs3eVL
w9kgEoNcH5nKmQSZqkRYEr9kQeFv58fjQHQ5ZY+ZR5KgCtFrxKoM4pCvfnZMllDs
YMiL1bTGe7/UNAziyNvQkXZ8aw6TVAokaIxAllvCZGjRXLOerBuPaNIp8g+gqHDh
XZkNeqL5nVaP1Q8QSgl0hDppPUZlNc0TfHeOYT1I6VUzERSYSNfM63FSPFsyCzCV
FKh7juE7CLBloRe4PiUmWRcDrTJj1sWpEkps0zLwcwakmBH87vwVQ17CufX1Qglm
SlJs8iI5jsxi5MvpBUMkt7V1g+ADFD7itXPKfW/wlXqc/EaEo0oh2zUkZspk+Gf+
tVA/CVbd7HvVFfXU6FYOBQpfXZIIjNQtPJPk5cUxwNfY6h03oy3jf2fo4q+NxgCM
1sJx0uJS9/3K6OGzcA0V8TJ9GGAvN0XeLexivnqg6Pwnn6qwmZcwFHFTrrIuiqda
mt87X0eEyprEfA1w3ofqxUU+IiLaVF/cTx5hmAh7FWEYKriZw/UHfHJeUe3jmc4h
5kmSrHSrDdA0wi9zc3B0DyHGtINjO/+xWz6TabShNduL7herVfD89csS9VyKAFLV
e5tm1JEEwDRdnchMpahaQ6fLsi22+VR+5Ei4jTgiz3o7YV1wxitwA3Iss7V5mnjO
qlf88TLC6u+2g8Gplku6CkBvL+lnx8llAmAr1WwFDm+RFedfcFZ4GupvmGkoEnyU
8wTdkYwt/LODDZY94i/otuLFhK4lg4XM0DvU/2vM9v43lbmAS58ilLd2iWCiSJaf
9dFy8XXGgT7W8YMra8yVWpQW4P3UuXxtE1iWAN9bCv4m2yU+K0E8QSMqKvZ3Qm7/
ju7HC2+CmnQvQBhCv3wWnsbyEZBn5zX9UC1hK+Ik4xy+sJwx69IQay2RCf6RV1nu
Wb0+SWv0cmxAbB2MnP3PPeVoKep124xjRjniWit5mww0dDyM4DM33Xpo+2f8uaew
ju7iPrri2Mfu/kyH/UOVV/h/bqMQvFb6vfyjrnFdYkh3xXluFYE8mVgYATC2yRrD
6Cwx2Uvf6ASHTH4O08ZkWy0TDQasBtTPYckkrDty+x07z4wUltiqUDBz0qHZuI04
Kfqq9FWCplp7mgiEgyo7//mGP+5bOSa9XjrkrgzhtTmqVvDEdcGGTyTaVqJJtCLH
KvUfepx423bC1iSQm2V0ZaIMKl0mLRN2qKBzWudyTNPLJzYOd1aIfa6yl/3cFXln
FhyWyywUlhJPDWwGeZJjhQ1Yx9JLChbIw9z/No9IAdr4ntCGUElC9SSQoojpP0xu
IoJsMZbmMRdktud33gf1a4JT9XKB1P7AA3V9N4jIAqjG0D2uHjJo0pQQ+AilmlKA
X1Jjwi24rJJ+x00UTTyvZYQ5XH+MwOExPawFnWhIvSEhWU4CiQVoPRTV6ZUdWJoi
AyAC/t1gyyEMloX4Wze7GYWxzVVW5JIdmgRiNq4JparKdsomJqzznZe0PpK+k13A
v3e1IPeOKaZSf0SIRzaW0VD6SPcAOMijwtnGUxFEdHuf6vteKfgMke3f/1X50O7q
SsamOcZ66MsY74QMqdIM7gemoqOB4nGI/pBm/RlgpUp77eNcSjxTD9McT21MSa2V
YGnTWvt/lREe/AJ4tqHsuaO013jr8wPj1K9mz4RqUkipS036GtciB++KieQulJSh
iF4zGXfKQzNbDCJm2iFhxxf9YLfSTnDqNvCTveK45bE+f9tHJ0tDAdSig9Rga3He
56BoRuZjSbo1/Pik1mDINnPoVPIiH1dpJ1Rr4sRMXUZ3hWvxvXd1NBfavAoKjv2S
ArFWn4fJGHsMO8hxYNWgjBmgna9Mt+REUOelEZDF/VjFD7QBwmwLWXKMeRtLGdL8
phioLFCzPHyTJKeyzB/wSA2fOwxTMS6PlARXa8o842GiNs4Q/ep6baEJd/O1vWfC
ZZHj5YyI41aul+YRQR8t5UdqWmivygoPO0Cz/9Y6ZCLGeWlUF4GWkbmRy3KjedZl
IKjPRj4hhCEG+rO4QmCssZVAUcqsHHw82Qg1d5tqP0gd9czpBm0YqlrtCFR+bX9G
FogS4a52eLpud4K3BX07GB5KYDysmhUyrMLOa+9BhB4nExsYEZYxuzIqTo0yKPaL
m/835lkPxE+Vadankz6CCqsWjI40BIR1ISkelQs2l28Q2nMxrC1q9CcyTFo1Gvxq
qZ0Tolnvh0lc3Nrlmw3MUHeFiOdkBUygRjYF4F7YW09/mNcYl92WZ+OD3+LxVqUb
m0Gq8OwbDc3Ql+oYNyZBDx/ZKFkL/My0jaln/sWlWdq3BfmXx+205eBMNpg7fABi
FtWKRLMSheNPzpBOWbxLTsTAM8kAxFFKCq/7VfTyLSQR0xB7L+LC1TQFfbeM+Y6e
/3matiVo5Ccw61snRP/Q9cUg6a7jXcV8JbWbocNsw9OkTJ3lhQdRCjPqYN/UBky8
lDwgJD+JOt60egQmaQLVK7p8tPPLbhn9pM/kXvvUWurQuqAOB8dTtx0kS6Lm/a/G
AXaroanEYfTExce7CoWXTiN5AyyHX/XK5CdM0ob14TIKznUDgA9pT24/LA3PlI7K
mHTWVlcG+VKdBu8giwPSLuTgWIuUuoIPdJ1nEMcOc9mZYf3n9AhuroBATtCZaeQb
o1vKxzRnC0jRsrCAeNZ/pKfMrnn1goc7OxGl3ktkFKMAg8mrFUVOVl3GjS+l50+g
YXhDFA9jJVcYVwkOApsquu0v8lLC6iIjeuyNPq898V0Zvz4NC/LvSpwa5JbxYOAg
K4SC6EfLNTC3Z2n+8SQNwEX6XB1Y/ieBwKEyAUK2x8aiXctvECgQnTNevgz5M4oU
QA+WgxCZHRx3pqzzUj4E0PHdk4+ZW9kcrdyY4Ka7LIFRP92JcppfLw28PUbLaPqr
xeC0lONDHJ/ndl+oyswyYxRx6aIBNDSvweKki5edAEgRZCuTSEnYL7R777ikzMC1
lEN8lN23I/BCysxE74ODglTI6NRCbHfyMLe5dnLwSEo++jOjva2/liF9uHwDFvlH
uvKGquDa0PC1UO6yGosydYr4MDQtZ3w3M4MC5tcqN1xkVG3gXx689o8XfJZ2WVkk
I0t9ZPVQwf6+kkjo/RbRaJzqQ9m4+qwygXWRrxESfA6BjxOxtLw3yTb/14Kzpjd4
6XapQqlVoVA9NOW6SO7To8xOyPGur0KiUg8/vPYyufXRGkjXQ846J2yrNXgZ+paj
KglGfdXaYn62v6F0jei6EWbfsdssjLAPTR3g7z+gKIJmSNG9Nwq59shJt6fQI8bu
c9o1+jjtZ7vxQo8ijKl6lbFubNxm7cf/BT3UkY+O2Amz+P3lqsDzNBF83nWEicuS
l5kRa0FCzXNTln6LMAqKhAMMseRapAp9qcF6JlB9dAJTDr22PPBh8W1YQpU60V1C
FuiY6BLHDM6rjM01u3h+2b6I+JYEMtkGn9oEXJ6nwFDYEDP+4wLcefFvXJ5B7aqP
ShEstG9r1vGqnpC/piPtqbHlS4IHTCrwdbLXKeHm0cHIpBjwMkJPQfRngscythWj
XbeFhQxu9w2uuhHZgrTq1e6PCSaV68aynNnIQSyjxrdmQ4t9Aezr3vKXHjWBqS5L
gM3BIgkSCTI1MqKYQl/ixcmxpFqwTqqUnrC4kpdUmwO3R+q2969cqaizHJ0c1U+S
EDMS0Lho5uT3EvUPCQhSpJKjegen9f3YMjyKKs+lGzPiLBEjcz6dd5UdOeANNBzF
9ttqxXUSDXaPkF4k+e+rI9JQzfVt92x/cFb58HKq5uhkLjz4RvcZ++SR44W8Dkxb
2ImCLEXxuFawMEL+xZbQaLhA2nUGSw3TJZpADLCHmHFTJT6SBQ9Mbr8neKmvi4JZ
ajTUGwUyAyui/OYj9Q8ko9pNLMTRvy2L0vrC7NKsZ+kq2/AKkO+39hZmIFuLqNPM
4c7HFZoEPQ8ZDYpcgwbv2+aV4gSTNaousGCOw6rF88yTdyBlMqt430a5O/peCmIC
ziiANCWqZ+feBw5uiQV3H5c/WLp8WMDXoDAGJrwBHcpsXDADb2swuvNtXBjXucN4
Xyb7Gz2tDVgo/wOZ0ZbxsQWw9Ly7qbmcO+bGHza1vO9Gcg5Z8RD65YUatvX4uGqQ
urd3IZ9D9Xf2+ZpZuvTMO5jy50GlQMsXTBl08IkWW5DKzXe1baFD6GQkTWsY52bm
rq7hC6fNgiGbKhCOhcxHkcqMEoDfYl6HRKy1afTZuGnwHcY3JU0YZ8UXL5t5QXYj
TaCOOsbwr6qHqpt6GXemv2MBje1XEWRl1t/jWnbwNQBq+cy7VRMQPQvbvwh7GADh
mQMJeu3UJv0GlngyODiw4OY/icr/38CyhM65qJP9K0DJKFqpJ/5hBQBxqwljtEMg
1v88hwnbZ7Fk3GWEKMOeDXEamse/oIBLLoaVVQ5hXpn8T/nfMgHCaNVwaySNXTFH
dInRHdSffwvll2toyK2c5qwXK2P8KVOdQfs/6HcDWUnOJTQqA78fXps/oWh94nVH
OIwx8TehdHrMla8LtBHYTTd79XVDHqYqnL78YExs3jJ4nsvQUlHRJK8EFuKq39aQ
M0PObHZ8ahnmLlgxK7pFyfAy6M+LclpSYrtapc8v845j2NBafv6lnQkgkKRgpjZ6
rSoHaz84KwCr5QiMa7zkcprhv80IGVLbMB44O7v0h3WvL1XLJ1Nh9SjxTbMJYL34
/bZEhlM6B6fy5NwydTrNRAGo3NbIz9KbQnKDWsS4jVS9dYCZ/ZC6JN/QvJraN8ie
Q2PKu+iOmw3wIMb65MKhJ15ZyS+f7+hyRiy3edyeRma4hAKPX8+UlCinQR+mYwwC
8fgCC56Lq3G2XbhIOsXZ3FMXfHt5kXsnuhH0RXKuDXc0Q5jb5LaGcHZuHBMg6FbJ
vZjj1w6oWfQTl24Tmdo3UtsrSNi/vGpf8sgdeCAzskHUhwrgvAVwoIuv6MWIrY35
Q3xDPSqIdXEIN4bVMhK0zEywne/cyElKB1vZViJ4UUDsDZ3/fElTcZ8IPtcdLAw2
B8xyoinv8TJj0mL5whnFWvmGBAk0F3pJTUzGrtB9JSxd6Re3FGxuUOeUEh5lhHzz
BK/Zt/JrqZy4cbICRTO8Dbnp0NzQMb6P6pCm7L3rkC7XKbkC90MzQhMVZGDZAyUE
5lReWjNZ2RjwjfjGXk/O/sQSr0a1Rs8nNeJSe0UD3LWnJsHjjaajygenKj6frhln
Q5vls5CREzrM9LzU5lcis1Jr3YIsmzeeIvnS3iqYuyaw7nacsfDuVz9FHO0Rx6fI
HoWLKpdoGxNqlTYeQUHyaHOH3fkcGUzYgsTduw8lutUOKcdq14FkkAT+ybpy1aJ2
R2qRUrW5TQexjGXQX+VMxZyAR+RWggFrXncGRJ0mH86r6ZJytnw539VGiqc5WZdR
DUDOK74PRZleO9zYKqK17qI+HS6/ER1SMzNPJcBAQXsy2aRf3b8BSRz6yvmsBb7W
yB/nPIZx39aMma99Ejlk7/sbIWxbxVjX2rqAE/qwmvlE7N8g9vTiZLn7p93FvU1e
+LNJjQdtfQy0E9D7/Uf9IocTCVJhwr5X+cmNT5wog/cBWRXbuAKfZxA1/x9ghseK
YV2eZOiKaIOIsV3ewPvks5OQonIEY5jC5ZJ7UUgdd8umCfvph7wiG5Tu+T//a0V2
yUu1KMF/fywIeFTfWg0QUa6KvWXK8y8iN/ht1Qsr6MK1Mh1Cn93I3wvOAQDvJ2RZ
QoEoPym25QsvOMZ0PuT3x3rSU6GqRfXEF7EyoVpok4nZVw28yHmS/ZOmKY+00bxk
80nH1emPV5/LsQSrrY3zE6bY7z1DRRCmQJkTok1M1oY1DaXPxmdoSQzEIt39lyAU
PWPUhF1LUHlkpsDiUvJcETedwYVHPU9dVYAK2leCcnQDTOHk1fxEZFFVWcX7ympK
RYkbcYMtdkQiSOXFVe5oNlLJXgmcjMg82Rt3kvf28KX3HafHHY0T9mVnrA2eu3CC
Z60A8V4sXuLLEe/Tf2MyPnYnAQfL8fP/7SShGo7WCNuXV1cK0SncOguNpOXqxftf
VqdSoWZvFVauzhRTozAQG3/A8BcDMQAXP00TlDcoNv2aPACRIXrNJO43YV6pt+pS
yy4pfeT6HtS5OVEJ1XMmBpiNmD/T7I8E97EvShD6YIwI1/X6mLC74bsbouinq2qA
x/6saJ2ndNbBYcn3YbgAxK/IK8//BKPE/e+5YO7Cj/V7EyMSxT7d9Pt3fnBkWOW0
4ZQh5pNshk+B51901KGyEd/GdPxWMeps8B6gNF0+CP9WmPCuJiAnpjwDosxxmc16
TSgP+t6h2I6PcABOSHxlzIqJqykeijmW9KuUW5IkgT3YJaoN43y0UNJ+2f+CB7vo
u+nnn2hu0TlotQyPPpxmqxlYKd8TFOhS6/NiA5rQ4zxWJdLuuh/uRdwUtaUxv7pB
ojxaGaazqI4BEH7wusTb24APUm/e8IvAz1zfWnHbue3sPfy+yWqRkQSLWjBMlJhA
0Gx4s2L01kxSVqEti1FSHHSIy9j0wt/9ZEjewlLcyP6eH+Iht0sjS+wuBCdF6oCi
ZSM6BKKO99t0K8rZg+kCO2qDQiWsF6G+VBYfcOTvU7cOQtuBWQDLah90yuLvTMFU
ogM4GDjj6aXwk35MY9OwQbcyZpGEGeWVS3uGQsSMObVxralmF4JJ0iZNdlpNqs/F
kuMkCCfaSVVqgXbGL9WdJMKE3cTXEdh8UC4cKDinkcG1gdTeUF5PIGfQJWF3BG7Q
f2m7n3uI9tw/KK4wnPjquTHJ11nFDf+E2nnnFga0dVlWzx1UBXyx+iBlP+wYiv9T
IV19bWiIu5Gm6s0ab99t1BBsAuVy34ZxZv0k9flvhGOQqkQSLIioUlzc3uPqM5UJ
29xUqNz3MWCNCEIHvYDlEkkb6n8dYRP6WDYH9thrjxA1ZJ23o9uK7zuE9TSqhYYF
G/hVhxGxAkH7idZERvmf9FTpK7JWX3LwFAVcJ3xl+bSajcglGLyYRAni4Wvvyef/
Gceyn9EJ+BC7fR+cHTeLEyiCHke4Iwvk9/EA+My+ELOyILdP4sazVTH56c6d72m6
NQyMwE3g3igRRenOu913N3zKLBJgHpERXn8mqpuc7qf8+QemW1H5FFThvuisu84h
AgJE+i0XMV21A7VhQ7oOTb4RWNFmyqBXEgD8N4yfJcaPrmFmK1pNhihh4ggQd5JN
VHtkbt7/iPOR5NGsPzc37vhy+lNfqmYGfsG5q/gMPVJDsfXPyTcdnK/mrxh//nP9
/dLuWuigmNIOkO3D/Y27kllHBqx+qBq4d6HV8G3qr1jsvGJBisE01wVJlG4Wtz1S
uTdQkwdYeQkXUUvdPhn0nYlqyOkfokPkbgW0Xdud7y4d8waM0tii5JwmrUzB0BqR
knje8qdZ+fTV4yQAijJExmmbuo074rqu3NN4dQU2HTBNiD4mN5E4EL7Xbt7YxkVJ
j2GrzCBw6iV2IY6DfJtYJYgDZtSzqgW2WT6si0q00W6U3tJs3lerPJ8bAEeTNecF
AqUcoR46/os8x/4Tzn3OuH63Z69RntTT9iBiy7FbHHAaMa0FAX5ULwsLhIHTM0Jk
xhjwzFkWpPEpN9LEUgCNwMCh99cpAIRTtVLp+vGmvvuBAHIGi0n36Bz083VGMPfL
sBxw7RCohVsJcsiNIWe8bMgYzjx6UYX8LXHHwrY3c/vkd4e0cX0tmzua/ryvsxHf
Pt6+VgrOx83a0kyQSdDaYCVX8tyUVdUVRClpBh80Eqit2Mc5h9qNNENXvrwKv2Q5
xc05iS1X0XbIVTI2ugCAPIJZCa+NZDdPUabAf2x47Sqd5JVpSA1Z8QYEFbYeYZpm
MLr+5syq1fQfzdxyNya0LMkFV3KvfBFvQubBnzPSp7BvootA56RilkmQ/XX6HupD
y1BY+TOzS27aDrLwOsaePE0eTdlozJPP38jxXMh/8vew6TfI+rCyNOmRzGYrI+oS
Gu0tAVFWF0fh4yaNIXmjyhGgi3E17s6MRgGwTCpo3tdTwT8yhMWyFIK/w6U56CPT
M9JxbWcaUbW+2mkqmoYbBbwuGxQ4el3oeTOZdWuL5vqKihXMC0etw5qdjx1xEwaC
JtKhmNkJ60dP5dVTFb+bjnEcmFNaY39RDDee+QuIRPqqmUrMUVHRvMUyrJVLoQyL
PaB0payxM5SmRL22iT7KMuPps2atjRbXbsQ254TnnJsEZFWI70YkmQD9RzD8JtJ1
+gXC4Goi6bd13MCYuBMONajKscXcKAvG7HfrK7HHpyZSQagHD0qqIJqjd8SY51by
5yrxmbt+l7YPSfTVWLo9AtaeVY2bJ/dTg9+9PlSK6PiUv+4d83YJ2BQx6zJuEuYR
t0pDebGXW3AribOMC/D9z/ECsKdIa6WBcMbQ4nSMd+FU4s/gM28A4i5Lt1mjChMR
Dn4yl5dVz+bpv5YzXE8DP82cstBYsDz+OjbO2yQQ7nZrRDwbsp81UWn7kuKcRGHg
8+mw2Nt4SF/IdaMmht5OoezNss6ZgxsCjdXEYyXxrho4624sUezUHedTfQdAgX+P
s6Bp+X0KyxmL2s1Z2koriB/7DvTxzQxo3uA7+05AEv9k1VJnQN5yTVFo05eGMQy7
NfOn6HERF4JO4SZnJb3cxeN3XP+A8zttuwPfiymRdGztFIEJ5J2+jJ3m35NUuHB6
YkSDjlrCVry5Qppy/vy2f/mt4htljVvbtK9aL5B/z0ekiuBtSW//ZEemFveOyFBt
ZVuBb3y0tR+8NrWKgKmS92uvQhd01BbIg/c4gE3FcRnK9M2sFIastigidosabkU/
9iSbtyZ1eArt2jKAearPY0VOcsyru7hroSiAFoUpClMpn92T0ZPsNe6QI0nhgUFL
IYJPGY5ECAn2vgjDsUi6fqDVUpW5YZB3M4s+Jjiuxa2ECGzmXuRX3dcksMUnFU37
oRrZGJL7h4qUO9CoxUnv9Z8xFJ48VNSmFTKVZ3bPoKpG5QhyA2k+BtZNeYOXokUk
5d1nnUA7VciuLPPqzxgBgggXsA6G8ouoAlz/jVoqz1jnGX23ZSCdxfXwWlsECrfE
Mn+VIpLdAVQ+7xQFyAQdhFdyi6v4el60ocVezb2igTFD5BGWQQ7hhRszDvobixzG
GCq43F37fItG7wF9gLaNQoUKIdpT6yVFYeHk5HTPmb7MKYSNhwfOUtnuThHfkNPw
IBecv4dd8JB/MKJ0sJVRbjz2f0/ZgBOP041n1+TYPrJHeFhd5bYd9HpiM2HmSG68
LGb0Wq/EdqKK5Vg+sr1bo3XtqtQGmhTsA6AGjVEhI0rBwCDEOVBMWQDEG5wPlqQK
G7d6Ndqhc+z5tMB4ccRrkKbrkY/m78D5KZHbMnQenYq0HaXCmb/lxx5UM6Avs0zj
wQCJgXui1DYpQMVKVYI1B4jMDjck6c1BdR3aYiVomUgRoylQCw8TAxW652WBVQpj
Mb12h9C7y07FX39djQVdk0WhoE8HJ8fTKLr8eeGAdsrUjROt22SkP6RSBbOmloGx
iI1rJ08vunOlTpQNdonk+GfAX2ST+kdXSDlvwWv0eLlcSvVZAmGcGETEgN2Y5rG5
dkfFrbpRxr1qEiIY0IAoSp2Nqr5Px8Fd5k2WbJrH6vXB9TbKyya2At0pZtuER/GV
9cX4mfev9D+VI3wP0DEeTJrDQA0xYGKwzzeA3VRa7OBdJiOldX12HX9KXqL6ahql
IoRxbL6VLzzPRLh6UC56PWLFFo/o75qIXSp9257Anmg9+IVD9U0NZAnqWJYKHF68
cesINqrNOQwbRCQr8Bnnnlcx2dJK5+Sztu+DaobV3v+aQ7n47fIM/JKNndOKqOml
nuAAWe+bgY5kA7unmwDbcNfVnRmY8eTQg/BR3jln8C1+xL9fsN11x0x77/D9ZH+F
yyFXmTzJS9ws+UhszvN0PPRnyfTAwY/RvqqHq5el46COYfqb3ZH5bRsyQbzr0NFM
OI0h9ETBWfCLzMSYnXhCdi3AOWmeZkCzYEkxQ0BPcXRom5B6cywUQhy5mQerykYA
b7/wCOey7GuLnZhAhPnGQVTRI5T8+wYlgu9IUyA/0oHqUk7mpUMZW13kwWip9G82
bfa/TYMKh50lXkMF8AM+zgNY4c1L19jadowiUPZhL0FMjRC+dM1xPfizRux9Ch0v
UO4egckLcv1DOF9L/WGNttxjp22BYM+NaKH53neXlcZKVycCSf4gICxkVK/c+R0j
lw5s7VffHhloWz0H5yJI9BODoqk9OOQikAU5T9BsAFbHeCTkxU8YWnBc/AV/SbPW
By42JcdVtCrAI0qZT/mes07jvPLXepE4m9aX6fLF4cc/KX5slaeGDs6lJcdtV/Ju
M6pgrbqrkBEKDojNmpKkNUn2LSEQurdmZx4fVg8euRDswG1/HAF5rDiO3Duar3Oa
SAG3LDSGj/a+AYy2QetHR6GoK5ehKvWBMsPY/j8IV9twTisUunwzVgVYCZPXMGlL
4a0oXC0fbN7Wb/ms4LOl6HzGTH1VlDu2pk4M1J1NLHYvJQtQ+XuvAiHaMmFFG3nb
Gf5nNAchdUfHUWjSK67PMwe3sowj0v7VpbuAf4J8ZxUH+D1mMj39eipn5fea0sip
GEK7ZTKROkmdymDlEdCkj3IDJxC6TFm0Z1cVqbqndokT1M2SeAHpk9t4QCpKUzis
FZt/J29CA9VskIPf4LpySvGIRFaQ+wFUN/8KtbcHeLb2KooOK85lp/19Ixh+e3nA
Yd2gpzr/yrTOPwKJq6z6eBUL5wO58vnDMzGWSLXvF7PzihsJG53k5G+L+YQogyqx
I1FANqKJyiXAb8ReySMSXBi1WxRekgDOgttz0S2oIt3cYwmsBDBzJFF9wgeOC6Wo
vpqDILNs7gqUSIf9KMXll8FaKIpBHZOAfC4XeJaVLxlVu6Du+6F5dfio1rxb0n5j
lXRMp4vgQii1w1OR3C/XU8GCU+TsuigOWlFJDj0+uIpRj0BZxNB+4aQbUdixzGkR
e0gV/S/gPiTz748VDLEHSMK4iIkitWHxDxtxzIq6KlaSkWMPRqwgB6RfpuSBTiE1
cKu/4Mr6V7NlB+5SsDdSCXvw2/QMOEvk4/Zlv3TO363rNRAERbzwyE3v27CjmkJi
T6kUmpZDSpcS5/xvxsaiRlLvrTovI3x49EY5x7n6/K0Mz/SKsyPRTOJR4hNU7e/f
Qkb0FK2qaT5jYllRE9060dkgiPx0nMwbwVZNfjwcCUKlJqGyX/HkQN8y1k+D+xjc
dZK9F3sqicnzBhAZgpb0WDYwkJNFpGtxkMTmA8tjW4BSII/h91QXQ1rdb/pD/bXs
7k+RKAiU5eYSXQQpYQJzB98R7tI5oAgZTphkfY4TzRybyGb8nqDv6vkpIvv/eYff
h4A/f75S94M0RkcHfIK53Sip52tSgemdUkrKyWGtybCtVXrDtNJg4xTpx7Sns6gS
78HaBM3RMVPJs9VAup+FSKb296lVSvATueFtxh8sGFj7gce2/v003SvQ1ELe6Wj4
rp4FP8cSNHjp/65wvt04/rMH8vHslYfC+iXI/mpwJRDbbJWmDWhBspMvQut045oJ
Vw5bvFk8O3C7uM9eyLDkKafgObqIEuyeLeXCFt6jZdV9ZsJJ6WuSmp/nm+oquUgG
e35i8n9D6BzvgRxIGNm+V/Lf3Sk1vOeovwpEhE/tJRAs1Q/TvtyeBZd8jcRci7y/
o4AiCJbuESK/2Rn7kecWvOZqpz6rDASAmQHDV0klbDNWCGka2HvN87W3SvCUIEah
4wvpbRrAn14Hf/dfucDX92tnZ7PLalUX/MC1FlYVhhwzWPegF9WYERE8gha7JyeK
4zx4Ei0TyPydXKugsciEdfwCSnkU98GeJMC6esSFykIEmrl0XCSpaeXMvMOwFOY0
SYXx0ybSdvV3TF4EI8xt7ODveR0VAMpBOTt+wATya1aiYU1vsQZRlROz/SKGmkrV
yFnFp4aGBT6BKwzzz8Rh9f6UQ/w5jweD86uIDthKRuzR8CnxbI8zJ9ZCZaknDzG5
qqaY6l12yb1e0mJztbJwAJxmNW+qgzW+WLR9S4w688TgR4qxztIspR0W5OHG9ewt
b3CE4GlpRt+liW+G0ecskHjfaA5R7jBo0GVSxHUM2Ft1pKFdDtbkNj0Hg2sv51a6
+Dj85yM8nvkyCQKSheTpmLo0l57eto35eBslGrK3Fd5VkBR3xGuLKSRE2nBFaNK+
1l+e1XTJpH/Wzp+dJask+43VrNJERRnK3HulOMu7o9tnRT0vOuSzwBjVBVAwBswz
X6FEWQ6YQ+2UqMSmx6kNwCjKdQCWm5O7cRoD4zPDEontbIWmSPGteSh0emT0qEOx
IMqLuj6uwG8XgvCzXNDvsT8cMZnneSlqkc2pAFPSX7zluANeKok6qd41Kc8QPgfI
d+O+VkHCw6gvw7rzDJmZVae97lYgAzcHC3uTLSxxhpLJcrKPNvDCt6uVlie820Xd
rNnPUo89tYbflvFYswZZf4CxJ+lQNE3qi204MJfjaKZp1g0Vgumcbn2PTyjBpjY9
uile/XGfkdgy048nIxYiBH4xYKgU4+FjPIG3AJm2Oy6xQRDp9chtBsFCmfO4kqFm
sRnTQ7eCqU+eRQvMgDSS7WMMdHJlro43kubxRHTvZB7ZdGReMp0iJ1pqvhj7RQp7
1gKVsdkBiiY4tW+j6+xJ2B73pk1F7HrA2FxoKq5x94rqOjUoPsTlIKebLeXmf3n2
V0/0C2F/v2CixAMjsx5Q90sFMcpATSboBWPdLUnLH6qDZfJWM+yjYF74MXf7Aamp
A4RBraXEW3RMzQCklds9Lx+WVDwFojWw1QaL6c158qmcD38/K0mkn6lnYdeqksnM
O4UZ/9E9G28/yfUU/YCs+I1nlpfEjZJ8oN5UW2/QfLm0kVhkojZxbbeqQf/XEHPv
dsdGm63AkDY6vIpE03sN5VlO7OpKTgPUCxqAhW6xolfDwuKXB+G2XmPe+QaCt8GY
0tR0s2U797asltC1Ua0eEgISXoTO3um8kZHbNbebNB8H9gDtsl8DO+RVhg0qtmRH
OElVw+BJ6hahfdyHvRgSqMCrqfM2UNCUnDhvDSsE1CdJhL+90Io98GHEKz5V3+BT
Md95YKt0SMKqZwfM7alTtWfc5wWxHtyoKpyJ6hGx33hjzUGp5GH8m+EHX8CWIL33
mjoeq2tyPg4Srbjd8a3FpnhFXyxf40CTutTCz0Mhhd6IbjlvBogWLQ0n4wt6/54D
6MC8zu7hVDqbJvqhaRBG6yjcHRjnCYQghG06LWWt/j+3NF4PHPHBk/GKsRgL8VeT
HPf5VeyPu6bW2vKggnvVvzQjv3thlCHO7w9BN9QF2piSr3yxOqDKbcf4nECcT9yZ
qjUqcPm1hvRgzQuVvJxIllqw0ZNldH/FMkk73N4TfUUkiq8mNVliGNhYQnjaH9a+
g4sLqtw9NX6vFJHhcyxj0qnd1kdjZOV7nYB4unwLu4dUicOKqRAdxc408nkwhMYb
UmB7LK0jlXKa53muOUgZdVCJQEuH9rolH869mBcctIalPA47zVAwx7jTNS2/Ksgo
5YnbTYShT74gkMG0G+gaM/+RW4ZKcC+Ys7ipk/Omf+6rYnYCKCPuRbxIWjZwW4cs
L7zKbglMKSJGt9fbj1VQmJQISN4n+kqYN2QhtzzvqwWnxI1T+zmUaptSOwoBnsFq
/p8DDGMcxa9JTkpYrApeV/Ex8LdEqge1ZfBcpH2Z6o4piyCHNQSu0dSFv6xhGQpn
a8C8hiEybda7vh8v3P80mQCguLkixLpJ1Hp0605JufjYF1mx8+EoA8SlcKuHHEFM
2bhIUe1MKv6Pg3aUJYv/Ju0YgJgbaQKbzA7xUZhlfuble/GRdAak7pwuwhT+mwxC
7tZnVH0rENt9M4hRUHPZY6Dn+jE3ksxk4opREubhlAFP2/N2iPudPklclX3CihN2
4hNOgXbp+5RqQGLq7vrOlhf2rz9ruZQ8HL3x2Dub6Jp6pEechPppkgWm8agBpVDA
NchgQt72ETXmr9Ow9aC90JqUIiekOrIFDwsn6zyA7gjjHfw4rw6pcYO19EoAXTs0
dW2XN3sQiQCs/HXZd/zzuU7f1kbKXgSyNGemd9L8vqko90IuxkJDlfHPDlP/+wY+
YX5vGJt+hN+WgyKrtwXOt/+VSaPBTkFh12bfvKouDzvuws/kFrkDY+aLOEDowfta
B9OAvURH3/r58If3wJit4Wekta3dJql6o4s/4LzCmT4b2w9ek0nkJor1PvxqhhEd
QTB1a+j4Y+r2yJD3i4TcD+MI7bWQzHa+xQ4ejbAg2kLEipUL5fO5GD9fv7xXqreg
dIYAVkrKkNVQ3KawDwVZ2WAmIV3RQVcThj3ij5TLHd4LNarxSN+6U+VVW3pZOs3W
ebXp6beCX4tla7L122Er72vYsNWMsJ4J3ON/wPzPYmrwhrgD/gmyEsdEQFZxPO94
aefEb3zQFH9iAddbcqUwQGQMV0j3WPG7gwd96/IfV7dUEmTYTM8sG4N49+3Fiv1A
NZn0CVwhnJkT1OJSAbqS9fvqHCVGhr6awhXWsNqKrBhntNxkGYQ0scpumP4n4r1x
qCwGJbAIYI7xyxvQ2S2WpBXhHCI6ZHtAHM1HaF3eWIq6U/T9EzdbmsEAfrTZzlzm
MfQ/m8YSL758JIcgJYAqcxcynGYlnY6pIg2NMWOoi11QbG/JD+P/iuurI9nPFW6A
7F49wdVnP2aS4eJbTjVazG68AqeZ1sME/x2AV4w6Dg4vm15nfL5VprBR2SW7g+xp
GcUn/Jv1hR54vpnRBu7/wyN9rvOveQedsjasMYaOZRG1ZTUKEy9IBOgjHYVIW0+C
jSTKpNLZL4JI8458PzOxeh+VGlVLvtFriQWxcQmsR1KOrZxxyHcH7h/3O2vSHU4+
uDahm9A5eCzpn3DEGzOYYzBGDh272WarZnWC94vK4aVqiscuwxA4ANxm1QG5p8wh
z17E57S7wEYvC3WzDjneyBXigDKWqH54nyzQs3HECdboNVIZOSPpSkC89g4offxy
qffH9Y8iZ2ndZWtu+qxtMUp+WBqvqVtBfugjVbfWD2YO5HBrS4oPSzuWtmUm7VwW
YtxDpCKOOLwtk7GmZ7GqGNJQs0UzXgOAhAp+CFXxH4OBhjKJvgBDJ9bolAnMKmDj
/NFnthM8xiJ78z6Gh3rsEFR7/ZqmoLhwLRNyGM6wteOH6lLvVV45fmCBnBPMT1Ic
Y6yTTNa5gDT2QP+mhw1e71A+Te1C04P2gMhX5Cq/zLV3lLzUis8oYEd4LkId5DXf
EsvirW5L7zbatJwI/YNxZJjU1lSzp3kfa+kgQrLDXSfwvMVZdWbrjkOHqDP3or+b
chL1K2NMK9B3WGcIMjPlDV5OxEN+tn3e+AVfDy5gnKzwMlo7UVVpcYbGt+j9Hupe
wS/8ifwa1AVGHyrLBj+ce+9vCFtOyiLDK/kaz7e6qTF0nSEQgVULl6JONAhM4BjR
+HuW1/ju8vfYNzD2wyAbX/KdZyg/GNlkWj5yT3nXd5bkrTvcdjpMpj54mW6Mc2rw
acKlMk/heo4ZD40Bs40pn5AwBZZop72n1bp4k49iPwVvntKvGzZWMSzM6fGbp031
BHSy+eLCynhlS/HWdIhig9x8DN0pHVqX7mTQksiR8iF+1/8mp9QPkJd8f2RMOGRv
SJ83ACIvS+g9aqVSlsp1dw0auj91XmIac/SRjK98CIozgD64XiaBVfu4C07u+UVA
uI4jLbsAI+XhxYNx/q0QOB+MPu6hCxfR2JqdQ22LDK+TUIXSnFIlr15YSkc8i7GF
AxPTy7MdV8AUEkcn/W4LsHSYKSoCa4/0e3zdCGHO6i9hAJwkE0xISykMJIqkTuLM
AoAo69rNxgbmMqbhT3eLLDK4+Rn6fHbCt4cOKh/hErYIB2mrf8DGy63YJ95QRMKC
0DAJywyWGH1Wbss1TPGCqw8XpUzbtQ4qboKZ0+s2MJOSaISvMfhQ6ZWXleet8cRq
8yxcD5TZtqGbDExw3wTXOqeBAjGDdQrqzwoHJfXOL49xibtzgx923p2GrbuX8aex
2pBDhDKcBWCXecWO80xLeirc5xEwzvPgOL82CHboXo+utpT/ZezL6S+FoPwd8iKN
ToTBYuSAXkCMg4Mtj1Jt7v3M4V3uSbnO01ejIzLh/j8Tk9by/c3IOVA59pWo4hfx
nFEc1rCgQ5iZkLOBWcVJ7zzmJPe/eQDZeQX5sFtT32b8xlVtLMkBdGNV3qzuwdLG
uRfeMxbgonzSND85mI+SzXyWak0CUQb7GeW9GLFGKZnf6bt4A0lhL8FJQDUT63Gr
V8J6aZ2gCZ+Pd01rw3g1pxJWvJOnCkIFEBm4/SyMK7dvq6OfRxtQbxMY9vR4PMTF
/oMAWpXFP2WvAq+vauCNVT7h/+czLx7l1aAsPUXONKBA7NnkhxHck6HDB29mmaru
YvUYez2Z9yI9QXRmxKF152+K6xwSbildy6gdMcR/sLpZe12MLuRosdZs+LD+jAN6
XM7rysQbcmYAzaFesVVkO3l6FE524uDvLjZ9fur1v13b9xgnARkzY8FiHIBEBPCW
sZygJcmI5YveH4/ernoeseIctrBuhu3WAGSpxNaEtvZvsEgM94FffExi2t2CmysF
WfknfRmTxY1DdT3OhcDdgQFxM1o46bykaUT/K9c8qDYh1Pyw4hLptr7JbYYPHirG
mD5XfqyJbqTGbw+/jy0RJIzqQe+2Y4H/oiLfxJlFahLO9kYQGPzMLygRA/ii+mW6
7zHl7mksscB2oJygSZiBV2IztQjgOi5h9incLXCzGHifb5noNGfTMlC8G3y3Xtmq
Dsce9/MoxIrmvcilXfEqCl0CTexU05dIB+dMN3cfyCPUbAshncxF2NMdnV2TGZe8
hPKJqInWSbSWkvUHeZRfLxa2SxTCOS9hMg4/rFQYXOceSCSJXBvTcjT0lAIGX6Y0
w3vt9U1dbPDNQ4cfyK3mJc+fng3WysBXPnnMHgjouSkXbP39yytS1Bbf8f/4xN/W
AUvrXcN0HH4qtQ3fuH/mocBZ8HSjTW/J4XROOFwQTsbYCLWl/xRENbykhhinJiXh
uIQnqb97P8KWbbH+p4ysERoIVIX2aCdM/z1H3bfA8f87QQ4Cf/J96Zz9glNLbd2A
itN3vXPtcoAZ05VamIb/MgUKvOYiZOuac1yo5CRcw6jOHDj/19/L7c7/w6efsadH
pvA0VmhkKjd23kXYunevgC0ccbXAS+gyx9HXot+YtKanXDajytEOpkfHmH/vgcso
jfBm4dPqx6JSaMXl0hnV7B0pVi+87Tjnz7zVnDp6xzHJvkKYa+xAwAndsCeHfkYI
yt6sgA/R7gbglNrrIQlgTMOG0iOsntA0PLl8X1quNGn9j/tTeqwlbqY1miY2a35o
IzPjRmfYWIsb/hrq+tbvK7Y36cRDcgy7Y7xMPUdwpxkBN/cvcW4ST7dMHirOhcf1
vUpq2991j8KNyLFY5NrXpGqEtRGRCpUV5qCGweFhO/PBZjFe7rCiyHe10ETunsZf
b35M3qyw3AmWK6rwBXRwWQIGfP3BpAzBtRkjmfuRABG3HRtAAe0Y76bxjkrWNuNm
sIdYVtaLSKfF49z1ttGZ2w+8HmCN+eWGZt8hEwkHMx6nY8rizbbJ2ueSAGsUU1D4
N3s7skpc83PophBpGl6EKebBymLwuPINE+OjHo0MU+C+oz49igtBjm31w88KVE0R
yTtkQ08voq8TubaeuXx+YYOX1voV+o19N4aIH4za18YnHh5NhjRXxJQ+nVHZBo1g
2apAh/fbZXAgymx5XKq/6uqdmhq64Xxt/xOMA/I0vxaK25K2ImGp+jSW+pNGpC6r
FOzPxC2OF4Ps9xxZwamJdi1kD1/S7HW77xMbI4pQmFvGIgqn8ZDayiUyHNa5qduG
1HfNKCprt7K8teidC2W7jL51EsegMxxQ45cv+Oe0P00SYQ3hdiUvYMbPXE0JRJBQ
iIIsBxR8KYaHZr/uRAwQz38kuSZVPc4QCtV6SknwzvnjLLJClk9MEy4qbgvNqLSe
0SWlZ2C1gbBsnjhQZWBmP3i4hvA8rxN3YgadeVgXbeTAx8Z2qpxb8lM1wuci9050
sKcaQHcXzo29mttyJrzAWAwY0u48ej38CxLb2wnfvLasT91bN5wyT9B4ujLYonwD
9sNzThFnntzD+CB38JK2phQrE3VWik9RQ0ARs7ygMtfqHu2PuEyiExCXSh4Badaa
LHvgM7TPpZiWElpA/i/eATGSGcfgM8ptF0QGpMMB0lR88wwzPULNv3nbY+PWz6/p
bEXHgzDtuRNXZ4yl6SfqFzvGn+0sviGgKyx8/hNyrhbd9TBid2jRc1kupSlzL3dD
QssfepV+W5JNsyMwAAMoZrRqu1hmAy0IyttSAmU1m4rA2664BmWtS9wNguhdSbJz
iAmFo6vMEix5RiBlRn3XKnsm2VL6NkrQR/w0SK8RysdElSxscFan+M67woRcMvYV
YodV2NHcL9er4nFugp0I9JJKMSz53jJGY9VeOZfDUg2c/YVyBzLBjJfS/GkQBWEq
KhbFyxLS4mFzP7B6C9lN19rTOz8j9CU+TNPwA+5MxDyInDxDX1Rx6FO5l1QACYK3
0Zs0nFzklqcdQWlUzqzkGoTojqlqxSi/23s2S7Sn14ArVsGvDO5MJBt8fhNCTFqS
ZKsO61D5zxN28oEbAPvgqTLKzBqUq9ToAi0V3sbBwrTN3qktoJkkYjnNLe6/UZGC
DiiDVoX35IcWNYHf5r9j9fNUELpIhOUtU2+zCBfWmzvzl2x46AfNsNMa6yCMMZGG
C/fTwJsgsfZic9tE9zmiyIz+bPZ1DsXhv/2ulvDVpClPRIiYrIpcdbUnJTLh9eoT
QC+kk92VASbhs3gRA2BSuI6KZFUHrubF7IUSLFd9tU7qdijqRLwpw6VPvDqNHeia
SjAsiymOLOH0IoTR/12/B2WJYCocSrIY6nsGDQtB5a3+j8D9LRIsC6qg1FDD2v1x
jbkbluwuRXnApIuiu1zpKLT6w+2EajZN47ebwVd7oYl1fmXoHJ78lhgkqjMuJqIT
7GwOD/P3Ar57mD05CgOi5Yfsr7NddWPPPcX9uLLRWEqgV4fjKKfwLUTRKXko9OEW
isv17iOFN285EH21YGjodPvTISKJMYBYRP9VeSkGT7KrFEntiyyHAzX4hyXQcpxQ
4iNgVWqAKXlQPa+3Hzh/BkRB3bj0XegeijGWdAaPxCbKFvEgsjmPq/e6mV1xGuTL
ICxqmonM0Z/+iD7dNzgP68dyDS6LUjuc29nxMrRrRYMfsddks5ShKCxxJ6U44QpX
76VCOvCNgpMtzQ2HxnyCgSPKO0MDPl2nS309cR+5YxmO3ulX47ry+64hn0Q/nqez
uUvnUlNFyMvsWswibqu3+9tD5QCMYicEUWcNxF3HUmCwez9ddyBNF0KBKkHewFNb
N7tO++cOxBYAcNUemsMcfYOK2BCF+JW0AeTLIXyJxNtw/icZ9IhhJbFT6g3fNpag
wafhwEOM95hgt5khbg27XFvMYeGA0SNxHRzfTD2yf7JVA2swr6yHThGnczgHp/HC
7pc+nxHhadakcTPVnqnlRnIVu6grIejAVk2hAMqyhczTEYmrvN0OBoPDITOIGclq
a3r4c6tv3783I8WFCjzs07BsNq7YUnUrKWJtu0i2oKy/UGfynFhsqZOXbAZ9v935
6ltlt4neT+zoEGbPldiE01mVKB8nVmHSPahVJTn5BYUTmYf5hlMiQHwnEroD9z+H
brVSF7ZxXxVT9dCyIfv8xHyDgbxxang2CGPxBhc+xsyFJ2L6TK0kMmvGOemqBRNN
5KXqXtFInA2e/NR2hKTh/pvpcwTQTuArnTf0uyNGFBObfeY6RNIMmQIpiLEo/yRX
p1GyS+WNQiPCmw9xwmxaCxQNIufCnx5ISPzzfz7WxPsK8Rn2thdjSWAqWI/UJ1NQ
gNOrK1hV02a/PP8gaHljK/5BgfiR+YmQEIvjaQFtJlzvYirAFq0KVXQ83avmCw1U
9f2OGQCYo2pAyXAN27MrHbojj4rMss9hT7WHURjtzIpScrmTDSsjk2R6Spc201au
zLCYsU6bBy9Z4DD78uY8sOZ4O+c8GqChQJryvHlDWWrbtst3IF06ruzvKWmtwEr8
d5e1LfDNGTxPmSuHgB+LD+jpJdb/2gVuRonDNfUE02Uvd2mngzyTZI6h1waPDWzL
ROvlKkwvBOYwJitURHxpBMmRLghK94WwgLMawherXIxFPkDJlyLyaILXqS9N8EeC
sW6scTOJzzQAutfvG9ZdjvA4yQh1Vf7no5i/+a4F0Zcy6HBupHnOEBoont6VGSUc
dPjsWSc01HXK9YT3Jl0EgdJbr/tXfj3BTLMmwGle5t3Z5iNeaH86VLgUCIzQJolG
HwAoUpUBT2NPZF+ibB1ARRFbA1m1SZc2RlmWzFaFW71rPvS1DWC7+oOOcvNt19VG
C93qbsGzMSoklgwXYHT8G28K++0ZkDvtoTlefd9iqITsGO3R2B28+NdCIdhQ638k
AjxhSCaSOJ3K7v0Je5M7ITd4FhhUmayrtNzsI/ivYVW6fHCjms+aGj5mJUgOdjO/
sFEd6liwvXNkqg0Kx0jKHS1NG1HG1MYbNkQn2Tcnf1mmAdFqFA776vBFHatoZV6O
phMnyPkYvOq9nF+2nkmkBj1TPJt6MzCyQo+OX3bKtTPpADRzJCmahu3rFn+XdwVH
fn2XRNY73OCVNJ+Q0lP0JBfFTqUDoVVVoanSQeTBEQK5yuGtt2G0oaH4Rgw9iTg2
CRic+LFZNEHoCLfQYjqb4A479TNQUWJLSiqp4kfk37c8vfOKI+04CEY6P9PoLkz9
cDs1sJHxA7TDE0xthaZizyT+sgetOA6Orjsm2OzDZIXXgDQRtq4sxA05G0IPsTWl
+KJp634f4R//9SYFi1pruZBXvI0rtqp8spIIGiegma8Z/DOhvPthMnDbAQ4roeW4
77QkfXE2h5kcFHV/OJL0q2yWuSRdog1YtzYsMdra+f862zP9M4ra98OuViO8KTVa
rrV4bbrcUlux5u7tuKy+9PCcz5OZgdhI1yG577aYeL41isZBwwhZy+/ot674T1o9
Ts3hwXSvADpi9q+LGlMzwSEcd9U+CCvIoxfbFxjMz/CtvmW8hHBFmHE2MDWbyT9e
HAr6/LAMabXrmWGUYAdu2UlXatfo1CIBl5oGf75UNESH4Vf/eZCSUxhJIMCh2tmZ
3UPTOCo4zzqnHTXvBibIkChQGHjdE/Z7/+K1V9JetShkY3vBzTUyYnipApctQYJ2
hapPNCMOwHJlttE0CPP8bfPU9Wts2pvWq3h6gv7EbeKXZu7BWtuKVooKEdXh6/kB
4Bq7AqIBEFfyBkSX87VRGXiwiiY471fNLZB20AR0u9BuNJZjlbnsdIKmHBUyANgM
DnmstpGM+X6+PwNJoKsFH0YRVRhkERnnt5pzMJkxyrLh+3m2Jcb8/9bCT71SHHJr
SET4KfkTnVB5aEMG0SAAos/Jxv7wOqRlUkUMZyd8AC5Y9npA4U9o5ykLR9jGml8P
AImYhRLBdhFvAcNLOQuBmZgg4a/l33hSr5m3yDIWKFGRArVZVjmXbxc4ITfB+EMR
sSFQ3M5teb0DOvFUTph2YuOeKZZAT63JOCsGbpGDjTU70KJTNpE6cNADW+XoQBPc
XDtmDyzgMgY9Q+sGn42ERRWpYJIxJT3L8YJctZVbKvf+w1N3jS2RiKH9Uzgg/D5M
8fem851KbwprSnUtNXvyZCoS3kTd9QsgJ57/zKBsjmGivHHkPafxMvkOuDq9oSXB
H/EbS81V73iPP4xu0aLvOn/IIWgksJ7e3858CFXMrbBiWoDmY4Jbql1jtIQ5TTTz
02ELHn/3FHSAmghet25oDxIwPEsDPDm6icOlUvRKaTKrj0x+lx1lBfz//HXiUYMS
big8mC6jfWBecjVAWkQ5lhzpBSyFIAkh4LPCs5Hgzmu5oEWEAhrGWOgWhZR5x5yw
YsZ7u3TjHTUB/09Ya7dnUMnkveT+XFsY+PBghKJlVV9nxBj92tPY7VVj2JtC8VIj
2dglI5M/+r58v+MpeXcSYQaO3xc4M/x8s4djU+pqvw1+3MxGS1CcnYMnPxvJtMAa
kyUouDTTzMBB2z/hEfKeE/ZK4ghzwpYMzttI3EE3pfGS//cybFSXKYJ6IJuXMS+q
Shg+79z1WmWYakYAU1CMH2BdMvsP4xkzNJE9eBlhRtj21vZkRYjeew0xhGefG1sP
SxUW4zqnWju3SISThEdl4/0oootINue3fMVb8IhumR4rhKSLOv1HCePsutCiglRH
Wkjp5FzHitcdV/UhPlspeD2YNlksOXl5YGwf82G4Lit8ggGzRVwUZIZFeO2+bDHE
z8BQS3nM2eKIewH/pdTl5+ouHxMEloTFaq0PwkeY/I8FeISblLTLkdsgkvBgBXjw
MKg08hbJgulJGtwZLPjehBBJULnyAlWgTCZc2AUQPIhC544wYPIBkv9VrYJmMyqd
rW9VqYEJkxfu8vIHifQ4SwFIVUMGqp9bc08QufbZUP1OoTcwbsXi9Q0rOpjkBRXN
Ce5HefWem1d4fNQ5+cFntYKRjgKA0QjXj08GP48qMN7j9nI/32RfTqZvViwLWrTs
ZUvlRTy6joGVZm/WELp1HxkQ/JExm0oC4Sc/uF1MVdb8ttQN5P9oaJBdMFtiBla5
Ltqgw4/gdHWchXv3393m9dBWuScV5UOi+hWXAUMhrZ7Q1bwr5DtIqNg4fgcR712h
2bUkuv0vdoKbi4oQZSPPb/TQGXf7ONzHHmFrVrlYVUoWLiMwsjmEfS1C6M4Fdb5Z
Y1fZMoISw4YBYlB4gHYor8qle5yjBBO8jhvn7ECRt+se2NHzuQ20p+N22hxsRpzq
1U4vGbXXpHKSN4RyUD2UinJDwiR9ofT5BwfBDuWW+72lCRPq5lk+r/VCYlpu6dnr
rcwG55JHbzjP58dJc8PRJHvFE25Fd2mP5PuBWPgudQMHq60dIS9oalXf0ZzBIhHz
FCxNYkmlZ/w9kbCFEmUvg6GCHBbYoQ3AtZVcuc6W5j/9gZD3DrGHOz9T+wHd/aTi
Xt8Z9fkeKAIQ14RygFpNRAigNtzwI+8T2c6/Fl2jl83jwVT8iIVgWyUXDsixvbh7
x3rl66Fr6zw3a5BzrexggHDsv4hkgnfTZFdnyEZxNlAQbjFB5FWGOa2qXnKXM0X7
UNgffeAQ3W8VqTPwpo1Occ1g4QNeeJ4V1hF81kZ8kV5oYoIaP7RTzxa/1BnF1o/w
IZEy1JHhhTAKWsfafmP4IiWAhWDlTAJ38w0UixkUBX4V7LBdQc134BDEmG5hq+Wm
zKKX+Zpl9FIfM3Moxlea38A81agK+ogXpwvxcpphU5SosXzlQLltlR+8CT8oYlZz
4lm3GUmgISyx2bSrTG/ALteRL3kSMoUGTR+WS1n3o0qeR+r09xZItsZqtqwFGJ2L
F1tJPnOSZ9hxsfu21V2OtZkHSvw18i7+LeKinwwp8BK4pttFLR70MUhBdFlJJevp
m6aBrfKFziIZlUSHl2RNLqoAiJ2kyLvvXp5XMY3+hD9KwpV8ecwF2Dny4tgRk2NR
AjUIVi9MXMuFTxYOZzQsYllaOHyUad/8+L/znbjtuvsV4wjdbrur2Y1dG59EOSZi
F7aFT+uvBas7WphKkb6pZuY/IB+uxu2q2J+lqc6tKnp4KVrJJMmTY8uwnDXWclI9
u3aNbDFyZcv5znnie3JOwJ9hOhbzbCL1fZTGITRwujVqq2Q+djYuGokI+WSM0KF/
Yuz0lYU6NTQ/dCJ54BBvBh7nS6eyzfy7xb85b4ggfyVtcKh8gWBO6q6rqOcCfALC
feUfaMl70Ss4FqqiL30AHNf4WG6WBqIomoz5yFOZZashBDU/uwAQW3NBK7+2fb9m
Mj5MXz8887K7N0OPPx2mohzmWGOjqStwWrWrJqF1UsJP+PinoLzsJzYYUk5ifelX
Ot9/l6daFg5kH3ELyAdtiYzr7STDGfzWqv0oFsvTp9TjY/vznD00bBTUnTUGuvXE
zKpAd98K9honpzm3YZw5PEezFDSR1FweKy3eH/cXZb/xxEXQ2RQ6lFMX/ZwvoxVL
wxuPEsq/UNzkiJwDi+Cs9mM2mF1a+iDr/726Iwgn6MRMnG+MJ7efIBxqRRfs6Een
+oUF4yE4+K65yI9KZXUm+BWQ5WXQFcNU5jJjTAu0oYyezcIbb1gpQwpy0bjeuAhW
uEESyzoDrFuYgsJhkVkyvOZUjaqLKPko1Coh+0fo1VG6DvkSzbwwk71IEjDsMDqu
/0yNeSelGj4KkbT42GSulqYx0RejfGPCN8xHLIRTu58F1ONeiawhpwcff4HcZRLd
kj990k8NzeDrl2eG1EbtkeadPB5vV2/AP0Eduo/2MXiphHRXPvSH4Nqefi48iPsH
ROdlA4LXCxUV/u1o5YqFL6aTzobkE9AkdyJk72doDnSYCImWvxTWQ2iSgk/XGn2s
yBzUaZwaPltY1lo806h2lkbI30l11zhE3VJS520c69AgESX15REP8INGY3IQsCk1
mEX9pWD4UlH/a13SVBc2tArHkaIll5IRcVvHZg75rIXpQAUOFP6VpsvakcgAso2j
y5jr1Dz6z57XBM7ECiRrJFa+isGbraAMTXMEX63rCuhHZubO1DsO8Xhu27XqXtSN
6SA3o8eglLvYAV8TYXCVjUrRtLEB1qVgOfKKOjkpVmCN9V4k9lRuBQu9h6mWaUjO
TovwyH/5FO4N8p6On89OQbR4Mz82761ZWjHkDskbz41O2VT1gP6nIvPYQDOrIVLR
a+i4H1UXdF7QJDg++CYXp4VEpremHeduUP1LN/pyVFnnQrO22aNKj2aHU66z2a/i
iFh3z2Fb1WU2RZjwBAJ3BzzqUyQGM+rlfpRUk8T4AFJGuZiERszrBe61BgMHR/o0
CPYVGs6L90uS/BhxeJ/UY7m9HKAMulW94r2AHGzGgUqJXPZJKzeOyerQMXSwVB+y
S4C0E9DS6/n+mqNMHcEcC5mmXN1nUWy1ISOGzn9YOEqqeWEPjFceE0Q51K9X6YEh
ZsLccY/tBpEcc+nc2/09GFfLdi2W0bF48kiXtDPHADs2AW4kRnALVA+T/YQMBfSh
5zqXTV9DiFFS4I78SAtG8hQcCH3pMIEVGQUmrWfFoDFUr4C0w3217XX3VKBOF0kT
e4naVMEhqvx6emt5mgGCdrNFgSW766HTAY/TXva2sKcaoLWGXUdk/8eZHeOnhaCJ
RJHghKDWMg+np7ut5DyHgMxDteutac4yaSk+8MNyxhLlIgivzsJ901OVBY3IyEuM
Hsp9FoNZvKc4yIZgKS7TnjlH3hPIWJTm28HsVRQzKBSV3qle8p1GX3x4wrYB09So
UGcElvzQ/qpkxpy63zojbJ7ALl0o4aTyApBnrPyxUe/RS6a0XZNZunqM80hWtnfG
bjtyCSUCZrhEwxtWYzPhGDQIsf3BZD3w1uElWTrjCLbvEazRUqouAxP1pYnc0k+u
k5iIeTHtKSDQJCXRI0XfEUdWhGJS++2orIWecrCutVfhKhp9Tb/xofcchxdv/O0L
q5B+UT0PpDyGSPl7ltJxn9yx/b2LLy3wMvPkpt+SrjdkiG4OECDlbEWJcOqcJ2Xn
x6b9f8y8fv1X3tmGuVqvR2vP95pr7Z07nYWc/Vc5VKdyvkCuQmxpxsqD9WYm5NJh
NOWgs05LhNXIyZ8ZFi3AaKbxNgxUoXt9moI1ui9SKDfSIGG3O34ZF/jZAR33//rN
U0jlg2+IMavOLAC91OEvrBabYmKAFaHUWQr27DIKB/6v3MSch5J9GYcRQX+A6IVW
0890jbJfqcwmMyxjc3glTC7Pg7wQ6plZxZkcyu70cEOe2aT755KPWeqKzZC+3D9J
I62ZuD9MBh50yklKqn2Rc6Z1JngznRjX5rznGAIdYZGjtZJOYGP1gjy/b6+/o66O
rKlN/piR5bHrMdboxiMQFO8dI/ILUv94xuXTJqvNkSdTV79KKV63vcPFh8FcnRoy
Ff9AC7+KRKoLE2t3KJlVH7w33rvDlEBTu+tE2F9EyI1Xg4dQBWDNCFGaBnw8spAn
aVh9i+yqEg7/IW4F3mY5kz8YuLdVC5B94sWQHvqoxDIKvzDXPnhHEFoyh7DySRbk
CXeh+CrCfKFavzEx+82ELUpwY3O5V1AWeaJuCV0BOfgk69sz12IgjrQM9v+69Boz
drkG7cXwdJikWi1zidDNj/GH7huFBJxENFqEVcRtMws6DLX3I2u1bIrfiRDHs7Hq
WHBOM7H/9IlsHMtn0EdFm+OIm3seGuIXkSH5+n0TQ3SfEte4vNceM7LcoIyCTCEL
FfQy+VbcWF4AXxLcrl5cbCSE/Hw07UYVy6ZRTELeyNeVW1RFJ/glNJ1z53XfaYO+
DYFtrVWFiYwXkJoFLpkRnGAVuMPqob4EfRm2No2MYt74wbqrh9uaF4LgUeXXZqRr
sWoR4x2MSAQw0ie2wN3lsJ9aRjPJvqcMBKGvux42Eo7fI+x5tvJ2GuxqOgQVK66o
1HrAjndOYR+LdMW6a4qNTB9L5OgLUfg/sDsn81gj/KOGOcOG8GZFwcS57cqN85bU
CU9uKWidLyIO6N56pbln9yuuM36h/nnVh8j1b7O4kULcvu2fwlskUVXM1JwF+v9A
Rv9sjbeRPPRTP+OF5Apb1BWExZNkEpw1v7mEyy1SMqOX89KU0ob1lhElv1goUEIJ
7qbt30HCIwtT/Gxr7iO6Rn2kRXYtvOyCm5lcbJRQ2lDpaF4MXfVZcuHLwRy+MBGZ
LMb53cWdjuCtPOFQWCYuMOnEzAEUWpSmy/ppOfJOvE2C9yM0kim9HOSPZdelkSmc
Uun7H5PfnFE6Bq5R9M11+S9Y/f+84fW5LPiZD5hoGG3437zUk4OGe40eOYk+Qb1A
H+08YKTu9uIzEtJUXCLmXDgxws8MjHGkaPjsHVpV0xb5rHqL0/IlWag3IoeLItjX
l2Vh4dtdUy+BtQfPu6xcjJSP2iSmKjJGQPkEke8vDFSr5jNJ5vlR+lprxRw4FIEL
gYMYlAYZ2+npaEatc9Sk8+/4vli9pYIfhbi3jr58KLrIS7ElWOzddsEB3yUW/vU3
yVSiks3mGOPVN+gpF3DfBqQsPSsCi/XiUqYTx201WXMpsBGL0h9OV/bis+dOjVyO
Je/U8OXRqC3/VQbFgfLShu1orKcO/MzhflqX5vJmIrAoy6cKCp1GWY7VzwAmt4PF
Ei3xyUoRY/yxgUFwC/24J+fGa6op7Aya0vS3dz6HcUiMREQEBVeKQotgwrhuQqoz
d9wjnyalhHbpYwQHQ2NeZlcOuq9q24kk7FKi9l2iIMxOEW15mP4v/i+fOfIADBW2
yFXijFoEzSqSDA9tuCTek0fQgsGM1cdAvON0+azkgcQrM/yc6qE7sdOnD9cRT6fD
+pfUPYvu+RYrLw4xxNDue+TeRu5iNffX0gxVDUNBECE/Ndfd308ciZ2jS7RhwDf2
Y/eSZfouOdaY3i3A1/ko+C54ZTMwVuBRlFuxm13WOPpADtNgxSuuMiJDNuUmHN7p
O+XoF7Ym70OoXLTsQz5Y5CkRnszAYNmFi0rmnCg8alVcxldIyQmoWsb+RjnnVGeV
044iqjulI0DfmTjlTHF8A0QXOXd/9avAbvOwgSnqPiNPemsegVDMRs5PTMSyVq/D
uOsa6hPijNC7lBnBnNVnPd2MgMIbeBV8nBqiRBLgjJb2Qz5rVhrasEYux2Uj/QUR
ESyu1qD6U4e91pxTAQm0ntffckXgmy5RKuwd8G+/7B7ZOvYl50KzHGE2OIvuC2KW
d5R0ZmmrzhlxYoTtXpRSP73OjTt75Gxn/maeu3vzJYUqmJgophJ4yjU6/EdG8oG0
Gxs0z7kg0hUFDjg7FgP0nX9qCXKcSZyWjFn1F75JfEAZq2Mr1G+6h/3De9MLdUNQ
B3y+vELcZ1gwIytNhd+5C3bqJs29TSqRDlG1srupNjbo0cexeeKlQsU99xvBvVhd
aQVBnU2CQlkHL3SSlh4a28VqGQCzp66YSG50S40pOkB9Cy/cKUTUVYb+v1GFIIKp
jn9MhaKy2SO/QoK8awpLXlsTIrQuWv80Ld2pKJIjkudoyauMMMXN0uhSxuL2XH4k
lcLgWvMP3ZB4PnrPR9Qi+Dhk3R+ITU3zhofKdGeSUFNdFA1GqXWdAw5ppUCNPHbB
AreDMNDmaOO3wnpI9ec0xNok9bglLIfcC9nawHxpwqfrD3ygmJK5erWcXPaIdUaU
iK7rD+zTqbrwRdKJRN+zlOhFZdOiw50fVHXlp7htrrJ6xaBcnd0N5Wc2B1mww64b
7cYJbXmMGUkl/EVt40ttKxsBchT4ynv4tqVs0nI8grl5TNb6IBvULNNOSu37UkRU
LQQ4w+u3LH9dCghfzOc+hTBb9fflywx/nXCMQBE+xNkj0xtgliXzUb5AsPfDdl9v
fKGqL/zb2rH8r1yA4XNvekKeZ7y6CPEiqaN60LbmIJZtbfRG1XP+n1vMqn5OlnOy
AgyJfRX4FIxfINSBbrHPZI6c03YMoxllxnUtCb3ceX+GaqBGmZt95H1yxynBJ+wF
hmVidZuo6VPpeQw9rhGPIXC4IhnfWGmqmTNMzmd+6QDmO3e72HGbYbh4CghCWiLo
BufZWUi9MYxn1HsqWSz0xLLDYFm41mjD9PRnAephS8oCQfkVnBZlXOFQnx9SNU1z
JBDCkYkELiPkxrykkwO491njtCzVhGCs+DezkT/1AUbzpoiZ9RJ+0rXXT+aIqqeK
RJGqJsA4Uq7lpU3LNRpckfV1WprXr6n61wkS4zqssOUFElp2+dTI2Nh938QZpB8a
p9+iZ9xTcRqoMvAed81qhLsvmg8qoYfo6lPWQNyKl2352fe0bdALDcMHE7Ck14WS
Fl3Cidh0PggTrVzyGEkkSH6owfGaVNFuPfy5dUYxQyWhfQD/jJ8Bj2VMu3wXLVGu
yy5NF1iWwOk9Jg+oAO5ypa/xVdeNu6bS5/ZIDL+7vj8jdFiXUR+HS2XD8FofrN+r
hppaz+4NLVgkV9bRdIRhLcDfM2EGB9C+MMxdDDBIxoKBcJlvbtIEin70wabKJGwi
+EDKGymEwsrv0qnkXIbHpH+5Jdef8nuCOTAuksC5T3hNdJR97Gr3JODQuVK1ZFYP
+pmd0yyeXMhlCssHDmM1SYCwHm9VEIT5Qygy3OywHNbUU27qeoQlXN+xH9G8yl2z
QEFodp+fvKknYsnOOCIfkqlvXE0EyR5MN+Fy9x72UvnQ3p4ggZarr+AAwYQKZNNr
zky9hiQ8e4qIRACIojmLvXCc1XkYfdf0u2FSiRlFUa3TAdkJK8+7qz6dbYV0OFkk
3IeWNBHpV4Q0/SsaJRtZXIA7HKNEeS014yHzexQomDs0rTPpFUyBT8XbnP+GQoDG
9yKVSrDvmR7ojYO+EU/j4go0vAK3RXf4DXwmpT4ameMoWRR9fULUCoGvLCW5MDc4
9l0fJdOMhxLtZ75hDOD5V/JKcGwFXQUpX7LroIoMvmr5I0L3gwkXK4A5DqEWOzaa
biYtKmlbPFysI3skoNuMwCO699X0Je2/i5ko6hfl9pivEY2xlVvWkSquMNQeB5KF
7eUfL6We/Gx6I6JnqrfpX0WrLg3krlbXupyoNLFDGLxSDdsahl/1kKCPS4FFXfBq
W6y2SQaC+e+CUGSR/J6DqS8jeN0K/sUy8/aYjfqqo5DoPZlFh4XhJDYdOYgDrpZS
nyMOvU3Irp4ITQ8YWQRG+8WR0d/6vAiMpt9uCVOj3QCRneB7tZjLBOW+xE13jShH
r27aumKJkNcyXphfiFVSLEAWKDss3JU3ySqHVfu1rjy6OMUbXKbQwDhg5Gjnx58X
NgjjQQZ5T/lELyEOu+5f/uASNCeBoDdILZ0DnyOiHL0AqzVy1rLTX0/nQnSP1Lto
txNSqdLEXJZv4hbVigC2LL5QZVh2hx2WwZUFAJjHEsDcRmCEbPKtkRjd0zJxLUD3
yjCElv4IkpvIgE9c+FCnI5z5mGHhhsSjoAALunt9OyOuMCIgr57God5xuL98csXO
B8JV8oVf4N1yiazgjQeEv8YrxRJUgSu0yRuYsU6MrEw7w9aMAfhtLcxGgQrygBg0
YcnSmSgnjhJq3ATb7NwrfU9Cifepz76MPTX78WwKCZwESwGbg/dI3iPv91ssFLR3
EZAB1jJY6lbe6qsrFvBTt9rTXKZtRpOsy2qCUNTL3T9pPaO3XnbqID2vX0CgnNKe
nN7gLOULQSmnerph2JEGFohseUlcp1/1sKrKE7oGAw4teZ00gx8Df/QOK9GvSx2i
ytxPUjO6JZrJ/JekatYEQLFCHcLiSoVaiomXQWZMGnb9YW650XCxcxW8w6Shb2Wj
vNy5U6GuRwdiYHQf52slMLYkivNuImVnv/Wxxtxp8WR4O5IWWnAS3ZkQzfp8bZp+
OH27eRzxdEx11lreptdCR7rZ4Lmtemip3dJ842G8WxECgkXMn3mcFzYviZm8w7xT
tpdmnp/l/nR6Hl7lFS9YKooPbjqhpWQT0/eJkDPUugxLwrLL4JMaBBMBRuk21/nT
QfPqVo9r478mJXGEdV4/HZj7DocacU4t6FBx29J0Jz3bDwXDv70SmHEe9voucLAB
bSjtZor6Zq5P9eOtOUlr9XWqfHqAycNg0d04sxG9vTCmNoNOSz7iV7AliWdcBt8a
yq47maLWmFyI6QD61fuCWe11TBf1ZtjNn2EymdD3+HFo5lEcEFevb/8QuzMaereS
skW8VAXpeV8DO8BmqSBtrsE+eybimiuwlflvkWa/axnS2GDlRaoXghiQu30CyKf7
6i5jKl3wykd1qGpwLNfrkkZYoRchQfstH7vESf8URxftwpjF2o4NaRfBMY3AFkjy
KTiHnzdTXzaxFhM/45oNfKUrc/lihP/y/ekXDsgonIFrYzOEOTLS2mG3eNWcF7rv
odzpMnMvTA8US1+q9irOz7chYnWZbBJR8LMBPElD0QvG7cnQgIPwearijnFGM6uv
Qb+PK/aLRKnkSHraeHKrKAvTt8aRdFUMbLf0wVhSRBGCd+Hseg3xY1VVheiQxdfG
pOJ6PFFZgkvA31hizv1mdyLlCE/sccqnYCaTuo9edE5ZSDIWyWZitf7dXfMlVZfa
fCS76RqN8q0xgMhbIyuZlEfRyfXSs+hkSlBJDev8ZHbmYFeE70jcpXAVIOGSnVHK
g5OUn5XdIsOCvRzNRSWkgnp8Q/PhkPYOgSvYCgHFWkDs6vFtHyTs33hdUYk5L/z1
JoWAA5nzKqURDAnk2didK3c6lMhobMI2kWcnQ9nxaPzoEV67cogUquS04uk87+tj
0BqkJ4a6DeG6U18nNjjCHMGCOBaQRmh+547JdFLnxrB3oLxEIj3JmwG5T2qOoOF9
8b1/M8rv6VycZaEWuGe0LnQW8c2kHmos49GgLbihJ9AdB65Hje77DVy0yojcuE7R
4M3FwKoBgrq0wGowgTBjOoW3misWrVW9qIZfbZs9Aob/erfnwZyFVXZ55xfYmRaG
V0E4vpJjFNXhNguO7TwNil0SiZ3XS+eHVJoxpXwazjdFEC5CLxoJgke9fXiMtXkW
bpB1k9jcM8zGsOVtS9S8g8ASkTLj4zIe5YNSp/UU7lOEJNOzpNbolkAod4nTdsiH
EOGnTjwDXKhAcTGPzskp00dIxK+7HqjiXkpiPb6L9hiTdG88lcSnink6WvUiWIQA
dB5tG0FcKQG2f7MvlVVKwKUEIMszS+I+8p8kYVsqVGo1Rd29sFfhWqrKRlbHHBFX
BsJF4iLgpFNb659oN91R9PEOktBwxtHkKm+GyGJ1zhRWluyNG8itf3NtaQ3xJcY3
X++WbU+ppO4x2LX54Citx8exIP79/P9l5zPSk1XUkCFbeubTXuJULtgCZpN0RcZb
GZB2O96zbJujjE9zm3rZg1M6w/OFJU4G/IbzuhpobPZhU9pkGIKiUHT/d6nOsSnB
HIiFArp4MyH2IcBRCs5Ws38HnXtSr8cSqsNRLFnR0jrqdq+0UHHlrtFEUEcTICGA
lWOguA9rzo52ww6AKX5H8C7HJUk6MVr8dapUXjSzy2IkfYKH6Jh+J7Viq50EaWIu
kOvJEM9phaNoeKqXuZoHKC2lYI35ZaochPFLmQLNdPnsGSVlGCaGIJyxIaxqu1k4
P/m3UE5qdI3XIyBCUCJJXIFoBxDrG0ZYwA8Kh8SJbyq74bHnKlUCs0FyzG9ra6Cv
RNUnWQeAElY9suftR5UTlalbtmUGryvn8NYCm/aCC1WaQIElZNazDWuQmep7BmXM
wSGJMnZRywxp2Y2XcqVInF25RTCHoQL3zaDX3NOR+l6tycM6Wv7M5H6+V8eo74t8
Jp8VP8uET9Wnf7g3KGCoheV0Xb9w+Ns8+/Nx+YF/rnuLuoMrTU7c9smNPiw5SS3N
LYUSPkv6mnx3OHpDDawjDsTAFx/r7YvGOYUXmu68lBnlgXLHo41qeIBaShi2sRxY
InWxP4uHNAoPkbzRSWrAomhQpzPhh4l6D4b5UB9rFj5y3bH3eIpOKK7PDBNPB/Y8
jR8RkU0wjh+J+Euhs+VZQYlkfy72lJNueRek1opAqLOQ131TSrpwuciBt4YVLv+k
2pRCqRs5ThTcyqCHTKsFqeYNuYePLAkqm11YP3uH9sjSD0xy90frtOr9/qzqPq1A
OEVfgwv6agjPIfzuIx9ShIHn3jBTYpXC2REsL1HxhTOuIBbkz6lULWQ5+rycWfU4
7bnDu82demL+brG/O0VdiPJXacbhaVq8lia2g0RyUgQZmT5ub+Xq2676lmKT0Vg2
hRi5o3SEOxXVftaiwSLgUu2/yt3vZ4be9XyUvPqyBhccA2htLtlv/MN03BITKea0
/Cf8zTmPcPrhjg+ax6Fh4ktLmnyhru4GYdHIZD86y3Ob+kb2E/X+T4UC8H9STrUV
0OH4jpB/O3ZkGL8MDku69w/Mmo/LIdRUBeDaWFFpl5SrEXPCqpEmatTFNFNHF94F
aDcsXxT08OlpeOyKaCSpIFm9jM3NRCIbveJ/qYnzFiVheSsj7tdjuF7XT/wB6b5y
XtMyNQetZYgooieq+3/MN3iSa5y753neTO/0wIfkfUGV/p7RHYf/OjQn7DbQ8RBX
29GqhKcdQtUDC4kyx9IWEWq4apGEwx+Bacj1r7z4WUQ19cR8gWi40HKJ7pYTsSTU
Ym2WB1vfB9BsAJNLg6ttS0q1afmOAEEtnGMViY5t8bFLZL6xa5vUpWaXdgatrO4t
pJRezRzL/nxEvcwUsl46a51VdxrnjgB4JrSKr/fnl+RjjQIovxxgWAF4mX04keW1
Q6VFYozdE7nIGQh+jQ75miPtfmzAVB9vxt3fW2hIHh4yRqAkTrUyi/xEus4U5aLD
vu9szY0UOcHzjvg1cLnEGH4O4eHxE6K+kDIsVQmOMvN0lHofPqEOzWDcWj7lNEQw
xK3vQ5znXloN9iKX17co6iXTsFREWXoEvlGRWIbgmJD7qnfE9lW37oe+5dFyZdxL
Vazaeyn2SUZeDK/w2T9ioFFp07MPZjs32UDPu7yzVkNQxshKN+GdW7xU+2sMQR8O
zGlKTtczgZFWiBJb2LIRukN4Z1kTiBF1NIodwurgLdnOgcI5wXXvgH6i3hc4BKbm
kJSsKEyWIH25i/3TjX2lNcdmyWh4RK4T0I0Nn28hKGb0fMkCFGN2baX70aU3ErmE
GZv8fst1O3LjjG9MPE1rQVWkr3xaBxOMOb0ODlyNhlk0Zh0Do/RTzHcha0F94md1
ki5IAoYX8QLFEJaUnJTijkJpnQ40729rRvvihDZu7SMA0/Q9Mm0PBElXZFFilGex
VAO32Iz+XpTWqUu9MxYWeYdcQi20VKFRjtmE2EYD5rfQ5Ro2R/ICyeHLTfXzbUFY
Fuw9h93d9EyuOXYmSoaVDa9gKciiJvuxxBY01L341M8Pa+ZK/jLu+km0oa9glR0G
MEsDxMQzVxV06y7qQCOlnmJh+bomgV+vLbSqjDuxkrKO6JMso0EjFXHfItz2rVNr
kSDV2VcMp5sk1iopXR/TnqQwBHq2FaIsJmuHYCqhExQd55rAlK50MDEI+tvYyhvE
Q5W+JUZBgUx5jqgvUN+XcaMI387BO6p8/tw4DGiKeVD3c3N6Vth42ScuscqfPPYx
5QsXJj9fJlMQVS/vy4wqwNF23bKw76JkSaGfzC4ZaSOvGJl/E9L7npvpT6TmuyfY
/gTvd1H0nus7dryZvJnzder7v+/i8z4s0qFC7/G//bcQG7gVEc3vAp8RKlL2NP6a
yPMynYT4zR6u4rTkHzrbkLbk1tu+Zqg0IdIxCZpLX7D4jhf4Yqj0rK4JT+E+pnCb
Gv18bV0AS+FJ+CPohqqAXN95ncl3BJachkBu91OFeymU7gEOTgtPx818Tz0pwXUd
5CBcaP1iwNtU0g9IQRXgnitfHcGlJX8cTZ3CPWHxfjfp8fI1N2yU8a9JSmSWYXX7
oFUaLcRVKGycVaHvBhqDSruTxpk8tV/p61YMoSGrYaSo/zrhJXusDnBpRLoAAyLD
kM+3mYhgGk5MdwBBkGQ6mWS7m7lqr2KgnmkWbksX/U5BlUxPG6JcEriamAzm4lVI
32FHOZeyxayVM8EZ0MMP0gQBYIaIpqVsgqEA67BuLh2mDePOn6YB+Zj8Vr13+9EO
ZVvs4CFWcCV4HdFKwHnm12CwUpcuGP1LYMM0RUv3JG+UCSU2ezKJBIq0KMO0wj9Q
BKno54UHMcCnoLVRovIeYaejzNuTP3TuZnBG2Mi1L9DGqKIG1D5v1cd800g5A8O9
w9/A6OEMlDd9CcrGESxDWWTAgp/LZsiESPqopnkSz9bzOVrHUAN1cb6NGEhFKJOY
xCtwSjnJsOdwJG/RRkP/eWUrywLqJBGSPZOu26kFVbUtGveh+bXp5lnp5P4XVwLT
EKgxAFnboV1s0zIzWrrRD7nfedNvmeVX1M6Fg4lOFikugzAPqvhIzHeh9KBokS4b
zx9cnXg35UJ3hH86awYl+BYB5zLom+q+f07KTPnqEgc5TysHlkg6aIa71JWyq+35
jXpGeEhjAG1716asm2MmmbJNV7NvzXC208Cay/CxSMLPUDFCS5kMkHTv+CGcBpyL
SgxKbvYmoezq40TojTVT4U7dgNDFzA8dqp0mTEHXFk7qY8+qlrw1DJ6ttmIqVE1F
grJxnv/a/8A2IZqeLDG09zWKDPnmo0Oetum1bbW+smONI2rMBXWGic3YgWU9j5aX
HsS05w8fNHZM7pZ9QdSkyeios/RU/TaiDzTUB20zoidGBotrApu0Jild+xcpr5S0
+GrUkJipOnSWrFrE6zbgJAI9m90VW1gNhUZG1TKxs1CRUPABGpylwzJQX8nHxz5J
zqI35U0Vl9jpJFssIOCKbDmz/suB8dQ69gG6ASDX1NkN3QcnKscuSDONnpXzmOie
EiDwVUOGiYPf1liqrQmhjYLNsEmn5pb4Xl17ZSv/kmA8UMHUWEsTXaFXcSCXlpIV
YppSVOMR8PVQ4goOLWvQ8dTVAafESRR6urWbTWZScVuPcYyxPQrdAWhKoHreW5/2
Kiq4iJ9nYLZnWU4/fZl16Q2iGKDySFortMKIYSnstZJWiP0n7/oDXfFCZBMY4h4T
9p6oOzEBSeNMEMMlFxLM6DumRFDOndiv5OdxV22Tbx/H7REfPXK7luGXFQxhJziS
xdt2YF0WtYZ/UDepvkpNsHIT1pUU/03/7arYlZoI7BFKPcxyCeOvjYtw2LP07CoR
ldgZoPygDEGvz/lX6VDKPAT0zljQ4uk5tSec9aNpIa41giWP3E9EzAHxPlVCxq4p
SRm5/TDNAIm16D8EPg9Kc++S+n5FfvZTmuZHZS0WVknUx+zX+rzI2nQ/EljxjEnT
+ucTmwHekmKDUzslAIPiVdWO635M7BJXpc/y2OKyrZ2KIMF4CYFDBFmA+/mepo5Y
mMVU0fvPUn1GB72oh9qsFgHvXcvBU7pz/jCqlFz3u7pO24sV87W1xB1UvD0MCX2w
YMW23p6lbl5bzj0z7kBqSSo+vUSnm8QOVicuOk7h3mJmTApTAP2EMqIquKeu8rqd
EaEYs68PqvtqRQ8WqO2Ioqt4+33ifCvyultmz96w8uk4qU+GWGaIz60mBMmEOozW
Ytb4AXkcG0AeLdsZd2p5vNNSIBHWmzYG+9U7TtDdqS+V9DlFy/ANM4AnGYgSFitN
817ftqrt5fLB5NUEvKzsKvtYoS8a3qguryOC5UH3H/ydtKHY6fWYTJVesaBG4MlF
BYsE/ogLCrVdchuJkdukYvrquh3Y1OHpgsaxIOn4jgLsznrHx5/tqrS9B/ci9hQy
9MCd97vLRgnNPRjL6x7h/B+Iu4Pm/DYvV8ZTPQ25KYbTVnH5ToUbc8B/g/HGv/5Y
szxFSU89ZWbhfWKm8D+nDGNGnTxMYVl8pEXL1RCPCRGPnLeQk22dcmr7pGUlHBjW
o3miaXUiXa8KqZC7lFdNdegpqZbnpGGaYScljn8U++kKxw5khsFeeQRpDNO8ntS9
XVD8X7ScIP6VXZqqlyrVFxMirN9BpMx02lEnEDDz9sCuTNrrltAgWG2boLk7vSUD
TCUZ425TEkeHDsJuqBSB95JdUvVc+ugZTO75EU1wdzDV7KBHe5SiMDnUjWSbqCKM
wgLnohSyQd7Mpl+yI7xrxMWil3OySuZsCqMLut23/ZIp7FTaBaOXotzf56Lw1JLG
1IaAZqLXtG9ZOmHW/z+pCRnwMv4I8DnjT4qXIt9s2LnjF4N/ucXNZvy+hlJxSVca
hc3DYOpyxpEt4zgR3p/fH9KcffqzkZGrr2nqzvIzmPBLEDUSVQ0s5dNUkm/Qzm7f
G7xR97Z7G4nH+rxpyxrq3vwJJZo7VRZu/0hK4Ts21VzVje4zscqZ6r3wTgO7gWoH
x3Gt+KAsDIuFnrwATDERzCXn08kklwGYYdb4lrEPgM+BG4Ef+Pxp426sloo3wKEb
rcEJdRJ//hjVqdD/zaCMPPKgbqEluH6dLlfE+kQ8NPccGfPtBH2Plz8s2lEywWE5
Yo7x9fB2HXNKZ3BsRBtnsnKt/vN6MJQmiqkmZz2lkMAt1nDmTLltS9VQDsYvsJGy
vaupcrq1i2rkCzuGMGzx2Ve0DVhskCFagFkfhVGClngKStANR9p2J0E7Poz0a2RQ
2sbhiaBRYHZe3GexI8mFbX232NT//tIBNJQuHJdb01DzkUUL78hDttAdEW07zAhF
9qToedCZO75g2J/E6Stcf0weOEVkLxgn5OvURzxvBbiFUDm6gN76YyuetvUbsT+s
0HgyzTKzvBqkp6Z7y5ld1MjMBZGmIhUjSn5VNtNb0TglBtmZCt3FmqzU001ljCI5
kpg4HpENVvvQ/NbSA7hkt+FB6/vKQd8etb0A66AUiE9TgMU6WvKzySKDeLqJFAR0
BC3s3LsFS/dck+SG7lY9D5sNXVbEf431CEm0uB8EONEkEvvWEgc4Na3zCumSnaPt
WGf1lEW0nqxSGj++eVY0Yqvnz9167x+Tx9wopRTH2i24C65+XbMDZraFS0utqX/R
k3cFTCphy0C+YkGV0gTUA5aHmV/ZBgDbhuRhGM1GhC3Et+Vn7qovPKT3SPSLZcYU
f1w4KKTHlZWPxO/yqoNrMn096DC+2SoQvSaR+nhBy1/p0fi1B5gpx/R7s8oDh0qm
naf7jTSysJz2XAUfgThK6kTEIQ3Fgi6U3cnSslf8V2s8duqZrC1P+ML+2sE/s6uv
cyeUjGOKWTfPZ6QHyYq7CxuOwXw7DKSLSsYXquqdLjrpavkWyifGIgQL7U+ZX0z3
f91jFpjzOHvnxzMXLlFesHLTMQEs6D+zr5A84w8DvrRniSOOYvuaVBKliTPbJQW1
lcLLH/Vd2OJ5tVL0kyM4/Ie76loW8u9bqe3QQPRnQKryJSJFlMiQGEhPZZXHVwih
5ahU+YONX/9YiaTAvttBgocnXYN2DA3KkOEIyx6PWdFhYsOc3TwPKblgvC4FMbqa
DjKTXYy4oWZW0+wplW4cUm7dE0y/AS8pKpn0ocEnbNRGcnlYeNR/4qZHVlQwQZ5h
x/wsgVHJ9PRH2RNAXgewgbSfSrccg7c8TitWwKrWkTDp5AKCHRVmmc3Q9ZM9ja1F
8BfIAhnDicebkdWGmDdruIdWSTqfyza0M3VP1rBCyh4D05LVT6CVIbuOzae12/VD
G36LInohixzA+2E6jocBIZfQt8w8bjlxK6384vKfQJIQPPXRIgYg70+zr3l44UDd
qVeE8cMXnCRqGuM9B6aseTYHCvYUaZx+MiqfN2njxb8ELevmSLCyrDCoAkk1Co1T
WIlR2iIZjARaeM+TA7xOYSU7VsKXTSyORUcLvZxRWeKA0Dlq4nPb+k6Xy1CosxLj
4LQ0+93BcHW/Aykuf/6CLPh5EcsDmihUJWO+p9LEiOHksNDdciaTU/B7c81CHxO7
zAkPohfYEsMVG0Iv1e31xF63pmA6xovqfjnd0suXJJFVF9cUd4qgCjPSB48lkpGr
EbqDXNCuWULxYVipueIXPW7ZVK7wrb2hxRRfTu2ofwAxiIgzYvrK6wBZxy5eVrVm
UgeguQalqrFPylRkvCNsdpUiyEC1QMsenvKgF03ErFY4o9ostf51I1JZy3KfeudB
EW6t4wOGOAVRLlVgUBwj2CBehzAQ6AoHViXUq6/FHi3mNlfrfGWZcH1aZar+C4nk
9tUZEG31ZDlsF0AwKdzrvsSEpffRzZpLI3P7GmdyO7sCU5q1U1XZCfVjgp9W01Zn
cb0d1bd8uG4+ZJ7ykBaedvnuJ82yYWY3+vujnD/FHmxgRlgJzM6vuVC6mLx/oS3M
qZ4EGnNhVyMlzqODympFr+TSkurxxfqaZH2s7LvyQgz0P+fReJO055lB159zFVGx
oB4rc+Fl4Q8WMKDKiwzLXYZ9igPY9vmUxjWS+tvqePkR185aECPPDAZ0wEWdgg0a
Lp3JzIIAIO10CAKqo4B+by5Ve8SgaCMeMjEUVgy1IiwIGBM179+VXXgrggG+OTFz
m4Cg/baT74mKWz2455ZIoaSRaO78zYvFbcLmOWQ5XqlWL/SX8NbX/7T/LFJOL7lF
dew0/zpzDFkwzBkq1esST6Z6d/CXgFJi0kMZCTvbnamMheNH2oCxzHJnobQglXHJ
0WU4t5fDppxRlGvFZKtSsV02+C5+gLrkaRBRX1lHync1CYZaVc72x0N722nmxg3v
lF/8cE/OOCdd3ju+3FPmmsSdVoUh6wTHDeP5zHJw/cY2ezruk+rSwXj40CLViboU
Sf+9HS8Oy/RExiSzYLpeYVbyL5FhsbOrZBmeEEH/OmVrDOYmty2N7m3VhgqEHxUQ
toBFccawa4XjCCF6CSBKBWLbQB3bt//lHwBNWx1+5RXgM4yi8a/MhaGzZhfgR+bJ
Ean+PLfkWzXfDzC5gyPuVU+XwPBg6290uGTLU6snxd8txguHd74JNd2SLXvD3jPb
/fgEaYnZ8vot8ZFopR5N4vng749iNncohQkJf/f+z6EyIElaHLpGMH82NAGkO2IS
hOK8CWuNBqhlIDfpCTSrE8gW+MbLvnW+ptZix3Hau/WiWJnbv4GcMySAyHJaaUTK
4J7M0GHhLI7Od6qhubZnIvhUJMYmE9lVmYIQevfomZQc5hLS9uoU+Fq3TOysMPqW
kaNdV9vigLJhkShQ2ov34C0SfHNiiPQBaKZF9Tv8fed17OTfaTDdhD8lkFFcfAHQ
wNi6olfcvrdYtiOKJi0yhrsQuiOzWyPC4bnMjIB41hBotGkhxkWjvKG/k3NBiof5
193nN1snLA5OZg9Lhbd2z0ik4FedCOrIK5p2SYG4GFlFcXWIzf1+1/W8PFuUiaNE
qJa5h8HOQsWjnLfcwiQw8qG4g5Sg00uHJoadKpAnPdwuQOhLX3vOz/puvGehi7hK
9gsaB6w/kTyeRN4Adj4vaW6F0FhEYmO6dqXWmwLhl4hB5bW3cOlgwVdVzeafXpr9
ABh2RhoFIHZPw9VWovm1zwXI8/nySZjRCoXzyDfL2QGHg1GwUAJp2uEbGzoFPMER
NelwgJ0B/pQriWDjbQPZEa9wZc/wRd1DfnxvaH6r2WdF8NDOqNlIsSsnqvnz0q+3
VmRcZd4y9yxx4yzoebBVCWI5cSfTxAcZ1FFU4al9cgU+NiaKCcaG/+y775sX1eto
cczvG4MwLpsuUD14Oazn2b5yDnq3E+vMnfcxdME8AIPNssHaEWDf9OhDhcK9XYrP
PeeRPkxKNalHl3X4ZVBzCOugEFdFynA6tplkAUFZ4UmAl1BMjpvuKPqUjC/zKJjJ
93cYimEmjG99DHbCv7HCG3vqs6YwriOR59hr11lzFdN83Y5X1EZiY9qZaEjRpQAt
PmyHPWTK5XHJHLGG1zIWYJzDee6G+jEauTwlTLBOQGB7FhHzLBSoCii98AbHJ3vW
IVNJ0KIbnZrg6ZY8ytqsWaQILxEc6+VizKpl6jxxpsEZtoMddYRK4OHQLlirSjte
r9zdxsMI7A+aRjIk98hraZ/nrJgLGiuUbnvLMT4IgTCa8XarnZa0jDElXffJ5mSU
6vVgLzXqYyVSyn43C5dMefaqPoXm6qtjm/CTQfSBtZK2rFZS6cG7603/Nedpp2vz
pN+kmcBVpBQsBRzEHS0abW4l1MN8QbhJ4yHDuuaEyyUHu2LinD9U7GrPCE3/bEzO
SPYhUqWJMHhgwGsVEd7MdNa8hi0hm86pLopvzRxGi5n8rGo4CJgBdaHet0MSBNRV
3dfIU4Aw9/Mz2lwhlyfy4cYv1THQvZNqP7BUcaa7k9PddO9B9NZRuD+pUyPdRhu2
xlkURxQpAZl6/sfkglFTfgHYBGzzsdbNC00HSv11ntZYIWZdCnGF6yALDBgiMEUs
hNCkXXvqsk+gF5K33FYxyWTynSP1QN00Is0xbBxvo1fz1Lr9vfuetJnd7kd6BjxY
LCQUDXs7uOS2ZH9Ej1jF33NK3RGv4EcNz6vAxsuRdzJTQn4ARlsilWc5on544DYB
BUkv6hp6bkoxEIVcVOulQ2J5tfqzIrekaekV9Nfhmeo8BxN2b212yWck0Lk5WUF4
v6UgqAFhbgPrbHshiVwIJKN4K9ulnK4DDpZZmQwdCDq7ePusYZ3phVSqI0qPIdRd
E1EqKWRdnSIon8tBrbjydjk9dtAUL89ePDjGclacf+Ch75pc5x/knLuXAA7l2B6e
vlf74ojaCTNQR10sIlnZlLngmDi5K3DMxfBslD4qjxI9YrL1jGrydwLUA4eYP1xR
QGnQ5ux8r1xdXf50zZB14g4NpgihUZFGYvNo5nKak3OWQOZ4VZGMjZvK0QPRaTGJ
JnHDgM/USgTZKqCjL6S+iV3xp3TN4SQl8DVsh5Y4xXrt6oJYGqtO+yTIDxtcR0Cm
j25IHY5iWuH2mvUzF7iW3Z1J3yV/u79hJth76vZW9bUODXBiiHTZJ+r6agPd1Huj
Pqu1cNAFeU7SCzAmlQMuWwKOnt7YdOnl0bPo1bCE5zg0qzn0zmZvhpgGlwusDSXY
QcVsB9tJbYOvsIx06cSgeKBpJBLkDgJlanq/1rbHV5/tESM6oUN9y3PmTaxdC6hA
oqW047DVxm3u12R90fPhloehkPp//7FrIlcw/OtpzznYCBGnwYFVudbKyGqQnwNG
UsDzDToIFYC6LSVoocN41hNCsSTS9rsfiJX49GLpZTr9eU0LcnNgZfD9vCbWtujx
dmuozwVRXtApfUoS9J+abSDMPKrTpxHHphkBKBxX0xpoRwOzJ4A11f31yDeiatiB
ol5grvyq2LLn5oauLbYNYwoLzlhtJlSJJlQO9s5Yr+il0Hc1EX6AB0NdoshFOkTg
5TPlJiUJPmgd3gQE5XkzCGplbW7abrNVGf/PepK22Z/jH4bNfeGoD1YqmPZlTaku
I4ILdpaVDMO8WmrGu6AKxFIeKOo4ReBkRjU1cwBCtagSSAiylNeiji5OoFQ7tAAW
MNRfyyYY8HPepRnxMl+4MTuXWLB7tNLZzL3xQ3zy7gaMh6hWYeGCqh8L2bOPXZF3
zWmr6QiJzM1GU0QOQNv/OHP4x6gb5JyJYOTDtKEMFF7qKZQP6ZYk2CiUe7ghRdIo
GPGHP25vWIkH4yU0SLV2n1haxEqodyHOWv+HcQ1t5Sp2eZ3cHGGz7SIORKkYg0Pa
j0VlqtP58CDAD5eSURm4A74Jw/ENFdmQDuW1pGJxsIHfII3WT++yfCmxO/LHI7aV
1nKsoaOivUo3W0HIPQ8Eq+iAPbOiwwhtmWYI1e2O+WZ+wUbTHkjWJlFTMqUAwlfe
kQ6vnGNukqLnEbTi+TrX1jfP/w8fXToVL1Fx5AT9qb/AfGX6Q98FdOMUMmOBTEYj
EPOQ1VCu+7PGNBxRqUWu38pGbx8QWjKpZUSU/vBIdgyFEECMIV9VowEZWIBS/9/W
cILuWhzFvPnWLQk6oLViGiw5ELhMyiDtatoOLeAoMncDh01H7oICyYriETlPQhP/
ltLp96+ZN6uEAbbh4Clj3Yvpxcy11OnHDQRujFJ1gQnAO4oV4JTeTaV2Yjx5SWfX
xQaZbUjwJYJ8PiLUklj/ItCHPCRMBzry8N/Z+a7nHu8nsthaa+eImB70ZWGFXqk7
u4OgTjyzhr5hQj/wUeiYfrBFU49/JoOdr+xGKJ6M43ondbXrG7at/icRGSRfkR1H
fz93a1q66UDVqIBz+uEjDqfLPfEAjWj4bzYWKVO2g0NKY4/ebEgd+JT+pRW9pBkF
uWw3MpG1hKl+55Hj2KDssv17SjHqmjUXDRVKFwH849sm5iojE+yOD98gjSQExprj
FUEX4FHW1LsfBO5WFqqFiL4alVAIrmlqKSb7qFA0mxB/v/8xVibI3N3P7TQxRJiB
jfl7CTjts5u3zs3XrmUXeuLRdXV4IIP6+y3CwckVbNioAaHCkno9ftaMarfN+0ER
TF0eom/5Yh9qiunhOSMNVSSW3jbv9e3Al7LxryWZoIFkAjBTnCS7UyQG6Vx/t+Yd
y6pwZBY7FV+3F+vaEzUVYxGuaz21cAp7UEoXgGXGomAS/rNVI42N2OJQdjPpO3UC
RVA7e7efGh3lmzjMReqCo7f2RnUlBqUiT07iKsIu/d1SuC6ShkwbdW8tgTvf747X
bpEJT1uwrcWa3WTJSynYVtu7AWz+IziMOUCoS0r6U+XMBU2951h+DQytRjHJdm1h
kBuv25sLbOj46MezF4yi+2wCTHyr0WBTOhGvG/AlWKyShMStLbSZWF09UAvaP6My
9vwFLcz7WHn6Ouy2iAAiO4yDDx6yjYjaLGrjDTRXss2R1O0QM8zdz7HpXFMjqTaL
inTOwje75Vi6km6+bdrp3KNOQ8KvadOYA2oU9P7iMti7vcJqJhtQoXX85zHzHZgI
ybJJ7Hh9erBwoYtZUE1FLCB0u0rcpr3dotjApxHxZGZjQR2k6efvyST0pScZh2Eg
gQaI/gAw98pmYHQ+7TMUHBDuv7j82V2SYsRDg59SMG2oxAWA2cIjB0FI1XxGsZez
yEF0lBSymxhJx+JwHtW7t5kXrpn+IOxj/0ND0zKQMpW3/yH7jVjIZWmQD5EjTSTF
hUDozwxtWtYWak/41uYnDL6rqhSnc4aCLQ20avqmJDGhTrTK99q6aePpT77zFyxw
pLLq3WsAknZQwH+JKY/7NWMC1MF87I3eEojUWkzf5yHoLBjMLA0t/dIRncQW2aq2
/9AtTZlM6qMSv+FjRToL03nCA9exM3vMGcN63kvJwdWPjW2oLCKO3GuYD6bel5Ri
BxcTCRepgT+7LGcbwV/7Yv/xVTItu9BBeJW05c5oxli390JchyxamHZurnaXqSgE
f3jfExcGKz/tCnsfpX4T3g2TU/yOTF/zAk4KF0qQwE74UMUpX4DA7kTHDaY42ToS
IvWyt8nKktg/4fhZ95xXsSWkL8NpyMx9Zs92/F4Mz6oRU0w/WP2qAXHjDfmKBHoF
NBefTh1fg/Ki24fI9jTQMvqkVrfhA2m5cKXkiKxvuw6d0Ec5rMQkOfFC0jLmT25R
+4OU8/DfR/TIWDPC9Hagfrt+PCaorw5JsfYFDSC6zNMsyoHZ13FhU0EucuHP5ZCj
ORIgBz+EiGWyC0IDL0r42Z1ublFJUYBnEgPXeouPYe8kNUIib5VLSY8FlK95rDBy
Ot+i2Zf2bYLx2BjkfmRofkU6cWBLzTEPGbNKPEkOS+6g7y5tdzsHCmYQ9KlKtWBk
t8ixIWftothzdBdm+Y/p6Y0U5D02+jaSWxOF30jP6oa80IbWWxFlcWdmwL0GlJ+f
l3SZvl0eaOoOKxOeBkD0YusnHZ9DEvQzLG6UeOb2ykJAQHt+kJLuGwiu7kXNUgTH
kha3abQZK+PaIME0IWlIdFxQ+9kUP7jPoYJ3lW4b1Tl7ul9CeCK6wc/VujvaPLzx
qpyYb4Lc2ViR2bNUMmW2LDVfWkJno5TYyDqnOEEZs8U7oUmT+z2W6zjs2Lcb5aVX
ZGYj/DJ8OJ5ONHQ6+jQlRLTTiwwXOMgAdvyjGDT/jdA0bvzjhEtRaoRlAn7LHL1v
px3VXuoXM+tuGaHqlVtlNDVnBpXrsHYpZFvJyTClLTKMG+BUmTmsKyJHozSNp79+
WdCFbd7wqi2YL0xj5jfGCZ+eDgwMXWedHkRUAhMjoYW67YZ9WUc0L0DrKV454Qzx
gz6kPG2pnLw7sFiiG5bHGOpq+y4G3EImGpx+xUe21717mUjJljnYFtelpEC5UyoC
HWbhGBuSa5Yysr/krqQTO2aZF2ZnZwKn38PrEHvsp8j9Pv7h28LlMg/Tnwms+2Ne
BcInxAaz/q71VOnfsc52m5SLKRh818y1UGAi/PwbhwJtxbxrLqtmZwJeVTbdBYdD
Lwl//Rjc4W021cogNUNQfJ8dkYvWc2N6+3+v53gRjkZYBQhC2mPTOu85VZUOfXjS
tMJHwkj75cSo28tHO42Cdg7aJ/N6Pu9B1TuefHsjBUsVH90q/EckqXJfyUwWHiex
oax3jxvNWRgPLWCrhaqMY0zUh1gVdhwxZ8bx06IReWVJXkeRWkqfDpSa4CVN7w3X
rMkWswPG3UZb6sbfrus+w0UwHOZmPzvxNYyvft3UAXuHsF2isFjpwa8ZgfQBRTRw
CUGpZAPzdTh83CH2uFdFfkFpLR2XrlxpGqNuDRF2QIvW8WB26zQbhWMWRnKiV6LF
/6/RCSq22jomJp8hf/QOORVodOTmDR+I1vjeJK3FFUGn2SHxvzHk9BbKUGMkvHGq
uu1iFrkXULV6VvofyyNMCs10EARZGHtGXA6nVqkfXO/ql+EGMHYsRgXnHRdzhAit
QKo3zYBKAbIBLRomxyCu8ME7TGkm2B9ch9XsoKQMK1734qvBJrGwkMcbjBU0Moj7
kiMQucFsTVXkHJZ9s7EfwkB7pWEbg+OcfTOUEIriG3aEPLq7rvcruzqhl3zdnKGX
Mo9cHCbcy5Rxd7xPOoRH/GL41ydvQ4s+fQj+Fd6RukltTW1zdjtgVixHJ28mVCwf
phKdMJPGKb6+MTq+gIrAeB9W+cKE65tHNEM4RkKq7o+0Lpn8QmCza+fBG50eL56K
h+LyNKzwJ+YwwtYLyIqor2HAGiIOncyoY92414Z8+CyZFLeHA1S1e9x1dKiY5JB3
0Y2ig9prLHCl7tB1CKuwEXCXwejEt3eDMK4/qkuVsjQP86JqHlBLo7hbyMCpbT5K
Sqoo2c3KDpXyscsdS6CCJb1WqWdRn+6L8Bq+UHuAPon3SLGUDslfzp0om8+AMuXq
pxRqk3/LaVOplZ8imHB2wQ+OW+KMTjl/U0GkGQOVNJ8rrNj6ijGaxkWMuI5sfRs0
R9HJxrCma7JP1icOJq2t8VJek24HKW7l2xQyBObReryVvdPJeHfdxuVpg0gEun8u
Huji2zly9nggjppWSw+6jZzu09mtVDXLQNMaSJcxFe2XlpGdk7eUQS9NTtpZxWWa
+/XAr2hJsfrEfPKbC6CubED6qBxMBpoi2kHDtuhwUSN4c7Iywm7WNOKaUQIiLkgw
Fm9NKCqpb8JvWKXYMMnpsOW6aZsIp1W6fDYAtArzS383utYK30lh13ZQm7/cSJ//
z18zRHneTUZDaE1MGgHH9DEQv0/Qz5QN4M6fdui8FAJ8BHvvtdp6keu5tWB0aVV9
hurGhN8y7hNIcL+Ol9d1/TKlcSna1mJwuIzBS3RxtmJ+Q1OczmSu/E8QR8IzxbeH
AMPwuHmze5GEf2c7g4PCVyobOacSO34Q04IfliMLagOqAfgmKYiKrV020ppELs3W
yVFJbh0Jwqfr+op2H+9Ne68jxl+pxV9sj4O3g9N59udGH8zvcAufUwFTy3tPA/FL
HE8TQg9bOQPo/J6/I3tA4BnnTLBtXXn+3eqb7vo034vontcC9nfgelFToWcwvmBk
bqYJpUkm7prF2VXX8qLN10jwjuJ8Hi42MIisC6svF7+t/JSnPRkpTMp/oJGDLgg3
SWPWz8lol0AVjSJRAM17hjMf9ty2qfX/tho0wbo5p+d/YY41lzpZxRfmPomBWDll
/m3jGIMjl6Ky7I0+PNiv6dGbSvl4Vx1tf9Qx0MZuQEEiKSIB/1DWRgDg4Ad174ef
Fdb0lKqTBY8ywSvwManB/LrMC/twKZDh8INrJb9USCLZogYoiBGGhCns6+jtarBS
tJIC+EFupsYrDD0nOy51Qf8Ehac65JE52XuNMpSwUz+VhSy3m8EgNlF8A966hJS7
3NCGODtwX72t38PmoikIrB2SGsv2XVVJLOusIV0ZyxP8ii283JdPd9mIEWPRWrmi
qpZYApDymZ3adybLNSAY2/k/nk6LqaWU7G/96esZ+jKp4K9QymqxvpaeE2P/ZoBH
4SUj+VUziO1lmpAtqUZfqm+OaHU0NmWJcNvMhKkDoC8hVhay19HXz6E7GfSc7N2Y
7Spbx6i6Qzbs7oboNS/HhAJKkYGx926ZoSnMex8Z4Qrwjm/4zS+Sl1jdXAR8R5HN
WD3mQtz8hbHgzACmR20fTl0bZ/ey2wNI7pDxWvwDHKAQy9myHE1SimvFACcqanhh
Y4/vCr/Ee/yK52/I1Y0DFmQ4Sv8Y47PmSgvCY1u8WSrw0l3oLvW2cocMwi4aM/uM
S76A4kg0kBUIGBNDYn2EMWac5pG0J4NZO/CsEtRDe+ccGUkqOPcBVsSB0cvRrkbl
Pa4ef/pCOQLq1uDKnre20cczqYyIDZZlVedDsSk9JhsmYgoidYKxSzJVp3/fmpQC
IpajvxQ9LdLKlVwVKo3On6e3mNwLfuIb/+cn5cDFlEfCvkJUUmPllulvuUvZQGzS
f0UDMeXdDSBxhehwoaupyRBdo2ooVcLnQ6Ixz9zA5lok/FJBGWZ4Zs1bNGXTA14A
YYDLEK/PlNWrQ179pBOkSXtdxr8FXhnKdKUczap56oAZow4yaV+BwOF+6OGhRdke
9an2moFw/3Y/qDI04eLu3x8xNnIZnug8hiQnWDWhXr7/9GHXYEyC2Io3mMubbfgi
FsMmCHIn0/xunP0vR4pB/8UwsrjB3tWazvbFrPa40+GMizDf0Z6hjJD6ZBxIQhD6
bqIncmJ1lLgo2GTglAPSO6sBqAfD73Ph3lpZ4ZeqjWv9kwRHancg5dU37UUqnwva
RKQaKAMCIkScwu6iaR3L1v8Ng782GONS1Ytsls+b3e7Des6lEd78bEkTsp8e7Mrq
vrTNmxtC/wEVvBRIZSzdmvFHstDJXO5Tk2sKVYROAPT3HAi0ZUdtHhIptIVPCnUx
z2cbQqh9h3xS6XBNCengbysPBOzcdIgErbtgJ4mvnWGybAS/ftnWYbWed6GU93CQ
PlnOyVd2OKbt9NjIC3zL+iaK6RZpG9UVhe7YWqjKnHkQG/7f6cA3UQcKLD00QHqx
dfTCIRd9bFGc7uJPwCkpZV3hNHcL3ClCJl1ysUIoQ23iVJPYbJ7q2SL2qOn2uqwx
KgxJAuQzMTwn+XICGBDuCQz2muV+MuVSPHsU/sn2KVa+aYlaEspl1MBxynM7mhn5
a7oQTE+OT2MRK6XR+vMb3Wm27Db9F2rAZymUX7goOEcp8fRqEkeE9ehFQjLM5f11
8gfdQ4iumtu0hHsMMgBpAq3FQgyQyd8fWtFDJmgYyeuGwmnBA/yZ9GYysSkWM+m5
IHvQN5r+Nk6MfW+2jRwQdtYsL1jo6gLbPSLJAC4z/x7XE0JDRqCRWWd4OuZPKmRi
/Ax73W4CJ9WoIO2aM25vJNRPyvtDXbqlSgj541N5/xgSZXKJdp0Pby/8ZIyBmMv6
To4w06R0ySqqUpvJ/Jpt28etg71EpqFHhx4B3PEikJ7iXIi8kBxV7d5WEsv7qo96
nxeZcKcFDl0zVnbEWN/mR2P1mUlooC5szuQJPVgIyI/L0kYBlBg3lJ19lAlKC4qq
2Go5xCGH/bDOc5+wgukmYLEevcHyu/OGJ2omMbhISbA9Fllx6sTyzxf6+fSfmzqw
FfoaUCOEFYr6MAU4q4owv3Cl6kC3+jc4fVTFWdnh0yrZbM4m3TcPuL8Eop/4cCwC
LPpjuGxgfZx0KAJlmOIhN7RXl1yhiGGPTRbm7Q1qlQDhjFafWpalMf3jZN64vRND
lNBKE0lTXi2ikt4mEvzNMG+DIMqy7f18imlibF97Oacco2OH66mh9ps3VlvB2C/c
7Ih1lhfghd3tMdpm+vACEfwyjpqV8MG/QJI4TXTUBUU4593h6EJtmIGHVGexbcyM
+YFypVCkjaeAnnclI4c6GoSRH96b18MYuZGZOIEHdw+HZ55FVgjRLloPNo/+WW+j
UTKp/zoKxvip9nL5p3s8dlAOi1lEMqO9g4CqeP80fhWH+D0wVHzvZTsW6mMCMgld
Evdg9YYXOP6ZF5tBHLUVOKWXHl5HTag6GYuOHcf55lnK1m7tWqjaBPPajbsHqpjC
81obgF68kspLNc3w/C79tIAetdrxFVUwXbdSy0NhDDAp4idpkVit3ntb6xAVKb/K
1DY7Z5MQ2/HEfPSYw5fGRYzYHTtq8UWET2xAG6jdymJur7+pU1a5SeXq6+1YHX8J
y1lP9C9d6pWlp29EyPITd7avhlFIdoWLP2EapIlyO/QOxbD8yFa+FKPL7Ti8h2Bt
06MLL0MzyEeU8YdaUr5SsBGAKP5uLfzZ5VxEzhJ0b7gs3q4ZgH5+J7e9oDmFD1zn
cGBCRjgXJu2qxiG8fugRURrKjBU4RbIiW2O18nGefC+WZXFR9j046Dt5ynUkupqM
bAW/uh8ejlx8qVBIwBnGmDBe56jcj+Diw72/bz8hOR3A91fqZOiRCPgRznNy0WI7
rxIwyIYgdYw8JxMqCdwzlFw68GGy7eVrPXG6cTz5a5adCb0xQ4vME+QrSTC/4G7q
0nRyJ17k55YfG41zWiiG+oGD1/KP52sYmKbM0mH3zVriS/cIhVBWjyZ5nd8qmNHy
Cwy9jDkSfrNmTBhe6qEFgo60bcoOXWW0B5J6gjJajk2qogH/RwB2IMNrwrgmuqe1
BETyZZ2Qc47vLg3ywr0UuD9LbIwe8sABvvtTXEdzgkvBfNhyQzFAaNk7MoUktEuD
SwAjnI4103PlQ0Z3p8yUAGzxs/hr7xWgZw2xfzwtDjzlOwgXY8qXlc2mbnw3C6Tr
crZlfj7/jYUSaqnmxQia97thJK94my861Ichn8FRgiSZjNepy7AGXhOkipshE91F
DP2jy5TLdNMYmFgUw624wr/X587nq4utndX+pdbBlgX78Yceu34Wh8Ze12T2ZgkB
YjQfBkkgOR2T+TLL8f8SrIjfFLkeyKWQ6yFp7A1qLlmGVwT1+EbzhuXB6SEbUJub
JwYv7e/Ej5WMnetJXOwCV4uEz9FCz3cPHKpTcMh1JML+HDu+M4GB6pAluFK4Y/Wk
uTBTetSshJAv9BNeXQ38Gbjp9bO9Unpljsg+DKw1htmnSe5vv7jHqwYLf50TizPM
oK+plKBb96XTTNnjyvfAxjQnbymCia16uq6PLS2rAVqcHTfs6x7eQcG6S4WjrrO1
lKAISDGtwMYpP8iG6Wqsh8TgIO31NAOAzHjYy0w3RiXIXlQJckwkPp/kKozY3oSV
zw/Q6jbOuoEMfT0Lx+bwQ4/uPTQfyiSqTt48UXGnmliJ0Ya80SLjCNpryf05hAwq
EE/4Kdb0x+0y50wtCfS0B4AcCjujcm81u+DHfehJT8QQ+Z/spvtKKdOFUVxnJtoW
Ki3N1subBvfSWCCPcyXFCtkoWdmZU8qnvjeAF7vHwbHMtQk1DJTA1sGl6ymBmkGX
SZMJPupA0YgkXV1gcqiTogaTkXScKqTJZUdkMp5ZmO+yMr7J+f/3oqXBrl1lADMQ
xoiUvgga2mYgf7ThLOnStS3D1eTsW01TYqA2d6ML/m0Zqd+uAObc+GiVBVt7VSEF
FowYtfbB4fFiKqccZ/HSzkb0WDHA6WEdYPqKlTwAhPo2K3Wb44CicPEaWTJx4y1H
cipZLT/qb2jHY1YcmFDQxbyKfr2IJVjkhGpWbOsaqJ5EkLLA4WF3Aen8+2dqiYnT
5dDh8k4UnirMJkpu/eiVZHEEk7cW5hIFAlqryK19DwoJA2tSfjHgumSXHrE8iadr
+x3kntHhcoOG4IolQJvFyaZsVkP50le0gqIH+MLPaUgJvN5PuTbPSqYLZriJse64
x3eKt+laVcCSywwLhf4Nxe6HXNQ9eyq/dYdMPKFU/vbfezCj3KO1TnZzq/tTY4q4
dXX3IWAv34OTWXKodl04QzpWoza4LDpMbFUjkKeQIO+oZGF80WXdUY2aWwtO8tsq
JNjL3TQqM7edoE32EJ8B4PnuP4R3nSykxY7mk/HgQhidwV3oLTJ6uztQVVpQTxYE
fqIIPC+ICChuB866LwQx4J5LltWazsk9oALpJptmX8Cq6NnAwVTwO/1Gz3i7GxuW
jKQHNqMn3IM5NEOgiRAjtrXgJjugu2sujiKRXKLEaCkKH2jzOhuzHiEz/acyebSd
R0k627LV0DCLqYpCBg9dFlgjGF6t0VnS8q0DqCcqL5ZLKHQR+tKx0nJWVgCEVwQs
pLk2O0vyKdotPnJMg3KwAJyveyYDQa/JuzHMxT0g8iUjnV03BC3sioCaXFKmCuNe
pVeY/ns+tw8PvgWK8lPRkqyGs0hXssxMHzqeLnnZO0RFDIZDdkSORvKtrsttHbhi
l9whuH3p+5lkzTtROsGJIivMei/rl+HFa2PsBg/6wmYNPNT+NnqOaXhXvnMeuMXR
JEYs0CcOa4RHkww2B72zg3veC9Mf0O9bLSoRKty02hORRUrsVSXI7Wyg/hn1wAI3
MgwxKSTJvHnynTVMtzBwiaQh13tqr8oz4n/tjXDLmVrYC7V8MyFgUEaYVBNvcqPH
v2j/BE57cPzp0jB92j/OPVMxT3rOKdxyFvhNP2QMb9q7ORxRv+bzVAILYeQfnBI9
fl+8Rwzi/0ZE/yjYvUrFJuqyFnshtS1X1BOLwF4Mvq2A+53hEgWo4i3Oln4p3lua
i0VcQkfFiMQbhhm4vf7WSVHyDsd46H/535+lPo34R6nvOFtZ4td5iD9iEcmzynRo
Fx+mX1bO8QosgFuZ15NS6UGD3jdF6yWVy0Vv5ZSKbZw2dNfMz0e9ZBI5kCunI69E
3+kkoLkVOw5DYkzL2VnEJ/tK/qje4RkLwDC99JtC5ZCTWvLI+2ArO+BARWqGxqsl
Za1AIzBt7Pjt1tbF8MCXv+oDkyJIauMc1znB/I8TpUkekyENO6emMy+O0NVJ7U+f
PHE8G95Yik7beLOrwSyDW6yFYn8a5IO3MkfBKeTSg8ZRweJoAQWkU56kHO/BwaI9
OURWWJbX15PbpjDdtQXhLbeDtIS3sZMq1p+Mrtk4c5lY2Q6qP+vS/9xalmvQV3DM
zZMuHjXHfDLz9kzKW5AHkArB3cnTKfDt33oZ306c6UxaiMN8KQNpgfaknp8MXFzc
t+b3YmS3GPjC/oV9rPmdjFHbU0gtvreo37tB1CMQmAheqkeSs0n2z86oSBi43UHE
Z+DcB3mb3NOYVegawFSLGayZX/eKq9OwFsZrwVeLha2Uv74AfyS+SHFwx00ZJDma
44qkzEedplLT6gQFH1wsd+uhCS1GRW7k4wHJ9GoU6k0p+bguP6KwDGJcIX5+SOhb
AHArpRq8zb/Oa3lPATVzjPIRLKvYNeea+2QEZ4SKV7rhjWexYVSJBQ4cCIofzi7C
5weABU3kvt/8CVqqNMlhIalNj5Fq6DIuGX2ELkfQjXalQWkL/TNXrq9khIr3eRw1
VXAJJoHeUVnYa5Z643t+VLwUH7rca2K789Gu+8B4gvZnORv08emlgsovpa3xXggc
ae9kqPp2wCygDt/kKN3tbzeD9KzdcmMy2YZ4tlhRKssVZoihB9UkNVkEAuW81GnB
8ffBPPbe+Sg1WvfmMKrSt3PZ6jNEId67sUeIogJgGC49tYIEl/dpts9a2MbmV623
9aMhp0i6n9RDIF41sDpvTfO0LGil+d0JzaklyRl08VfbffegHIjJiBEpET1XOhmZ
pDQxitHdO+bHFHkwEVS0rPAs3bCdrut/WScLyjvewk3WpUpOLUT8bsawZoALRX4p
v3v15LRv1oy0audZIs8S2bkXf4h86JaraK6jbNTFqB3/7o9zdMTVewsakefprOm1
682TSKvDq+cibKXPktfxSkZZCwS7qYnD4bQ1uHou3wLlIh6sfj3DcoroFlnr2vqe
2nlGpzotNQJWhfPaQVpDCgW1MwEJGV+0GX3BoKtvi67duKZHbXo05SYqXHHChNa8
8b5RtGMxzuEAD5pe35sGDqkwegOdBRXj7mUMl8qiHC3H6R3EpOuNoEWhy9q41Fc0
SMjJJnXzZVa988Xf189V+0nWYD4EIAI2ZaBXtpz8VS2n3CiH7gZUlQI0XuXih7+t
CVmAlsarDw/8HRQ5RjHlFeRq2x02nobKHp84monzyRUb5dRIVJq3/vzHXBBkUk9U
lm6LoiBa/7UaXd7taO1rX5QBLer/qDmlTiW4kJ3Zf1MztCznk3W/i6XHiG81Foxt
s47nxdFNBhIB5zMFPUlL8wdPPCbl17xvgOh0iXdDXa2H+TB2RkNXPim4/b0plAW/
0TuMVj+uModojoZUcyJbEOwDO7CGGkL+YuJK622h+HZ68oiLu5TtK6i3CgxJId2R
y3YrJJkxQi4scCifkyb8UaFPl8XkErcp7K7SCrVXYWYSNqjCz9T9LlAyrivyoC3g
JWD6T01R3Xk0cTvWZbrQrpvc1/qvAw50VG3U/XUgLTs9+W3CEDBimYkW3Ckevh14
q9i+O0GMuKdyGwKogFN+1QWqav3CbijgzqX3vfrY65E+RPidfrA15Z0y+g1MCsUa
ygDttKr008Vdg1kz4T4gHnaxEOZE/lM5KuPxr9nzxUYnHS8BZAPOolrY8WGtK9yT
g7LAC5qWWjw8OchprvRfWuulSfLRIO310hiqd5H+5i22Q2HQiDQUlTo1rGbWnNtr
TaDcaCEo+wzcgJ9fKPbV9Bs9B2OQCFXr6CJk3az4p+slVccmpXM0WTao6lH7sTLO
eyF7Et26JXBN9sRfCwK1bFtKDBLQmX0PpdycwDLONXqPJd5APatCLmWlFZlWGe8U
hGSKH911tumS6JmWs2nlMhXiyip1p9vpun59w5aRadFqVJNF9BmnNNiJ61EEzaMl
Yf8UfiJA0xZuPnpQHx9AbZlctudx1bRr/EEsftRRrtSlCJhea148JGeWRr6UZ4j4
7ZogrgqwinpWOnG3hRBbxdR8d1vFRdTD2bLDQD3ThAE+y1HvYkrl9e/lVDXPEdwx
+jnbbfNPDYBOeuuqF8bCRLSkUmrfT86uoslIyIIyIAi3hsQJvB2tTmuM2jxaRRbO
Y9ATN5mQuLn4E67b418dGZWK7226WZkp85sV59UbQ++c9KhI9ZFJ8eof0UpJmXWi
Q8RK3/zr5Q8HAgcekQsFXk4fUBmxZHNeKGzPwPmCgWfzCDt+KWPtF7TYEqwqhatx
UEX+KkgQSkMHuPILmmZEt/eQxZTrgW1vwrp51teHGKBccAhbTJETCJTlHqnDWi5+
zBtCftIODW5nsMAt4ah3T7svHvUNWuZ2XtJ7K5COWLyDGICvvxvZnihyf+qhSMOW
ngZYcm0MljvOvF5BeAlcWdJvvgG9GW5Wmtncju5wPTsDSabM3d6k7BekpJ7+bytN
/kpwGovU6/S1+8jI8hdc4eEZLlKFoCNKzuzZwsF0n9iEciAX+4v0YnkWPW1H4W15
LBBL4080iL4GYHO3Vq4eNtOc+PiWeSKok7ZtNgh4SJ679hq87YdFCczdOGBc/WrV
X3bjnIeu7HL2ya8Er29M/XxJ4Vy15nCq0/Keii1lUtcY+AV+POt4VEGkJHhTyNUw
ziBavMJarumxaNB53a2zJxX2l6jDbOCBgYnRJDo0dLd8AUjdPd7QKrYLs1xUAV9e
or3kGOv7tXaQboXrLhl+jvsLAkwiODN/eflXioG38KUPelxs9jaC7hTnXUPvWmUb
93ETmPZzERSmiv9U7pbpWlajciIAS8sBaxGNu7/jC+VN/W4sMrgGa5EPEPvxNwi0
u8VTGMfEJerXoLkf6m1tAt9nxzNlOcmHpZN1pPqX/nTiTYNPYxcD6IOp7gnMeL7B
gwuyw0yOKv8q4TdSg+yuZ9f/Z6tpkmqFX5q0wY+6pCizmjcXlZCK1NMI211a2Rfo
0f9FW9D+g4ZUHLn6n6lWX1Ex746aNG5umpe7d2YSaRo955jNPW7OuILY43DvqDkJ
fRsjaUFk2J8G4kswJVJ1JlefGl0aD6JyHa5X3B7E2vrLrU6sqBqf1B7AQYLK2JIx
H2wvCN51qbSUpgciMlLbjUgsYhCfkYshqbFbMNvy4ja/NjBMc8517siF5kSbTxhU
RnpI208vmRZqeNWT20eHE0Hz2b11jHiHI/cBYDpGB/qIra5QO2CN6XNH8mIeP97f
UHFpa+4dZz8uKJ0UUIoQHcysUGWPVfmGpqq30cCaK80e3XJp0zbLNKqp2/cy4eMu
Wlk94BO0pRfTYJ2QiwoqagyT4z2bAu0uUDb/WjXHQGRgVbDwRCMHFQ5lVN5opqv7
eJFYFmFVdiqEekFItOX0ISR/Ua+W1uGD1tguzN3LE7BjRT0IOizhNSQdrGpWnvz2
7uzrhwqDzAKAVH2aaF9JBWCZCLKKBoqeTWz1gPqhE8UMu3+0T4XsYVgK5zF54/0r
0ylOczQuUXbbCsid8Cgddtk3Ahqmk+ZSwL5Yk4XgCA8qaVAfl4Tl4hiDthoCoH3u
yYj1r4TJ+q9wct0VVZruz8rEQ0ln9DPKGqpdLuMDSXsqM4e9YTkHDkZ1E4MNKUJS
cxHWd1frfH0u9q0Wfmctg+w3kw50CoNYzcLr0GnEhc+ewI07wLrlmwMXLkPL5zF6
YwpQymW8hBtFaW6BMpIDCjuLA/VqDskmlLJm9MMTaKOJIoDaSbB/rMM+/d4tiPlY
b8yb3PQsdp4hx3d5dNRnUxUU3Cj5yavCyM4ZRW4FipBqJDYkeCOJ68pViXB1RRgX
8ETPVjIitjptsyWd7loWcRosQRexzTvH/MA3Cf9U1AhUNXSPpZ+Hl84orEOSrhWY
qR2INeHnjQpWUElE2rZ95lCmXeeOTDcDPqIIMSw3BsLlpXkij9/lQ+hyL9k/bHNz
R6acwNOFOZd/1DLA8xc0kjJOyvreLg1xcsU1VHwfXq48M7/LaRbAtPXeVWylwEI2
OJnCyLYZ9yBXGE8I4hvyIwkEqjfM1G2abiIv4i7H/Kw0h2xBqop/N2bqbM4z2tMi
wKkktmGgKSX4M5SNaUmZLCXc6izMHE0CjWo8zpWxPrPZfMXDmoqyIGUamLnsZchQ
uggkVJcg5Bcx1sjFjqzHk8T+x+akd3p+peBBww7lCk/3K1LFtWFwrhG32FNJ3WT8
19kLpSa8s1UQ90X31luiyoSEi2AQ6opJonQK/SO2OV1tJsmNg3HNf746cE5Bjf2B
cSvwek/OmXRkW/x9ve3XFnehFwQ0fDfVoHDgIBupUanp4PaiUpqAhVuhFZY94NKr
qdQlOm5kg5XlA/5P8ydGomq0UGqsx+M7V02mXYsM81n5yhHcI2tgPYV48aYkMmoU
din5ovNysl7lTM+QLlK6nAHqhIQxI0G6X3BkVII28zCRj2Rwy4k6nYiV05YbGkqN
KZumGByH5nD511hX+S5RFfH7j6G9JUYMheZkArqTAPoWkulhOoj3W3a8U0iQDEOV
3NF5DCwwqr23focwOUqnOl2dxEX2AyKECVn7A8kPoZEK/y4L/5PHwK+bHhNzPStL
J7LRAMcvfnxmkkPMh87QDSXB2EwGdAd/rbf4t0Y8LzOjeQi+gj5Q3S50u+5UekGt
fWcdqPrveC+cW8TR/509NkpEHgBY8RkFjFREp35p4NLVujdec4xxjnfW1tWFR8mT
wLdT2MPi7kx5bOtqFZytrHP+Ey3K6I93BOdMibdtgbkRzHSUyQ3ZBWAWY9o0V6C5
A3Xf5CQLtQLTol2MaNzU5h/HsLWqbaizFer1/18AT1z2pc3bbzPjiyvu57RcmL4u
FiriOXtJHL6uzBLvlmTooxWVlbfIdZsBF6HDm6OhVJgdA5p53f4l5mwtkE8JPW6X
Tx/BKkfneQUfysWdXmNT2wpx3T5/dWUrQxLSTc+vKvsm9mo51BY3TYdRqvMMA7O+
FzKJmrf1CEk1HySuqWn+A2Kl9bwvS4ANwxCurXUS/yVkz7/iEc1QUP/J2ogcVlP8
sLwurkXSPZkLmw6T6zHgXLkLkvaAFtKeIDq1kFeiiTKTQ6xJtmSB7Qq1YNQsje4T
1GiyyRETi8eePlIO/yA/s6P2rqgl8OnMpekJrLg3eFjRyaQZsX3C0D+J0JLFsxGC
lI9ylvcXRFk/mQUB539OLGGI3BI3CDGHp1EvS+5zIpi0qALito0SVlE4LBlxMFSR
07Hr3SrCV5jdz6/XqkYkK8RAfxUBQfl8bWGgZjF7v/UUTNTbqeruiWBf2ntscQyq
DCyc6ev0irb0/5w9DkMgV9ZhP0hk8SH4fTpmj4G5BQShvG+Na4ymHth6lDIg+Q0X
FVhd2VWjDvp610p03Y+/Z7Weulvn0wXylokmA4SJvPKNngIPAqxYMVzEgMPVGnRS
UgzoQB06ONVgMXVhFUz4/kaG7Zpb3fy80amOUHCyW7OttLNjxMtDwM2w3QXBVk0i
36yEw7of93UjxXNKu+tkes1/xDEMv9Lcv8k8HxkdH36so7X2VPw/A8/DIdpL0LE2
xT8k2zwASdGTwCSjIkN372O+wdZIoCTpCv58pO7bNqM3VAx2Rr9A7GyOJRHIRTK8
RvbuNTQSHGF7j1hGXr43Cif29IBckDXSECV9W6LzHsYXHWNtfAe8c62SXKD2H9V9
GuPSP7f75nN1ll95dO+9vDzurftvwLAJVeG7jYj7NFxVZDWMVtk2/nQObkEzUgMU
65FZneP6BAoTWZXq2WZvH1vW5aIbIWG2GPeKtZWIImJ7rm6SAu+BgScc8RyUFGNR
qR1CohWl/1ikZWWymKuhBRUS7tDPV9K8RSupJ3otbIg2DV2RhBIJSmMCCrDk5dc7
UrqmTuZx4sdsF2kbq8cuBHWMImLrJoPRtJ9u4x1RN7ff4LzDRtGnxIXQlO5FVghp
F+IjV8fYZ37nMJrkVGKLAncvQ31hIOrNnuXjOBYDOItagzkuCJZGPt0rgyXihYxu
jgSO/vmm4KevOb7kjwmjuua7kk7CVS5XWoOckViY4Q1CtBxEMVK0KL6nIjuom+4b
nBdN8q/6i8x/yW5593cTwlIqsQBAgmKvh0QxehWOgtl1DtyUCcC9x2+eScGIpe6W
1A5kAWj5W2c1J3OQ48UcoZpS5DG6OvPGB0fXG+IIG/NzgURg+j3xtkuQ1NmMzlc8
OCUJTe47kp5aNGxyDD6loHvlhL0tXvk19nAnSC+JU3jC/t5e1iSFM0/bzAQiuyyS
OSlxFYsFUwlSbkTlpYDXMuzW3HZlvFrVOZM45uOpxunm2xIlaHjU3hloYKTWp8w/
SJysRKKKmPJU/p4QqnS74sagGYjULumfWkCRWVUbVxOScHTvxQXJUpNkGWzZlemo
mJ10p/OXP3/dOiAKxKzaXRPyB08n2v5UcWoj0EyUDq9dRe+zgukUbWWHV7OSP3/x
w3W923F9VaJZg162tgawgo2fPJCcR2OL47pS3oUFfCL3EhN0uiJk1Qq/ita67i8n
szWth0+viKukqpW8OOhu2pSyScM33ISBzhWHsEoeCZ04sCv0g9mwyikFS99vqVYn
jqFk/jGYdUnJKH/pINMwdUoK/ByuuOvl+FofQBnq600qIKRlzxsFA4uq5QrtkfDC
9LCVWGJmbWp4GCEDcAg43ktbi9CCgb0KrO2iApcxWJ7kS6InuKCMMPWihTCS07zu
GVBkMIdPBukmZaROOJdUSdAv1tlAFXTp1+hntPv8FA/nX5RGWXGVqnj2DL8v9DSp
v6K9pBRwDXotmvZvUu9znx+BMxh1EncqBKOY/UnmuFLJ1hTC9lTQXLdsqgsKSLvQ
bhdTi9nz0+huAgQFd0P4gmPy75Zqc5nnmXp/2f9UjPJmFLAVBy8Wa06GKWbQDzdT
jGq63uJJNJYPXSTNxc0GOONto1Iem1J5X9HbZEYnZYUWTor355twsQf64IjAKpjx
1ISBXsnqJn207ySjaknapR00j4nGRJm40/um4HQAFMsw2AJnSUvfDSrniTBEd7uM
ttoIUpyL9AOoUMBE0dXdtUr9diuz8NG1RPoJ5uIioMraockThcF1ZV+JU0pmHVJw
Ttm44IIghCkNtF3O4kKCntnOnz0XDPfGDEP+93q2RXZWMjKcixuKe1mOXRCfFOFf
UCylrlKut+jRrXrRruZCuydG08uhCVCLuruMPiXnEI6I2mYDR2N26HV8Jq69aDAl
fe5qXExX72KwnPvrRbdfU6Hx16/2HCh087yidgClNl7ua4zD/miZEsvazWVfEaP4
pSO8oVtmP9dV3g/9+AltDBl2nQYeabTdkX8R3bspui6DTLjyXk767Du+6htjx4RZ
zT1q+s/S5Yyck+Ho4t/HQmFZ7SvQxHB/wqF3xh/RBvlgVTWoQVr1TQ9m+4/JI67a
TfkXXYX+KuvhjkAHX2Yzz1Bi/2gw5I/Q5EbQgSKKRq7xNjN4R26RM/R1w9QEZCGE
tuxfeo60/dHvNpDfCwZ2Ob+9xQmilfjWnnx83I0qdohim5wVejXgI0Ejz6aK5WoD
btMCqJz8/S3LoMDnzv3nzQbkta/lRaHxqexOomwt/3spsblnLzyJMy7rEUMhOplj
Sv7/6nowaGsnSdsIENN20QFdb3e+K2FPib9giwixhLSo/ZznUSLednj8tTMBXP2e
+L1Pp3U+Zp8zB7y0ChQs0YLdLooLBJ+QUW4giXTGjHBzvKOpMNl4bNtGoICDVy+f
1MLgGw2eKVtPtghUpDgRWKl5vd3ih6NwBtsphLe5YNvldYDJyIBm80/22rf0xy81
vM4h0k9JHK/CaPLyfZNexyTpkXk9mGFHubqC+sJhTJ2k2sjgHsRqDnm0k5NHzwv6
BGKa7LrvS/gV83ZaBJ4IzBa3Rtwt6ZJjpP8XnimfDrVmZOYACMxWEaGoc1m08dHi
3KmSHkXK3W8XCtrpbdDx8LivrCN11Yrav3YVUX76qTKxWjv55w0+R7W6oTxSdvD/
Uk1I5blyXUSnz8ksDZ3/yXhPhfHfgVeQ/IgyRMy8YFB6e3sQR17dofeOXTt8csFD
CSN3U0jUAjok63qveRSd3dYXDvJPtVDeS3O7Eh1i/SOZs3/zgxtyM1W2+OICkgHq
NBzFnZyO4zmgKL0xRiVV6d4hJp0JEXjfbNT7BmNsM6zKCgOe4FqsnDgPb6DGs8nM
T2Dz71NcHmN3DjaXkSsslTlDc1l5E2Xi8XYxvWhlko7fnHeGpBkyB+rOeTPRsgKn
+/wLj3ZRka6PpDkizUJWZuIJNZTE7wg9dw4nHuLvKkJsTySVxpIPMqBIRyUwpFuU
OcgIwFX/z1Uq45VHx/YBQuAqxGn/+6ujBlsuvIpNzBjHcN/qTF6fpsHFOmh3F74u
nu27v/eWMooFk4sTuDcZmj/bk9hwq+bAzbV0OXmu37/OQ3RMmMHXhMDURNzjZpPz
woQDqXRrzUG2qvb+Q2lGGZVLYz3s/Y/nqZY5r0lLyeTNgruDaXXD/yWv1Ny7Bd3d
z855bIo6Sw+i7hi3XvrFPW3I0tEdb82dqQc0cr1U9gNMsiYkU93qq6k3FzZxJZt+
7baD/sOO7DMJj4goKAfgpR6Ul9VyuhpT3P1orzz9p04Yc4qUPhY4yNqxuGCzHkgG
V4scGefge+V2iuPYVAogAOQaYZLoePMm5yGTB8c40Q8HrgAQJ/F1ozX4xPhIbKyG
zwQ+xcnx6U8jidhhkPPOzH6s3zd7b4RSmD+VU2d+en7ANEfMHEfbAZj5TowxJx/A
zEEWaGxM/Gz6Ne/SAl6D13iarIwkP76NW9uKyef86tgY+25xOGXcVgAsR2PStI/o
2lvpPYTlm8NmoK/HZ9e1TCrUIPXWxn6Zi696HgqM9/OQenOg4f3jWP2UrvBO21Jt
zsCPWxpG18v8cBRWTslcsvhRBRIPFeN13wOwq3Z8X4/vCzU3qqyoE22gPsDwvCVP
6zTGs6qcfMXnweqKfqvqQFai6bh2igSiOarkji4hg+jKEp5IotymEBMmWTuUlas8
B7DaL87fNmRZw8zcM7GO1IN+PTfSfYUEcUJU77nAaCFcYed0/xwKdghqFqFsCCb1
eDcC30cXGLcgJSs2k4ZT1VPKlioKK/r65NR8YIj8BuHwSq0KawvQmc/tuV/hWtUt
4qn5juraIfRnFcD4Rd0wSpJQCg7FF5Rwyyvtr+lda2Zb5Q13tZNCm54FOg/i6Snr
iNox8eL3dEVcx2pOzLBTJRYsm3OnH8UAc2SowxbHGENE6bjU2SwQfFX4NmeH0yr6
cs5c2o/SWTd0DFgAAWO9I7WFxlEJdPAwU2PL5vCP2yv/K9x/FtQt3FW9Asz/vFPO
nSvteNP5L4uVYQvR9CgrpRb0pvvYoRGV0L6n2BFfARWjbOZyGcLHlzaAF1okMatV
c8kKGc76gDg42xl2K2L0P26kxAkCbfSVxC2N687OZ1MN2pWB8Tlt1377ChMAdktj
9jcVap3dRFvxsTkrVLYWFuV7q8each9bz3Agluz1DxZ4ijkg7I2l0tm0fNk+XfK8
w4Msj/0WUs11oNHpMtYqYmNKr6yCy40VnxLrNTLmFxfjeYiiCjrLjnfcuYsTAHVa
JMyrWqUk3VekfPrMsDHyUfQayelqU/nWyCfKLDh9DcantkQt8rQVTrtPmvioImNs
pbHb3prLcc34wcSd0mYjEMGlysw2za55kQhNnGOb+/xknE2IS+WJna4oi+U0k2E9
LmEVAG6uNz1gN3Cc8fGNqIzhPv6ZatWUtJjumgd3jfWch7xQhtPGh3o3u8Cwzw6e
fFXnvW6ZTAspd9b9QP3ukJZNwK0F0YdXvH9RGokOkUjeZqEYm9kQ0RvxWYPnDkHS
SCIsCb+BQ5pIunh9PLHQZNdzaaxaQZsRXaL7XuBD5a69y7IKvAczFEQ6RVmaqAcu
hvNvqiRzUWdND2tzJ9v0uBDrL32RdxsXCVGzXQLgjBAOHrJjs2lpxrAdBTfglP70
H+lnARN+TgJvXfSKHgAfzlM5DhnCCVuec125hujNVDm3dUle9ONyq0euvgWcWQbz
6VTulpI5Z2CaI76BV5nSc27/j1q2LTtmwegF2b8yj3qL6bSQDX2aN+RzsBrM//6q
tOmh1Qtpj1r8WbKIxJWvIKyGk2Tf39ojhVLTZYXOyZBkvYpUF8PAcMhMtm0fBdoS
tQA4UBj+WFQlhJXcqh8P6/Afukil8zpypdqcQ+XmmMr8FvuZFHkGXliA5u3snowT
qOfU8P8VP14KzzngoJC9/py8zqwV6DI1ECdOk5U6m69he74Xr8p0ABEQYRj7h0/N
3JK9jiKuRw7QWbcPC266vCjHVus33NYz3xEhvVdRmIKi4ATwOZCC1+BTvkK2JDeY
akkO3IhjLAQ1q1jax3k4GRRsg27rbOHHC14g9oAfXn59dBRVpj5bNa/oXiBRuEvw
R0YEAKQFYhaegNSZ74b2sdQHdUvbnGN7hDw7A4LcAmCHQxIeq5JaSiNjTKQ0q44e
qnRJU3qaTBoh31u+SoHI+cfM6nQ9y5XzkizF0Rei4lqheGd0Yj3KC+nGebO/xTeD
IHH0/Ab+Nlf3vAMgipyY+VAAWrAHJqbl938Qkwn5x4mRaPg9/OgCubPRxDUczNya
Pciuk4wVfQO1wpW0CR/WihZO10XxibgRkI2t1vGTh/7BF+V7s2PBzV0UhkI5oNwn
AMeBWpruaJXFRKt5hmn1+128aVJic2x2R3LLzyDrDvwpFBST9GeuuiwDa3YDo0Q2
tMQm33TRcCr3DPl5q1Ox8MRWlN+1RzlmtnTeqxNOsiPv8r4wwpk0ZTrZjOtnGfft
U5X5+gxgsB2YATmaqWz2iDhi/LTDb2tPQounula3lvMEAgSFjGIIOKpnoErtWy9u
2fG4hwQvAJOixl2AuFzQGxt3ndNTfJwQGmme+DI/F309QaX20XTXGSJX48EWD/XY
0hCt81Wewq9FS02X6FTJQKCYuwMxSENa4+61jPA16TnYhLYhVaoJngryMqprlBkU
9zNhT3cI1BKY3bQFiz+U400Ao/3T5x0QkJFVrZ8Je3UrLF/VT4ugvQZcOTxZ5FtE
nbJXJG3exh7/wX5JmIJxXv09Dqoxqujyz7foa5uBet/Gp4397qlbh4nTrzdSw1ll
gPC8DoczGB/eEXtdv9zMVyfbfSoyxrkizEY+d5ezEqX5p8tLMK50qwDDHb2lrgmg
+b+Ggd6rgViEMzC2x1thdf/TindlFFwRxuREuEGcX35+GRsItqCAI/vh/ZSHOVNJ
9rM1IFL+pIyKQIx7iHxVEgErbNx7MgYQFV0xvGCVioq6De6SZ9an1LGfMcUNC0l+
xQ3lXV/ZkNpqM1rXzIrD63eV/p3naSjCyb4+M2XCWv/woINwuggafM1Kikvus/M9
ahPUmJ5BFgexLmzV1sUjQBfsIPDcMeJYKLA/RznkxPtYmXtBUDTzJThnlt5fijje
fOzzQ6SmYKfQze0LD3FenK9i9hODuxIlX0OOKvalOsbVuypP6khzraEftkjuvgxf
loPFnB7lylXmFl9ZTiqWGKgkyf0gsatSHy7frSr/nAjQeWPhX4IgSnPYXwJ9Umqa
4rpdPJDJsX42GQ15TF0MRva66RtO65/QNfKQPSdjffLK5E+ljruWR/OjLvo1TJLP
tycsWB3NOz9a9oRYba6glEtFXHw3/n4qAeheJ+2VB0pHEVEMahz3+b2kmqSOjfkZ
aCocThc1osiN528AM/IDm34qLaNuL01yglqVR9GsUADoVETG1qrqPCxIWCumTqWu
GuAF/Y66keMak5EoPcUu7G40lGSj+onYNvFjNPeHVxDKQF+l0usfbj6Ce7B+5inr
itvpvjYsYH6IUrASMH4VfopIelm/4eAxtVyLEKeUkIYhmKZD/liRUGFIjV7Xlpv8
hUZQIKIWL0wfxIgPhO6obIt2/Op2prBJSwDKXqOPhZWt+1qdbt3Sm4J5nhIaDskK
CDvzDsGI61eDClQByEitdBVSI8LrVTVQh+zL8s2wD6Qgcin8hxRhnLzHFmvnEAA4
Fcz/BRf1mHIc6jsxSoNqbAr8W9YcXqZx2dZFPkPBYtPG9wtP2uktLpM/K0ncNrRC
0cek9fnlt/lhInpUB/ZpPPx7PXX8maESUy0V3RXaLN9Sfjz8APhycydmpYiTRgHX
l8b+jN6o8W1rJAqXvPLxmRK4wG1x3PSxLkcQAKgthtxZdCN/Kp7wwPR6s3W4ibMh
8+thlj6sVkzl+L3/AtrtT80We7FYqdooBaF2HlnOzakr8aOkoW+MwEXYFrH17dJW
EQGGLxFSlIzAZZK/pSluf4od4D/bK8CvaeLTjCaNayVE5dh7dpd2j8RYBgu8nuc6
bmiu13CjlomxBTAGWb/RPDyR9YQURIDTWu6XVzLx6YolgxzKalcKMvfp2z/7hivQ
VDwAaPISYGawHY/imCLFkuyWmuU1kiKogZt+E6Lmh2bJLGVZ8e6obHEMRB4+UkJy
B6/Zk5cAcn1rV8c98IcHtF0FZC5guVUGxtOEiTFa7SqAiqtCir19IDA33Oz5n5nw
XG7Vc4kYVJ77O8MRtPwK9bSlbAY0Mt+RAW4prG9Nc6qFS2KOpk6hdY4Mxdu34JbI
7AQK/8uKHNIQyI6I2AiUTDt647fiSUUikWNC/1K4VNxX4kW7nh4b0TaW8JyXjd89
u0HfrGFoJgyQtXZLbQdYWPNy866L+wNugvWvniOoHN7dhlXbE6DP2XAvVkB5lE2I
7GETZiH3ZsOwVCcz/DXXOdgQDUAmyQvhDbnIv7x+s7mWV9FvNDEfmKPAoFZHvCz9
2cS3+m0Hv6sfphS6nS8Ffb00umLjgH2gqmFwc9YmVwozkOF97OjNvqDMVWD1fSUR
5z8eqR8Da6nz2FsoRZPicnliEcjGO6HgskEdHhTJy8BbrqS4+r94tBbX+ChkzHOs
1WJrHulvD8pXKPfG91JNfWpoWOUarl/7ZK/O4qOIeTXZI7u9cvhddQtyOIweire5
T9sggTC5lHkIPboCCeQowHmdwSLcOYKdJnbJfpDWcnSvu+5dmiV+m4krbtTdQ6FN
drTqsySHF8flvTVy9TB91H/WThO5Sh/6a+znKnE25s5E+BsDypDSXPcqNFoKgZxL
Q/I2/Y743+DQlAGQyeanDYzFKSOPcXXhjRFJMdub1jlg1RVW06bTRsa3EpdM1Au+
o8d9w1FMS+kaNzg2jJHsKTIqrmiRZ7IwWz9qGQ0YcPSA9wbx6qX9Vu8Joi7eMx08
M56Dlf31509s/9+/9q2wvLVaNbY2b2Bv5Zv6zuZ/6maFyUHi7QOKDPay8vV+3Mar
xod78YElps9Lku+vOG2i6xpoErSIBTtzVMM4TDHFHeaUVHRQDk2j/vxkbGICzH5w
wZFCNu68yvizyc9wFhFKyvn5CkMGnG929mAsoxLZno+sa29HyXuZdEjRXV5znKWa
Agfvh6QX4nQH81L2G+ryFgbZ8O0wJUj4Dq97o7AiLAKA9e/iCU4x1FPnxaWl+H1i
gSUJ856aWghC0QLT3BLFUGbbfe/bQLc4dpK0CFQxkbwgJCIL5IgxeOndoY2UtNyN
fofbnAmVUMnKBGShrKd8rfNt80KZWjzAvCJj7rIRFPRlYbW8M31JLJ3DsX9dTkro
cQFx+hCYsiwqXPl3jWK3CwM9cBUVbzlfdW0O9AgVIJnDa2mgY2lfiXOE2UyD4rDm
0sG0HJb5xpQ4fCTMGNRtUXEir64E5XL+cX62bt+hGT1y4VPjDLbjY5IJHAGyDakB
EzVBnrQdcqmwJ91vbN7gahE6qz3N9qmwJ5E1eNzVJgp+HvFRh04TbF+nZXU7WigN
eEk/Ig8GpSF4IPVLBjcPAAvFwxpGxcLcmjnmjfxyCu4ML5sE1K1Kuv4EbiP/8nk3
cpHhF3q+dmHADYnboeDSvHdFfpiHCzE4rML3Cic1/qHRga8HSAVr5RqN+kI/0G1e
xYY+4P7K88OSiqdYlLcg13tJWLkJCQYGeD06+khjFj9Z51ZqO6gTA3cI87F+LSiX
tMaizbXo9g/ZwEiiE3B+5/QA/OP23IwgfSNU1c0Nqf/18J3HZijwZLG+DQ/+3OPg
LnBTC0Rxg2b13YgFzvtaE5axllr/TJmSjRcDu4IgyFaU612ihJn25sM8bxQO3Wri
ASIIoVgjOx0ZaXqk0u+oYh19Fbuxy9LVUx+lsfHh1miXurdjoJC4/ztCgdT5IUkX
eQrhdXHOG2Dea6YkpsYw0YrtYrR/iapGTNftKY94F2mFwwGB2PCjaLaJ3rpH/P41
ThNbqaK2/RygXG/zPOadRt1C+Fadwo9x6S3CEstAvGcR+xgFIVHqoRMTR0mcvLAu
oH2aFy8ZkairesEowZ6XFw3Yq5hTYhetzICVg4C2an+1zklRmstlR0NKDQGP4/n1
L0rYlbMjgGoRN1mG4IpQ3tQjmyqeRs/oeAZiUh9yCGZufIlwA79MZ4gH3PXxR2aJ
THd/Nyp+H45jdMmPhZ5nEuUSe5qVhtB7R3CC1ozReP7X1AeHYZp4z3WPwoT37FKJ
nTLrSpqrH1vWRo2PUkvvFTukjuIJkMZvQWToDMFaPzkrNXDVe693ZvJCSIa1ZzmS
J6GbOj1iAoAosZY6kKoKnM6uFnemNbTHA73Wb7F8zcsljJjF6vE5nw49AMLnVQ+N
bTzIx8dJdBJ5QCpmoe365eSrP7eDvw0pk02pmi/1iu6jVEp0oJg6kQrM56GnwSMS
+fO5/kzw8BhE+iCEPSIluK4t8RI1q4HGNKkvGB+kE6jB7MO7OeVOeS7wPSx6oApi
TGGwRdB9FEGVrx9FsK5t+0cPxyJOZzcU3qmz2eUWeFOLIgXC1AIb6UocdPwSC7Px
G5pXcV6fdfHY6TfCtlZ1700w+z3WhXlLH9rmmLVq4b1V0qBuTxtv2+NgyBEphCjS
Ntt2wHB3kG8aftVh26+r7l1MuDpD1DKDM7GK3MsljU9R4LUgXTJJ+InfXE5PpX5I
cDVp1hl6hnEASMuVXB7JCqKK/ZIVYLmBv+UlPCTbGVXGMzoO84EKNP9GBKjUDN0Y
us7JSvnN7ag9Y33GbbmwxTlv6MRgZsvsDxpZ7gEToXIbV6aTr4yj6mMrSsl5e7WA
5C93JRb75hR49WLF64IDxiffdKHBfU32wwaBfcnMCPzPgJPPOigHL4k93k+i1YNO
VomSI58u4jQtuv8lHhteJP79lSsF/0lIG7cqh4uPtUw4zsg6yDCLlYhoQNLfxOQg
ozqBFj7BFYKZ2DNQ9OVKLWpHMjMxKvxCDZTX0rDtI2Oq5euJRTm+roUT/90pew1G
nSGcWHAszoeLFQ0UPX7cFcd9s73xY2dfhW45AqI9NkMhI+d8UR9ISW0+mdEgCFlA
PstLBiOV57AwX1PbEKdr6J9bijDL8otz9EqCq9KNP9Jga/CPU4pzufk8ap5xbLbQ
F2G07AnRTsv2oNimfGJckPOJBb6j7fP/NFjJGo4jMGOA8QujB4Gxzvq8rJIlQHe0
tWd9dYmlQZGRnxHkVZf6LTodg17RL5I+cUoVSLTmcVznA0uoZ45HU+sMZN7e0Hnd
Kz2S0zkYl1CTk7mupiSRjBEK7N9DifoeecaPYfuUxp2cfv1tLOJ+YIkOCVA4i5jD
8xhM+4JL4gjQv9Cls1+a0KyCN8F/KF2/gihIzAN6KMzqPX5Dq58zEs6DaAXyfaJw
QXnV8QIOO0AGOYfaRmGpo/ufiQ7GW86VZHrKKXJdAxImj2SWHuEm0+DQDOdko/BN
q5WesvTK63Hbrh8WX2WHGY+ZxkajiEUHMkmptFmhWQ48ZVLkZYzcG/tgzVMyzpVB
wkUTzPERBw5xtciBjpugHNaGCKiRj+9JCMfbmgsHkZzX2aRrqb7YNH3WL3m6TOAI
wLQ6HLAXD9emOVfb7DUmxtzDWjdT3saegnYvZblkEd0ne1JJUSkVgN3HvcIWZ9RO
mGB0E2qAeW1MQAdPq7gd6h/hgZzRzFuqIDq8rkr5f3J2bLOjXWHpN6/l7odCYL3j
qUCutjq5EHf03GddnJaDcNNl+0tqkZPmew3ru2PdDgFCwaOXE74gR8CmW6qLCUmH
ya+OttPtIZ2mdHHmvv8xZwUVceWvknp+DL7oNI8A+qdYSbmpf3kDCXMZsh77jkkS
zrNirEFbk8ZFW+v1T9g9fCOFeXZhGS8+lxO9SXKc5Z+ZeK4azlezfV975K1qY3Ip
8xXWu0+CIBeluupsfNVzkiiixDXb1FEfMaebWTSkO2moPWvyDwMvkNydD9fPgRLJ
evaWEeVxUZpOtzxSDtSEqwsj2cX/LYTaJvSyCLumroCITEDED1Ijb8tBDS+7mSEe
kU58MMuBooQn/IQm4bMEq7XTRz0wRSGkvN3+rUaXR/QSlw5HA8hb1qvvV0vvzMiL
LU816M6ZT5tSfWkdMST3AK5zjVp6V1nRbVEbvNWjsr4fOWILCTbGHXWU1y0EFQ/H
J9LspEx/9KO31Zw19V1cZeM1MNehK7zfqXFTocNCUKGZ9RhEBK28rI9ze7Y0a+hG
ZRQAILm1+csSR42PP/vQhPcDLb5cVo/CxE8j8jJ3r03epm4DQRWPpn2QUihj927x
2eCf5dZRVuG0yUn+ngyYT8Y35NEgzBHyqbDAkBSJOEIcWsu0pt7EUHjQOt83Dj38
deqqz8sOcI/Zs2BSWYgxOu2quyK/IQWzh5zzEezsNMi0dVqLTzmrGPczOVNDfm3Y
88+BsV1Yu/ahtoS0jVOQEcQ7CBOM8RnirnzCIsz3aQYhLGXcS35ArOpT982hMnXH
+aONH+uLvAR+UExzwQOvMJ/G23c0UhsvFGMFk9mysJVZom2HoJBTyvoJ2dvZt/x4
h4p1cHIQ9Tv6C7HHiXBtJaAiXKsTr088taa7kG/OPWUZzc01zfLNtX1orw0B46sX
r0QGK8Rw8JaUZ7f9McVeL3AKDhDc8yrup5Eetso15TousxCNT9r+pYRbDAy90mO7
7C/ZsRmoH4hqQak2Hab4V3Mvbj8pi+N9l7Prlz7yHYXotvRP2hIOWk9TAZmyQAct
eEYs4DhR7clFJ/h4ZJhvWXAVmVkSO8hEyDSkLhRybeCosSTkLdt/wo/GtIawqbqS
umMXxSyIhmwkB2bfMROQPGsbEEMjtxxOypl3qzzlUU3IoIRi0yO8+APHRi4rkbbl
ASWtSHsZACozh5O/Yy/ONy9kCbOoiv54hdQfFpPMO+bQzP9RsONo9tzOcsjIKBPP
ttrc2+BGLLlFkc3qpn71BReEO/quD6nEiyQnZXeXmVYV2v4w/rqaA4ZRWBKZ4/Ij
kQmMGNcn/Kb9z7F4vEjh3EGoQYFIym0764g0EpqHjafQAH7SEA8bmBpJA7UCv+jO
SjBgRA1X+AdrbogsucW8lSSI5nN51LGsMmwdqonnB8Hv69O5o9hzgwPPzMJnptlx
BJBbknGUbLRLJvZGet1Y9irpVkt6bSCTnmku6JNo/Md9VdRnDsQG2LUk/EyIZnWm
7FR5LR2mpPsEP33SUycB1+plsPui7Mhe2gwx05VeQ5j5U9bnz67Y3Q0YL2oGTi4e
ptsI69Mtwpv7msmG97kZizHWV05z2JFji+XJAw0L6VFyk9Wr+iZFxe22kHxNrHEw
qa8fC79Qdh2a2FCrDftS4AYssaBKbChaQ1vn/D709zUeOIWNt9MCA2B9RYKD6y0d
WXgziAC9OU9oIHwbR/ms1UDHvXXbWrbsPVVuL+USn2RUg2923aqiulbvlqhChsHo
cX1Urt7LEIQbdNvLfygxS1P8fOBA6oC4Uy2ZRvJXRsSL+JZGa17dYx07fhPliD77
T4HaX9cBIszO+suKX3FvR/KdXEXPoGB2yoGNfRhSo3Mm4h1N6Nqhr+Lyq9dDkUGk
y/Rj9VxxMPHsJcA2jtnZmig7T0ob5nhIak7Yl96KgUx/ZDzL/7br7IlXHjsqF8eW
uhJ06nVgFm9xEF6XEh2+vuTGHf89YyvRGFaMgyBnY2ghbw+SgIaEp9Ib/5VrsZmd
kiDWNfxC48t2WZ62gC3gAjhBxLi1fhJjtiUwXbhjTVUUmxshYwofNJV0bAFqxl5c
OCtcK0K05u8jGdUbp8Cmu0Ad8qYY21FiFoYTlIkfI8RZKMM7AMzTzbvIXnwsxmwH
LypT8KNLdMsVKiv8xJvjNwJvm7yYNVENCZIsyyRrcxiRC37VIcV0TgOtu4GI/hhm
uL/MjGuUVrG3ykPDwakOqR/A8zewIm58O0NZ1Mf0MIPKZ/akY9xqWyLq2oD2haJl
JEx6BUi6efx4mubjkoZf04QkaezyEjOTXDGItMRE8F5dCVV3wGeCfJA6ZYplLnLS
rUUB+Q43YwS7FJVkvvOFwBzi03CH+rDyJU8S4RSX3t4/lgJ2tuqUk2eT1qQzNuvs
ieTRDHxFVOqaWPxBWkJ0PBlKKlmbXLBQwkZsbTTZgSn0tTCkxpd/iasqLkqBpnET
Pp0L4CLiGWPByig74EWzsA7lqqGg395qH3Bk4VWDHYY8IyJXTHA3u6YuS4524AOP
WVgWbsLHT91FGQHpk+lyMA/Pl/uigGz/4Ro2De9DUzQssWVqp6nj2KlGjCOP36mR
mWNKNzY+Lj9OmjBLkrfXFH6m3YO1Uetk1HxHm5j5KXndhQK5lR3uHkdWDUHxOepr
c6IqessXSC5QiAW0vg2VErwsafABgTHQ+kjAZWgSs/dmr0J7JRm08FKoY9/TZKpq
rsA04qVieCfTg1q17PKmWfzIsYJsIKxv5VvO8+uu3OQO8NX7ngKkn/HAvlOOJCLs
5TMKMaGMpq/ZjhfmP6JigZY/aNfKQPZalO6e3536KuAeVv++EvPGMYo+w/MEjxyN
1w7p1h9ovI9e0klLm5B+PLSegbTKaHiHI2cWpOEH6w2fDIKCQJ0adQLX7av2pYcc
S6yGys5g2HmF4d3/vWP/+MQjB6HO9iIxMERkyNhu7ELWfG7DgZFUJHERtk6ftpAR
KHGKo16N0sLPTNi7oJ5c5EYuvvCuVsNOIWdlickRyf1HzU1w5clk4gPKkmbt2CxY
a6W9uqPg19zlENJej960Tz+8Z9RhqIY9PjsJcRnNCZISfDGbt/IXlhtRPzyd531r
bB03RygnknM0BBZ/6hitNhhy1bZwR64IJw6/f2Vhtb5Ppu8+zbVzSJ0FKLi1CoKx
f+r/M+DqLktIGJUD08mZYsl+IEMcrrf23/dTJwoJtGpNLpXP06fDRlyHvAGKaBPJ
RqavRLP1nhwAz8A0rOOqNDcJr9O5f87KX30IIWnQeZsVDiNX/GkUD+4uXYB7dcx4
CPqhxYiYJF+I96isea46jGpJmj5/wC6QcBAQH34MYyvAOolNYVtFTjPg+Fx3HfGL
o9+j3QGmMRsLZzi1klD3Xf8S2cuZpqmSohDWVy645UGFMOpDWeDxq0/rsbPqkJrc
tSmcBQMk/+3tcRWZYEnJ5sWDm0g5NhOLMN0Z4l2BLckrdvEulzyFHHCQ5xIooPwr
+xWxoBK7sGRj825iUuSf6OsKhAJz1+easirM6pjyas7PmRiyTvurDafd1EnkT4VJ
9dHIo5GIN15a2rqHohtRctxGzUjoQ7rbHU1NxvIbG0kJ8lXZUVkjuJbAxN06X3Hf
oYWqXkLYmFPBX1gzk2DGRLvWdyuBIcbfrjO7kqEIo6Ma0ckWUcCRX+L+s34NbNoc
cODSmKEYvd2EGY9zToi16jfwnrcy5OaAKbB3f4TBpFbqc07jHUiMoFB4Bz0B8RQB
VKiDbgvEgnbpFFKYDT8Ovkot0UxQk0dsp/UkQ7swKXReoTwgibR9c/PQjZzseow/
j6H2MQdyhC3AmE4boWYuBdhvl+6ZX/htVrbM4G04sCyKCyCX1/xxmDO/KNZJ7cgQ
qRHQdjxf42mSoDqjev8bMSFHlF8aKbRCYEB9Bj7W6SNHo+lT3Adc3dSyEEMFqpGe
OhxPgcS2o+gVhrdaS2z4J6GRT2ia75eC94k/Ay8D20LvhAEG/ga2VWbMli+4Wb2M
UOZSOqjJ6sQoiGUJ4yCBVznTaX8tSGofSTpxIZN1i5dLE20nxIZTh8jmINlec/Ir
+q7/AhCHs2N1aG7vksfvSFxts5g9Fg8dQXz93pNwKwzvykMTcJpKomi1q2vGce+P
cdznaW+OdSY7vBj7aYHgXmSrHvxLGRvosGP8ScSiEz48j9UIaM5NlDSNTHMOoIaL
We2XgCM6fyO2TSIAEAvC2FoNL/uUy38tA/s79h6Q7MY5eVq36bpOX91T009Ioy0U
Pcdawb9TGvwXU2UdlvysSNH+R0UApcEBy0Gb5bW7FM9PeNEbmVeDJs5spKkmbkwv
OakN7IwFBF9ktANDQ56ySnt7+1ZUBhkbI2Hb350a+CFBOQxe+HSftiabL/BUdtNq
fvQiDCdXr81257BbKNC1hdrSjM3MqKLhDZOcjH5ZMqplnOKBHEYWh4BrlHdpDL5i
iNxLbOrAk9NjtXIi4mVLZwmWmACe+/QvIC+i1r28KXmTExYZWX+lsJTROj5tEy4h
M7cn1MmNsz1XuMlqX80WRtActVL+U93nSShc2+/rVsrYPZG0ylBFIoygvmBMToFD
C+Fk1pcB7BTulYoG+jxrM9LlN8cbJxNuEf6jGQ9DeGAi2LyoQQ0KcAbswyAwtnZX
mPP7jP7W3ugDeiTl4av1GVG46d0ANGJz0HGRX97kf7hMZxbOFQYHNpkT6zsFnoC6
y9AlEw1BHHWVd9pxY1BgR16q5ahwjidjCQ2TzOu8BrCCEPYWAgi/C7TvqdJAn45I
olu2s6qR8y4l6+9ZQrKMmYLqPpmqSsfHp79j2JViQPTc7eMn1tK+c9jjLVAPwF7K
+HIwl/4uXpuMdl/WbZRO2ETQoV0Ba0ltXZQuk2rFpWWSzJn8d1EDGS13aqjMhnD6
xjIkWjvfehuC5ymDYd8i0fDP5RjBeIFnB+op0oiYZJxU8ItLrtawFCqu0TApmz7a
u7ryib8J0YSnmdlTEjhqOtB+JVRJaC9ikge8uwGXWIA+8yJ7jE+iICQIDbuXMoj5
Lc/ZWMaRWqD81312zy3HfaZjJI7C2UJEyJIkE021eg91/bHHicr4nXKxU614Ijw1
5Kzndp0qGCagFZfcna+YC6cJUrEt5+fiqdev/jzbojumtsRCkEmu/2eKe30AEivR
7x8pvvD9f6QOfVPjP+VheDAJN1P0uy10RvkIE9tTKKBEEJC5UTuxaazAYx6uy/7s
FullxG+2+lHcPhWEPgVCBxpALqqlNlC5jJNmJL/PY/tL3keZ9DavxN85p0LdITFv
OtbohasIb1hbveTdyxVQU4pZX3tDge6A+ltYoRE19+4qZ/5j0bE2wOcUB4boLUZC
oBJLxR8sHWrzwTuBoP4gW16MOIsftHg5XnYAnrSWExxgH7hxKNPOsBNLRurnkupL
fd5CEuOHxNRKmtWW/7EpBeoejGuVNQNKvXIvSe2zqcFUR1FHdk95byMlgfnxqBF1
M4DdRwl7bqcmBHbmOb2EDOHTJJMWsnddPzbxD1Y6B+CAbmKdUuwR6H4VBsocm19V
Lkx0tzVnbeajHIghGemjQ9dAkFhXhbkeVqfOwvBm/X+5PvHMlg8dfJxAvH88uKMu
xyeROq3W970GkTpHxdAL/r4kO05/58YUf4rCGAC4gEAhXvNJP1shZZ0EKTyGL2iD
Wrs3ECcY4TQkFMsVoXm0MPVDvVtyyV+yzwzT9CcsOs5HUJWG/e9TkCGyTqe4sqGB
i103ZJlY1Bt9OYukT4ScdCr5JoHojtOJgpsefp+H5KKr52fXhavQ0bptvhYoK6SH
aCfYKkZKpPeLjIc7Gk3sy8+h+UUDN2ndOxnrJmNPMgQf6KTNORK6kP0c1qXJYt58
8mutHBq3Yf4I5Z+QTVVtUzIW6+CUJJUKrMdYhQrQ+isyP/2lALP3eoIcExacHcHS
iYVrt9O/teq8BOdFfClXqMEQISbRA/mL3IDu9qL4OzLKaAn6rNwJqpjoHPs7gjEJ
fYwwCrZkegYf1VAUccDw8CxPHP1Ib7Yw0kNqqY+FMLrTumulKC5s4S4oYu1widfE
0yuhMZQ7QJtaacokQIonH1cdIh20y9zlk8x2+37b5F/cDX7PjGvxlmZkkJh7D6mZ
gxyn5xmswl9lslMAQTeUBc5oEeV9TwQTJaJtsRDXpOZzGgDYMY292yCGhuB9X0jH
lbvK6kUyjipKlPgR7fGsWFQbhj10Pc3hrizruQDVDGKwAsAMdBiE5cd7BSFBno//
bk7BV12LveA4Zz+5uq7N8vhAcKOKBEmFkpVPaYxxx3BGb8Mkgdj82aPSLn7KWIG4
XjAxYj4zZQu2Ux+L9UbGE4vsw1n+l6mhfjil+qDnLYIaLW27PRsFyER+f6Oj2hPI
hYH5lKQX/TgkYlm+a8Vm5BJMQQrgXaxlj1bvdjfC0onnHQLze+Lc4lmjgwkN95nZ
xRtRm7cV+PKF4mwt3Njzbw4NnuL1LqY/iH0+H+lg4yk1HD0x7UOMihc59td1vM9u
iHx/aSrhJrigKCFgwfHCf5ukmyLwPqB0Y7OBBKzi1WJmJlPenxFkn02aBEZwR5qC
C+1YnhFa7LgPpzuiZv+T7Qr6evFv0y4SPVdQ0lQpWvRVmWBpUEppyDWQfYbNjfdn
m8RiNpnpQnT4EG+zO0vIkiipQhZnixNYXeA/V6eV+h9Qk9HgACclzpGKDRq88f1q
l7DpgnnVe39RYiKIR1PnUKHce4MO/Kczf88/yl8LX1vcwoxPrpis0ccurr6pTA4F
1JF5goO9+dsD6ApGQn32KsFe/AWKfx6v1t6FItpoAyJlLqIagOMRl0+SjtCmYa1e
lHcG1VfmD9ZUzroQdpLOuWJKW36EHk8eBIybOnTvKJdvytTA4H2ioggX/i3HBhR4
kjZXu/YPID2eV1Trxp5kjHR5ISV1TyjIE9lAzccEoUmC53ZNl+W3t7d2DGpvky6w
pc9VCoh6uxzbizUoD7XlNPWuYjZyBgWCRkDFXNsxaqh7RqO+w5Rzw+RkmHxhvNoR
PLWS3wWEhUsjkam+8vqc65m5lAPJSNKbohY39MeKCEc6bbtZsLN/tgiXHO0c8Zeg
ORR+Yop04lfKcfSahTisARJ87qS88G/Zarbf4mw6JOLHXvonhUsd5/LnSxnK133q
xZgWDvHFeML1syRLHq3vxXZcQzCewu91nlygSFaT6nQCHEyZsj8KlVXFkveSUo2L
L7NH/0E2d3tLKXaTbfV/++1jpuQeXqVrLpK2XKGQmuhnZ+Ht/Yvggp71BzwqmzMi
YLTcno3s+HpNK5tfSI1fu7WVWo2QBMkKGhPUuViO/FpViMrqDrH4la/1exOMst//
RSOX04gMtLOzcv+fQlarahrh8QHyvoWRt0EtihVyQahoV1jVNo2xgZYXlm6URBKj
foauTm9/TQ2CliHhIfBYuOs0iX6e6tto3YomGkG0gURQIow7HLLrjYjsjz6z+Y1d
1NmHGEQkOvOXA7yHqli1QYp2LUsoGq+oFSgyEmVpL1YR48xPMcNaelD1bQNpyWWR
TmRvwXyjMDNyAFvIzou6POkuRsqIKZJwCjqG7wvCgEMmcX+bb+zyD5l+Bk85ij78
yQg4wWUylyxslMLvqSZRznqnMI1CNhBUPX8qQPDV45WO6sAvOeMQU55czg+48gCi
WLLFcdhoXwzrme06k9fUm4YrJ8CIRKFobBz1hQHOqRtNKj4oWIFXRoSjd8uIlXbQ
eh364Ib+Qn6djthiBQZwqhdF3MmBVHhaEMBUeV+g5Ly7obmEwGhiGkq/UR8qE5QQ
+amq14WE6EnPTDtJ+mOKNESudbs8CXxL2ldOibgx5jN1e6eCC6h8OcBGLzAE/sCb
0j2bsXXvznok0RTiKa3WwAs0EcDESN5tSjx3D9C+jsObitSnFGAYMv21R9ogvqTN
HVic/ZeCT4iNF0zEtH+CvQPTqeMk92gJdZceped4BKLEuGqKqhRxZa9vVUZLagry
45iAGKZ1HWlUjV5tGydA8zwLNJ1XkXBmxVJk1L5gEhQbaKHt2mLSIugonme2m0MR
0mC51461hSCFrx4OY6G33XGbOhyIj6rSKQA9Igjcbtx+u7g8Y/Nl08OOuYJno4cR
zFSv15iRXZ5PVXS5sqBR6jxnNRnf1raCNq7N27Kp9ixoh6OCTtscUmFbKNyBA2oC
6DMyTnrAJSPujJPfO1t8UEzF4iCV7DiSu3OtOwjEKKRPzWwzzzRiqCaOS4XABKG2
LjIOub9n1iSknZdFa0f47htSBDWFzBn+tvBORKACD0RTNs8NPs/r2guSy5Ks61YO
7wnlxjITHgEhOvWXgeDAhSy7w1b0j1O/q8vrTnFY9oAyIbHXYj4POpdGEr04fN//
dNHz65Wlt9qYRj7zZxW1iEIyvr8UqbNCKv18HU5SxM5JmvBZ8CaHwd5dbi8igk/o
cZ4FHdtok81DmlDZWKX5Xu1m0fCS/0QQOeUxlfpbTOmlu2m9UwlFayNz504yeYP0
pO521zW/hA7I7PwtBG6xFqiIA/YPnUraZzLllAQK9PV1qGkrofARwu3UTtC1BgHB
hUtRS/AIPuhUBWt8yXuG5KeHri31G4fUmlqD6bLOwNje+u/4deBxYn3QXyKdyBfX
QqaO5X6LDWhCbyE28QqYCjuyrB4gSHAmV8O1yJyYhN0v3jw5+fOV8JVF50oYNgRs
C/RMbj1B1E8ZrC2+k/n9AFbgBUo/Jg9hfcAKQ1ZQIMu+k1zZAtGcycoyXenHvFiy
sHVvTo7yQmSxPAFJ9rxAiWoBEQJUkk8MXGqHH1zjJXIv7C4EFFZn/V0ncRlCOKMj
cNmZUxl0grIdiV1gUo33FGNk7ATUZOvL1nkjRFu+YAyrzRGS0e9EeghlVG2xYLxo
Lw/ByGpsj/OsWjuZAYvEKNv9mHfBBy/C9iAi1UDdkK2xDSng//Wsls8NKl8KKpe+
UsoQcdCysT8QQVHgjqsqR3ZA7ooDj4DlLHBfVQd2LzukL4KD1rn9R4/mcn3yZbhH
xGIB7UkHDI3M/hkBAoGO+PEPnbRLoJef7C6RMod6Xfg5wlGdKCIuwN2pQUqxE3hE
2eaU/y7Z1XfkjDQ8QLTrnfGM/mYNFhvgwclad/Aj2eD+lfLFg/KCCb2wO2R1AU1K
T6bXkA7Tv59twyciwLTzn491O5vZVf2k6+ChGuL3FM4Djj6cDQUBixuLeACFn/VJ
mJo8zdhtJA81U3Y/7HWMZwOCWlhfz9JONvHiRXWH/2uy1gyuv6bKPo1WtBqQatQY
UQ4fXO5QBHYvSLk3yscHGicz2HTaU9KwUSvu6NAJ+WGAXMN7ajK6rjcTwZfXzkPx
2VGRrBw63j8bW0te7jJNtVhhW5pQUXXYVyMMaY5tTCMDOai2ui1JqjA0nTKU8MSw
r2roQIdtkzZUIOOTI/TA0yUtRvze8v5XrhNRric/H5cATBtAWmBEwpiFVmr//ED3
7fevGVzZD5QPhIlxIVx8lUuVISdH2itJ4Cy496eHXMHQPZehWvwX0gzO4Xy9VDdV
EJruNOGc3LKtiSG+XHEbmSAM73aasqo5YvtPB3lTck/33WMHyS93ThwKIcXaTdVD
qhwtym2mBxVSWmTPIjK9kiSOkHgq7nVkB6Fb541qYo0f7EvytC5LxCeyfQ6QNE9k
PSo4OUi/wDO6kp5OQqoQygOdJRM2xIb7trqALBSnZQlLGA0R56P7aeVq20BHKXio
kMUAxQbfT7zSFYGCI8fYQN0OU5MQxHHtrYg8L+dBJlD2MuKRKxPYi7kwoVYiWfPb
gWnd+IaIlNTEnuqIdIgDT5ZRJXxhJ305oYxfw/iPxiY3zt4I8ziA/JOvvd9RudwD
Mo7KYvVr7qxN2wSDBX0ih9JyMB6G9IZDZqqzHMrfto3ElBKEcwde8jaBQeEnbwqe
tnxindF/1H9aWCsX+DZSfGvcEcLBdCnsIjiOaLcoRQSUQyDpXbeCZzbMJh9mP/Do
gRnvhEl7x6dH5aOO6UzCGB7lbWj/mltMbhWHTcxfydLyvpImJ+G4qxxk2DWNvcx0
mj7uF65gdTclBPnAW4RbRUKE7/UIwg27/1g1U9UQfi88TW05OAcWu8oEiFyqybn6
Wm34RNiozE0yLToocgX0mxmws095kNNyIf8Wps82oqMjBdPNRGpDhS0bL1h6mP+/
3Jd+9UYt9J8FewNJzAN0YZpJPsgG84iCAqrWuGVgREtTJsa+AtZboUzXcr+giTD3
Kj29sYrjS0lV9tS4iWva+gC7ZvLByqsOizkxAaAbttCW+cbdBJWc7aLt0iKavuxC
u47CE3h1+1rSxifed3Vtc6cR0EamL8cX0i+Qq8PkupobpNfcdrglSaOUEyh/OZhZ
JbFMXvrX7PrAOO3G96BQ1gleIt7s3Y7zDnDiyKpryuhvRQMbZOvjlrBcFPWZLVXl
zpFJF5jH35AsO+94Ao5HSPtcu/0ojG6SBmASgx85ZKczRW4MeQKwAf3MiBe3sQQF
Lew0QCMneEYUkOARhOj5XfkvN8Z0/28GJA5PiRpPnLM9lO3O3gLgpoNxhb11bXwE
M8N0uIO2ppDs/IORRA7EDP6I7lVlrCpV5WQM7m7JydusC+zBflcULcOj9gK/J2/X
qtwUqVSHsKzCd197sxH5ehocIHJVCeNVyJjq3YNeJkzqLC6UpahGmt9iR0BmZIhU
sFmkV5asGoYpLLpVNYxFpZKB7YTiiDkxSbubsNCYLEMmhbSCee+g9loIwjeoQFUQ
XWFCkhnw3AXytLb639iWBv+YGcbBk2Olz3o+tTJyqXLQ9F2thuMu89QeLoIqVYvp
ueZNtc6lb0DdHb689cNLX81h0Z/rpgm/k7/VoEsDdlRWLz5+8zxbCpLC+twQbi2m
4hSFR/QCZD5jdgVpimhNfDHocp64enEEatc6bVRgPxxA7CJlRZQprFI2n4MhVWNm
xtX4q7KiexRofLwQzOPVTjjDA21kOod99HO99exo5N3ZZcJ3geq92B8PIwRJ1T+G
Dmh0U0XRCeNU3+UioDWfdZceZrRaUBnmkyelf9BVLyWtKNJVYYlJgJ//l8dbt+j3
/tXqKujEnAbzQQqsm02vXkhrMRPD1WpDL62jqnpLMEvrJNclw3Zf/Q7yE+CfxaOy
yfMpKjTJgu1vl/3XYeGKQiG3riJsq1MNh5C4iFQz0K8bVFB1pq40p0sRJe+fHihV
md3J2a/PwmxbqOnAK+eyRhPs2tpmAEc7JTioZ7DWEYDa2ol9I63Aau4zBOChs8sC
6e8Z9tsMcOPYooAJjS2Tht9RrrdjeY/xXO3C92klDaoVvGTsllAoY6/iMuWAOo6w
UqFrHtI4BWFea9KO8vmAsBRy+WxiGt+qap3JeVogLwf8aoVQcoPRwdDdqo5ROAr8
IB5guLLzylBLscgQziaTsJ2ZJkItBXZ96cM5lt+6gIu3rFgoKcr3k5cRZtnJ8A+q
HmIz1AlSj/pRFojkGAU6bPQarBhfuqsTsaSdXo3OooePuwLJjx2hNxkB0s0aE+gG
VZgG2vnIa8hy2fZejRammGKePN+ZWF8bQ1FHSmMEXj3GFsjidprozpDXA3TqrxE3
Uy1u6IK9TR3s9rr1r05yZTyRqScB1tIU+vyJolVpP/ztRd4aLEb+h63wP+at0kBb
Gu4HRAyAPXBxMt9TlnljvDpfm2UIsiXrlyccM9pIb8a0ge44ilXwb/dO8tmIf9OE
3KrxvpAxZhMfuNyhoI/px85B2QthNnIoCN7DQdiGAHuKyG+4Cslmo95j1/OySJvS
B987sO0ViNKxB6IS8VxQAp2kGTYy7qmUw6J6RRjEM+TxrxZhhSlZd0Q/MMv3pub8
loO9NSTVtR1GuXE0b2fmhUy8FIgajuEJ0FOnvfxl44+x/DBjDT0o53NlcgAaQ1CX
LDJxQCm6zlNjk/y3AwwTCXpxYcPfqT+ZDyDZPBBvMQSpM3exaTHjvkc2fy0pPbel
XKVZQ5NkSmiOSSO3Hi++6ad6K03P/7zCxA23EVV7FtoG1UAvqMtRwNV0/cknacNR
mIdZSEvGbmq3Z7wNTKgfkOBlVfof9uBTK+Js9OIHgBpGLxMnMj8UGDtxbFWD9W10
UyujMhvjyNIM/OdR0yC5fJjKWUDoLjEs2l+eGo4Ijm2idwjo8jdWNX1ZHGwJLG9o
kzUQnfB2FznfKRXAexoNx7Ayf1xvsqCUVwyJVY7ApMoWNdmIpHmJLQHbTOgnstoP
pBeTodzArn7oFhR97ecAvcYgH9G5ymQnkUDegnVkngYDRqYopx1Eg5f3v1jN/B77
CdYnahM4Sqtd0hbOEiJEf+AAR/qkAlUeSKRmAIOTgqPk2R0hX4nkcrOK7r3BhUa+
40QHTYnR3nsCQFcub4+rtzEBPhJ/RDHvghuGQzJgKKUURrfZMqY8bkQezTDriopZ
KU2gPkeELtNEzqC7sRRtLjC8TCduJZcSKrcNJLR7QlAcu/27eT6M4ysMQ2EC0rL9
S2DaqKHusfXR96F6VsJO/hFGMjvKbG45NSaBDCpTz1OO0jl1d6hPVDgv+htSQFxB
bEE4qLEqjph+yFVrreGbQA5liSmtNhkBF5+SUNTNHzwHl+3tOgovaHZCdd5+NqOv
FVPlxwRPHY+q+Pjvm32J9jxFbH9k/V/riLva1m6ZvpmYXs9R+c0yEGHvU9SrDZYf
vC6zJUg6ELZ953DAayeXjwIcMOMZ6PU6GBqpMk5w0kRv5lq/m0pmaWlwElXEvREH
2BdiIGHE03VMhCTw+JmiA/Z87CAspYnpaA/h/qj4TzKu5HO/S2KxQhObcbXip6RC
Kyh+0ly1/vw+5Nj6VOG84D4a1Dbdl3UkYeQzwIch9BlyB7pToykJkMEfVB/1MbnH
XaUQNKueo8e3ms9RjfvCd96tdCw2WgkflmOyyJFxSwhFCnzLIf/K4OnT48ejjjB3
sJ6wPyO0Ll/xlwO5F6q0jPGJb0XW1pegI2hn1pm/L6OucXQntPkZn67lsi56Jjo8
JnWKvpYjAzAypq1zbYY8c/KuhdI1gU3pAhs1mWXJT3U89nwQP8JqswJB9Ly0Fq62
6lmTak9j42aFhqYtl/KDiqIG7P0z+GWeyqbzjJJBdYrQ7/fh5qvC9PieefQ8zovj
QcJ64rEeqGZqhnELDHgEWsdF+x7SgaafPvrZJgd71383lnQKATje4KSvLvblrhMA
keOlraB5iqQvHEV4vmaOyDNnZNEtyLEHlX8waHmgnXeMVp8pZUPOsOd/O5COXTZq
vjQGYeBYtqnaMInpqnqCqazPyRVhErFlY+gczYpX6hnzr6g/YAWW7Ordd6+rjujb
H2xt4giFMoWQAXQVfodhvy+s/sxk0n3ejIRgXCbuypeytFVtX3xVYw0odF8m6rMR
P0ts0T12iRusxuXREOZynAqgPrl8E/qs7q0r8SnldVyF1eH4IKdgzGVP7xLabfg1
CTjf1+73ZR4nQssGt4vDyvgNm5vW3lrYLfICLFIYgUCp99f2nsVlbQGQVt/2vmpZ
fCLWZNFIR9CIY51DrSnNPKmja+iup2hD9H5ByH6ap+gP2LISQj9RK6FzP5U3v4pt
eEVfLEISqaj+bcnfh7D2X7XjiwpnTtiRGXUTB7fero0232yhFnP4+KQT8QgPVCGk
1sJWUaO5XYLJ19ekacUavlgfIPqYS8HS8KtUfBD+6jSChC7pq9H5bs53JdNJQ9pR
43CnEfO91bl8CsIt0MjcnlIGiSTO9FjZYl5Qeq4Erc1PTIcTogNRXjM5VMSTtmUA
v4ZA/6gLeSXDcZcObHKdvI5p70bUDrqxozSBgyp9moe0L5uYDYg6GuRy2aOPpYmg
Z/QN0pTFJBLZfsjhNyz01GifqbO6FVxkBTHNasLVyINjtKF3KXfSxC2an789jjwL
FuXr96k/XN3v328koEtFYVlG79lBAKRXpgSbKLcMcIY6tQquV4KTZ50KNl01XiIC
IU6tq7o+Q0d5+OKdvvjIelaotMCOmrIjOMGIzW8DYE3hZd1KeZ8cdPqcXXF7Wrlm
Lwvkfyxd+hkZhNa6anLPGbhlDvrflmenGwJMlRRWwz56cpxHdJe54yuJjDg8KgLt
iR3tdrxH6xFo1DXy2caQshXu0UB3IzNHmkoI9/eHPFUB/NkaJWcCVpAewVg7acgV
M9w7wRqt4l0gUpqmn7xr9CZBeeWF5wg/9xCdss3oPgr5dLpO/khbPkRGBQ5CK4HM
CNGWT+2kkA6T1NmtdmbZDC/BYT3e1JIMIXpu9ode+uNEf6X27jvSWtjOlqgA+3+N
eLJvNPMSNWCg+LnVZAO1ZVGDBlXpFfRkIKsHfUe1idEURYcbplszNv7JCfCAz8wj
CPSbKDXA1Kah+w4ryDQz7+kKo2mRjubKfhwqHYo6k5dq9YQDwQ5Gv+DT8Wr/haJ/
2d+Aks1GrIOBn1IjuMZHz2ixBpUQjzffxBRUiihk8akr1KOaj3OMqCIxL76TVzzo
vfbdQlfo0lyyc2ZwhLd3UORFT7SdwZgb7H1XRWb6U5fPkA1YqMmXQH8lQ/lCduEI
T71wPp1ixV0/DrNK1BlQBBZSocbboEF5SPBn4uuav6GuMLWrHVcXiFqfht+K3iq4
w71KJZJHsSJfPPjwYppOdNtM8cs2bXiU/qP3MH0MxUzxwRcHadJaZ+DSuB8QPdBf
JSSUs1oChAekue1BSvg81nfJNm88IbwSx0s3Cg8y0cHZadI5xxYwexV+lw2O9e/1
gwNp2Wjkf6ihrITdYkiIPqMaJvDy6ReVUeoK51DhbNdI8Kb9u3WEDTw9gcoNp1xu
Skd395YB01LU+gT3MSYULWE7L/E2A/vykviYYvepZbfua00NwOfxdoU6DYyvTqQu
Q1bqBDtoa2zBLX0EWImDe180pwJosuugvYsyUj9LLuxeoGeRMJCpEp+YKqIJVulN
oF86EyLNA/1jXZG95dYg0SQ9dxrq3PgVwxPMM7xWGQCxeUqSztlWxO250Eu5xIdK
X0OmOg0pnJ3RPFX06Bo9hQfP2CTmwDJEz7w3MXF4w2E75KZtFqIp/V4UrsM3XS+e
GValZ5/TiiMT0zueyrrd2Lr7Xf60JJjNuPAYlsQ9H879vlukracO4wESX/JO2hzp
zAUPFLCGQ4i7SZIGfDlYwnG2qcENsRSrr2lpvVx68a5ka0znkbosaAdm/XxoCUnO
trEuGACrsyPsMDqDhU1e01eLhqO0TmmXwlhWNMZm8Z7v1qCBuIDHf5sWlIGElg//
zKnmT3yNBSf6ecfgv8ntSDxTFp6+eW3GmOvwuIVbAVJAxqXDf8tVNDW2V81hG16r
o2EcKybTXrVGScBahZyw34zLxKmzjHupw3PvI8kOXpLPMGWnfTZh7kJ6+IoaJRfF
rDxPD2K6f12xsP9s2ZjFIYO0o/11gHf74I413C2r8xbbNYEIgqK97X34ysUt9slR
ju8K3uteUHvepAbvVhsd2MVNwry7VQtzbFZFWaNZIlObNxRZjBR/HoQalg/Z+ScC
Zdth7TSXHyhuMcpNhewUI175dIi+V4h84wSwxmF9jVlkLAMeLjYy477RWCunQ4Zu
UVLHuOiB3ASClaYHZfzGLflwJDo6VHl1+2ggA5eNz4a4ZowQxdPawYtAFEbMBxKX
5GDNMWCVnhUIXpcrZWVCEgHW792NiQjCSHfrVD0Zby9TCUERMB29k6uXAe+EpKVo
fORn/MjDUzBeguweN3IeEm+WPBfgXHODVK5mbQ0RuSuI8sTTwMa/lRMxq13dDpJS
RlvuzNm7lFa6NB/yMYfpYF1Z6BkMajlCIYTU+kL1oBfOuMgrpJGxabOT43HBn/EP
/BLWKjhP+/5dV76gfu5BTpdIVRCyZhkRQKqVz/1mlZ26XJDcoSl38QqhtOnAkpNC
cYlap7PtZv5VxTC8AmG2gG9Q9+EO8HRZE0YlQymggu2th59gZIZ7owP9YTDpPExN
R8Edohe3mEmOVbXTB81HQvxQJ9f/q1r+mzGnBJ9vgzoiWiTsN+4kYM66c+l2Dzf5
zbqFpwTbD9gqYvjjtKEFbiwkLDqCjPV8VMLiAVOj5WzYBbO8fxpAYZPUkt88N8+s
hgUvV4et1GIUmj5274tWMNlWbR001HnmSRc2pw5h1FKjLGQkOFaiuvnJ11GF58pU
UJlxFUgXMgb8HanUE/TjD/dmn24doc9B59GZ/ohsnal/0pNRA328DjlEzHRBN6Og
MZYD0U4fxBcvLCrStNulWBHwkmrLDuaen+3R3yYcUFMMZANi27n9wUqtzk7TUu35
PQYeQmFvNY034PaBuPPZSgFl7KS6NUIJQGC3cHLYyoehq+MZecptqFg2E5FTJMXV
epHsQSIzlnPLqB0Fyx88G8BNOcyxNw+nCjnUX35E5txxDVc+GoSsexfOTiFvJ2p1
6/jS5pX5b/KqEpaGhkdz3EL7OVugroSmNBWpNfZEdaKd7fkweaw6k5puWHF196RH
MZPjkNDHotOFmAFZDtU79oCNjJFqfjJkhqgcivpMIHpej9JEnL6AEMyaLx6iSVfU
/tzd45VNb3mJfZMn4GqO8WJGpMP/h8pqK0n+yGOZWxooiDdT7X98d13Duzdd7ht+
3kHTX4lKhtSrZ5m7enZvn+dz35ZBrCQEGFCoxEyNQQAt89+bPTSCFj7QvL3mhjkv
GkDz6ew0l/CA2S2dGTPKbfnUI3GKR2wUrLlL+cvWs+NJyS5czIiMSYaSPZjwjSgi
pTe7Q3sFY9yqjHlgBzG+MNT2ZUINESqyeJ6hG0l5H+XTxMOh/MNAiy/iQz2+ECya
5grE4nNq2LMnE2FxJveZirQhEOYy/p8fTRC0YJE/9AlW4BpbYuMAoQIlqi5SL7cv
JeO424w1fF/OzICfqrWUzrBhOe5rIGMty1csHdaqz3gYmcM0M7JqelzXPyMllvxD
DGNYJWxBLFJWzs6kyXfa4MtBr+7jIfbPo6oC1/rO2cQnaXi592Dn2KmLemM1plsA
CIGPnEJ3b2b+11AYu0LaKgMMmbsc97pokGQtHrQtdMNJeYLxjofnWdtWRkCWi+sR
DYGjsn0wcQFXltHwesUWLoB8syANXI+x7eoifpqbFuB3feUxDTBXtk0VRDcbr9hV
XyS1wk5bwW11tX+U4oPzflACg6kRD1eYM961B1+6BPetCKsZSPpb8ZGkoZpBWpFz
5Lu18Jdb1T2Z/cBkxx8MwIuyezKAN37IwPrtJPeJdcqdx++PZdz2Wqc+mkRjtxIK
QZJzy4h+s3dMPKzFu1M81sf7qFSpiliOA2jUw8tBPyANBSahgWexBqCAaHCodgXc
0tN80tzfRhhDXx66ayrFzeunBp1ee/xcy9ABq3aAngXKqUN1RBAngDNnbVRqWo06
3jrQ+9pvaf3IjMUK+fUDEc1zJMl8sTFZQVBX8b3ZwXOpkFfxlw7Es2t8xI6AruyJ
Ua+F5h0eBg0dFL9GbJWBHecbcmFpzZvspM4wJnLR0vEXnUSiBfZUDicsxxX5k7Z7
LVuOjpcGd/s3p8Yz0wCRO2NZ/LCgHPjyk1H6rrxq1yLtFmRdO9qNID4w40wECD10
FqYMgsFj6Cy/Qc2heTae0LJltqJwuRCuxjF9+uPEnq/nKUPQ4/N6Jv8yL87lMLxu
VlDW8CE4yyNF5+6gCxdXJjK9oRrDvwBKOd2r3DL4UWNOwlTDFw6B8snk5MzqqoV7
uvTFMDW0N6gZHincNGwb+5olv9oFdzj/wFDM3ZuUDBeFtWWdAhlRGMBsLxHbQlUS
0rIhCtTx1elRCK1w8dXFvcEAWKt7ajlk10yWnm3HweT9B+OMmI6ER5jcYEXWfGwR
NjU1MZeTAGkEblNI+sOCHLRUliKKQyKIxOcFREzVjqoy3dX/wxmJw9I0WBIhGtU+
7ec95Y6/qaXSUyrmJiXEJs3LWQSRITsbqd/egMt8+EA9NO2yjxqvJLwxgp7SEQVr
1K/lTWMrFkXEJzpjSSEj1OnaOalwmakmD8RMzf39W2J4zP3OAlownoDgUKDTwqZP
C7eT88UQqotsCqORHP6ufTBtcl8McsGkGxMgJO6Cgogt61iA+ImUuX4cVODuFqLD
TejN5bBAPCgPv4loPcX39cWAgDzkU8Uftpe5Z6ghBHcOFLfwPutzXTbMFTPlTLEK
X0kuM9LKYN5TYLTdtJzsvrzphhL4O/znFMS/sqaUJfnK9B9/6YSQ/rrUWd+tgZM/
jGDh2Z2q8qbJhLf+Q2kz43n3SzE+49CZ/+s//AVt/EBBuz7UqAyKozQ8RiRIqjsK
FIaehklv15HpWuGOEBImP6xzryj7Ey4G1sAMj/CQnVNYG0lVn3r6KedrxHz1g2lz
Zk76sZaDI1Ju59pqbC5Py6praBc49grgHEQnzem3lnAksbieHtCZmbPCM5J4SP/F
45ITnXK9JCZC18OWA8bMQfRQ95XDbXXKWFc7aDvuyQUzCUbLJ4Kub3qQev2JlZHp
+qT4jGqW7ZiWFzlZMSlRiUgw4p6fbnWiwQ6jAhk4YOT5AsDH8bVaJEKn5jucTr6m
erEJKs6rjz8VqIHkjIOSYI8JWTlKJJyl9XDe8L88WUuKMVipPLJExQbQY/HKk2aF
9YwencE2rrLzGJIiufk9yBAjOzLk1ru+edpV4dCooWcygwo3JmxOI665Q+gz6DS5
v1PXAv/fWoDHV/Ta2Lq3nESbnK9iFanAnp5lj8XbEPui2w4jfzTTsa7ZSjBcmfov
qt8TbU2zUcD2qUquP08hSgj0Lr40x+ZLOEoWnGZQzAF2v1N93JOFwyHCrnSbMmXu
g/cdmPO5a9G/w/lUY/wl5ca3AkaPVQqKo4JWaHrhRGbv2eM2k1yylA6XkikJvwLR
vw2xRsySKa8FKCx1xo+nbAY1NlWqjGGN33TZpsGetQL6UrLB/yloA+QNInYMplnS
29Z0Vtn5fIelMbNP64qmcbXMS8bt50P6oQKoGw3/STwP/y2icyMu0DdWv5kyhrTL
1OA4/pftMaOaPInG+EPaXxU3pH4msI3vF6RjdzUi/KQbZA6TJvdAkZG7Df1eWVUU
rXEU/6Waph5RmTlnZuLFwSuCzJx328WIq3Pe+NRHpjJTsaZ5jxRy8hzoSLgdp9s/
tPzVypMrPfJwh1fWrSTuMFax11g+6QiuqLwK0Qyos5DV152SxDwd8ll142b7lG/T
9/XvD4Q3JgNRxLr5BEwq1M3clFuYea/N9cJ3wklDU7Nzdx0w3rmgk5nuJH1rDyMj
N+PKiXdD9OlnnbZbKg/VLPm3x2wprGnBhgdUL26DfxAdlzN8Clj1A+j3ia+gaq+9
zMuSWMuqo3wjPkOn2p4VndDIyXLQKvKuePSrJqmSrVkfbFfheUz71JUbEWICZZ4H
RUW44+PEFNsK04v8byA3jVLSP461gEynIvcbcx/OPKOqjNWP7pEhFFc10sWKDDf8
UY+AteQhC2Hc24xZxKzEOj5zUoDeQGqVQa8I1IEcuOEBuj7BF9C5j4B7K57gpVcS
ULx+GY9t6JX7ILUIAM/ImSnO/eX0VkhpPyMHk2ZIlgysqiyIyIWeEmLQS4EsLLCa
O9ixGGa9JGUgOPpfilXLa4XrNsd0m8Oq5JFoWqrMBwqt2+4fKKMcFOZEr4o4I3JO
iroFEhkjtuQEEuoP7Adh0ZtpGXJOYc4cwir7PN6iBY9FpPT7T00W/nfIE/3GYbTN
hO1+ICh+A3Q1MkTywXBlfMsDEFJyeEWZgJsV4Wax9EMYYWj8pa224H2MBcE3HhZV
Kt0Wt0jO4uis6KoYjfC0/2lSgo2p8npOnIfZ/DVy3/Ymy5tgWBYzR0JHxHHTrPtZ
nbrGNC5NLNA3wX5Lvd8x8tiL8bJPTSjk06qw0dZ7gc3KpYSXel/FMbZj0aOIr2E2
+iziNAiwmkMq/3WQFU4Ykt8LY0eUEitggacjsrkJYyA8qqvrT17FV4zBjETCkn9E
qrAuzRXbS25egazw6+8eWTVoieA9MtpByFKY+aa74Ohx9p5Rdgx8jW+tSVQtZemB
tjeUhrkB+CLSaQRsIjB2tDu8KybYlvTKUXOIWMXekd2YZAPnNPuKIUabr2KAVWUN
MthBiClRGDG3eebno2B3pGmPpvykZ1af2Ioax+Y3l5pk9Y49pZJgr4XVLlDzFlpZ
6F3bEgyuqPEbv1jxCXX7sw5pik3NeORSkQvMh5zScr7cMa15sKxkirmeC0NdwUJw
t6Fyt7O93h7ZAQLiMVcikI8DviG1TnZaQ+LDbYqR15U81P1BxiDGWC9Oar8SgqQJ
wP/omQelrkGEkx7+HKBgkzdv/CZ2ycYv8eYEJzqHXvYb68lhlO0JeZ8aE0HwLu/q
Lnt7bM84sA03VXf46vfrIdlfrQKaMa6ITKPVkijLfP0AkpmRgiTNRJml/gkldvpL
P5HnJYvHCSkj8tTCgf83R9mIoODwEbeW4KrjxmtKAjW2K3Kng3OPqIambLJ2UFo0
KUJ5nR5M0+k2tnzqWYUJjSGF22RHGKSdJ2wQNLkuneOec3TJjDoRlXr8TaiIRXY9
KxesYOpA1RbdS79A14UqMZ2CXbykzeXsXHrM9R1ukG8oQQ5mj3i9mMk+sq0xoUqy
BSACsuy2Mw3kOcIY9BFXOMyCt7z7BslRsGNzq8eLiyH5PUUEVa+y8JOaGlj1aCKO
mUUKl24m5lxaXKumjh27ToVUTrDY81kTqqoWr9LHbVy9V+8mMiMjXAwzc4Vkodrp
xOregSvnl56VPEeU2/l4gzo88K7L/kjsx6pDPpg7nocRX86fazuKs4NwHlX30kJh
h/qLwT/Do65gKAo0s+CdXrDazqeE6ka+xfiX6Dkq7FM7oKtYqaECCxSUN8bcXeMy
FZpVpaGdDDlSGeX83GAxGh5uZYmDvLOMHSeBnmpeKwfps310i628qx6v7s3NaQJV
W4lo6DedxmE4i91qThzCOQ663OPbhz9vuqVeiBAiuE4UpY1skaTtFQWK8i5yucog
M/rKbyUK7cNVw3jQTUb/lZ20jiVO2XlmxgHSY0qhcJ9OlY+EFWbxzOKATlKLo6Z4
NnqxHkh247DPgFf09iBgEzPFwUd0YH+HmOBHPv9B7bt9LEIXEUDev3O0dQMP2gb6
QYOsqe1LgqELQLAC0y1RhXCA/nyGPqvWxnKRe9N65uit6sMIMvMNS3qxnM4ruNk7
jWTfRPUseCeXP4JxVnV60Y0yLX4/m2kgM8zbuSt7qHx+U8MGglhPse6rsk8R8U7Z
3BwROPxsDu5ITkEwKp44ABIL2hmdRfRPLS/J1JV2j+dx0k2I9IrA2jrWY1FHUSwi
OpOCpOVDFj2G2zDfePlR8s3PuRKHnjJW0dZe1poV4XAtxTucejTTaj6S+Geg225H
kFJNR+NvSfvIsC2//2wnaZEDe694Dl/jUy+JUEzzZSfa6GIMhK262XDcHn1k24py
uo8feiyqQiz4TNznNvLTJLYXmCeygX22QPFhY6CGxk2BcfafoXtMkPFPP3pGeAMX
yNOxL3GE7YtyFPpNezpFXGvoBItCESf78TKBHPBA5MpNckHmEK7GutCgpGHXT7gS
RkNZ2DXGWsQmXJsbV1ufZTZHoBoqzR7uLi85R1VWHuRu/WXY6JjlwcNWB+nb0fRN
szLPPsBkSfFFV07mPc3SZvyONob9T0YIoPfLM4fmHtSl+H3YHorza7R2vDXrlWqa
VMTXB+KocoHU7CQUtwI9hU9l/vUfF15R9C+OkY2Id4BJS7EfvZ26LNPwuF5/vYof
SD8mx6m7GtiNoiz/eCw5HTFUHTdc1D245AgfOAfUALXNtHIsTPl8O9MifWx9OK2F
/wExu+EVh1te09OaVnEgIVlfiGbi65DRktNlC8jWBeEswj8H2X1AtRk6T0gATALG
KnxiPdUKw5/JFY0FLWqCTMdBq44Q8nDtX08hWnm97AKxfgkjPNtClNnHX2eU4i99
7jbm1Jrrxwo9jDqMx+y3fTdQAmxvYtSqu6CQkJs5ynVKOhokQoc8a/S+QlfoXHWf
714s4hIp10LMPqArIf86zrpIfVquX3XzV9M+pkdFbSPNgOKRkq2tWo1H5t7yL1Q0
VqThSJhpFDngefVoD18TC1TTjF/Pw2bU6YibVX6SnYqalS482XOe9bG5j13aHhYc
NCWizshsxQroBoQepK7nCzz9bQsVpSfv2mDsK979mwvhtdrdvQZZnCXc5F5i4ekB
B2FPaTjB3Z+5w7ShDy+JdQBS12g0SowH6OjAuZMUznphVlK+db6lMxURv2BPA2vl
Z36+e5g/is2agxfq9sQO3jMnhh8Q5ZBKS836EozLx4QEtrFgFHfM/y+BilbFBf4w
8vvg0TRR6QVzepJIU4ceTiJ3wQSZ4fsFC2mTlPLBiyYZI49A5YSewUltpHNBIrOz
5STTx5jAXqVEGLJX6vaWMJ3XB2+A7EWURxtcqYz2Nh3daPAqZzDGsaeyfYGfTnWX
CI+rcJ5YWREAD4eSarGRysQDq8K4F4h1p8cJlf9St2xdKldfIYUnPzFgq2tjA0EK
IlXQYko4qKPpcQOWJgtl3bbK3Z6tQ3y7dbIePuuM+UUHFmwAD5NFmyxDzfd1fN9Z
CMDN4z8YN+PJMGL/wmSLLnNWQbcapX2D3oWu9fc3kjBPenmL1icfZa42UFCMCkyo
0O9LtMdO7iSUHnuPxAiLpFamtzKcy+WXTlnAOLfxW7vDPNmufKc5IQjqiijIxBt1
OuthPjPdUEo6GPa5iw9Z84+roQdCq5vrY6qtKa9VhZDcpJ/eeUW5O1/qD/EuvmnR
cI0oLXV/TYf0EgJSY9rUbbk3yAy6LSWNmA6OwZN77iT24raJa8uw0wRyra8042ko
JHgJAzOn87zqLCR3jH5vfEkEYAf8c6brY5ZgSUlhgWZjkb3Pi0kpeB34tYDzPA2K
bOyTG53u3kkBYQe7ubKTFfBTQ4ywW86rBnbrwuW0Fcf0Lv4CXpb4znbYqzgLCcqV
ysqHpqCnWXw8uYtHG8tLoWb4KfuuSArE18Xv9CH9XFBXhGS2HJKPwDyahJYnd275
wRpPanXs0xy3oajcHaFhWUfmre9bKGVH6NZZhwcxVrkYW3dR7s2eAIJqvdHgSwNw
bftGwQ/LtJlcxaTN/GETqo0xBZxKInhCgID4019hxKZtw0ye4pa5GHhyM3yoCROs
NOi5V6plSJZwxv80K1Z8TNPujKX6bgRqcYImTFkUhrvQDwItzVcvlMwHvzZWgR1+
wYaVVtifK3OlDqaMrgUWd+4SvJg+n8wxQDFvInwm07qRho30VSgvuMb/9FN3C1Ui
XhranvtmHzdnvQ/Sl/Pb4FEbu30lNyelS0UvwHtjWr4bFetUnHUkU0o0C3dMmNbf
NYLg7m07QidWg/EYedr7v/8SzDV2QSRVTkED3sdGybUBaMtaC2CocWNSee6FftGS
QuM++o0KoF3EKLudhaiV8A0tI8eSva9Q1bpT0E/c0L+n0CzJp8uqOcwbUHh8/af6
Ls6T+JRgRDtwe8hc7alfrbpbS+CdmNrAuhFza7O6J16c5cgWD23vqvQfj1V/1XR9
GvYcAxrPIjYsIPofoUwYaxQnt6lmKpb/baW+OJzo1HwXhxKdlgczDmTPRRTIUMQl
UxoAqTf3kzmKM8Xfo/mfOAs1Dl5TG3qwog5JB7hy47tG6ajCmjN942zsvjP0mpUo
vqL9NOMQAyNAh5vSriN7mW4l/3OQfPbUBOVSxMGFwmiXpu+5j0gfYTRtl18vkzqc
vFeURRHlt28S+RCeHGjkahAd8PhXCjm2cFJCcExadILXcVJFL6sHZ4E4uP3I18eS
FNYDeBeKw/3LJ94R8RsSNln40/40TBf4j48Q8IcblhqgtTTvOSw8vF3MbzQ+k1VR
mXK3Vch6kZ1OjSJsPg+mf7Tupd9pzjDtU80dmbnotyLXNV5sWQdqg/EfavgXUxEE
INZcDGhG3bTkzis+X7OXByvqX7Cogkw9wvBgUF8KXrqX/Dxu2+LNgT1geX0efSxY
imHvvydXRZ2JzcsJ2eDGng1JURhrZkdO88IqpoU2yYqyhN7V9nyDjMgwtncRXVrc
ufvrQZhSf/cdO/ZKNlFUfcyv0BBqnjrAIjSBMHTmUGZJE9OAOfeuFnrhoARoNHGK
VAi3Y0BLFpnYtYhOOCpVwKBuJL0++bFF08IKzmdLnwi2e7ChjI8okwuKZ6ql6bRc
OKW5yrXB+bRsWpvb5MDGiiPAo5SVPTU82g8lVAFTZ4kIoUP55MuGizGSc9JLPKQh
3P4h89+TDdszdTeQMyTVirrJ8JHw6jC8pk4S6TG5AoXIibtDafsjXNPrKGMRuF+t
WR1xkrVBRJDxyFWbWhEpRZhPPbGesS+ysvKOpy3p5w8hBGpG3AJ59YVkLDnce1EI
w5SjHSt8t3r086RT3XSvvkKPmRN+9RuYhbrXKT45tU/EKy1xfNdPlqmhVTtbQItU
nyigF5flnpBPFv9sl/7fkXdYMJSLJPXFxwHXodDVcbRmtJwiz2uEGZFeASqIZePA
PLbIx+7FVXC2gzyDD7M+pqOb/1eu7afWKhUE+mgK9nUXyzCnQsSJLNNLVqUnLeEQ
Zkzm3tE+j0kELUJjnsIaCOh8uq6f9lSrCEQrDZKnbsIIeEwQAeFiY8lsFx4rBhh5
lLmQ0ouejq1q7w0NX4/p27JAq+VrZFRbp05ugAN9s50PXyHTF17S0tZamtVb0xvP
tmncatfOIpoZnY0MhQDSYfKMRRdLiT+sirqwhHriRvrpp/VVH14DAdWWyvhxsPDh
lfso85iFZHBOw0LOo1ygJzdASsBtpGl1Be/aeKlLqCvhCFuyRjBaALMqay31svkJ
zFO19gVeEvk7ApWz4ZAGeW4gf1mG8YvKYf8JV8cMMs3rMs5Udw3kmYmtrPH0aicP
FvSlV2mvZUTaTMALkYGoNvVvPGs26CScA8/1MM4839ggy2EZMMPkPt8fnpNYuyt8
6z21zD3hyzyVjuiBOO+r/jyWGsDGFBLLlUlauuP+sqULicyJI36POyl6qwpYDG4I
H1PzEObD4vpVLcbmQgV03na+gQjY5ws7oSJ8PegMad9M+xqc9Lt2HB8QFCh0LlXe
0MVzgBYWNoLo767JU2tAJr9f6D+xbKQ4SYbIPvTIk1jIW8YI1WSzCCFWxld0jTYY
sSHI6NImigoYaD8O6ae1DuYH2Pxq7W1JW9MonhODs/nIqQAAVmefZ673aBgDG43U
ueN1Q6nPtsxwfjo64goVU+uGreUWTP3z+rxzcPrkNyFL9yoarBkN4Q6D35K/1LlA
NGMFBDoPdLnBEijJ0FDNTFe9s/54+gsy2IhT/4BmWmsvNJXzMlDrSozYXrPOwJCG
dm/nSNauwyZ5wSQiLiWOYWA/CQTNFrlm1J+s2h3CpenVfAShZYXAgSJyfc+st1Rg
7QyuqRkS14ocaL2ICQTdOpS7WRUkLi0OeP+I+c/THPwY+98w1Fefca/EFe+B4Y2H
HNEsXzvxCKPK19HkEXhvVezGiL9NtXAzh5ra3vxH5o/wcc7KBymLDdgDFC7MB1z0
EpNYpsHkO+yMfJheb0l6mcxueXisYb47Uc2e2ppiaKExF3FvKBgN2l7U7038zQEr
zfsmuMTyHGUrz4cA8+C2a+Ke6so9Kt5tWpOMkICFDJtRb3BcKrjIvyFQlDeuaF/l
ZtSk7wmes+ZwTcsipT+f1iCfDgxOmHTpGbdNPzhKnsSfsrZJd9s+0lLtByvJz+HG
A3QGsbzKL803V5rXjcOqVgM25ddv4/of+FMRy4dCbXHa+kxKMLrb14Bnv/us+iiC
FbGek5i54ICdHL6D4Vdd5an3nr6JUPdznb9zcnq6WB/+c2WdKTMPm02SBbBopkQi
7HmqD7ehUIJBqPG1mArmbgJl6rnv2QzrCmCjNijwo6F61V35oGECOIripbEFNHbF
cgiTN/c1/OHS141ZNQgrMFa4738uo6WoR4DDzXwp3zyAaK3HM8Lly0Bptwj9BvJu
GbFzuh+gxYV0zZ80otVQLiKHcKzfsxVBhyHhP33mzAaAAaTfoaLjcaTNSQx37CCX
nPJgJayPpTkfO52w9OoLe+64P0VOggyYQJz3R8exdW0eyI4RrohEtbZ+sEI/S/gn
hhqVaMfq++D8e13Ydfp0Hkvj/ggEUUqaA0ATngamrWVgLATGywW7Bu/+xEod7CoO
eeA8fL7wBBWaedJQWzUHzpPRFLNUH2/xb4iJGmVVldOP9j4L8ns3FRELdsh72shb
jaiMifdYpElLn3QYiwcJ5qtDHeIAfgHcko9Mt0P6CesYoW5q7988ucn8ZCXp6eA2
GMTZ07dDd7/8OZX1C1SlUaNY1oNtvn+m4je+oHlYwaxMyuVORGqmtuCPH/ruH6E0
2RmOPUpHRTHwEQhunxsEbzx4CvjGnYagUsmTu50i1da6MgBZW2JUN0GGJw36sVcS
5B2FmKXo+obw1ccLeXjc/NoRUM5OOKQPhetCQ5TsxDRPPvoObBIKZOU/id/bybTT
q3dfGqQsLIA8Azd3SIciG1hpy4QLaQxRqM3PgwsMNmoFl+kEifhupWcwtyr1vg6h
ELD51k+ZpsZsINFlu1DzhdvFfPfDtbL4DfohAqCQHbHYmTF0LundKQyyWr167LX4
MU/XTabQ5dYQlv09LFXJt6lVOvqQVTN2DjmuGM0QINa7fB57cus/fH03tunotdZa
E0OEXSEu+JO6GmvHmVoFgPeSWjtwDPRZOkhJW5afWr4XCryhNv/DhvZ6hRB/zYxn
bX2BhNDO3rA4SCNMfZR+mxZP+qp33Rhc4EGn3tv3l3l0Zl03KQiyHKm1PsVmn6Sp
fJOwrk7OhpoQtuqW8gwK7qz+dpxn8ETS9m03UAFh1nEnawecFDQa8jWomyccpzf9
ElloItt1T1FJPs0fYmxtjr6rW3XPyqfBw0pPsw8+PBdkXs6DT5TANdSKn6q+gHzO
KtLUyEmTpsym8NeE3qnbOctOf87+8ruuFg+5K9Fcc4zoavcnsJJYMmCdNadETzPb
+C+bVqmvQodz0UZ1Jnx7WnuVe/YKrv9qxUfxjaPFC3WWfgtb4RWppmarZKN9/0pi
Ewjv7t1hJwuqP/MCv8YAf1JqzixdgF56OZ8GN2D3mpH6HojV6EHlFenSlyLnWs8B
obbvKTxx47D91/i+QJolXjn07rekQz79MTilBFF+hsCSTAo1V6IDrvr3NqEHYPjs
jT5+JxA614p1YEahjLZ5eAuCJZ5jJmeCqB22gQVAcPxnRY1rNNN5gAjP4l+L0yA7
KdrXzvHMXSNl/FeH4++zOXGXcq6Alx4b1eEF2AY9Mzr1wJnU/r5Dp8J8tFGb5njo
nqtIpkOjE2xGt5ej7ZJVtixtdERko/daeOxMij650bs94De1BrMNaZEwqUXbXahg
fC8jPAK8Y6cuwFXLVCBstdKNhaWxBUrzouthuwteYY9d8ylSOQjg8TzSrqefROLL
+siBTIxdjn1OOjUR4W+Pn9ScQKCtCsZ5lFPB24U+9f/difnnfppVoKrFd37071GD
bOAZTDA9QlkNuoSg8zwyO6WDDBKlzl/zaeu/EcEKAcu0bqk+slflJ16Vkxji/rh1
+Wz1EF7VB4gUc3QNQd7udo7u2yfJ9WSuBJpe1uojgrqUCd4q5HoxsK+spxeZ07nf
TY9L8lbDZfY5N/ktBhEHomn1ErJRBj+m5cDQekRQhiBI9HzUzSISoZ1/Cx99BFGA
U152Pa8H8R1qtCSwiGBH/6bkrb4fsN76XkR0tadQIdhAAJBraipD4ZG+fS6alz+T
jRDw9n8FJtKQcakNaeAx0KcaZoHYvxPJ6qxvIPs6cKV+4gKXFs8gqWM6Q55JE6A0
FpZly8fBfWGW/kTo2YPu9GaWihgj2x0IDblLBDJn45svj7OIxM6hOVxJn9fUM6u+
HuD1JJezkPxJeWOPWdPtuBunUGy0097CEPOgpSOpfUeQ4KWc3sEmKvmD52cd4T+U
NqlYVw8yQm7nzo7oO2Lk/3g0ccjwXn5B/nsQOhIxDBZYDOQTxJywmMiBdaAm/R/u
dtVubaIRFU1BeQbT4MVk4APqT+W+OsHT4aKfg/4PL7BQdz1c3iTPOdKxFCwTi8pA
znBaoQA5fDhNufdhT73AHINtUr1Fhc034+fGRUxu/0SiCVUbuNfIKRIiBTjJ9w+l
NLu7WIie+cqhY8PjaHga76o8wAAC5I9lFLc2QpXL3ggWFGYNOOOgZ2yA87fDBGx5
thZCLLeioHhyoalaKylAjayl2Dr2ksv7BDOAa92kyqVmqw+h18AD1daxJUcx3nKn
7qr+6uP6jeHmw8yKr47nc9GsLq1dVtdPpC5HdmLTeY5Hgkh57Ue2VFfy2L19O+D3
A3huHIrpGPvxaMz8VMOhWWybjlzCoRtzwrkIzQCX41Nf/U4V1mljY4eetUw2/0VY
RdTbMMsU0jcmisHXW2mN+mUo5MbZTv61FLsD48en/fcavnIoQfF3bFPnItc+QF1d
eUIIfosyLjLQS8hibpUxa6HCo4DTGLPZk5R0j0IATwGAe44I/VvPn1VKQ1ClZDTF
5xDScMwVuNXQ/t0fefBTeq7aapk62MtvDoEiwCV9Ez+1M+MDNM2F+aMMCt+WF0Es
tcSxchrFJUVS69Nzuc9fSA6aH5m/ofL5iMa6vlRipAeIZYomCvgOGhxtM9sejIcv
ngycTEh5A8ftj+8mJ4ELjnIdlHAF13ciACS75W14BgN4rRGyEsVttjXs1Ak3CV6c
NT2U/yYz3MpltZA8Pd9aNlnZEQ0l1DOYrqj044gpNcsMtR1Fa0ZoJvPUueClZDBd
YZRXx9qiyZ3k/m8TYkk8SZcDLNmsCHXS+tVCrZeGIp+Po1ZecFnAjObcfZcxdPEI
ZIGZteWA5y30wFDpytjmr2PH/YZ80GzNG8KLEE7NemOO4RDcVZxTCgA5ziGRSrJ1
IEotne5guhPpTzIuTOwt2y+IQnKTdR1P4r4nGpMa5h5nrm1QyfFJcC3BE+Shaism
CNklm0qBwgRHOz1lnSCwq6qvEb3+ZwFUebdD/i2ZJNSayAEOfShby7XzjRFflZoq
13tARm/G1Cr4+Wq47RI0LOZ7TncOxEIWwKwzssregnHHcefk5ifIqPZFTfJ5w7Mi
lWH76R6F+qBOiXEa+jNKhUp+ZmnmKCzEJBV7jI2mlSdSloD2mft6cUe72/hvmO2T
ye6YGV0QGsOh2mZrA83DiubyncnlESAsBztXeSGRQaMQJl4GuOUKgGUorHocEWtD
1mjrZVa5LiiPDAkDGFMfRmOiMCs4Nbi/dqxbH59C1c3lRjZTfToogSOK5t7XteRv
WsFn4DNhGFmbdcmeTxQ3A2qyJoc306oW/C/FU8WUjiTqttxZL1G1+Iav1Rma/L0B
JvwgX0IWckIR7xAFx4/12PvrvpFzBXXmz/Ir0N5fqAAnx/n+0mCPpxpndYQQ6ho0
UBv8sSl+hG2iNsCSEveEf0qMso2/bzh3W57yIM7gZ9EId3L57LyND3t8mFXoz4Ao
MOLlAW+9zzGpUFvdbjKtOlczekaKGwC89i+RnMU1XVX9242fnYhSN65js6ho58Bn
LjyRbINNDA4l2WSHhjAnm+B6PWql+b0fMKRJ43EntRwp/Fc3kjMfy12STR+jg4rj
SIUO346UD1KpGx0zoixFh3l42W6Fi5nykFLgoqWLQNWhhQNYXPWlvCyTZGTLMWKc
nppjGmiLiDDgglGlPBj8k4esRf+8yCdjR7fYZQdpnCW81ax4YkiEFQbjy87m2UIk
dGu2YiS/hkKi14mzQHrefgJxnJu1c9Is84V2LQOF64q42pnpwBfNycAQzeT28Lxw
c3RV6IKU+gW2PD4hxE4Q+biLatgiL3MhmOpHLa874kcFOdaqbLqtrYHpEZY7Pqnv
kEVzkn42aVl0Do+t2YIjpRnlVSp3+cGlc4SXXSWmbP8TE8r+xneOiS5DEEORfQOR
7ZkQBWYJsYHIqORMBDCXvsFp8TJqzxT7rn//59quaPaMuH5Euyf8auMM465Wrcy4
RlQXAStPhSechw5zajMusU8CeQu/bwQmj9YujIGeIzKdyVrm0Css+D7gtbIKRb4W
1NhvBPv9jZjxNy9hhewMVOvYSjS7Nawd9cNkz4c6F0jT5y9YqSCRR0xGbMmRst+/
Y4depn/dMKsZ0hdPwO7okl749c4+eJoa6EkYjrV9xDytuIlpkoEhKtSo9Vxdg+AB
4c+PtnjoS06rZDXjdPzyU/oGbCW4UMfM3bP9L3t+FQZustNk1dw5nTjiZTbSiXHm
oP47lAVQfh/uS2Cl0LcZmbOfBQa5MPWfQGYddf63BZpE1zQmqe3V+ZTZsRNAV5Hg
N+n1jRedbVosJvVbIpmD1UFHMXznNpMUJL2O05dnWzII0XALpzGw2nPRIHym0XN/
SQp4ZRRmKfWccc4C3dkeeULvrU08s8HJ57R6r9YXxuYNSWJCS/bYZ2OcQmzMNFUk
F2xJeDMDTwWCK0xfUeKGu0q6n6+duFI/32K31XTgyiBNmHZGHxkHpCm7LBBNkCDv
A0KaDvY5TAYmY/FmPrnAM9+HoMZEW4dkzyfpxUZX9XSzcekx+5YOYCyDFjLVqU+l
qUmDnKKdc/1XaV2McLKDGNJWBIPWWaAkYRV25r8b9k7SGzThvNnishWd8+82Ir3y
X+616/F8SVYZgiKEW5GjQd1lci67XWjrfRBHFldMl2RKXhEEiBE95LnRMkDtFXAe
Jvd/G/bwCOdwY126TI6ge4LYH5NAZXph/EXnt9eLDekqYJhPWyrVlcTqXyST3O0Q
Iu46pBBLZ4J0K3ONKjebIMIuXG4g+Jkn1lqEhg2tCTTh/y2VSdYkUU/z+SaUcHEX
mp3iEDj1215qJ1V1v1A5z4fsM8h66r7WENWd5iiV5hOg1N7SDfd5ceNR3Av1KqhW
KcEfPibpQxUZGypXgEFJl2aXurNvqBCvWjv9k+rAkm+r6m2ej9V5mTfAUYclegXq
QyyKo2rF3+FoskMqF7pCH60Z5i7EbqraEjOzebxD/PYcRKJTemIhncRfh8qIkEvc
7C0o1vMfTO2vA+C5agfaA6NpdNjxLo/+MKyN10twbkUYarXuhFlW4zOend9cG+Dj
sVW7O+WV1DYEh/31SAe2VnLODtDhrXeIJVHaegRY6AI/7A9uqsGdmMVYlO6FZNB1
0N6S0Dky1p0tJTUwZOgNYC5XSWlxHtmUj4Fw7n/ckqDkPWk7LjUpUYmGegShMDBi
7RSky8SHM0CgqR/qLgcg8pXjrS/GGLQZmiNGuEnk8gkJhDkjfdXt9ykZbFKHTb2e
L4Dqx7yBVJ69YlcWD0NP+SX50I9h07PpJI3HShI8K07ePegP212RTcPiJX6rvAg+
6/0cW53S3GMm4RkfgwADXTfU5FM5bQ0do/x5oKAxk7TVHzbsKA1TVSr+i0pwBA9F
VuW1mlKgSh3RvXISB0bgXB+u2ncpiwrtzUce5IPFQwNzymDrWB8NtfQjvTWYzoKf
qlM/LcR8+t1wRJGLbSn2HFFaHxRRzDc1EMMDZLTIhL8qTvQODtxuL2KNi5I2H05I
BdJjS//MR5V2cJ1cPS7akOe0jl75pl8k4QHYRD9+RQBPvy/5ykroC5jBFuAKMvTJ
qVjA4arQ1rPQxxcnNt7xCR9/owTOYWKfSAuswMRPD6wDIjdIRcr+V9iC9nuIEBHY
v9IudpwflpbSvoEn0Bx0wIqYPaewkhUCKFuGuomH5A4iLkSzzGzMoDlPhr1ZoluC
AIkD56WHFWXY/AJdab0CHXe3b6dIslO7mFcUfkTwjJ9ed4nKuqootsjOmM138t2m
EKpJIElkRAxyMp7I4VcfxY4ovK0h2efolewHgJ4FCyyK2Sts5wxVVANCOcCjPxSf
Cj70nx3GeE8/+5xOVWrDxDCML9zuV4AfrE4IiLG9NsoYf01fUvWQX4/PFvhGizoG
ltJidgDVZfCu5dA8McAtazW7bh5XM980r5r5d+bXqSqktTthx3ywePIjxPnn+1xS
asf84DKgs4EbJkPbYD6XvdXEsZgGwABIL5PL9QVCVbSu3MhaKUvtF6oN9TGXmKlO
BmdxqY+n/7iX0qwIptEdZzAkFAA2Elpugsf+uAVCsay6H7soWBTsudQsFwyjbdE/
maVbd2BFCI/PRBjrCNWI4jB+00XSm0br4Gl9c1EsYrcKA7QLWhFiiO6z4cGiwUMa
dFYUAjHQkUPcFrwi1I5UOQm2nIr6htBlQLXgHpoFRYSU0LqERX8WuCKOXLLkNHAa
yrZVrpSR4J8StJXEP5wk+v5oEXNLcqHvvVm2tE59n6k5S4dWrn0Wm3hQnivDB//P
72yN93Wn20uvs2pVioOzRGUP13LZvI2XFHg9+ZySx/sxceiPRJHQ6j/t9wdHsC68
fLG3ZcEtIUxi2SX56I/3BfJU+hsBBwGWy/ZfrUFRLm99NEH5jslVkCZSwhHG4k26
uuw8uIyEgmV3T6COxGL/FZQed9BSlbh95qsDXs5SIdzxWgNBa3ssw1OzHgYXJerq
sN7e9jH/hCaQ9dw5btxeJzpwnTvK8KE2JIhy7RQaSdyrxwnQtLxFO7X1anIhG9Jk
7y8keTwjagZg6Afovqcjk++nJ2yue3GrRU09PeMC+Y7PMKmpfD1p3OGp1Og36ot6
Q9qWjSOW/FsKlfcTKiwx30Uln2wihu3ONmf0uhY6VSoYBZAHLsahbYZSzSTVqDI3
FUo8eBZcK39UKH4HgoZ04Y3fGPD7ibKseCVz4N1WsvSaof2CQZ1skGUT3NmSlaRZ
IhNdE7Kx2FzEgZz6a9iu9T+Lqvq9AmMAsVXFmxBAOveh7ujZ2SCYBtdq7lPwGstv
DsItREtAkBuZ7AgiUPykSYQ0fCaYGGLn9DdrtWQZh64z5gBurRiuPvXg5dSCoKSo
XCYo3/CSAIgyfVAI0Wlyce6SA6PjjSdSf8QIJdLWuq9xrGESo5S7u5Jc+QAPGeo4
XT9GvRcUrfmQXnoWw+ZA1xWg60qxoxn6IyY/CwXemuaFK9OYkBvKM73tKwJCVx1c
85MZHpNSEDOeqksxImSIq4mNh0Q9Bcc1/BvzRXhgCKNBi2D6TlY+gX7IGA82KOka
QykVpGO8decNGb+AlJCOhL9xI5ZCleW13I787mwoCMJLCaDhSu3a4nuqvjYHH6ZO
Gn3Tc+dDIMGn0B9Tl1aqGrzR0vluLcpU2tOHHGA5+kkV0Kk0u4YC//UsIqdmjGSA
preFZRTvdkE9v6ltuND9SieXu9/f33zUySpzuG+bq1bwYsclnDrjnPBv1IpGZgpq
aoK3bDuwVsBL/a6uzWtBXyMTG//Hrrd70r+0mdqt1CTDU1uej0lAutwA+La0vtnQ
NbrItQQkDOMouXCykReuWOTTdT8tFQ0Xb4KEUAHU7PxIXGToqsp+nY9IWWaTggNF
Ynrewhc5aku18GdqagvV/wcLmzMoQ9kGKDxeeQvwxir8gEr75Elm7P24bU1+gGSS
DhZqzlGP6OauJabtT+aBV5Z107KYk6EdJ3Pa4mEVho5NI5RTq0fcOkZeJ5w2qrBE
Of2eIdbgZviFNEJ9XcX7qHnSwTTxVEqbKoVapvmOr0tjMB7NPtnTkvuU1L0FKK6O
cp64xBBTCjXLVeRKzhsD8ENajrYCG9hIhqu+Dv2sGEAIeax3+yC2Wp9qzrEIbt4M
YpzSerl40XEaO5V54r0vLeiBRjQA5MXMhsaW7EMWw+XiKVhACyKOlxOMdf4K8LVO
ylCxHvRT2Bl7AXrGWkDOCmxqS+19pD/ykH87zXEsrOJqzAGsUKFG3IlTnLSZvWVo
JqmTYBGBGcwU+egKUQE0skL1CvlGJ3SnrVsCmM3o2+Eic6kMDoJ3IUUPnoriP4bR
8ZZZMTUqHsDv9jYJNH80CPma98ybFrXfTNXiCh0q4arKxV0THen83NOjTFJW87Ht
gk5Dc1EfvwfBil69JNdlpQzGdOlBZ7q90h7HcENwaJHglHw8C8zArclxZCAsTOZ3
8caWc5tAtwNNLSggl3ueo91/pCBQAVeoi5y1QA9bCGHydyC5+gb/+CYVFHHdYvzl
vqCZfmYs6yQdXDI+Ot/Qk5ezXi85AWnkWlaIoWN/uIys9F/Xd70X4Tl4ZisD6IYC
5y4ybrvKbj+o4J8KxOhKAHTF6/m99lUsaUEMcjl6BTxhVKDfVpNxOJbwB7K1hMnQ
FDnoOdDZKEfOsb7tuwyHzpHrXcb9nf/yMBAzKrrajM+IGlgO7v2P359nEZ1Z3ugb
8BFx+AmzVmP0pP8W2SmE//h4gJjkVL5UM6kgRIg2ELrJKiNXr9vmtL4z37JpuxKA
fZfiEhFYNd1PokB+InrSlC2R9duE5uKrj5jhh7P8ZLApdED2ABUAZUdPDOs8PNKk
MhcZxxK4mOlWvIK47R/Vsl10sAAA9Rqr5xMsgfOJDvuUmqoH5Ufjo4A2+BQonJtr
4Mcdfp6bjHG94qhtqG9DUmpfDPHHw/c/tRCRqXmMD3nqaSFIiwpqZPIs7Z1u5z8I
jviifkScujLAck/s/872odKcq6294/LU3LFpuPfSlxIdnGtLQ/kWapJ458GR97/l
BbI+pR34vFDmo4yqGc52Qes+lTUcFZxSi/VnXg/AA1v/ojE0ZQvcndBNakdud/iY
jIxD3hrXwLakHJdI9fFo/KPmHVs823YHWR18Lnn4CrBFnuZ1iXHGGqoqIP//RSNA
98KlYBI9lR0PcsCSXIox1XG/ghI1mlz3k18cTkOA9Yr1JOM2/xVN0oxODakJH2Uh
ZYZyfNRdKE0ZcbTdzaQyM2rRrE4z+dmjciKPyqxzcvquiEizE4uE14f72pfqxPff
u4AVKRXOjqlwbsuOMmNOzXs2e9HlbDCeVkV4HhkTnotjcv+77M5khcygPXpxf0vi
v1j/+jq0FpeOMixWvxE+cgxhqhdoHAykuHlADqfRup375jFm5l/N3+IUVqgjk40Q
XQkjXiAdAMuqe4qKPWXsOIdfebXciu+MCH5uJncn65WdOR0HaclGZuLah+raOFHZ
BijZSBXx3LS8fipiHZP+Q00arDfE56ASIPgOk4UZJh6iIb02HecifgBsovASUY7P
KvpgQZ8caT+MWNLLo5c01ifW+EWUul/vEXBmrKuyplD8gT5yc8Wd9EX6GIq9d3Bd
ETSc5s+1Zvuzo76DQueAInLAtYt+JW3sOEtCfvUqiSyD0aKpok+mw09h4YvHGW+t
6FNL/0qqySq4k2rGN3u/zAmICV9sdSnMAJK7JH6gfn0MVLIl6GKY0eDmFk2qROQX
W1sfgwScdVxX8sm7FyjOAzxlnRG6PVSA8u9+EcQEZ2yfSqgCsuoiNaXUEGezFVwL
mCREOPTU+a1xMU8v4Cbe8LuVohZCEwOh+nlxVydf4oB7C72N1NDIsmx5ZyO2A0jA
6jLldLTaishc/D9lRi4W8EKJ1l4GEgwBaVxIpsBKrob9fglgpzuEawqW6A0UjaTO
1L3Xydt1Ej+Aqno6Q0jI9aWsca2wFSSE0N2u71ZcBY4V/H8Dzk26b/ITtGh+2YHH
RkHdPrCeMuUmOdczkK7YpOPHTByKztmOUBs1x8Ke319YvkNBiws8K+o5hMQXKaYe
Q6pKm5SfamDb2XykvwyJeg/xW8/qNg1CHTPPGB35ssjfBzNrBinCsKv+nJUS1AvT
HkxDwUX/uZwqa8OTyC6AYu0NKVWKDFkG6M24Dh9BFDnHC/KNlq1snW5Bfiq0FL7Z
fyfWFJ5H4bEBqt3xEtTqzVScDY8gRemQ/tJP6vAz35V5H7FEzlh6gKboVnZga+Bg
IA00Zy0Q6oh6Ht4nELkl65ZyuwWy4uN3Oa1q7IOcDeQ5Ntnhby4bK/KfkE+jj4tL
QcE4k6TipguI2SOnYfjswUPqoSPul38GkBjLs3LG2xPaJa99qY6Y7vXGNK9KhXbq
JH0lkCPy84JOvD8Mpfhso3KJpnB/KfZZoAitki/9pbCuwz7ffoOwsoqPZDl4n9jr
73WWUNeiaD4FZ6cgWaN+RUV2Dez7B0AtK0duXlC4LrqT9iwu3XPlAnY67mMut3Of
wyT8IQQEDlAVOrQq6m+bLt40oojtkz0ShdUpXQ//4eGkFU2Y+9pjP2sjj/gKwKpb
TwV1RMR6UmkU1Z4mF3e41U0n9NwpPfKwkGYm2wX2HqLmGutoWNuzLVoGiYTNz11A
0uk8YUf4kCPjAN9gDbjCXoA1rP+LhROPxDsLDd2pKKKPnkIix6DVCFq5DkWkG5PD
NzZyIT9F9nntT8IY4UZMzjGOqYwl9V1F7HqpIxHK0XVzaoQfs3y3OLhvt8BEzh4f
mjBE1bF4gA6qiAR+eGQ4T7Kz2nhLUqmQ22/7v8Ra6SLDUuzKJvig0W15Z+mydRMR
y80hiUhspF6j1vf9QYy81wHaOFptM0Jd13Q+57z7lwb8x/7I8zn7Dp8e45BMAWXu
2hJYwhSbVn/zY3C+ptZkcLYhDcW0qs7aNdDFIbyvmsS8SADzUBpKRbvJEgUYyTnH
DUjhwb1QMecnpyQ7GymM7RC0uuxdk11IPFtpgJ9hWpF3d2+bjhAKY8AtlyuN1tQo
VRB+6/kw5X1rnSAqTN8bwDEEnSSmZBcxmtVDsw9pDOsgdJUCZVUWC/a7HfajJL7X
GqU+ae9wPAKPRxrFje2SSoSR6m5mJddBj2rRKCeZy1XZqiQT4S/YQ7Wnh6XWDjMO
YV+/I0ohTPmb5EPtOqUlWqhE08sTKuEdZhz1mVK8ghNPXRQcR0tni6+1kMLwfkc3
sRAQpq53mTdROzSgtWkK/LiyC0I/RrLXVFyH94J5vSgnZv87NE0NZk9CgNK0L+VG
BvsIQ3DDpg+xO8vhyVs8c4T0tBbhtVVRUJpJegggP1EpHanIE1tyABWojGJ3d3Yc
rEk+s9VEbK/RdO31FT6HtUFNwlWolSufZl6kJZJ/FcMx3RXOiCcxFemkkq5JiEza
/NJUMNFVz5ylHjv13CH0BB8kTYqlGIcRSYZFLST3KRVvgKSn00RQIgBRbAcvZeC0
wJJ9mFBhWbGQvIjDVlpZqlUGvGqBHkD7GNna4d54tSfyfHOfcJucP0EhdbQfw53P
4E46z/xsXh95h1UDP7nefEhmYmL9Etjrm+dPGmEsqnr2iTdF9HV7d4UBXMdt9d9W
KvSAVSZpzB1UIrGoyrFRQYRLKONF98cIcXDMxn0pqyp1k/HJqU3wv0lfnQOwYWbS
dzgEvLiBorPXCwLFnBaCQEJmavqFcUYbcRTTK6gP/ztBH3KA6wwgHS8baiHK5G4G
IKS96xmCjR+K/Nr950RpQny5PbESHAqbKJPQQLtTp8Tg9PgaM3JPEGs7NXX8huIN
VsskA4+o8cYY5loTAND/raSSgrpvSDmnopkqoT3DLIZb2Z7vwcKyRLlkqPkZHg+l
oOsGoUaO102d6dk9ea9LTrtOoRdHjzF+rFaw+E0QQ8GgkWXodhCjWS48918mFPRe
15mmQlBfrmL/3mO5NS1XD0r2oKKP/nTnfrCSEAVoM7lTXWKblnTTqRwH9yr9H2oA
OVd95M1/aL9enaNVCR+H3mmevr2BPYYUCsV80XzlRar0f5/6ZbjxuCkFvd89WYCD
O5Dok0XSre3OeVX4u+f+C0XtT/HteXrOsJLrf2R5xZNIPua3nI1QIkgv1Y73+Pea
vJoHtoAvflFVgDP0N79ESpatXnm0KAArfVGiGvU1W4fs6cfB5jEeacwTTmq81+IL
d9tRU2Gje6D6uAQd1rtWiPlwwfvjEm8ngRB5rDnIakPev7I+1JirlEaInoxU1KIb
jT9a5Sb7V8AHUhwecWPQUXsQRn1FdMekavUre0xwM3+K4t5BB+7VzE5LNSeB3fcC
28kIcfdEyEHUEzdEJfXUD3LsGEiOOUYamxlejklbrM08B/ivnz9sr5EaHDVGnF1N
OPgDTB2n+1rC5d32jXp7PyGT0jxK1nNg21JWzQ/Nofv8zveYzAmsi6kCPIHuClF8
Nz4oFr14MPMnnCiHYhg9vx2FQ3/Xl6h9V2jlRfDPQQrQlpckEwKQ05vDWVThFU8q
vHf/j552TzTIGGxbJFMgLWGYNlR3WYK3PwHTD08YykqCiWqW7V0QIm0bnBpZE+7V
+u+Fe6A30V3RIRhjIdH/cW/PLfLrDdfuEkFXHp16RF3AWKTyPvU0s1T8DJ1hvXpT
DheMh17ZEseoobuiPcjOv6eBEqdSOfVKUagr+ddLEHyHWy75vcsatx96vwOILd0b
m27ZuSmCCYozDYzocTyt/mAoAMwz+FOkqXaKbBAhg5aeAw/rqlQwFd6ezIOtOMAm
XCHuV6MU76m1zLF7UASwS46MhgxJEfUgUFkqI/xnoFWdpfM/TAA5kDK/nYO3y/tj
xMsd1MXp2Yxfzbpe2Mxhs90LsHXRI1lvJKxFX9mkDol2HAmHWp/hRYRRu/iubodn
6Y+BUe6rFteh3kE1KvfYUN3BUxzKW4grX2GePCDh0Hhu+wrAWVJ9+obr7p6AhjFC
Zeim1O+1nhdfq9buVmRsh6VBy2foZLjZpM0WfJy9Qk/F3xVQrDIYr58vVLK3N+cy
kgC9qvDaSHAyE0a70Mko8UrK032Z4qF+yXJARhDPpiFp9xQksph4GbqedhmBoSyW
stu4ScD4QO8CnozD5gLrwFs62+X0kkc2ph7qqYK+xOliYXi4o/g8xMIuNNwltHSO
F3UQTVp04bZkFAUXtMdUQNhYbUSP1jbeopyU5ZWIc6q+l80J9A90ZFTOAKd3942z
VtUQ+yatDtbPOaLYoiGcJ8pswc/JG9S3j88h/RKVNSbSNrgPw2hQggKTOLARrmHn
HBXo2q3VX0S3oo4GrIKv63ICC2XUCtMAdofats/h0pnu2EmFr+cNcPrOrjCCgGqm
wmPouS2CyxOzohsWhjpDYwNw+ZH/z6zeyP0a1+6Q36v60imn9vv1V/QnizOKzb75
doLiKnuWZM/WrvvQGzlivx+iInIQj/LS2ArWxRWlLt997XitIC7S1l0MYlyJLL9U
ahwyhmLuSJAgZyIU0mxaY3ONrOCEL09J3XEFWKRZh1Dcim1JCjEiatveBLlX5G6s
viGffmLD1A7u4dM3ajlgkjmGjnARoxrctdPkFtEEpjCrzNzdpiMgMjjXMnrPdmrf
giuMBDmbMq0eJpkHBZybouUf4MMla+KcYCJOIAvz/aBeEgxdVjZKFSGkqdIsYKVB
7/qvY1upQ6T3ORCUupihJkErCLCVMvLUl4M30f9+BOSELiSiIkbvaBt4rntR2rVb
394HYNC6sCAR0zvKsK5Urg5AcT8eu8Vwrw4w7/va8scPHNsnejLYR9xAqi/t7dKb
eWc7beMPba2JVxJCYYYRJpJTGAVgLzqEUbeQPDMSdntsZqLJyLepSyDOxt9Lg2H5
YWygpcfIjwR1yUlvQdXkWfOIqsR9QhoyWxloVQ1o1aFdtk/NvV8TmPW++j6wRNjt
7z2yy28CwA2+Xg8Jdyzlbe/NEJN34Nl/95qyRVJcV4A07FMKist1QeRdIBwfvU4Q
8NfndkHNIe3MRov1wAgqHIPXkLfV8suj+5YTE1Iv8ampXy73M5oyehav7YQQfTSQ
SxAB5pKePiNdnve1Skj6Eq3Wmpztyy7Lc83hq5joZrFjjyWZ6aJhbkv5BqJe3JJ3
r2cKnl9CkYD2W/z1DW6MeuHyyvQF2iXTMZTSP2KK/JzV155ty1ACRhGMAAVg82a3
eVkJMmTEBlVAbUYZpHRyMrIIPSyh7LVCiaSu8TqRVV8ZI4SdPypiXtbfYvoTqVo1
hTwuUTqd/JnDjW9qz/ONVD5SBBWgBYUtqIOqhw51RlUf++3nqNNLCLq86x6FGeTi
3RupsNMUNq9+znOV+CoJC+3UePlBOR8m2v9uWubs/L7tnJy5iyFt7R8IDtz+Yp7Q
Bt/QvzweK5p0AIUsrzuKUOkU15CxnhQ8bfGK3FOsiy9UW/uSifJhtOJFg6Iu719g
5tDcWn8aaPRGEJuMBAEu6lHDY/vW9S+DDtDKRh71XdQQhZat8mcDDyxZqeHZgff5
yfR1DMusx9rYnNaSm/tLRipf8SIMyso5PRMbWX9PZuji/NXH4frjfVvmUb8brqj9
3v7MrOU4O8T5RUV80yv+c3bQWrVfgxlxbliyRqJLDNGPE4Pa69n24SacLIadMpRH
gT7V+RMsZlROqfgTvyuOtfyOwT6e20qPd8blm/svJV4v1l7F9cUvb9EuOA6Gd9Gb
N9Q9h8S1WXlSmw9Jbqk18wNER0EgrAKd33m0rAsT0ioSbkIBr5Y+1Q1gg4cxBR5b
pCNvrARQgsi7wPPNMCjMx5lJoxLLQn9GI28UKGThSjvw5QwgrJl+ueQrDTlVQlaS
hhdQQ5erQoTOL7ted1IxWY4MaUtk+6uf1jr5d3lLTMRoTWSKuj/INiSQjAGiLxXS
9ihQ2SGYFusLwOzr909GisK0I4hhQS1k8H4mT19uG63EMxcjhOml+PaBcPoElGhq
fwogU982HZyQP2H5dwnAo978kJ++XPtr+O5R8Tox0QGtQsmGWtDC88APzodOwq/g
5OAMVFCaSE2wmfkS+BJNxcrz1/i1NC+duLl2s5FZ90P6MEhNWmPUy3S1UzPeNAc0
iBW8KWuNkqQSw0f14RhRZEJQ/DxzTvGyVOrGNpEqwTr8UB5bd84QdNV/prpztAMf
+E5iyh87SW+VTc3IwX5ay4O83NS6Pv5j8q7uuQZFy05+xP7K4w9T11Vo2VxS33RN
vdXkxSEqD7IbZmhSrNzgeJ+peKRaargsgyFkxTwk72E6YnrTmCp6YKkUL8kZ34P7
hs+Z4Xr9xnz0Dlf9/KkCXKP6P2bsH5zile4Hh57+KIUVdh2qNJkRjq5Wg366EIba
B6xMfnkqk1HdCsLaTltDbtq2DbxooDRVPwTkXslkreVf1Pf+yGwBFNq0Y35BVLby
i359KOmvhogIWYm2KZLYpq6J/IeP0essd1l+AjHn5KTKBh9UEEbZ2sAUX5s3biOy
dyuhnncOTJyL0KY5ec90xurx9nF8Nmf3pjBBtw5oHraZfGR+y4rOHaCRYHrN4P3Z
DoTwkZQt30s9KVm5Bvj5dh1T1GtzEERwJ/gnnjdI/ZdGLJ5UED7Y3CNez9QB5KrP
pt94T4Zojr7DdA5IplkgvNHAmzFa96fFn6pWSzK6z2NdGKwC/HKxf5SPV2YqQbZd
om1fLXqsHlsZTeBms01YFLxJyDYTguQckNTAWi0sIJpmKXb27W4e5fwTthMDM808
xL/ZB9lg1GIBVMAkxhowlr9ALZeym2x3BUXLMga1XQ2LaYJaZumPZW9/8fcxw/nx
lpEyYq7x59qFbCfQbzGXelYeZMcYw7EfCo/h8VuLS4R5e9CqHvRGJae7tlh5CKkU
/kQcoPniozrCXhQfHiu6l0LIJWlDs6/loVhdEpwaeE1hiu8NcI3gyTfXwPMNFN7y
Rdl2M7XMZx+cfPHSoTIb9uQL+SLYP1eWyPIqWVXYP4JmBludBeoPvVvy/Sfzsddd
23+KP6lIlDYna+T9f54I4ZtVnsVosEycK47Plwl3JccwNvORK/NIkQm7M3CypLNI
q2IdJis/pudVleGP9+LXKnf0D9iVUktuMDfj+SZXYEa3wVO9qFisgyB8hUm89sbn
6tGEd7Qos0TkCYYWhSQWH5MMxz/vBk+Owa1Iax10kde3Bvov5uzQJez2+gRxG/0b
rXy+oBkm1bLwWB9V+JNxnpnkJ461todguJtavNk+4M7FaLWneFrNL4KJsTpaB8As
fgYAQ3KbF5gJLDDLIxFw5JQG/vOdTT/jLBgvTXCQH4OVbCpgHGrEYu+g4ylwPXKp
hWHehQ09+7a5ymudNqOihFjTFYT3+H7LfTtoOa5ON1XVFdTki2vCU7S1DOfEtMiH
+Y6iE7Okd/O078ski4wNufB8gLlgW7pSugPMX6k5y4a4pjMiZMLN5AQ2DJ+hgRdJ
K3vu29y0Gl5bbtxQxjPNPATBVOs248D7dHbgv2lRz7FWLsHTI2aHHjm8SEnTa9z0
g3BVynq49gEZj+I7uCTeL+zup3807/0p/1b9B/3tcvVcaxeHPoTC9yX5JED6ecIV
OlUgM04IKg8hoNG5nbOAOcjWAzgqDhnc3DrdkI7hVuybIAr2Lur/7G9pH76STByK
W9dJWXZxySq/0Z5d3VUmzzYjr6vL7cdcReELzukgSyJFJrAV1Lo8NL+VVEYyw2VL
qfJhrJPmAyw+uWX3YHAmPW7IQD6s0q6xsgIMu8eerZiY2+K6AHh+WS6MH4EFqWvS
4M6zer1Ysh4O/YoofCBPqGPi8smkMPqz0I8pnu5GFzxQOd7asiZNMA16OZ8uIFZl
djbaaJ22EtOtH9l/+j/2ovuxqMBwg3vUVf+Zn3l/CZK18txM+2YXWDXgSoGfS7mx
TAujDALFhPO7IavDxoBGjDWAyz/4iBmy4FuQ2KpNS08rsPb2QKf1Kg3BmPuOtRBv
vCuncF/HqI3i81zkG6Km+M8zVozJKVWkaTHtaAYa5WeXKLopNK6dOTWgCBccZRcg
l0298eoQpG+YRxBbFxWvfU/0OJ+46z6dBkzQBJ8kOS4oP5VmKjLEq2Wi5m6gl3HW
Y0sYxB39HexdzXV5E8DmOlDRpvwyv/vTzR3tjtu5PHVWVanPRoslv9m32GEqkfnR
3hVde/IZe7R48B51fEaCwSjP3Hg8G5aJmgm6bsLJvbN3UlvZu26oCFQ8PTOGShXX
ON+5RatT2TKLkyyBOPNhncGdm6aSi0VogS5gEGIPqIk8/OylDkNEYlpVR3ZwsR/K
78SIYdxdHbtnNuKmaDayOlISq9f6gieJn+koH3cXckStPwzPugRHdSFCk1wqHtzf
SVnnz2aRPAz4N5AMlPD5ohPKkw+tsgw+D+1x2vOWFQtHp9musgfyBfS/8r2D/Ej4
DGGLVbFMFfO8BU64zNpYRyuo3RKDnVJXTcekgtvFe8Xx8AFudeQXJcLeTPf6E502
bcHjz8+jLY1EWIR5WO/pZHv79TE1rnkM6gQzZuqr0fx4MYnAgJ6itjHQvySBQtfA
r2xgltmcUeyUHdWZayt70P635COH902lF46iaMzG9mLi/8A2rq5eUsJsUA/GqIbY
tkR6mSTmG4Q5UAvTP43DtyT0KjKAXK89j7zfshqi4kx9iVLMz4UzFi022u9Ojy5e
neYX0PVHyNP5+sVx3RucHMJJPeuphyIgvu65bHWaDxgKCIvP3WMGHTqzkd5sOh5K
v973Eo3MuSZ6vlLek5cIUAzAMCxh7IiRP2gO8MP+p22huRyaOsAH58EiKRy5q2ly
YADENq6x+5FqxEc/EiH1aNt0VmYMTqoCAF10zT2+kUUF7v+RbJIxzRmZqfiH4Vkg
eo1rE10PwwYeaGOB0DZHTaDWn9x6plOWN6w1UcjZWi8VX+I7XCQIi0W1bEdhfLeY
K2WyN0rav8lmtS7if0yyF8w4cl0gNNDpAks8qGJXhZASa5ylayVCxkqEQhYUeq9N
g6v9C2FHC+vdL2xaQw7baVlbJKEroB4sY/BsseFmi2pyRN7VbICQsFV+gAQ0kQwQ
nGcmHvQSJbYP5kNdm+wUAoK1lB/zwKnegHXSf2pJAx6NM+YBpNwboPEYUBBfK8zN
IWR0FcwA26C+CJppWKHW4NogZ5leSKhIAqiWCB4hCOONXdqvXMB0vX+RTeMm/xnp
2L/47t++vnAcI3zGrt+S7dsqPb9xQ71NE+Klq87jXbKLiuGspeXZUrg4B0XhL1FY
TMpeBzeITJ4QqzBz6BJ5+SVqOulrJmUFwOJlmwKH9PKrNRdSOL8nmkU/90lSTFmW
oZiMCHy5sDHGyX7IeU1+PPHd0JOMYa+NPacvkrd6Nq+6SH8/2t9I8ut3Fdwq13oA
whR320B1TCoMIgofhbVKTQapyKi3udasJN8cANqXDddzADGJeRAlq5syN7+vOqWS
ATgO6SD93XxDfZRQnir8ZPTLa+Y193G/MtRgJsKlnLft9ce8/ize8CsmKUzTkwBS
cJ2A5iAJi86t7yrLQt0rvETPyNon6QKSYP48haItclq5UcnlYsOUCq0q/UZRViv+
t/tLw2YBS4ibiYv12PAGxfuz7KepFsICMkkTDrAbeLKXes2cy7mCp8gduWpQM5Z5
HIzRjMfvH/MzIQXXUEaH0oDP5MRiodbNsLxpyZSoiKTphUrxvBUL6YyK8C2Hip7P
ZZqUpLGC3IPesvVfZhuH+SRgXz1r6tjYWTemZs6RxfsMsbGBYxxEaLws4fKcezPa
E3kPHPNUH+1m3Bn4PgimbohpIezPaqJPgSEF9wN5ob0Eh5KZ3k4oA35DKVeuqpGx
/JScEDsgjfHvawuyCctygd1yur9PxdNVolRT+virv0NIQ85NeSREftQkYZlySsi0
GvUMvsO0F/ijaVcSSPVzD6SbhLvideVKIqzoLOpfINid9QZ3KVlCl0O0Ozif9R13
JOjZN7iZ6ewGcDToxgj0R/fbpuLM+EGNe/oQKEsQIdB1rEHim9iOK8a22sCodJvO
kth3e1FlgfFg+Bl3oFGT75Hg/wUHP79TPc/JzVBQOFeWAYzJZZK/tRoVQlB+XiUu
wrofEdZH45Gln7ikVCR19OKutuWI8L7CgX8WL3LCBOwJY8+LVctAN89BbvRQGzpT
bwzPJmRAs8WVYIxca/2dJGXAfdvYcyE+9eGR68FvoCHzcL1uZeWKr4ETN2cXOllr
9TWhTNHTE5vWuNryR94VkhzYktYu2O8iDTMTicGiyfEG48hiFbPxH7gnOtb+0TR4
jwp7asGWjYsDk9EZkGOEUg5qSK6H3MWBM67IDRoNh8ka/BHLDkI3WHuydq9kuEdw
SP3LB5jeIz4Bjov0TqboGEUhegqia0Gq6+nphgJ04KsCYBVCmekfiWkWBAGuQhKl
l6wl0LvL2RakyrdJdPBdYeXqvwN/C3MBbd2/FsW0KbnB2NZpRYBx+oXrv1mB5JwT
8qaZFWEHthRP48juF4YpMZNQirsHc+qxz5OsRNIfjnpcG3P4y7DhR1Yq6xRrBlqg
s3wEuMb0YzPKfoFSXxkUJ8r8nWXKeffb9zCfH1Dw1NPRAiZvTDVkh7CzKQJMtvr1
VH2cw3j0ESPwwOadgHYtRuXtjv34N2wdI1N4L63bFpTo+8jnDH3VhID6ubkO4t0M
SQJw3dEg5GkIbgwIG/z2drbTIgGEyvu90WvuppfseaLPkjbsV2NppgcCoEyN+q0I
1L28yTboqHKudWqrW5xrdI40HLVAS+Qmp+XHYsWBEk8t0XEccPPFLcadDJfVUvA0
h+EGKEMA8MI+pkOKAaX7GkNx8k+qOCw2fnkhj9q3IqQb71t712Iq7MqQzHtEBNtz
DkeISA4jro42BUIqKCP47NuQX+4Q+LIF6RbtINL/w6HHWvxyEKSLoCKU5r+4C2Uc
SlWeZMa3MBmWA8X5Jf9XPbivDsCjYn11a6HBDNRhuPUbrDVv9Qx7/DcLRR7BUKTW
qEgNGXWo7uI+yVYc8FsLPItJ+SckM7A+e40GTX6d4EvJdbJy51ep9SFaekMEUG54
mALLnzB/QxIcJQtleeFuJhCAuM9rHAzP9BEj2hHT5ApRzlmJQ0lm0R/NdzgXDWQx
76sSqL4+smsovGRPxXjBhSmdm4g4aI1/amL8kASmpSMdXF/UMpTkSQPTH0RhjaLd
1MrsO0vePOXbPifLctKZxD6CHU0Wyf285i77oBPOhru46FExpt2luvXq0UrQH/H7
BdRdj76RStNQWukq1QQFx+LIWLHQMAuYX7zXgFBZYwMIyMzjNcQREjMGR6llMfbH
+7+XJjW6DLVrNd+V75rW4eWx9ytF4TTtPcvav1ilw2ylnYoR+SE2IBQ/22QnFZ3X
Wqrf28FyF05ZO+H/sk9Kg4WdvM5chxpSLMzllr+SOH4OescUjDJDpREGWpLGIvcr
2QAGw3evPhKFlO+QZe0YMnUnB8s52Qzrnfl+5Uutpd2kfphpx1sPZYieTXPNCcvO
CarL1jNv+8KecaKp+nMrVFdPyNBG2CUGFKASa8OISZegLKi4r31utKFKwlfQ7dWh
NRzNwB1WjKY1rS8LvHCZu5EJ20Vcw8fWau79wasy7HbYJowAkDYUHOdRI1moW13X
CkmfUDF/r017cNadpdITke6fjimhXh4m++5gjOWsBLebIUKDtUZ6mNWGw7yBf+v9
Nlx5X8Ayt8tZWjMincefp0ypPd9p73c2SbBAsN+nl0gmpITRVOgjmHsikSAfq5lp
xSuENC440uVPsUA4c6aSo5CkMum/wQUkivnU2vrZ4yhJh4ekFbzZEJLzZ8njcu7S
HMtlOvZ5pZXt+dpOW2aP/OJR39GZrJe6BJ1s7062TQBkWdW6Hf08XJT0tGx8MSi+
yauzIhwUPysm/PY6f1sWD/tM18EO2EDjtEt5xOH0KoqcVeHdgXwHlIiJe9XZmu/F
pFxYRowgfQVeiBpzh8FQ6L7St8//b8GLHp/Pmpxf5LSj9nofUfhHNaa4SSbYyYfV
TSg647+nGdAoV7LPpmbzeYBDIAO1hw7XblMLO+jXYaRuHcqbMGbnIYzRlXauaXop
+99MpqCSoUyJ8ShFaAV4uQHFulixKPt1nK6PVanWjJQWQ23h4GSLTl2joBjIspco
5MkxLTA5BnZUmDWxOk9cGhotDh5ibcH7Vv/IKbBBnuN8PIvO3mqeAJ64AOmkFxNF
p7Qc/FP2jG3r0L3bq3RHB7uFRPBNpWCUBrUIdFIs52bCYGC11beO9lSLK3pSoiKa
CZuOkvqAXfhutnugomn80SpBHecjU3WyzOcdvRFTc5pi/Z0pImeSbjZMW6xUKw72
MMkPz0jzwxhPCXYHlMCC3q6S1hy3GItI6dRlDNM3XvLs2wp6uoGf2MqmvDSfduXB
Qm8y+3lYF3LdMZoaYj2pJbGm7wXgpfFJiey3RgrOd9S4ZrX/2qnyZ7h3xWqEPuPM
Kv1iwKinW+dlqw4A4ALOeR+C2PgZ7zkJojbMNHAld2wAev5RKmK6Klt4cDVUF4fg
yVUSEwFROzgXk+DREJOtf5rV/FJEYXk2QYszXNdOZ5TDkhiKhY9/+gaDNdscfrdr
2E49qeBc+C8mXdx+oMvZUkWHHavPx0nEna4YgVU6Fly9i9wVbY2wS9lDmjlPcdzT
+qR7Q5EqPSAELHsrZIQqwQ3QxICVltHgbCf9lindhYTJNkoU1MCxgJihPiLTBOBN
Dx6e2wh6VHQMXgavzGAXmd6BMRanxjQ1YUBlEHPCNu+mfv9CUUF52UdjOYDCHYiQ
tqVkPaPLkod8hprytBWz1/lN7UD8Z3NDasKrueiAZL/l180Zu/rCN/DbdjpzFixX
dcSZ29QKQKgeHGhcYuTzO8/1ziMe/JYFowD3T6YxgJ/yeL+89Jx3PAOD22bQv8NI
mk1osqwdM9rCl1qzGleVBZ3WgOTJAuEIZYXsxR9mSlRx7srXmaXfAVq+f0Ue/jbA
cUBOjVSDCCV5flMuUb5u1TDtdEx1ETrTNXg8ZCBu1kX8qlLApPjW4Xtj2W2wUxjH
uI1zu3XL9w8O1jtMzaAFTEj9y/1SIiyS3nkHl0TaLP2NZE4wwiAjKyd56XVu7Wmz
w/GybhMeUePwMFlEwoAbUo5jm0C9bKOQER34XUuelyhBdZGTGJMhqfWBpiF73YPq
al0XB+ifI+DHD0Msonx2GJjVazpsbI58AbaMmyDzrgdnDqPUGAxEfE4e36qCAh5P
OqDheM2PKAIrRirozT6zeV0eh8GTgy6+32PNLZrXcmJc+jgigOY8k8Sq3GpoNSUo
lOgD/cnTs6DpqAVcYL7jTt+UwwNPxU6SHVu9Ew3uspWC59WPHjdpnWmpyB+w8d/5
PyqNUUkF+fW3tjtXvdHHEklUVtjBzjKcTS9naXDGK4OrmJjUgi0yz0vLWm7iaoBr
JYgC4U2hiReOlszqcGu3qgl7cC08GGUidkf+Ytz6AfefbMjiZhnuuDZzIPlPNlYq
/59gklmBYaEiYKACQWqLAzDpac04C/9HY6W9eRvX6+IFVuhud1p0+OUJiN8juz5P
NP+KvNzjfgplFKUuQWpmZJaZBitFCYeJmelCpTymovMJhSVfw/uxRiJZU1TKFN8Q
4h32C8odk4eSahF2GvocL2SooPK+FX72FYy2SzvcVkYPsYUHI50rTYCs+LzLGwYi
ph29PdPiAlRVJsl3SdAf6ZaAbGtveXn2xAbDcqV72L3etDcPdm/JO6q1jOrF3JJk
5Zdf7hmYhuUsO+ieHUpjor7040hRj9ECEeT/HPkmiTwjUwr8RyP44FP612Qzb5Q2
h1/kXuBkQ2BXpg+BMVljI2+6zepE6ngrwLioxxVubfU/aBKl02Mr+4ChiQH+k1xG
4liltQh+feSbrDrd+sQgefICzsxFTNizy3remASQ1gMPhHqvWFsDL1ApjrShbsHV
wMp3U+ro5SdJtvecTWiNAq9IbWIRrZ9gh4+G07N2hwYm39aYP9Z4/hci+7OFyUru
GrEhwj0euUCNjVkUf2GpuFUfKXHQknaEkBRWEYUkDNFpLb3E1v5lsh8XHCaFpSrp
qCCjCArEfJBty7C4yAXWhSccaPRFxFlBZVSMx7olq9Aw/PTGWI47hFbHTwgawqg6
Aq7E8mZek67uCjjwSmwwqVn1/L2VVBRbCj+FTNOb84feP2FFT2gk4YjcQn4SS2/+
f39ejM4GQC1PJ3yUOa9DZQ8YBU6n1nlHao1dqiR3MXo20CLX1buWqUzH31VhuaVN
EFxlmHCPPRBPPRb0OW+lvRjaC6FCOdvN7A3+Xylt01vlP8V30XgcrdsMD1cNFdeU
4ZXgLGUtyb/xfGoLy5/F2CpnFjliihvoEC0qsg5/wWD10PiiaPrsei8uQdBUEO01
drnIceXEU/ipymre0ZuWyT0MGO8gZp8gqc1b6jSGHKnWtvvAtkZiOsZ0P1EwzLhU
/pLfvA1f59+YKqz6SelgXgRcGAMOQ5VGYjOfvihdq5cuhEDTZ4Bl1L3+BmYV4qYH
6euaUwlSL/uSv6p7lZoGuWdeqFNNQnpC8drbf0j3f584IknEYD8hNzuyLbwOSZ1b
QjCYr4up0avC6b/Mfh82m+xfXcoFsMMnw6Lx/gb77icVo4kmzM2HNy57ZDWlWp7c
vsdUvelL6f3AE2FGCHEL9VinpMHirgBU1ixWS/zheEmpfKpcn5gxQKAgkpZQfucv
uKSFpNqLumxyXMuezjlBkcU5MDt66QnxXZSaGL5v/VULMPnJhuFWIM4eRmNTOe4j
abA6bqaWxXXzj4dg4WTxAhcSfmN4K1umz2eetqNiYwhioMFxt1PXYFhASQ3HPOdE
hqThKFo2smbmTgLiBId41Gwv95TWsKq0HRSD7tKEkIT2k9rbTPJ52ECkFJbaGt9b
dd0hb+68hS5//8jvUaEzBsla3lLuBgBFzm8BNT5g4gBAgOL7HcEDSUAvPPrNJOpi
HVersTkbP0xFa63N5SUpBntVFsYI8Cgh6rog7cs/BryWPlYfF6tD1FQr2se+7xy2
tJBqc205ZsE3duTN4RhRkqLGZzKiJpBluqvcc+GLT1Odaj1BXvW++Nu7eIPOkfl7
j4ZK6EizEQfh/o8E7Sx80Jkyfpt7wXFOcPlvZmj/spa/W9SEj6SkTMBI50r5Ryu3
xifTsZZomnkGPEga2WcRjgLKn8ssZdCXcSXIjZehznRWOWbPedX73Jmc8Vkn0PHi
9VFJnNTabExlsMYXIAzCQ31Lcysh/Np4IWpOfMgslJVjKi9VI74quLXla/VXELJg
uLm6EoMB+EdfySAUr/o+AeRYalzYumtqSddeuXPGgXRKi7cmcQq98l6aV0isfQiL
4IfK5uEdulRErCThPgbmBJBE5gtgfSikeWhhdqMKI87GsKc2W21AHriG2rCD5NSK
wwcPyAgpEfYzrTNKV4SMZJy5CMTrKUag6TlABFEVRl62wHfpT+L7DwJC0jLnIQgM
Pw7yM9ZbT7EG2WlWQnq97Ka2s1TDHd1MwcU5dYkNT2tsebB+Nw+F2+yKIq7VMyeC
eO3gDaRAiefiT2d6eLl0kp2u7uI6RT6PsKjBMqKQhuRU7tnsqwnWsV0KtY3iW4xT
lsILQpETfVZhGVo3jp2HP2d1nKIMurVlcIeDubxNHGjB6MX9q287KUQHRRgZnevZ
0N8Vb8NmpTHw+iUiVcc3gDD+XPf9VaxIkMrgqQ7rc0C3EjCt2xKQNGkIWFP/Xq77
Y5wcaWRYMBFqvmYPRDLrHvzOm6VS63HS3APRJ8LY1OcJ7UQoRsslwb4uIv5V7MJA
1jRgtpqNhbElt5cpO5O+lnqbufylFFiH4Qjr4m1EpMy4j3wf+TIhg7vQEiFGFtEd
LAzNt1RQyofyrUurdpbfZgV8PUhLuqKrJA5FvutKWUd4y2LT8hzzRKxXAQ4fM4TJ
1crl/god0JPdSfXOFwQ/M8Z4AVRWdbtHvnVDxwaYcOVRACiWtdGvvTe80eYIn8O9
D4sQhUnXTR4ku64p2OgKdK13I6DPg6ZZoUGxDbFOUjsxQOWq+mYgUevu5k2bF+w9
OztuHFzO3V2VTsYGuTq3bISdYsh6XpZvFghcY17GWqUGIrn5Wg4A2utQxYVBpLCz
NE0QcyfjuwVUWeL3G/aE90H0D93YwC6Sl8dgCM9LYWztdFmpFXXI5ysViFVzv2Pq
/NAGoLiElXuwsqaASmv8quKpEJA4niKvYv78wy7eHGNDxAKPNPov97taRq6A/bIT
BzZio+t0KtxMgE1GBL+9ndeKaUt7V0lfjdOpWuqTqosLA/xnMu4vog5dJRAo77+A
KJHDWZXx14/ORXpAXRidAn7IH5IfhVmjHQ4SoHhKE3qilZ28g0KD9bfD/qfDNx00
SnnbF85IGSxa/Wg+XGrKn5Npqv8TZLpIdXqhkS1WGIzm9jC0eV331hJAlB5XNk+n
1iJVHim7Qe0qOxiroFqBuMF406JpdHKe7jQOyP3m57rpgJae/IQa+iF1c9uHflhB
htp1yGF6kn/IxdhSp6sT4VHHJG5fH3xSkqvl++AAEZbwSBhcMZoOoJjb3LpIXFxs
uar1zpATb9t9bUph03uJ9klBEeBXU7d42FOHjkHZLg+WFi7wzA0m/pNI7z+L+AAy
F0hTsEiJj1/RG9nmXRGUldWCoOS1+DspSc/W6epYd6M7JY7HWgFkUDPqcpPgdAow
8VyXN8s4FV2pCtBz4pU+a/nc1mZKvoWs1tsUkxQOtBqToblKQcIQEGvcJwVSGuYo
hNW8ZOvYjeYOaLjQNK+4W+0k/JfRpfqOTaFAMwqPUu0b7A0dMbfIGvppTtDYzr5B
0T/IBhJKt4wkMGGi6E0I2k0+KkT4zGSQNv+Nvmc7DN7gdax2LpA6ANm2tiKsDArH
XimPqHq5Tx4e4bJqTpMiPIGZ3j1HUbeFvLBXV4cnKBEXTq405tVDUrFvl8Y2wGF/
7tDhgZVI7I75j9ze60mztNLhzABiodM4ElXOJxaVCvgefI8sqFWgWGlhn7PoRPuq
MLbGv3rWFla7xaCyS7vujSn7divVxuPdSTTnRUZy+qTTjou0+84FZ1J4K/+Ze6ju
U9fe03aNhpdzCHq/v6EBMrHjDxUVmeBz4QQC4Mz7KdS5FkAC9Efeidmn+Mml0m9e
z7m/aqJ1DTGZbNAeeBWd5lQ0OjEGUkbJJ2eDAh/8nYg6mmPQJjQD3WGl41phTOM/
kp+wIaXXRzNw+N5DQIy9zMIjXo4qeefQXPyZPAclXjtEe3A9j2PmtO730PQNuYMF
APIrXL3/G0xkSs5rwA2euPRNGWEEEpuvvIH7264bLkSm4clXKJ8ZVVapgDEJySVc
i2cEKnVUyygkbKokAu2VfuRkNr3Q9rzvoA4svjy4edyZUz13DhZoq/lRS3Pprj6d
xukPmDB07MLbHGs4N5fLersPz60T2D5BLsIe0i8arcs233uMRBc4109JKWtEOsbX
qtGw0eWnIki6JLukT5LyiQn3i3iLDpdm1iCBlK5fMe4XyndJd7/4pGe3he5tdLEv
AVzJVKwbyqJoX2DvOd4HJPsbataJqWLdHBFrzwQfVhD+an9HhhlOTvps0w4vVtBo
etLB3ETds5hrtbTDitcySm60oLoo+hBEwIpUzQTSPskIfTJeTyRMtBUAX9rGHANF
8lZsibi6aP+ChxYVQse0SYcY9BrHMVM3hbCSN8yRAhK59/AZMUgc3/Ulozl58EIc
1s59z4Vh3lrUQmuhiazK241+p43qhmc9vkwMxpE3JQ0rqAhLQYd5trzZ74AEUYrz
QxVhS4GB6VvxXu5WpHxpril/salUz7a6qLXFXrEf4jRiIVEUt0zcL8DLEkMOwG4u
agxRmxufuLKPsUfrFFXjK/hgruBJ2rm2LAFYSQprTseL/gExRu38OMsVScG4uWie
fpKMfU3pXr43ZRFW8p9oFESQcxbMS+pT40RH625ZcaqDwRqBvFGnoNEqRahzNOns
QpnEqpMBDaNYz5tZS5laOtjk3mW6+sxBdZCZD5crFTGhDnwizcZbFpICjKVytESa
KYnSS5gl48KFyEA9+PNIkwsBwDciGe9p0je6QoRUS39c68K1vl/qekYPjAwuITzp
du/oB+0jBPqyaohMRZse+gSc1EEyYqXAIqh4EAjQRS9FJlxqPBaVFKCUl5B0GT1K
+IF/2vrOIJLLdCTemQngUnjYITAeOTw1qD9nrVnJmv2Caq7yLmXMQOBSHlOtg7rZ
2oysEmFkmXNZOriC5nBQt7vgRvNnD/WueslKo47QLujnVJ/t/9KvBYtQOl0gYVsC
WXYCCEj1R3O6EKq2XhTGWgBF1S/5PwUjXGCS0xby1P7qSI8lObLwxRucIj7+7120
dvofGMTKu+Iah9ZhySavmN9qmgPtXU0CaH+htQ8e5krwEZoFaoafWqIzcDLwanmA
gQHGqQkacaTT/n6cXN9c2lNTSx+S2POgXCxWlWmau4KDEc89ygiFCdHKfmg0z20t
Eu1XOhYx3l1zhgfvAmgQrd0WiO8EiWKnIOigT1pgF/3Dlh4AGDzNzjITyxl22AvI
C3itTlNL7DZ+dKShFDPwzTeH1FJkJW4e4wd9OAnILmbnOqSGooRaRc1cbuG8PNv+
mCkLRVg3a36Z6+bV0MA4ntCsfFWvJbiupuiZY9SeWxhL5FmiFue0X+WItvEuxTsq
YpttScmLwCJC42bN72Q89V7wEDxSbko3yuKCLAC5Ao+F9TwjeJJoLO6yV4EW9O6R
baUO5EusVyEWKQFERGGJ0idq4zpwbdyuysXSYUP7bH3Y/0HLdiEKebX+a3nLlVoU
EUtwCbaUQfkt3UsByW0gbv4rGMSoKVPxuNLO7WoXXpvYSzdKLfBBOB+BPuyQG7aH
0gz6s+X34L4Lt5cKIhs25Yt90TuDExCmuS/2stZ5ah/cykYBVlHRsTE4XCgC4hYf
ertVzTu1OGG8twNxMgiRGHxT3bq3vPDK4k5m01Tn88MnsArmqSy0NsmoHjyrPtJp
PHD2T684PbFzoErEosGV3JeyoXELtzJUDFrhLAEDY75akDiQ2SpzBKmiTxeZjhJt
xWkBcwpkJxki+Ze4IEoFWl5ECV4fY+mWY9u3pLYJyT7IYqMIJLmu1leq2EKZWI3x
Cpm4XlAP0tVDMYsI7rMXh18v2KrCN2bGlYm0lVKZaCNNkpzumfJ4eOVzn58Eiyin
RF+DXYbr7pBtWvmZpmeerdLjm/542z20btH4tcuWmnubrKypq6MThTEV3daQyVx3
WMkzLiUkY8f8F6BCsjT+48AnwAhcpuQ0gL6Nn/RDHASqgksp2ZIuo5uape8v5KX7
Greg6bje9aVPQ2UnrVkFHNaub09umZp2qZwJ/WbwbPVJQBV9+F254jl4wcHkGOjz
LjBfFuk+iMXaWJ75IOF7Sowq/CitkQ3HX8SRdIlXZvCz+oEY5pVBE4fgYAulWjVu
upEGLth0UfsQoeO3F09zqN7VUifDIH80mPsJvfugwSxxlmZ+wxf7ALmzn3odTwrc
XWot8lQgVNH/Jghiw6IscuZeyHlBLE4RSBqJz9nkaRPXs7UFP90LUtUn6BjqYAkd
wwaiBaM9Ap9bsjci6ie14ZtKu9i/XLx7mqMgze0CpS8W+eq3zmZho4O8YNTWOMLP
JFrGo2aZavlGaGtzJafFjhBbbBoP+35o11f6Y0FJk03oYaakyQ8wjb+mrp69egJQ
Dtc69hDcorNOCULplG70FmGxxKmGuCS+fvgsbf1vbfXi8iclyXTXpT9z7wOivY7q
Us4TYmVSq2BkThT45g6W5bjem/TnJUf1+ONZnaH3AJoJHr0LJEihJQg+oJyyQwlQ
q1u7paGRytgW2EdRnKsCNl9pxRZzepmgxIDAECDq0c6c+rqEfP73CHj8wwMpEtbU
DC71ULdVHZYeFB/uMS1+9Lj42Z5F2Db932F4h5Q0s14EsLi72GAo9eFSwUgPh6sw
KZq8+YHVv4r6zgC3R49VlshdISTYg5++Uor5ct1afHypNJNVjDORqc2z1xFrrC1X
V52J9zQ4gYWz4swTXELYjkWdJ2T2jz6Mm8MQD/BH/4ysspedOcprpQdtD/7mSEC0
G3tefYy/62ba4T6JAiEnSiznfO9144UXxJeJJv4NCkbWKgZh97zf6ErF+ZoCQbj8
w7hWMTtuPJy7tqA/Mzwg7RVO1fb628nzAhRWoNXFnyT3Ymbort6sofBC9hjxZ3FB
6qVnSYQsoB3ryutCVyG3PCNMmjBsezQXF8hdenOdEmIVhll2TkxZzprVdi5Dit0k
psZZGA3+FgpPuacJGlTiZf8yZNvxkDIB91ykFsgAk9/aYzPcnNycsBKGDNJCdsFT
IgSHF1ylR3QdItoDFW2TRCDcGfVbFQk4tIQToLOQCSL1K4Mccr5DyoxjGvSNZIvt
bpWNA2/CNzfrOh929Dbqz3bmGAKQw8kcX3BTkIQKH88RypFYwyKZkNkNjjoF/X4X
BR19qgS5oDJeyVTHeppCNLx8ZFkCWK2+ULZvQkWXIlLPf4ef5IPS5h4kk7ND6GJm
dw0JO5nD033KROXO1Kmh7a4GIA9XnqjMUfTAedY2dE7ocFToE0hZvpADarSXpENg
Jo59eOyy2YCiRoic28sOZsIH7yTHYUVoArzH/f7lX4ihpDkXDx94zxGQ7OhiQJqe
tmcmbrdZoqz+WWqTktZnBYpBYNd/dUovFOmPpuM3XU2g43Hl93a64pRqsiYiAwYY
0CiB7yPqp7be9C4i/YtTvXtL8/oQdFBHLrb27PXjRiHwgbL2VJRqQglbNYLtkRk/
z5xnXfJBQSYMrIVJo/kC/palAjmvXHAjklpmliu6fMPfjXNg3P0dTu6E2C2aeVhP
WuDzoS8CL31CtX4EPigPQL7iufvzV0qa43YV0UlVhg6p3p/wTtorjF2Vpjym1lY6
9dOk/21VizRI1BJnFrct1Ql06l58eWn1ce2CX98lazFGO8r8ezWtfuNrBBZ/9adj
q25enZMnX0Xyy55akdwTCNzF5ssCoR+zIw4ZalyQdi+lXXURWBb+i6/H28Q5oh+M
BkPI5P6/uJHU9qDqtxNjKMQFq79/0ltfc0j6lGfPia9M/n2nfLydF5wL6bKt4cKU
aEZ5thXX9nQCLY/V9EyPTDQjZTb8RgR4Grzy6T0ZFOYLYDIc0YpcDv3fFHlbkVqR
lkDa/kRAFTfDjoTcPiOn6NiIr4qv+C21uWinXs2/sUIg9B7azzFJjV3AftU7LEeN
HbQGevO0IF0t6VOwPt6BCg6ECbDj08gpZjjeU8yoSqEomWJIPcvOS4VYtni6x3mK
7DkEtI9voFjNGpE4bi4D5+5vLPBoGQe9/BcWiA51+A+QOo9rRDdkSL+Pw9fcYT0W
8U4vfzy9OYTK2GZ65SR12bD5kB4C5SAg8/jkXKaGLMI59LAw7EPf33x5Qm8wPHNN
QMG0obTA65dZJu0II7Btku3xo+kYwGAdDU+Qt5a37Ny2+eUORSs5jX3c5S/iYr3a
Fb/BznPqEN2fGkmLvN3fqNWC9ll90we903Axr41EatIiWMsaNxdWJICfG4zS9NFb
l4zfc3poStzCHg7aDJrY3AMXooMSh8KkcLwQtCjQmUNgWNtJPxyw61LJdViwdE/7
mlq4is3BwByg1K/6JqxG4zOYRoLMHlBctZWWbcQrJQ19yq0wA2W7/k3IfD61Ga24
y04ni+J9OIBi9Hi71vUfmDeWyaKtzltsqc+eTMdV/D19RLmM2m0S0QoPqHl04bb/
a7s2rpXhfg7FaG4iBQYKYNIUuGdc9gh/K1xTLbbrgjZLLG5ZXe0pCfAbPpImKS1a
9NGm6f035MV8rsS8RdsCoiVHEtz+sXKY0W6atNdqO0C27BdKQodn8BFD5gcdBuZZ
BvzU0WBstPO3GFnMOvag5BvBFy84CxopclhGQvT5xxI0EYe/WFsFiwWcFzWjC4Ha
5zBQUGAWP5p0yWy5QMbSg8M0q+8dpJwW9b2GZYjBeHWP+Hxdlt/a3A5biz55rbgM
M89/T5lYXv4FCh7PNvgHzHaWBkFB5ZM+GkeCb7jec3LXtBNRV/oir8Vi2VJSJUrs
A4PXzYHsN3Lm7LMpiiNBRqpzZsLltzcjoXtNNRguPdp3Ex1Re5PITJHz6yYYc7ud
keKioxRr4UTpajvR2xjsw3o/HJC4c9gDNYfsYFqIkU1NgTanv0cJ206mj9404b3U
U9Ufre9+7ZfFWLmzG7P7FI4v/Ku7TQj2HRHvljsmLSU7kumbBsBuL3r8lHAwK/Jg
zr6LE6N6h+XRVfVpzV7x6dbe8Yqn92okk0YMiSLKMAvKFgsuaaZD/D6pt/BpWN0U
dDAg49IzfR/Phc2U/Ir/kSsURPhCLpesi9QzYQNuV9FFfWgnt8ymxHXrjaYvHwFO
SCeixi0VWSrpNIsrzoGczwIyU0Q4jEjiVRqB5mVll0PCOL11pswF4oVLjKuSdtoU
tz7G5HMRdTD1vza7YDtgBObHbElSsADzBT3g8tBs/W7zjG1y/ATImTzFf6SIjJ3I
E5XzQ7ysn4JDRabaFVs2PDoO3Ek19JvJj6+nMQopvpAiN0uB1T6AXbZKrJz+H5is
GVD3Gc4F3OuAuFn/8Jses101xuuaGixVi2gZvixFmU9yCAMNxThSSlmNNGpjLeV1
BEzmnkA+lT79o3MOKgtka8GgbPl+INnEr+t6UxsyVcXjfVhPiNfCuQjQ8SEsOWam
degfFrvoFP+WCOW1JLvIUsZAwkEPXcLfhgTg3mEfJbIBdn4Brjy1hNj+OjuEaQ6N
IsDe8DDhX+Vx4oJDeU0b6b371JRrQHRx3JuJQACpI88l7q5EEnnL4KWazPeusrNt
tOhGN72g5K7dHsBqhGUfK8clnjptG85HM13L+Pzed1/KvG3w/gY46OLDKAqe17ro
twIIuZjm2xo/d1GQtEHSxlXXPRwQAPcHDyDJB5Rq/HIVbRgSfQQo9iZWPhsEjkdO
uHsTmR9X/hrRelznKF7gjSY5ha3dLJFLRiVAsAEzXsgY6pR6h1TEqpZmCdOGfEW7
F6cDGZFhXe2X6ngZEeALNmGk//f0A5J7KveALUVz+BQBrgcPKOaOesdTrfsSW7V4
1RFTuytiR5CnA7buBruIUgBihhtY07feqQuQg2mcJ4RhplH4FNQ2wZEBs5fWI82l
ZMHf0kaq36gxDNJsG/eJuiAHOzfPiqu+x6mE+g5POcgEVbxVjKI2hQ6YGt55V6wl
Q0JK47m92D3q4d8HKhempGH+Gb7KqNywYXhi1c3kzU0LOEQiisArpZjtvpIaWAud
vnqp5o7lv0JP9LOzFyuxu63WS0bRQ7RfXoqU7j8FK+0/X5TkgPabaRMUhe5ErXdU
nvKk+3D1c7lR6AlgQOVsljoO0Rv332XqkalQ8qF8zk/m9JkAoO790pF26uENnNTr
eMorQCnAJH77cEC7oiRm9vKq8+nyC+FTOUkMQSXxNMcT5a9pYHIgCQgQk08F3G9j
bxZvWhW1NuR0ohloWBUVyeBJZo4tfrKIuuSBS/6IkZ3jJs32lX7fIMM1XK9DQ4AP
n6BLBm5GFrq5NwOPP2hk4X0nI8w15X02S9MnFBXsj6BBXs8JBJz/jyVsMI/FuUX2
SLXlhdQHnGYw16BktemWDcBdf91nGyVJIpk2OvmWfGbTndLPXE+WTKANRUlJ21XF
FbBghpCZSFnhWIdZUJPges3OJmQ6cfvcsoursk+3nRpwlG3LofDMc8+OAstQ2k8+
SfAc4glq6PDnt/qpVlZHka5YV/9aGCYfUZKiePmB00854L1+L+QgY5L0bssIEV09
v3RHsGBWWBaPXQK+Ym972WNzhugZ3S/50yyvAsZeadau2CMqq6qH0PflKKdDv/lp
eKLJ29wmHNVBVdoAA77i4u1mhNU2+jIblHnsKBwpKEFTTMCSokYBj+yqFjVHlLaQ
okwsEjfxw3I/2tRzLKv8S0v4CV0LVaYDfEJi3gw2E/jvNAiF4zR53jceyowtIgBd
7I8cOpat1nDLIjOuJryzEbOZh/VNcU5jkY1lVDW4kZVgZ6n61bTVhDHP/60JMJEV
0aGYhGXkB+FSCnAksYumTIovEqUliscgDQJDicLbt3eft39Cpjibjendt1+MNzX1
8SSHoxhv/N17vYB81dvdSheLp/KCP1POBqvSbvqJlkzflZOiKsvV82eCVTgSXfzp
oQlzb6nSb29gjWuVfOkY9qe9aL+Hvp4lQUNE9Whb8Kl83gLZ9l4vad8LzE25eeVn
5kqwGxmowuifIOU71UVWwKR1NAaSip9Fc1abf9C01EIjHHWjdxnp58b4A2yFna+0
H03ErC81JCDmrHElx3Ff/i5Lvyoc/kYH8EognzNsLdqvhDQQr+jmGEMQqqUm65Nt
jbLaM8zFYVfAP3iBD+hFkbGCeFAPlcCABe80wmCjL8V2HqE2srbx6IV07NvbeOjm
Af63EH7jIwJpzhZq5IYagFVrgojFelFtJSzBz1WN2NulSHcuBbIBiOD9LqvPZdr6
7nHwl+6itEUWi8PI95JAj8RqhF8vKw1pj0DXaprcNgIAiiTc47xe/McGffMbE0na
R8hlOywY88MN2vedu+hbnRXOa9HIsFFZvdscHnseqDbM9xJSL0jlngW7eFF/uBsn
H2MdGskg6VnFDdlV/3YlLUo9uUoZyC2IRvPdY7PTZS/il1YQncWZPxirsCv3bSeM
Jf+ZvsXGwj+7ekILNbFPp8lH7YWqfMZUirEDANTIq7JIuzayIPQhtWUev9Ypt7Oz
iEhNsQ4OReuhu6VP6Q8C3aFDHqzfm74GFwYoMt3H1X0ergPA1ggYDevS2VExWof5
N2fcyAh3s8AJmirS/jMkaP7byQZyZ4ubWxhit3V6TYwKo7E3kgtsT0KkGwnIn6Ro
+OFJWEGsQHqdLo32+SGF2PbPqgiX5oD1Qsft7m8yrtytzuRMYf7XbeHGwqXpoWor
Yc/gpwFFUVUWewFMOs1lKmcPX8X9zzNTuyMvHe8htZ55SHpIiXoHAb9nNZYfeUgw
YP1Q/xERUW3qu3NJdq36BDT6bXWfzvg4xgPF573V21PSitACsE8R0qfSPN5eLsUK
mT7GVaJ7KKWGzZ7iT84mhglKvRxCWbf0exZEF8sjW4PhmIEUtmPEGra+gG+RXHmy
DTlVQXN0jMIPzE6F5VtUQruBRU1usIehfsRXcGxX+2ZvIIb/WTEB0Nsa8NesxHyZ
seIEYOwxHgS1KME0OppabRoKnywNLbSr9rHaZwIWNMdZFDaOeH6XPtUIsPhOYjqj
GoFWJy9wDv3o5JhzpNjTIgqFcJAC7reYsFWbO6l08xU2R4TfAz8HLRoJ8PM71tio
/nC5uiRQx5t+GO8q2ovmFmKBR8V67PR7vJRXRI996p5PMciRMPeN13KuFy1bQIII
peIuAvsn7O4utCl1n8oetg3QsOFER6TU8dPs5W/GhjvZXTzW5VIXdqILz33ayBYu
gzOuWXFIhh6b9ypoPlQY1zSKl11ivolSV/NmXyApIYIvJe6aaPs2HGneS9eIcIP9
mwrVrrOfuhVijaR9Ih3eUq3r6BiBsNenyhxCM/jGM0voozXN6QfqtZ68fv4Qk4S5
iHFXAAe46vYt0VXuFxyonWh7jP6WFnWmw3M5Yw6NF48MnTiYAe6cNYn1d6PzSJQW
9mOHNFYTRicIQGYcGTpjt8msjkLcjSRVff/zXTZHJZWXxtmJbvVmE/m3QJ0G+ynL
n4fz2+xeIuglVGDXTixNCAVND7HL+4I6PJ0NA0rKk3PU5EIpUvCoFXcazfPqgVUm
9pXJ1YBqiw5eZ5BiGKf+qjNljuRsT9KTUXvVaPBphbdaA/8kPq1zQxDfPk4tTnST
Y0CdJb+vGS8AWWLWArUGIgvXy778lojcxF5hpl7Gs9xbrMuaUc0sk6wEoM2BPiEL
p7oGRSvPky2WrOdj6XK44ugOIRK55ef5aat+fNU3PCGz54U63+tbvXBiGtL//Fmy
Q1VJ54lGmvH1bMT18zGfkwqOI7WbPauG81cC2Y4evNLXqOfvq8wiPRz1w9Jbwdvm
LE50M0d9Nfum6pFaHCMwLeUSs5P4weE8xeXllQozWAkH8crTYJTMHPXwbOn+stLe
akrIPxwht5b9PiJBibIPFntpNQPyjUUuD0zewk81Kh1Q+s1D8lXWRtqH7aqP4gOg
pDscMlO59KW6wlp02ShSVcmKIYFfRr2BX1A+spn0Frznkwyrz7ZWstEvdHh6xbhj
kJeABOcF14FQPvo6EMUaV5hm87imKGeCSEEz/CWcP6vrIpq/jaJj2ggMsiYjEKMm
E2/pg1gGxdC77Oe/NCAT+Lcrcw4r1EGFz/5NohLZLR/PEdfrVvE0CZa5y6nQcLe2
hokcoo6mBclBYw79SZMRvDNKW5uQ0XwyEozXLmb02peEB4+l0hQ+mqA707pi93cY
rG9c+AJWAhKDR9u45MaQSd3+ovN0cBjsA3BzQ17GxK1qs2YRgC/j96O2DnHxQwU/
gBFs6O2E/ymA6eoDBb0fKQ8smN3lT8rnOQpBdXHURjFMNQ9+ZaDuVjM/oZHmIxIt
yQpUlfPjw72omA45e6uhe3x9y5rETBuZvK05QjffV5CuCYmJYaWh4ux52jItC0DK
sEk4yKUFvSLItVFkLfJeHvs2bEvlla6qfCGM0Q9zY17vLTRjM0CCAPV1sjg4iNuw
2GodhkCmNJ/1edXeCq11ngJkRKkRtK4l1GIklCPs+XzPbq1AcpGuQ9KodkIAD633
twwPOOn7rljA6Ex4XMBb/OO/FOSifKQvmmYJd+yEGDG1ayQmbrsGV7w14VxCChLG
LYoaEfeJ5yPTg93vbfeDCvWTft+FYzbHmZasINM17hc3M43u0YbM5/9eQUAFNLQX
lu4IxcI2bvXPuGLgFV5Pu8EwGS5XR7n8MybguySBxktK1ErEN8PuBjPvV1RxZzcH
UZNMET/QSyYH4MYQNOTk5DM/uIWgwf4mSiBjaiNYHBmqBZDafJvR07eU2ocR+TFg
rGdYsXALUJOQfcgDwstbm7sb8fcMG+azvxP++LnZf68kzWG522vDQ2lQbcp+Q9Cr
bo2IClN/VQpFZFu/DGnOaYAECgrGZFF7rMmvjE0RjdwFb4pcIVYYZjAy4SPJzenL
zLbFmVTtyt9iqxZjXrvqNHNempApJaswoq4oQ1QF5GlHgPJcLLRoDXlbgHxnQ6hd
YAVlpzOJS1ywwDKLk5o6rvBGiaDTAp0yWNO9g1zyNbI4e/xEO+xnOpl3pBOHPLDj
L8GgPpnWw1bkIT6jSqlqB5PnexZoxdLSRfqerWQLVQpEa4DN4S+gI1cv+v5GmSmJ
x2xkDdB6cqvnu1Ujtj+hKg+ghIWFhYg4Jbg1oXO/MHVowtXMW4uLluyqp2X1sEMk
cKrKPXo6qgzrsfDC2k6uy4ai8N6GScSrFAkw76rHmkBhZP92JFs9oKJR3VeX4aye
GwGk/kvOEhCbmUyqXEU3QSJBdXz0t6p3M/gdb9WxvkqenH+ziSpnw55+OK72qr8u
tS0MxrSeXeE3D3lEYn8HCQAkyus8qiQMdX4fJdRCGPWwlmcJemdIoqHc3pgHa7ov
3SslF1RJ5nJII4arlLyQdpDDUG9kacnGqG+2UsaVwQbQ/jK4wzD0Qu+eM5LZj9xj
Mp9xdZ1ZtJzl3k7HhYvbxDxyB6WYBbmhaKerQQG4Ltrl47UgtSPtDofjLsG6It6u
B5y2QYMlTRFRdLO6X4ilhaBdYkuWBtv25irwgzj6qf7APWaJjM/rcPO17F5oUM9r
B5QWLGljQ8oxm/efCjV52aXK8uPRiqyzKkJhzH0zLkYDHC91uzwgRqfghZfg8y1g
mPd/9d5wKsVPUI7qSPbBHSGVrOBocrFlw65m3kpR/INcgM0jtBBhff+XtnabSv0c
unEl6Ro3T3ZHWlq0rB7f9aXM1zMwmX1kTmuItvbRtFUK0GLHzLVI/4j2iRoHunSL
+wCHj2Fnbfa3UWlXnnj/asyFtY1xa+1w3AQp1+wM42wrCiE2OEz+zF2bqA/Ios6f
thIRip1eTgCKuDXjavhcWD4/Chi7olMX8VG9qc1MmJslojwfBAQCh/+h5yIXe/Jb
0/0kBxVyk1ReKi7NhjHDIIDQ8WT/IPv5wRmUwuNDpAizCkOQ7s0PcTQ5t9aO5V7p
2MVG9EIyQ9xwfYMr9qixIfZTmKMeGd4jd7B3QAOGWmu4uUR9z87ZRwZ+eGJuAS2n
USdALWXCgs6Lic8O3dJFKm0i1dI9eqyvm2KGP80wZJZEstVGpTRRDhwnQxqISG7U
3n1AgBcjY68JGGREXeUAOjJjQ07+TucdupYyG2hMHAibv/jo3Qk41pCB3L4y3kF9
3dJMW0w4AAF36IUYdSaBrUqq4CCqEtFLxWBUgLdlAUaBRwhBA3BlrohdRPh4qSn/
uoGT2+of7ax0yziKAtJXf2AgcNCJDvkeNtqC18edK/R+euQgUIYvkZ+HlAtpkP5N
0s1cG4zv6L60G93tzJK9btXXkeAgC7yQQAyxTrcvfc2iDrLgdvrc6FqNr8u2h5Mv
IAVHjxrKMBljAKaCkR9oApa8GXHSIdLt7M2M4D0zP7g=
`protect end_protected
