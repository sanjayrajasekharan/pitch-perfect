-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
MM9vZxU/0MSKkwABBS5x9SOM3caSAyasiaWtS4PAGlSiet7Va+Bpt52Xff60dJeb
yYNbWHNH/9QVJmwQRi/TNQY5VXZkarrnFtpTvdS3JDRpOmZzOBdJOYSPcl9Dlg4n
XZVo74UsEDRKROrDvXtx8T2CK7Gpmwl+z3L1ab85iao=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24091)

`protect DATA_BLOCK
lbtDetuQ9hwOFP2LfwzV4n+APlPCM5NFjRwnssimrBuDF/3GDEAC822E9euRv6FU
HtDhHqb2M4AbdoB9mIiFm/YozssXWTuEMr+3o5i7cghDH3WrvS86VN14G2DCe6L+
CVz1k0s5M/UixOabMyECz0kfjbV/cVH72WxjWvTL1gSIsaCyPwguStYfSFsI0bZG
v1cwu2yFrLYFwTiP2lrNof3Lexn3mdYBdsiC7G6FHnxIHXblKaO8dNr4OjYH4EEe
K9XpwzNLqHpj8GjklARh+DRmEZpX3t+ps1vrMoMAxowryTkXSwK0VrpZHMLLu46W
F6/UKuqtSqClIcvV6cBhelAAb3hvySlJgnf6ASw/lL9kiw5DI7zHZSg5+PeHPhAp
9gRKEnZjgvnfvhoVAoUVUq2tUl8V1fUAgcWp3oR+6z94YXW/VToG2v9lmQSkFO4o
vd5NycJiby0GCjiBUCuAJCexL8frGDH9ndyupbgyXwN7cutuQzkNQyNHa+/siRQ8
Z9yV6w1b9WAU3a5gu3LxW2rd5M/O1XHXoihXvM0a3WoWnrQCpcgUQNkTU45kNfFK
jvPbFSNU08o+yjLmuLWir6qLcc5iKmZEXWCgom1WPDu2rX68tNovoA237ek09mji
/0/rwHeRzVLkicBGUeV93mtqu9tfVAeqhkdKgrV8TSXmtqkCecAHTh5qvY1nigEM
JVcAqgtaN0bm0MWW06qVORIygqpex1VaYwm7QCwJ5fbBFlXcJ9M39Y1C0qkHt9kX
dnRPilKpNTO52K91fITn0Prqy9e7JxA8FSG5kt8/VoC2JoTsD7uIz8r7gF0mgUEF
0ZwXohpkNHVeZ1lDSiHKIQctqRUkourccH3ha5Gbcl/hPROfCGtlfKtsrhAxIZb1
/lRRPjuBiPYdei0PdHcJDwMd6Esge9o/GdcPa6CYuXL7xLH0nwSjmfGQGzYTjMLF
9BHQmnMS4ny8g3cvrmACfw3bzeGvMnV8zHxuw5XkUODLEGcJxVLCCr4Nl9OU+MeF
QAvJAdY7BWwOehsYKGqhIRQ+agU/OPf09FoPVTHkcTwzC9tc+ARoSsIY+AoAS+UF
vQgeCck9m6HcfNjpc6TY9GBLSsxFjWrE41PvZLRcFmgFue6Q7MmF983BRyC1oeP/
7MBM2VM1fOOjtGHZIs7q6F8pU70TyyxMsqohzGh14UmhsJIF9fhnxliMcqXDMCi/
JOrgTmMZTTI2m/MwPaOPKWWIuso43uQERIdmbW2DB1z9iKOTvxs/mHMEG70VKDz9
xylKpGLjzCi63Glr6xEZIaBSEJSbDl6LtRWqTm63oU4Gz6J+adD+cMBKdLt8K6I9
6kWHHSCHA9c3EGyx0uSP6iWToS9GAzn7gYzJpWoMYLJeyU6uycZrmpMGAwG0/N4c
QABESYa2yexaWGSd4wUEiz75tPEVxtJNUNK/WvBEdm8T/NJxNf5hP1IBGDOJejO8
U171OF4RJ2UL+70LRoUIy95Ib5qGIj3jhSfXebRl2RqaOCqax3QFH2Hu36bRVkxn
C2IF9Jxm2nt3dAK6RyPbCBMqWYHVBVF9rvrJnLazs+kmOA0K+QpTzPli4zGlvEjw
UCiCjAO+7fvcv9VTDiSRJCCQLgFxxdtKcCSQ6YyMfDy0QSs5f3GYOAGvbmxj9WCC
0mpsYLUGDckxnv/al5Q5pOi7+6PaK8YtvjWeb3aQtAeLW5qlmDXgFPLdtYYzuTMl
F5OqmSXeUjqfWrCSkIg85LS9AWOANIScb04b7OceYlaXrtqag6KlLQP1W+yS5lNS
bBRB+Mclm4fH2JV1cWtIhoSEY8H83X5MYJ5ULxBEbWjmugudynUBcHXmhT0kMN4F
X5N/yufxFl8v9dURF/FPYgZ1ZZjOsD1s8JQ81CN8fW3arJPadqEeLJiWZuButdbq
KKGuJ48v5xno6j21/KwB3Nj2dEgaD8Zs7xEFm1ugRUMkXSrt/Gn8vMfihPhmaA7s
ozuoiEqTXowxI14m9yvUKKUtZSqyY88BXAEg3VRdKiXev4lbVZpPRiffauMH4BxX
vlSf25ndGF6EhUCQhandtMq3A5tBFMibUGyesr0WoJKqFqEwaECQ04dxAfyI5rf6
33QIdIOnwI4mkrzdopW7JcQAnaH4Zkpp3atNtiaaN+82sOdnKJoUFa34Ssg13pF3
zokujB3eZ2XBpUAUSHgF++C3rObs4ZNQtHtlmGiPaZahu2kqDf4e8dgeaODKNKAd
12M1KcrHVMzV8SZB0M0KEP297DyiAo8mdrRm3Lk9EG8+7dRbyplaePl9Re9JPYeQ
E6uQPTHpD+D0woReuWJyOUwubKcfrEluWVHqXXDWXaJD5+c8XmEd2O5msHGGHV81
rY/6qkACDloYzqfTFHnzKncCmhLzfV/fpV4IAETabDXGoprLWyS5PKcRr+14baL4
FgoxfzTHSlIlcuWl7hQ0A+yGuaUmV8quq01eTJ2+sIOSb1iNhQr+fR87/Fc8fOqw
xTHFAe9R9AoDNQV9UMTL50NWNITLVil6kK+HFDOt3hoVQiZkrVOu5cEH2IOOeOXk
HthQWLVXramG4SvHrXK+a83RNnmaO8P7vTij+OOnReTj7L6Ul7Nm844GhI9FPN1p
wR0+61S0mslSNm9/N05cI5Zu/YmUbpxloD5Nxzk0bc0DLAptKAed1Ts/VBKAP/8n
nRvDcvWrD6fXnJBwt3HFq1OrIqGu+9CfZdNLJBGccNUo6ihW/j80MEPdxy6Lqlux
Xh05Yeau0AlclDAt5+CFy4p/HgvigjOt33zQQpU3fsE1ORhpw8KU1OKdOq0VxBc7
AtofLLUzavJaiFhfBdXQ+cXbMqzfbrxbiFt4jnnwsB/ITNn7dCp5yPn6+RMm+O6l
Jk0rlB3yS458bmAEoRgbDaRo5B02J77CPY+mn3FZWLmXIHzvV0R/DoVZNmc4LFiq
qcwXt4f3bYqnUw3dbbFG0pWj6wl27o5mcFjrb2BbJJOWwguI7s2NsRaOYo2LsTPN
tf7iym86Ws6Hj9DZumbAwtGzh6T0vcIk56Ig+7mPMV/gQLbUXUlq034DG8yjTuLq
a1vv+hnrl/YFWu+5cxz5VutDrDsIlcmYwSizTaRBo/sseAawhA553+7r0Ts7lRQw
NBhcdul30hgq9/o9yQhS7PtRgoOYUCAAR/sTjpMGHeMZojpmVISF9rsz4JMyzvBw
6WCU6CmDRNOoU9DvqKYC0/r1B2GvnwjwQL4QAoX2ECq+ANiSrRzsAd+xcITtVuej
F4Sl4BHbiK0txIhTfd4A7wRraxuOGaD8Aexz96q1LoAf7vPuJCG9b/STZSEjrtR1
lrhxm/dzR0ZjaoupBtaxMUz/qDwJjghCdrUmFTcAbU402TUWEmgNYCI7AxahZKS4
e4ZF/hevvwpnR1QdpVFyDGFcRwg1ZIMAqo1+wP+MCSbxSmRnW59ELFp6vHCtLhz1
1nt/wamN70GPAJ2hBR4HO0s2MRCW40uoc33RkCHJ3ltQQMFIsYsQ40gidT9djbEk
+Ep6Jnv7UBncMHpOvkNS9Hv/ReqcFWHn/eOLT+jnFjzOH/fwxmGcqXNcFvvsCO4G
rqiCv5lKFK4efXWSLbHydt2nycfJUgwlYa6QCHsTkFstQYqIPKxCLEyvOshXBMg7
cEwdUWILjcFOOpdVLoxgce22suJGkSB0EKzVJtnwgMTV2kXb+wb/q+Qr9Y5cvbVO
Tv+A2GmCG1KX4dH49I5gZMm6nIe4nEdlQEmWG6QBRZx/qELmTlFWChIlCK42lQRD
bWXHYBPXZ+9hg7cgGLRdGR9WBw7WZX47nGIeTq1J90TAgE2s2ZjzCIUZ5sh5RbaP
YuJTnYMDr3YgA0Ks6NwFF+na7Hi/qkBsIkYaVVt4ge0xcz+6wBT6WnckgQHCtlLo
D7MwSnXfLrSHu4LcPbcVj4EE9okZhqIfPkMrjMtPllTceN7BrZv8gPOPz57xcfns
AbHbpoj6bXNDo0mVTrr9G8Btnw0yfnyuyaNYC4oU3UARa+1O3wXcy8aj7G7h2DsN
ADH/IwJ3i5kLozXDmpuYKuenVU4SuYv3FbkSz12XcQARDEnh9DTABbEDVbTTN4a0
KEkg7pqUKyQcjWsu+Yk82rcn2E0au+16lMhNLD+PfaQXOtKNm+hhjXANVPM3Vp74
5hfPqJ6bAe9vEwWMw5/aQJngu8rs87LUZz0vS8eD2js5BSeeET9NOyOc1uZoMCP7
czAw7F/RTz1sX+Z6WL3WWRWsfuY4K/K2K8iQZYcwuGqoLIbj6OEGqMgwp1snlRH3
RFhe1wIod5Z/h3f/+cW7WZ1GQKvThOHqqfppwsoIaLdyzzeyS2Q7l30D6avObBNb
qmH77Gu9q5TdpWGoioHUQV9pdJ+fEwTIimgAEgLPX2TGMVOsyAmgzeEVFmV7ucGn
zyPEjaiZ2KbwabhQDZ7ITA8WkZNeryH1Aw8Nex8FGRq/bnRk81aWPwtbqZ4jYYR/
By6ToCvsi5CfynXaiyInWVumiVCIfqdXzeGyvAbGLLZQi5R9j0fP0TiX57keRiEC
zL7D1Py0tcQQaEvt0MDJZohiRsjfbmDIWTgVXe4Xh8VClwM+bsEVK6h41OCYFLrP
WZFhnKgo92l9NO6MYQiRwo0p/AzL/VSdfkGZCfNnn94Wyq3zLMKf89DO3S7iJ6fF
5qs2X5gbwOvA0NlkTUg35GxWuP6p1sTmTOJu+FuA79PiwIDJq6SMy2cuhQ3CsatF
YORpI571Q0HAum8E+ozXl8DKUP+Up9pMStLy6A+dsXPkGGR0ZH5FmozNECzaEfiB
DK5Wi799vEXTjV+wZipUv4VHotKiMIUqyFZ9a/56ULEzQ/2zUdC8se/YUulzx1T/
qZ31GHR/7SPIsyLrdu7EDPMIkZgJ3umezvf/jIVB8K9QYQDsfHAMXE0RbuZAsCKW
Da7iaDBEGISLZmkOzqC31p3r+37wkqhLopMESRbQ3WKuuv96c2UKcBtziwxktPoM
8KZLodyDngsUeYGcM2pVdp6Cpjswzsd2x1zbSXdUbQo6pddjVqS/JuXAbNThXOpu
/eiIadwbBkTkuJspQypVRcI1V1hoZYA5yrX2XlFa5VDuwWeMvFb1lP2bLLN4yxHs
AX9RZJ1tqcUA37v6pd5EeqFEPQptNv0ybGriD4v9sheVFImDQAMlA3W1hxpTnB/l
TDsV1cQoVvJ7xXQQn4FGK5AuatUY1yJuVphYV8NlMouoHaYTlUWEFE1HQc7DFMr3
ASTgRVeGPHPEoHdFHpVvG1uA4v4+QCBFHFYNHt+oafT/D+iUMF+BAQwUlV9tjvWd
65aKW3coL3hWKKjfIram1klgvH6NWsv8+2lBitjl40fO7cXY8y/485hdpThjaEpp
jL8JZmshdrU+27GgVHVG8f/iOPE1enMhbsEDlhLJ93kUSf4CiaNbSumHeWxGQkCJ
+bX7+LtQngNUvfjqYCP+fLodkI1VHUcIJouBC2j/FpQ8TlWCmMig7IO+DJPC7U+t
ylvyS6UJH2G3/2MVZD22KR7zDrmrIIBMGU8L6/btrPAucd7wKALT2jszeGzlftUl
ZfMYc08eUqnPbKTFAhwLp+bn8IXEXE3nLIgN/WLptpMZjC2kJcwNNQ2kC6G6JwyX
rMIpdTwPq8sHFz16/tVjBdGAdpFkdIA1PPNImMxqf9vLYjmbvOlNIs15+hZkBvBH
ZW798KUtYhU4gk2vjZhZgBoEy7EACzFWyn9ks6Y7XyHafmAstM67Zxqxu9+0ghb0
BkK3FZxHXnzaRnERDv8fiYfiePDHyZiaG9qkj+4czDeOjFAS6s2bXLvYfdy6yDBB
b9aRAk52Qynjc/Wjts8tImkSgZs8sbHlNpH6jBHDd+0dDy/unBdh7ijtpJgjoM5L
739BPSVT1hWchzYkghtnuqLKSB+3Elq3A8PLiTLNn2FQvzdU6MvYfrG/TEYaQ5v+
sTiDk2wO58PeYHAB76QNXEYHXs5CVg7EigYkwSc5xqqqXFW5xi6kcHg4t0xUytNt
YM2yBJ1jGMxESuP7e2slB+m9Jlw1RuxfidUEca9Uw0H4k//02AGyBBxDNPL4F7IM
yY4ZBa+rrphopYGM5yrc0fRl9ETSAQycyPHpdlBj2OiNer2lKguIcwPNJM/KPXxQ
+gzIpRSN/UpZIWphxePc63UkKLNXA5Dlhub7dWbPf0NBgp80KMJSQKqMd+7EhXBb
SgW1UNQQv9nxcCWJJ8xqfhh3UwBiSI2H+3hEH4KRxr/ojjwaZHeV2jkrRygRyUKl
5acpp3au1YCQ6q36jEwUFaI/ZbDybBY1EN5zOuUXP6eJg+NCem0V5CLPeOmjpwoJ
D6MkuSqWVl8HjN6KyflpwMJY3VA+GjQUBSMU8a+v5D7/295ZOWQEwvJrxO9esz0V
VfzUrQirzSJBqhKbLvHNQDXrr9NqZyxKUG6V7x2tEDH//13FQwxYfEa1cKLSv2gW
wqg4qDgxXPst1OQItn7f78PXWYTvrGwRIsAe97iz/T9VcWDNq+O2uZ8q/O1TMEfh
mK45w/GzJuLM9cC4HpajBXx8Te1KuNnb8YfnFwcpl9suxap22j9zG9VF+1O50eX6
ML80svJ/g4R/CqNtGScdhuILWXmJlDK+J88cpGcm/N0VaWsDHGn61we7nEso/QjK
tVuhCDk2UaztzDQg/Lkh6kQ/ObFizgoGU338aChvJ9xZzeUKqlY5PoX/sJbOKB6d
dfaGC8/2qEZwSwgr8Y70tdsSgieYJpIeBHvB38x3Z1zJ7fLaQst5Ml4LYRvjfzUo
WlvlPyztYULhTKygxAAp+NppCkfUoKaR+ngYqK+fuxxTF+VmWU5fFdjj4Qt0xO1F
joteEOjYsKxNM08YVY5go6UQ9dn05J8DzktbzgpisflngIXFy7x+yjDL0fzAxj0u
0oF0xRUr3MhdR8mnieLOGd5S/vr/+0xWFQq1v0KPvEFgGhuPWkE0WWflFrSAJb1+
STSWG55hSQiEklwITuo/vIMe0ZwgPnmTYf/b4/0Pex1c/lqVo6B6rAo+ztnWvcKo
bKUeQ5Efkju6EGvvjek0PbZlzYBX+ad6faP5xRYd47QGKxN3G3yoL3h8d6RWjHxf
GBUydpr/1r3kGWTVjt/LsiKwMltvqKy6V5B6iNDNRMgi6FIQNjqRMUihESr0Y6+2
gP4iuQUMt1mLzo2EVmJDfnnLrWNvmPoN0mYlnP+j/iqkNbFc4RmnWgeH0LFtVUBC
SSFtSdC/X+7JX4LK6oF3kYLB+AH44Dwq83UApiYf2YEhUCXtliZ9bQwXZQ1NWItP
h68grTrubmMuvyTIyMVJx3c8SA6M/ZRWO9lIr1Mz2ojF9jmOKFKewcDYUM8NEABu
L5mJ9LH3bNa0G5L+qVBfRkBXmBW2Vo+ne84qXi7WnFTI8jrLz6ryu9xMhjqwOAn/
avByKliHV1K68JaZ2yrpBias/dQKsZ7fgEsI9Ql+2TCY5aLRcI4b3obKMn36FHQn
7/Edws2+54p8DA64s6d/f+l89V+BUP/uWvqNyz7b52VVgJJHcCWatKvyKhb8gTZt
MxmhmQ40dPTAPllKL3OrdSFHB68JRY7Da14d3QfXM5eT1TeAzlNouNrYkye4KZvk
HNar+bETmJidpzFRtn2k1CqgaQABREISlZl8ApcKxX+U4DarL3MSeVITPI2fFXfu
QYDPUKZqqMbbcqChHe4qbqrQ3b5BNRhavUz38zhElJqcUSkPTVrbShkgrVRIBG/s
uY3okF6IKX7Q/yPm3MHZ8WjRXoS3mEQrF0uuCkbRUajoBpaKp5CpaYALTd4jyGQb
9Dhu+CsEydFBxyjt5+MCdndvjUNy2FeDLTT4uvtdyAXwapuI22J/0H3VzWjv9DsF
pjv1LYZ9U6EzumqsoSgREzPoy62W5W+ktuc6dIZML7jyYZm+eo1Z12W4IPdhCzkC
3Eb3BLJTInEWYEzd/ExZbnW6Rae8T8A6pO+D5ansNEp6sqZ7Q8ZSAGyDpkwQ3aGc
D0WVgTRMeE2oGOSOwPWipSx/4BevZ2s8zmlia/aIYggnW5kdDNoN65dmbsaEbo5u
Tq8ueZkjYSYXJcu76iX0XJS8WBB3LDVkE5v3PgHYNyD27a+ROo+UUfD0AmOAWC13
8/ar9YBEIALyqUayCAV5NXhcoCtWfs73TUWgmr8C1Yj+h5kTMvI/tBUF+MCBN83/
0GcyfSsNcg1r0OgHhM7O6o/qPYmLogIugWEIL3leoT7ECgixfM8S6AwceZXM4Y87
K4PxFBxlq0zOc66ECjm1GdcFPEUT2xv9aMBFdNTLT2pys9F8as+5Sv+xvkRalBmT
39z98YTfAneLwgy6znHGAFwvKbPYcyxfogtD3HjE1v66ITY2aRb26EHw8xNvZ1gI
ew9T6DrU44XPL8OrOMZwfFvMsA3vnHwC57ZR7RYx/HeWqW9ooRcAo6d9xiDqFe/L
sFSovvLekVNhcbw1czyCSASD948XvEC4Y00Xh6k0eFimGCvWBFOaZvzlsPY3VSmY
vIKQyAzdTNR5bPxTpp5W14e2AAR3mW3BDXYhR0ygsljJL+1X2DnLpLix6s2RWK9F
Wb8gaacGEo6VKHo9i0tVOJ9g48urDOkmPg2NVGuz8soC635TXXs5pinxQUUQjzMC
HuuRnDSyMhj+AjxjKqDclDQMeqgE3zzhlhNfn6/bEMmLAGJ/ksZdXU3VBs2zLWIX
czQN3ELKLkpfyMlLmNAuDu32qM3i9Oz3DpI/DoAv1KaeMv28KHfrxpsdykS9B79e
h8sx6IlgCGlodUHX4jx85rIjyOwrrZXaEnLWn9sH8U7GOWY+ORvtTiF5zJSPjT4S
/dULSk771a58hdnAs/4m2fBmQrwwswfB4I9VQ3wwKZj84KvrCiACWUFgs7loHNem
3h2fJ08KdvIAQXvrwHnNY5JG1m5Ej4sDnooE9RpI8oAdErfRucag4OPkBzNuYYMI
kqLD7I7aPNlnv6lGPIG9MDbiV8vDEknn+9wqRPOTkC2J15leaz19ksy/8/xLQjns
Oy2k0MQtA07Og6WaIZeavx9DUYNt1EHlt3P+jG83Hj5F1yY+I/KKpxP3YgeANSPE
l0Z/YnmV4MrGV4XGJVvmONHq9AgsOyNIkrKrAOsh9ZoDuybkUETW2sN9fiA57oz8
MflS17q0ectQhrXQEWvinu0eQtDw2BWbS7fKwbqG2iCY1m4R4L+pIo8ySuHIZ1SK
zu8o4Ywq9+RWLzcczuhlX3weTazM4/B+g64+4UKfsJlKMAlxJAlfU/4uRSt0oNwS
mgWC9tt9UAeW1eMnvHpp6NAy9NnzJ4mFTpjLGXosDBZXRoUanCqXSkO4deC2q/Jn
BzSAazUjq4scaZrZMptY1M2rZncSP2+JslrmxipBhqq6T5ne7v/RciLlRMS8mqS9
Sw8fnVHl4zzcqmh+Axr9Vnt/QKdjadtcFVHz2CirUDhV/dCzaJFqH0ZFlaOMBe2b
OEQkGlBnUIIGAXg+XmY2t93p/rWNuqFGrEedT+n85819zj8g7CwdPkn3BO5TBxwg
QNmiRBwzr8krcDUVwFj/buI6x5Kw+2Zj+vOJTxiQV28c8989XCAve+8MLvHeog9J
t+lSyuTRrRwNvXo1jRE2a7MgPn6OLxNJbAVNo0eeMl/dFfWzUTT7R8CduK6EsDTN
Z67uNkP+ktgMXQbfXFcMSI5Dq3NC+PlWSpBaAvvCiEfJlZilkDVihfGe1fpc+SjM
M3kLq7sRMWjXLWVsVIydN8U8W+MpQ+typCRi/FcyANvcKFZ9yCMISxaw24O4hT2L
QIbnHnRta4D+0lxXYx5hDNJeo27x7PNdNMCebkv9My244u6B1mc2kwne8WPBJlxM
UxZ4bw7EJ/9sHun0Re545qazpmSezBoJBsghkhjTzQrccvtokKQPkYUzp1jw7+v2
jiVYABQG1e2QXduWtH9as5eWzvVgY7KCrJKECtTwtdL1kYgGk1WRGF2dSIzh1ivu
IfoDpoAEj2wSyPkJs7Y/zm95q5cluUu1sejYJWWKSyl58R4ZA2+CC14zWjJNE6iQ
0Pgx8FIAvVAJKi0vHNqWiGfhryGRJWDcO3jN8FJkwLtDERuajEi1fD3IBR+C6S4k
MPkTDJFUAT9JPLVZipS1PnRWkkgy/OrvP6veVkt9hOzK7xCTcgI/qwLZOflCgv+p
N9Otl5lztUMGtSy7XjfJWG9KZL2eXFpCKgljaX3a7zYDnQX3LKbHNIxQkD78NAT5
ofziWZOI0mV+ii67Gtel1JetP0NCG51QfKPSDSkRvIOrBGKWUMs5GBuXXxNTBOGY
RgGsnCyaYhUO6n54MVpsqZqVTbuEEP1sbJZ7F00rZ7swCyiMkaRb7kmaRnk8ErlP
wRXSmCK0HGSArLE15VsGXO8RJKZQ+mqwNqjYMy21yBkxVEM5gst+cUPy9U+j/fmZ
MWi4psnV9a96NcRY+G2B/igkwqMAFD3e04sIXLgyjm/6n8FOGx4bbEiaY7uk/PMz
k4fYpy6q5x+5Z/v8Z73Kr7G/ZrShqcXL9FqVKm4L+g1LqUilgrZGvJpZv05kEMJC
dAn1AqBYLRM94cfI9Bx+6HrJ9+eNs36pAw4pCAXkcl6WGBt+KWjlsebRV34a5V+3
SQNo+YsYez/B9XoLE/5WFVy0uuL6+KPI5l6y/H2CYxQxP8/RTDdXrw4HE2QxCO4t
X/AsaKz63GcgeFkGGuryeBA4b+5V90J10TaoMAk41NTU0Htehk80U9+8+hX5DTa7
AzvdVsadlEQav4JPfXYtnV0XOWY/E2d1zz+YwfwGGiDZRbTJKvzhSGXwKd62XPqk
df/tLGx9yO4KoS8CyzUnuWCuuH5n3u69C6BTiKPdVSF1+S+KCQ//XSxIiAZAYFfG
r+hlWAT+oUvHbUEbOdSRP1hIvfMGPtJtd0zmKQT2gxC6L4s7GsNT2HQmcZ6qFCWO
mEq000CLzksbRuBQ9I6njlBjG2GgUaWvUZ42FA8aqC/Hqo1g02Tqdxj0NbjZlKl5
Nw+e82wwRMep06s40mV7AHNfvXTObydsL96LMVIonwqx8sUKVsntCTmE0tDu+IFq
UjcWSCm+e/4H4rscm0Bt+SIUcx2nNjrRoxjyClgUB2KEXVVVpWzCRF2xBhLO6VUx
WdZtAYLB/e7fCbW96MYouL7huO193rNNb6klY+sbH7uX9+L3ZWmHGkaVmY8uqs2t
Z5OVX+QvTNtxRVxfF4JbGv6kTOiyckmY6aC6gB72iHLI/5GMkCjECZqVI3qolmfc
sW0KCVCM0xv45XSEv+Rqf84HYrGULUB4G1avr3nbpwP4dmo/Pf8RyO5qyrdL3qmX
KcPBMbHm7rXmJYKhgbKGIh2e0pyB1EdaoOv54FcTa5M8yVw7wbYgIsAKU4si5n3j
g4kr/NIkgRM3msSNFIXvFLHfg+Q9JmBmVam6GhG8x708cs3Dg5CLGFqzmZ7QO+dx
QBO5MbM5hTRIUoG5UtGBjWhgk7fYZ4ky+f6FvlBTzbfslmi2ODTnmAI6qlYkGu9S
IAz+e1b90zAqYltGjVIcKen6y/i8UkAmdkLbRRU7kVWtAjDHWSTm4NQJdkShI4cN
MWO7pL7tp8o+Z7yuBezsmSz1nA7Ky6ZHay7jQdrjiSic5Mwk6NGjk3toJCcuj180
JPWdlW6KUfHfE5bFDYpjDfIrZVSENxcGqBnfuWqoNDjcTKLyHvaTo4CQvBPO4aFk
Bnmn8dlWAfLDrdncnrae+nW9rErnYHy3hre4ZsRSt4Q32DslB1YIAcGlvUwRNpvg
sF02BpZhMbEa/pDASX5M9RD0WYaidSvzrUFgkSdV6XlgP5V5BwR4PUCPGQLL/d9/
fj7saL8x2QCPZnsnUUyrOItpOvW/KygZ9++PnQfS5/DJEBNTSRnnJhR52jsdTpv1
cd5ujtBUa/TqtCyScnn3LSTL1Rwgd+ofCW3Tdn30xgRoGW71VTXKFMR16aSFUSQX
ZfVBIK4Rn/b0iKbJwei6ZZomADqq+UECaKu5EwDGbiH/DzahCntfqDa0KfkRWwOf
tQoOCz/5+x/dgdnJ5BQmskK5H8e0lN9+idcEA4IFrA0X372ep1G4wIvVFSnywIuD
0EUwjiex88fFIqDsNZYnc6e+K8796HOba5n2ajeOnq2oAIU74cakoVS9XHMuutzx
OMQr5Ujj//HAdXp5WtZ0FJ8cE6it+N4m1BNoEHEHSXQYwEz5gLlzT0Z4Nds97UXJ
szL9fg9l1R++a9H6vUAE2QBHHuxn9a2n0/sWgWFyhkw3AFvu0xb3NI0kN/IFCa+c
seFsVp9iwQaMpiYAklMIobuu/NjfkkFU9/Hjqjxxa8UyoFcimVMV+bCBmcAWdTdD
6SJIiFRs3rrOb6bF5IeGMvnrvV2qdCc6ogAwOIYI9mDX8xC460oFy4egRG1f+1vY
2gN9PUz7glURAaz7+AQ8oDVW28k9B0koAd84pE6yrTmer9m+3ItcvXC6DLgoqDbC
6ygoYBYZIQVRgCAxO16HNx1FmR1yTiWUXKufxC2nOws3b10oIPnQm8XAlSOdULCt
lDV7FGSjPrlIf1gRcylJ0yAa3QOk1V79EcrRQbo6R19drY/PVNFnAJKPg9gXDEs4
ax+sX7K0v/VQSoBR9JsSMAYyrmeqgk1MkAVPqpLeqpBOzDTRcTUZINNpaxmDbEz2
vx8LzvcFQrVTX0hqqjGO13oZwrHZFtX8bl6IbbQvCPtxIBQpWg/Uw3nYcWGZRk4U
G+FC461s40gi0EyOC5dveXKc4xARBoFOkJMU2z+6o1+lfQwox2opruWBydBUzMY/
DH9DUMVIjVJRgvDj0XqBf/QbtHG+wA/WC+QUN4En0YM86GAWwTmg5C6aojOp7mMG
WrjrCuWBqJYf3XO+dg2UpKLdku1ne32YFqxUsQ/VizZ0XzYyVA/JBEHag3zBzoxz
v1HwxsKRJFFglWJnYqec8AV6+2w7GnusSeAx0tcGhjfmUv+QzXQ1HlsIw1hK0oQc
YNWlj661OB7i11aBCECYavwZB+Xwxrn2LkF5MEZvDuhTBdidcyL12y/XV3jBZIIW
Di10ynodiewkZQhJv0c9psIlKhkMka5eSRk0EXYRv3GuErZe/gBvm3tiYFXTPqhO
IJt6KsJkpy85iqFwdHniBMsU1ZRcAQdbjFM3QwHiaDimFgK1yvAMi+K9NnBCmTTh
MUSe4cl1fR9/rfmmIDHWPMAEBZlxuYQhOHd48Be9CiG9rULQIMe4cqchIsci1he2
TGSfmQgXT23tI38IgnCaAzhfYdp+9j1Ct2hbud9OLlmJBP8FvfPRW+cWexcSMjtJ
e1wp0NcWw5P7FILeGdK59ZPS8cpgCxO3DXg9+NdK8ffvj4Ptw1VKZKoysRAYax3L
kTHFi8mVXDvOBn9VxGv1TbTLNnBPEm5IW0HXPtIXWN1/6Nxj8EmrU0AbMqwc3fBq
qyh0/x8drBLrHdcLFO7AQ8B5Cnb5BFEoTFsGmial834NJwxjWFivjnGa/8F7RTeb
epZtR3uhEjvVhXN6FzA/pIT490s/cH9Q8+4qW2krPXvzTNDJmRUh8F90eNAcUYdl
yfjMg7qY124yiFUDg3DydRGg9MrlSFrm5vdqdHFcvCvfAlbCn2heHOZgOOEpI2A/
UVi5kwGD7Wxh8psqyDGZWL59nKBgQazXMvguK6escFBEueUWk95dn0zkG8VauKzS
EmUP3rOrvGW8ORJmqCWfpvOCslFzaoxtNasAtH99nsC59w/z1Olv7tlMjTs2o2mr
nM/ZI1fwBcnoGZ3p3yR2VnK1bGdNCkdbEs5KJK4MXlbIDFcPtjOAdCfs8AO5kDNL
wXpvb9N2C/E3cdjgsqBNeETivQKToFQdN/HosTDKK93sgum6p88jYe9nFZIeud7F
KF0fjWUS+STuoq0ei2X+NcHJh5GvY2GOjtRbQZSwNZnKJ6Nn5n4dyqxZjqRBBWlJ
I/6edXM4OQwnTyvcqV4eIyRf+km+AxyfBYm974SOg1RWClsc29jFHswX9kumw1ss
x2J4uY25UfWBwQMO07+HqaNcRzJwE+yhGIlsf3lJAj7Bq7nxpPzGEQOhlLK+hQc0
olWkBBP5NCa79nnIeUqn2FU9+9nqTJE60LoopJs+5cfeWt9XxfhcLdouBtSQlBGL
KXyIGdJms9gHMP25wqY3LIBpnPCYMD593b7Gxn97o/AYr5srzM0tFfdXwYaHJCLc
64cFuN+x8HGvT8thfm/o1N6UJggSUlDCxq/znbi47LQLsPXuN6Rq7MKNieSDk0g6
DXYXeUACTybeUNBMoxAfn5YdEwyJmWsBZwSKXcDA2wG0zO9gGQYMh5RmoGGY2F1O
OwMavsgids3n/GORnov7lqwku2Sh4ENv4cVlLDl6l3fjzrEDspASBk+5DXRuy1Mp
QtYYyMjfe6MyROawm771co1agyvR5DGXi4HxLCs512fdE/Ecp3F1ghJq2Dtlokv/
0AIIdUTe9wq5OWyJGVX2N9c2jjPV3Ur6ZrM+8ITWqevgOBQRsHiuS3oTabYmYbn4
HYEOn881DFQ9Svf9wJGU9NKporEKKyyVMQbBQ41/VK1bXfcOrrY0AAnkAORcWIfo
SqjMpzaPB98VAtVFGwjxXQRuknLb6sVbNkaKcztauSbzJH571/BEPp8D5QYcZ2Xu
0gD8umZA5wvUzhv47kEAzlFU8fq2iU3QKkkmOrrCzrrPfIRzgjLc3FbsjxXn//4z
o/4MkhwCg9/07aSsVDP503j5I0DE5ZnYwBd5Zf0mhpwIaQo2kUvRbuKEXsdhydd6
sUmkd/+VSX83D1nUDnp58l+B/aVE/IEdy4bLKLSNw+wm2RezSYiZDo984eR8/992
dO2twY61Ju45vxhQzwb58U987hAWo3wJFJSQ16NhDFgKi049RBG34lYciLF+dKBC
b3HMrD+QUgzWyBzYh7d6dULgF0KrduWFaXtKJw88Ukx4sC0xw7BemppzQrJeCj84
DsnElMPCpZA0mn0qHBnSFz/WrS6pjwD1Wn7xARPdXEESVdCZWUvoYrYs4gw8yVoP
46g9/9rWC11yEXUV4DglmhfgAq4B8LhbnW2fjfwNqKDpnsPz+sEChmnkCM4FqUFz
xo1MVHhxrxQfPN8fszLeId+HqtZ2dSKolFAnSjFIcOXBLAZizt3G9tHHLar8PYuq
5/p/PZNt4m5SOLY6WtiZ5XhtnDv8dDx5JpI/Hf6ysamV1CJbX4k3HhpRE9+DhsCF
nj8z7yg3kuJodBeu8tRe1ukVWq6KLTFP0sFta33fMpf8TgHuHrEnNbMDm3VHNwYY
2DxUvjWojmw+YaNWc+8DbaJHyYBPiNZib6qRtxDLRZRNtqC0eZUNVk9Ii1jx/dmd
O6EA8+X3qLtLLBaM2XTp+VsA6iNExfbB8w4oQfGQOdI0ucog1RJrBDjvnSc5vSr8
t5xDu97EPK/mHIl3FrgAilh28j/L8pkqs9a60kN8qSVGczZYZx3UPqVOAU8UqfwE
Z2md5nZNddEsQa4nSBNrqc07/nj01//ytFkJpIW84GAuhQfQf6MB1yjuMzmDWiZ4
i5NhCiXqoiaxEVnbiRTM3fC8hF/5iv7hHYtvTUQgdTZrI/TTPzTXNgZ2YUFzH6SC
OGReNVv23XgrQwM6RoYcWN3UHvqYWlSEc2/Y9+3USjv2xhSdEnDOm8htIMj7sHN+
5DoiQDYnI3R1DKAzYRzZz85i8Q5n0gJ17gPCAhf8Swfd1JoCmvQ7mwaAXORG/hdj
phXiHDff0xmoRsDuilBj5papijWCgck/PpNqln5ToocW2Hz+5XwA7mdIaLaMpzqr
/ew8E8E8hwm70LCqJRFQQf8+UwcXxLNcb8bB78XJz3Zu2v5cLXX0Hsjg7NChV72n
k9cpf7prCVCP0JHR4161E/IrCN2cH0jXc3MEFUWowwcklrTSg309y0zJEgKjkT7w
ldWBXyGlKC33qxm5YNxVbra6JJ537IPi/3xoSIRvjNjPojIPlzPsiWpIlIri1WHt
2k+yOcdxJBWp0o2THfIJSQTIWL7CyS7gN7TEtPlmB2tUwlr5y/KpqUN7/l4qxIQj
drH/FEom++qDHNTB+e84XQdsAlYX0NWQRQ/v0FaKwWyRbFl9/ZUxCoKBHVyEYZqS
faHNxoekPaL4M9l0ZYkgT2vudsyJlwD52OmwKJXl1Cldeq/KWzpbO3YhLR6A2vWQ
QJpBDN4GiovbcVfapVeDEfLjZTLLqDRDKJsPjn4T4b9INfwEYZ364MKPmDrNapmb
5DgqID3YEtiFVvkBwklQbqvvixQqkrUYdRr090bxo2fX363oOZId1NvZZWuiaYDL
lZsYb9iIivxlYQDHJ7qtvtbtUl6Q1IlV0r0PtiORmcApa/zkTlCD8uAuVs8YOry+
BbxaxUF4rIPF6dSEiQoD7drEKlImwpmgBEmoRI2t/07TNqPjd6iFK+7h9qaW6J2U
uXl+6VO1Hz9DN672FoOvRUKgKygVJBuenQTFuw0eOOCW6aofvFwsi6UDCtHNy/Mi
TPK/B9nzr5qxSDvK66vnoe9hb5L3uCJITHgArapLGBqTEW1Jf88ZDaMnhQ6pHfJW
orD4PxIASmr9CcN0pTUyMtQdPMOI+aVmrIbrlrYbUijMXIgEDRmpz1FgNk9KgvIh
vhinALZV7WHZkwgDJ0jdh07PUXGXWQAF4QXbeA8bhbJDJ84q2Ued5JaY60sMJ83p
dlkiSKWPp4kFAR7zl8oSd+N/JHUs9Zftp4HdAvCf7WuRUq8wtIA07Wat9gRJuNYl
ptyQlzzTMBKmU2jWdOTUxHTfXBiQC8bkrgM5WTr+32164l85fr5s4QohnUT61V8Y
frZ+qut8qDBku6sZ/PKcP9Iahu4vDQpeDbfls9GH8IvLiA4Q0/gQ7x7/fH4355yV
kO/BprWdPVzJh1mGiEcChv7zaDBQQUzSqxlnIVC1QELojkX+/rfk2LnWWOgHNW66
xIzD7s0NR3FKLJVyNDNXQQ1XgBCh4x5mhrrAvLy8AyuGiIMyVxUYCH7EmydoI9wd
SWJps7yvcSaX9EVeEuSy52wEnB7okPqEy7zZuDaHw1YPgq1mp6oINTHFERsjkFWS
V1KvJT7DpjL34HwPLlyker9ByAtWDWcMmOFIh3m81W3ZWtQgKPvNApGRRX6WFeMT
g5pH+xG/xXBTGo4reHx/ItTexefl+nBbKJZlfwF16IbnIJ+3zIXoeZn85sS8O/Ma
+R2AXyomQ3MR4gj462YHoy6bTDb57RRG7SeaQKPTTddgwwq9BgVWFVl7ZOBiix9Z
aMIYXB7Znmg9MHKrDkg9npmrzji7Zlt/aowdKjIp5hLXZ/kzMCzyucohRU7dxHWm
cg7aUy280ADMGuMAaqpkCrPSrErql2bSiLenPVw5B9gTAifS+580B9ca35PDz/3Q
vCfI4iYVhv6T/owFFObBhOYFPbEEmjhSOuv2gqBwNrI/sK2mnjNjRdhkRbxMWxhS
dEW0xSKOMuIpcSmACsDwIvy8musy1MZd/W/mSafMu5vN6kZVl/RfRGARF8CsiEsQ
ytFTZEeFkbf8qn6vAYTP3BzvEORVdM9cRV8qyzGnernqSTcUUGLfCb0+eUAwoiNI
ajGHYSoJglwXVJt72zHdUxd8/VYF1NycuF6Vd7LXEP0V2IClzJx1SsssbGFacx0B
S2r2mPjBVsalgX1JI9YJxVsWDzVOvebg/L7m4w5dm25wzWBjEZ/wAoLMdjoyGdUf
Eugrn5yDv7v/kiv1JSxOp70uh22echqedUYN7oODN2LLVABVmImnbmtGd3GUJC9C
UwFeag695cuxFWHMklEJEX2Y2oJqaLqhjELB/on+/4RQc/HZh8PM+1iM7W5bWkhP
A43Y18LSkxI2C+HLXvnI/MSMI1aOcPeBnXifSv+QdRrUt5pGh2IkFt2CUzZpJKN7
+Z+duUiWKFVVKnDwUv4500mhyt/tenAjjSQIJXZiONJoIxT07DIj8W1VI0wzG+xD
LwXfvjHOkzbMJdVnGitcWbETUotnJojakoA956ei0ysTQXChcH/GRe93RoKfCfWy
4oUm7rUJ+wh3exxkxIQJqO6quIQMeg5DswucSePEyqFHCbnDJOcf+KIty9icONsI
f6v8jazzbNZWKcw+1g0PlgNpnzhLn46pHHDzW8uX2Sxg0tcL/oqIh5xnpGjYrvtQ
MZ0z+oSVz5bvGEAfYyj3DFdZ4i3XQcdtx+iN3onwemmj491PC121n5NCJYQlrwLg
5S4a6a1SIkOqhJrIFH++MwF456j0tu5f2thjkKTITumQuWSFOZJh/2/eohn7gwqY
Ooz9GUTm9Sih2vIHmx9/1nrdkXqvi6uMU5lNn7HvLPkkOaz5TRtcKRz04dqr7kj4
axpvXFbvBJOeqb1Lpg2MIp2Q3AJr5b6NmmpopZ5GvbhKpcLMNBz6QNRezE78mloJ
A29aSJ4NnPY1MyIC7EnKW0vzqAcHSmU1m+P3Tb2yFxylLH0LeGJkoXLmeriMvkM1
CKL4XLEmxmL7gnGTv5AlQhYIYxD1+hnEBwbEDZtD6Ro5qSRGPhWugZGzZjKnVJ9N
YNIGoa9Zzu0i9ndws25Qrz6uwRyPrv6eYu6P3pWeXdUQg5u1NI+yo0vL3rO1VSVS
jiy2/YvlBvDlpMtiSVpQ5oI7e0RaOg9lYm/8o16DGFXfPLdQ1c5wTHha59yKOMvE
tVB32SbOINu8XTViQTGyJsHcZVRwGXLB66sHhP+1+eUUTUVJRhFGxcggjDa/JITG
vepEysXcvdgEwIRMNuhQlyQ1waKSRAqRj1lcXRmc5a60OV7ql6z6t9bJV5g/S4UL
NvCKy2ECN0ws1FvhhjaHXl5/Ed8t10GECNqATysmdtJmbJrpBcK0D6DuJAVKJkch
nd0HE+O2JVUfmV21C8TfJaoWa4IMjIRw+CMp/FwjVCZtUvKLOOC0EoGNSsRRhVTj
rzuu3lWQmftbkPMJcCfCfYJFfol+EWevscpXlf0uwb7uW71KmdDAdC+HLbPcQwkp
K/X7j5RsRpmUBN1jWdCwX2CoUuW2U9nyuK7FQCtpD7RtaFyAN+S3NW2Z112WesrI
IqpoPcQ1zsSQ3iYBMa9AE7wr9TAltbkPv6jEM44SgmUMFo3LjdlyXKS3VyqmgRjv
DEyBeF73pZAEQRRnb485CUV2Q8a9PzGtc9TXsbr9gf/2c0vH+jXPZ7CWC0rIg9Ql
9XW3NUa7abIQYnMN4XbaqQi/oltpYWCqWgE0QEWETWSdXIAezMvkGgXUmsAkOU5z
rXIZ0qR3RTxyeVsoBaqqYftv+m2zJykaepC4ZoNWUDi/r4qdFOBXX2xqDW51i73d
xxjo5g4wXaVLlxJEtzCMSscsU5fZEOMxYFe1dUVSnV8Q/eFvceDwT3QctS8q9FgQ
z69eftVWB4s3zsQ+dd1FtQaH0RvPRqjjsRAigyM500Sd8GqVuAJNUvxef6fXOBc9
8JopAtV/AkaoGkxI0pP4r7LRcKSOL1DNJvqeIdH1xUTs6sT+f/6n0275k4feDWKq
M0c1RzwhiC24ls8GJM7eEroLkHgGNMHA3s2hoW/ijI3di5ujvVgrr9Ic0M8tQvPL
xCtyzTCkMpUZHsuAkPBig7Flx5RTHURU6+eFe2b5gZLLmgkrVgo2DqFGf0jkq6nC
lIFhszoOCcEt2/nE+uD0B5LbMabkNrerlyZ3fAq6u1mMKXRrwynSmWiwHaTvb6wX
PPkvg8lzCLlqd6n5QIWfAoVaz8AQMV55zc1ts2ZdoX8qWO1M+AdaZT1t7OIUdKx4
5sIHF55aWM5AiQAKQqSpJhp1wrrQmTfmr1xyjf9Wfm1lkq9uYPfHIPYxYy31yGRE
hoF156UIW17dJbHojufj2l2qBnDmHf90lFoGnkw0xH2DZ/oaHRhDSO8I4EBH2nNR
UIZ2z/z5Wzk4mlnS/wDaI1pVH4JxlPVvM+fwbY3Q6CqtoGffi3CcwGy+yAcNF9LU
hhtoLF6+h70rW9QO7Uph8SgY/HAxIPyf/zGaHHYdhhnWvHvRatJsCmnprB4mlNjw
VpZnkj8Zeza7iqlpovqS8bgw3NF9XWL5tZBS1I3Mmv42sp0G0gm+h/xH7Eo2GMRe
BoGoTn3r5Adff42KFFArVU0Y8cqphBQJo6TNMtYdiCe0s5bZvZ9iqIzKwZGpnpgS
9q2oOsaBeiVLYSqDrBOzE5d4q8xDKv5XRp1V/oKMKVu5nd13WFGpwjVwneAdhZGZ
PdDHNt4COVE1mPLJWSamJBlfB/wKiFaPfoFq9A3DCid9mPbQcAE/QLK/7hfotgPr
FTvAwsWa5+X5KqkBe/9QN6grzdKcW9GZf0foOdYTUA0DxjxTgR8mirAQFY6hCQWw
tKDFqSLx4QEeTwTRu2S5JTU6DCvHI9V1JOz/kxdtsOTXP64TbArRNX288O+EzzyH
W2jOAOQ6pcUWJxiYzz390i1Veer5MoSMaZZZaNlZ9b+q5CN+YkLD/DAFA++aqTF6
ZabqaWvNL82yI3XL5f+EHsiWJwhnqAhA+Uns1shTtdz3syA4XvQIi2qPldMCflx4
faIgIZPj+ig69EhPl334EPt8aJVpBBS1O0Vb6iJbiYIlBqKMnkScmHDDlDUrrcIv
Qrwx5lOjl8f1mgvz5WGzengPppcyGykqE4Jf/wSJzXi8zXb/kZTEJZHTuQXHwB9B
r4nlFjF9+Vg0bze4dqY37zSNZC8Z6hHZqpZGvyjYt5ASwxSF2bD2tXjTjEK/iMt0
Sgnc5u89HY9lXpHvpNxcIu1D7rGxFybysmHxIQdy/rRdQZumVCrevTXa06qgknEc
k9foAQAJ9rve0JcWpV04m4pg+bdCy7U45KOEPxZMr6XC0iZyRobSU1rKmqiEN4C/
WOeHBYjte5777784TyCmSEporFoXx53PEWyrl2ZxAFoknT85f2ku2L876XcqPUxu
moBcGxLWiRjdgHsVJiMbJuoSKTRHFlpebuaEy/anWu2vKgH5AUf/BMTig/Uq5lJ0
ElMHcB+SjtzG3qfMqil8514b7caSmNzC2hQwIArAqFZk6+z0PNySyyQNGYDxfbQX
XDOXUMyrPaGxA0vv4tAz42oqF0gO0ZwT4R6+8Cv8fIFV7Z3S7iQuthDi2tRWUI1N
NaNihDwOpKpcn4meu4iAPniwcKaJuntzkFu+F29Bw+wQE8qYwv/8uhhhk+JhfR4H
HNYdJKaTW6MgugswCZgFVDCJW3PuEguD0SPAP2cCbC8vZOH+luLtY1Iz7VolFpzz
CHT9XdpFPIHZAG366CQUpgJBIyXutvr5LvcT/d0y4yccVS3a22SMWKK7z/mq4JI0
W+sW4MSMNDMcCdFbdVomWKKuIruV33A74liSYv+bYcb/15CPzKnvb/bXxctXrJHi
cwJh+ZGQ8Xxo75XvAoSqs7/71q2/xxwLMyMNigH9oPgt48W10L5UzYq0OPdngigQ
7APM1j2be5C3fyvkIu5RirvZgqZhCecyJYWDQTFySaX4pPMjuF9OfSpQX/H9nVUx
EYcWEDqFVGe+l/eXcuD+Q25aIKk2FWfPEwW+XGFJ/zYipeLgx/K806UVpSLj+fLx
hBzybRWBwy45hHgJK+07AJJHvqntFD/nwJ9v3SmjzbfXN7TwPLGWqMUu0vVKBAe0
F6A0LnroTRKudXHF5PHOzxCyi5x2szX2TyFbtrbgldonGLk8qnonQLIr6WMZ9o5C
bs05P0aXXbd6eYHQF7QEkMpM2o14bz8b0SK0nJH7T5N5kLVxAJvU0eG60a6taMBE
XlH4F1pY2R7L5xMr3NYbu7kBmExQTVl29ONpW24POE4c24GebntPQnCad7+WpzBq
QFo3Eq4Ny2oOlkj3c4YDgEmL/ib3OjBqbGtOBjjtgDar9QdYdJk7ZLQG05hQlldx
AWvFFK4Z2igh5HMpzDyQVZxY9teBuzFtjgKufUJYJkPM1h8u/qavECTfynVZY9IU
G5YJzXpjcIlKeb7TKyUDN0eojjbFHYO0zFIli1apHrAIkyT5fKp48vv1GjiUZqYF
JOyl9YWFQTHPZrx23UFAu+tBHl/VHy/jYt9zHLJCOGlAC1ohg9k4TGwfLZKXhoNf
1fH281FHx5AdoL7fdtm8ST9EWiE97Xlfx3CFSdAKGa5sLM7AJxZ6fKdKU/m9WCeM
iPmXlHkDsHWL9vqFmwz9bhH7JIwNNgZNP4KWX7y2WYoXcqoVYNG5BbZ/KlVGBGgB
TxMTGtPlZN+JMS/m98QRm9k4xFnmh+rorcyhCXXiuGBfBHSO/6F9SKJ1y0CFuRJx
fpT+udgzqaZm1zV1vFt0b7B1Xu5NASRvuuKeUJCwkXPXQAlm09YaZZjY2Kr8aHy0
6TT09dgWiBKQmKhlxTV+6EiaKRkAzA0hr71In9zZ8XHay5SbIAcgJoiOsGWrzeIv
e0a6ReZVv4fvKhdB6iTN4GwMB4auPX6BRDcSQLWpKw6NwBNBabidHcwH8bs3N7nG
UHIIgOCsVbRHxgtAb9xURp8bhNrk0Y14bRzv1akm1S/NpL/EWcK+XJXiPNfSfH5P
b4pr+AP+lXgV2vuaeJeoT8CKfYMj7zOp7uFxLRLowHWtHmZEyjSvtz/MOWgumAR1
2gP1DS1/CCmydMxlA55YjQNd2ICa9e3XWn5AR2oP98rHL9hIIsgt4p0/B+Ha/Qr3
lXChahFCE7tUFovYSZs5UdVGvf7dLm1czMGODSG/BhQ3hGv2LZyvejw38OGdKBh+
N/Jboztfy0JDVVBbH0VSpQmD/yFFs/JVmo1KE0W+SroxhmShseLPPmDI8Cszlf1Q
J8oEHDEN1E7siUAvm8x6zaSspKqR7XNZIjy/I0XP5CyxYleskTBHNxwbtmiADpMQ
6q5W12MZX5ffHdUDTtN6wYVqpVAGf4rzhZV1uhoRDwXgdcm4NpqenRVjj7OTlpm7
uKSSo9MM8KsxkceJ47rg/fwNNtK1S3Ty4plnI0gbf0tM1cN0DDqE1wJW1LAawP4m
NkUKxbkkgxHFauaH6gCKmPMeD4EToIaKzTM+mdJLCx8VUCG1nblJs4ulOmE1khvL
C/FXazeJW3ep9R4sW9GdLHBa43XiYFGCpeaNqOlA02vB+EBT3C4b4T097AnD5Srb
oUzLaIsni++XlGeKNaCVsbPVM7Y/Q+VIar3z86hgyYiStnoe6NDKv2Z0Ypdaq9h1
19BuNtZs8fSGRrvzrni/omn8HN7IylYvW2daBQOYhOlynEAsozRZVt7NErTkfrqE
DhfDBRdeIvlTHdoreVdVYsxhZQ1og/SzQGgqATWVO7rT3xfiWVRV2gALhTaRjSc5
vVfcTfTZ0P99hntq4tdjzILYkSJTlAczEL249PTzOGayLR4SyIdlf7mmHxVw/6EG
AdemaoDabfGfb8FvUlLQB+e0vCN/BqokPy749DazPk8mepvkGfruyeGJh627dvW4
QRTKZ1xtDSnWgfDvKsxLSktP32aX7fXrDPZpD2oNAC2WAAayVjDV6RCM0BLGePx1
02KBO8bgNRRtoZ31XOjmRdUpFx3sMcc3LKuBCQQ9b+uEB9ZRGaaGMoAkV+Qwyqz+
9oLMfU6+tzJA3uQcjNUpf+emevnmrdHSP6rUe88uZ+6gHGYlF7X0psuqSSlJNzwB
ZYCqTQ0OFK9xTCrUd7TjA93ok3VTTBioqnGg+PMcNvnVl9X2DQ9z6hIobnDWuWac
h9DeKdxLS9tHTWoCgCu3jGyKcS6HW5z3LC7khwHXHs3+IcfYaox3Nm1BcCkgkBc/
bNkfLoSEAXrwg7z8uA1ZPjbPd8alREEwRzPgk9HNJuTOtJsiJV+y57peEcnCT7ZY
vMRbRSew8CiR4MHNGDWp4oOtHf1SMXvf7edZNN0sXVoXbZo7Ye4tNZmOozN7i4rI
zWx6Hzu0VO3N4JZZCWXgbGdFCM4uiUcWIMM8azU3afwc5sj8GyuDJDTVNVUaTWeQ
u3JRMlw9Ce9VLqP8WX3Nz5ATKFFRnWpbDjkrEkE8B1aJbrYDYe19SzfB2y4Z2CdE
zeqbGfiQtxG9O4jcgTtRiIxzkSBbDbeg2iF4l3EbqzaPerzybF5AEHclmASHt5id
yrobvPG3AwNickxangsYFQ//8HI6KBEWVTJ6stun1Vs0LfCGVea3W8iOZWHDHZ5I
Q3DIT6KktJJmKjBgrgTN9B4VBDbg8OHenjGUmKaifxa2MM/xkZ0B6qa0/sG4Db5i
Ow/dCtGThpHK9xGpHwrlgUuf8zm33DtP6ey+AR9P87weMA5CMj4dAtQKdD09bwiH
hRfeS8eTOiytRn9cLXRDJBFqpLhqlM4QhPhjAmL6Bp8myL3XLlEI6bym8Ys5U2gF
wP0R03FPaCDz9xweIAf+W9tsReHmsaxe7gaehJx4svf5mSrxDu5Kd9NClAjdkVbK
bGP8PUGMirDVwsYLh2Nq4i9Cu5Htu2GbfwNOPfDwo78bNqALKvu+cXfoYs1i0ECW
wYoufg1EdIL3a+0bEb4FrS2v8IevX/nrPqNyg8hLD+5kroz89QIMR061v69rd1ZZ
e4blfMlkkV2nLkGyrHB81N1HRoQHyxE2xTXfcIt92ho9vC13lpEV6s8U8s7uJE9P
C9OChRwEt9TtI1IxvYHO/rpu4z6MYCpUprNg+ZxPYVcBOA5W6fInFloCqeNcPJjP
zFmE70CE/8IiBEwJndIrtcKmFaf0yebLDp/iI4XCsMVpsbBVpYl8HPX+jSLIgYRD
pM0Rbxn9dcaAyGLmAzZ9jpNl6w82qvEslrdqGdyALB9I4bLDpJul2TldqHd4u+Vn
wmAUHsx2jc8E0Pcfg36OfRbbcHsjz4J94vKbFHTxAM8/U0B0j9poKFNJ2+x6srG5
DblTS9rAa42vhzXXKQ1vfp0dy5pdo8+IbJ6gdfQYSJ2DgP3wSXSbxREwokOKf5L0
LqPkJkvRcUUBpr6+7v0DxqVXuueXp+4ekzIE406SosFeryqUBCaO3PVLCzdhHy76
PvGglbus/vY9ZBZXUPWtgdlx8b2rF8jGMjHTgHM900tSQZrpE7BCUSk1AjuYWQ3l
cubM5kzd4EpI1bUQrxKjDGqcIwkodVb+PSUmkwi56bxdlzxveMehkfWMamMrs2Js
sYKHs1WhlLmJ8AbPnNcrDvpKzMx7P78l/V+bUqYPLb4KDjrwzhwkwmSNOVxohj1R
YBfe3vl5+W44GaBYZj03kU6ZoyrS94gCXhQEybvqUodLrh4rAWNrb5As8W1JxBwE
1++jvf5YT2axUglo3MYVCEDaQRKLx6UVlOoSuvKVkqjBHBJhGVHxpYEO+/tc2lPB
srACbilEgGQxk5bbJyChQgRgNQpw6hUFE56OnMuUPByP8zixNwvyf4xZMcbUvI+V
ZwfUXRy32NOdiceOuhvC1iiCZ9crskV0t2P82YpN9338SX1iciswPGD9J71Duyd3
o7gwCdZYIlpnZxH/OUreMr/Go7y4P2ZKfbAG2nl4y/nPALMhohMllLPnmRoGIeeG
AE8uUoGCVwggH1u2bhneyOQ0Xax02qgiD7l0xiqUu5zYOSDnopd3YmEpPGibJprZ
eRHzQIWiuMQ6BSnQcvu1C0cg4EYrwKJTr4HdpV6Le23s+veT+lPKyhwELnwawuKj
oh370Y1JB4KPCBoudTM9GARQuSG2yRWG91J4UYVcsOtLO8lzp7ikC16Ab6J2N75I
lsyUUv0szjPhSmhJDyukFkTteAuOpQLW84Vc4QbRs38JzIl5W8tulmkFQRHklp/z
F0TziQ2Jx4JgtLnWuMjhA46Od26kaCJHKtq0K1yMW7y+L6KM0MmUbVh58iG7zhqh
/8RUUpi++hxI4D+9XOEJQr6RlvVJxYV6hJ8ytOmSf2ksoe+0sezkhJJVVkU59RIY
2fVZHXPbQ/lBVbleAJRKGX7I/5+SZY28kXisQfQf+3tOVhD/q2pBza/fMhCWyFWK
pUw+lFz0NYwNtoZqIubsyFOvU09PxGZtpXClpNQn4YM3K7OM9FBpVbz01rV6Zt8d
A+Z3yO4u6EC7h+S66/XZB9yP9CCve38w/6O4YtqfmufEkppi60EON4liBLcaZ7b5
i2pNfClbvdJ1rO11ZDgBlqbr+DOMmgjlreM4vCansiz+3GrLUqxm2SATQak8NyXp
j8r2Jntw/IG+6M5e6yR9Qi4rGT7AGPKXXHj18WxHqxBU6hT9ZpIYtfJXDKKDwN8f
iB3eNryUWGczfkT4jUu/ySc7AeO2C2Iwt9ItdxdBTQS5IyY5UzWsmTI0XnFfuO43
L4Y+mnykFs1SMhnV4caT7WD4QVid2fUIY5Tv63PquWjqksRbXuDBFI3LXXDLw1Xf
ydIpf8q4otf/EPG/m8pOMN4qVpLeNeYxVs3oY2I7QKZdZ1UUS2jHsXJsuBoK5PDv
j3+/7+uLWXasOqqjWAAJZQDp+9XVII/qM6YzIC8MeAMDWtBI9FOsmufoCvF+wAst
GvhUfUhEMy98XVystuNMNOJZHR4cSh/jKXDU9wxzBGdTcMMJJCZEnE/HY8Rwz64x
9yH4C5DDPu1UGKRTWdlwF5RqyPw+K+pqYGEyryGRfIHUHXhqpt+EqHsQEp3W5i+1
0PWQ4GjLr0tkSwYzPnlqfH98ueggABn+vZCBEfnoBTm5RzPn3tkbxfxIQryoxIMQ
D1xhFouF1goB5wd3pnDyP/nc0UtfSKCa5e37PczkjorM8YyBAjSAUa0k1V0flk0q
a3+Mpdm3jSHH4rl1yoXxCOKsn96C4cTe1dWkNFWSG7OfBdlHaSFB52R3V7p2/cAU
Qj11VFtPPi24ESrT5Vi+4cPH4nsmmv1T3rpAnn5+/KKMMNe6ug66y6rNUVHSmJDV
RWn8V12+kx9ptTSnrg0BGqWUtxemx7KQS1+Ic5E1iMoK8Fvzr9MLhdYxZZ1hiS/O
4HRHZDVRBGdbipbM2quujk2DHfOGfV2WL9eJ4rFjD7O9DGmxC0oIPpIxdCxNnCYH
Oe3jxwy7hT+ktosCc9gEss2JfcR65JpxN4ycwt41NIDggWDxaMvtaH5AL+CHI1J2
llarsJurm4mrxIerJ0mNjQ7ET0fxEXukuBrztlSbG4pFpqtQu2llo+qeAMSFOqvY
CcIQUXVsfjtTWlam5S9/brZFN8SiWBWl3aPNB821QX4T/YlosrNTFYV8T56inscf
qLbSKLkFsLXHQ0OPUkRBTLdQbK7SqgJc3bERLdj1JSNVjmDRMHF+EWC1P7vQljT2
IOEv+Aaj7iS5DX2HrYilRQAvXP6WhpeJJueAB0DkhxLxEtfhdPw6dMQp0endosVR
jsvabLuRXjw3l55dZFRbXtJCHridMyPpuVMxRJmcnYNHdlYCgIq7HjMq5UHOM/ZA
cWbtz+MrtBErNn+XacKCARDaU9HZykLOM9I4TDsy2hneMiUhm7xfA4Vt9NQOG5bV
aai3x1b4gEgPRukbRdl9nJQdpJrEtOS6LnKZHQuyErjfv2nWGyVsGeOPcXtfOeAC
2oQS3GHpzMTHGNVvTZmjB6GY9ystodKMY3jK9TMzo4ItsGmXDgzFOckUP8wUwbGp
s3mgy3VY91pC6JzPmlpcgdrWW5NrBx8aD+bnF6vrKanIBAGLzs6VAiqv2Rl7Bk6q
iYus0pdcPUVt8vy2C85Q5jiuTKFycFoAMjZ0hBzyMjnCjc+Di+vs3Ymnb1XQe/Xi
xRJcPxveStmkz93IYEA4TLxhapYjwWeP2s5GwaVnZRRbgqSSxxvJkf6tSpg0TUOS
C5DTaVbewCdYzpUVub7y3Bfrtv2AVFPnEY8hd0owVw1/f1YBSyu3xHzBjboMwB6m
OklnuTGjGjrlLVfv8JtRdPNkGp5KkTLIBtFBTG01+YuLDYmNsaRR0mG3hUuW4to6
3UUeEhuQOymyDhaSbxGR/K5CBsk2nqu2Ff1Ldnfr3QT8mFU+VApCNEU9GsuMwzHv
v9UzU4p3jYIwvLLP8WEUGFwHnLcK60Mwc0bQm4eQ64tPdGIt3prPKl63lYqDoB9A
mh+fWVZXpbcUYEBylSMgIHz/t62ygSSVs6MbNbuLw8YlPKnurUhOWs4MtTe1yJXH
lbZcRaaqOyUd1lIrVBMOkHluA8TYNKDbL8s2vQ2g6UA/NLmDOOHg2g8oCL8Dh+h3
JIny8/OfNkM4ZnSdn/qKBT+TarNsE+uQM9JupNmsS+jiyNyxcUSG+gq+c/dvTxZb
SHcVRNG+DdHOYHbN26M7oJ+La5RSCewJ1RcctVxCAk/ViaI35j0/pyF7BEQFswL8
HH8R73opDF5qQ83hQOyXD0cgjlvIjWhKv9N2g9Nn8d4RNUCIHR4MM4QUNLsj94KF
UuzrKiST5N/xnFnX10BR+qJC0Fx2JxYnVISPZQx41rzJRiUWcaRwP8lJa8nKn/Kq
kqSar3gfHCPgwieUQLhW1NMIn+6MbDo75LtjbFSsy4d9oi1CJ9PnyaouDeAC5gyh
3XmhKjw3PF3Py3lcQ5FPLxOrsyWZR5dQO2goEFKJgEwkFfcR2+nvmzZ5t4mRIccm
8FewRv3MsWgJVEHKkOSRfqOZHu6fG6+ZGorSrDGJVCIDdudLwommaF+QAxba2sh2
7kSpRzbImI1ps60aAVvqWb4m5M36kHTC/m9bz15Ge/hgryCUy8FuDPsTqRPDBxR5
cly/HxzsNHk6nH7+fV4q48zJf+lcussuP9jhzbfwNxNR0rZB0AX98eyl02WNldHN
HpECLGEDBv+BWj6YILAG8f7TSLHhIrN8ZQ6ScBF+6s+HUk2DbJY8OGr/c2FRr6sP
ytlZcZLZ9gdN7OJ0q1bkcEyF8y2sNrAQu9fHzVYaK1aDqgs1hUkItKsVZE7nrYVA
xEWvWpa4RocLWSoQt8oLaDA8YvHE/41QmHIpyTiu+PIvkgfxXq5fYS8BhJaGdzlT
6k0Y4p1CcpOIg0OLBESb7ZzRD/pD91e+d/+bM3uutJiVdw40/vcyA5AqUDCRN1Pk
wnHd+om7cRS5/mMd551cuLIsr8z0AEkFkRUj5TZKksjKFYL/Iri6gxtmZx97uKNp
0zDJJuV7XSoNjMGFQmLwMzx6kzrosjghGI8QdzLEfAkzv4E6raetL+AOf0Rptuyt
mAQa5yQlmDCld/NGG1+blb4nSUFE0T3jeMTDvuOCgAgLa7PEqSn/3qsIWZMuW11W
BZpqV+pA+QwU0pc2i5CaZDefCBtFMFjLKmksZs1Ic+hmUrnYHP9EiiQ0mK78pd7j
w2bhFbrGo8/C3mm6hhBLLgnOvJRLI/Vo9IYwt2v/MCvrUv9RNktdJlsORsIbj/DZ
+l7uOq//sGuHM+cP+6jBtkuhHOawLes7S2fRJNXqomDvA71R5nCeW/QrVqImDwHf
6qcVs7U66J15Gxu878sC7VrYsDBRF5K+tHhjlMDiuEjIwEAvx0wQZTjV5y4TXvLF
HmZGvql7+i9PfRntig7ZefXqMd6WYhfqO5IvEhu3VZIs3u41sQQ0KZ1TP0rAvnxa
8WASCaSe18BDCsZQ4+g6OCZzIBwpLmzMWYx5FlrTY0ZGsQ9t71KwVsO1WxNFa7Xt
iS1KSFrmeuFwr+0mho2Qg3fVnVszOXFAoL9sLJJNYMZU6ZGKRj0wjfXW9ujaItSM
mmq5SuK9esIhWlNHlxy6v87W1b34S+P8hFJNxzwkhGO2L3ZqcAy/19OwcYdbPCkE
pDfAp2ZMop40fgHIips6QZ47tSGLsp8WRFWqo4cGYLj2G70un3ECH0JeN6RbDRxl
F4oZ/cZkLTOnLjiy4JTs7ATzQ/xRcoLXXbLz5CnNRR3Ua+1AY4d3vZwxmJQNFPUi
1ju8mpdxjmNExQxVWL4MTJs2bznHwmdHEKdF9LbCJWhMv2HfrereD0k9n/PxpdQP
QBZi7kIFXD+6se9wLvPn7WXu97QiNCzdNWA+z0K49Zl336heMmJxzl4NUM8h/7pj
ek+/Tqrm+ZZdLLevb37vIsErhHtgXJJU8O7uw1KiVfTLJ2j9mdAtAiBMK1zAgTzY
TmDNnLAic8dsGGU/GbsbS1zOYxRjTs04yoEWFyBhN5fzkXWfg0NkknyPzjARMbpT
tqTFvEgtLbQlHtj84FDnoOhi8feigRnB5UyMXA+Rf+Vg+UO7ESZ+JGXBGODO++Li
mKSiIil5p999H43QaXuOlGV4BXj8GuYps2qOlRVLcuLQSzPchQUKigX6JGYBRU15
lzDm9ER7Z1OSehCVDAsPmltwBvLTSNrhKEIF1Sd7Nh6MryWxoJHlDzpWtfG6xAob
rfT+wVYhokHWBQF8U6VhkgwFGQng2oS0bKMb5jHg8+KJXcSU7FWUTRKiqt5QUS0G
Sw2HF887rRGKKlT4z1vZpxJJ7c9wc4FCMGMGDBaUa3ZBfdjYdg2HO76yscHenhlB
gmeUA0D9uvu+CO6oBDkQ4qbnhaW8VUiBBi0S+tOQYZ6c8OPu9DpsfaYG1Pf1t1Ng
GjQ33ZaFvONlUEkea5LKS+oAznDx20PVYRROjX3zRk7rI1Jgfvi1IKOQ/zlINzF5
1XJ3uRHQe/V4NDr8RKQXpmtJgKSDD9wQaWaqvtPQSCQg9tLkIgvEjnpehThOpIdK
4qGOGR+LLw1weoZvXYidUZPOh+iWInwKQ2g3CZzyCDS+VXTjs6glZAabxrS3cSn2
J8l+jAMoQ4TFVAezp61V+GgRizjPkeycIAll7/cAcw6EUxut+kTicMNSuFFK+VKG
T1hgWAYgnNDuYkOBjmF5qKAJI9Ceevp8YM/4DuxS6Fv4Ypn6zjmrx4rdBK1Inkdx
JhjhTDGwB+7T87G02QwgJWighFS1g1J8eybfq6D9jI9kwTf5P07VM3BlqlB01g6S
POvZCN/EEDFou7PLRqg2yaMfrBjH5ToJUM/UNtNznHYkwCgtF+CHqWqIND+MITa6
ypd3B03EM9n2ffjL3Ym+wYtoUPKaBwwjm2ryzEHrZSPJEBaXNt/9F7qDto8WcmoG
cynRcdOfwXSXaBCHP1MaO2bn+uD8gqqwp3D1owFYBmQHNZCEBsw0cq1TXQeMoyv7
ibq1KAxi9Mmbn0tqz2Vsnsmz3zeLGcrCrU5gvaBIne8uRqhDN7ahzboGETf47WUG
oSdKy8PriqY6QXjm2fzvQ1Dx5r3kzotNl6l8aiMB4KzH+TbSvWIU8Rpe2zdS3uuQ
dMD+Z3ic94Vcg8FsU12T3A2x1SZnd24B2ARZMAkCnXxdypAiSFqayxWM+p9PVFTl
YJKkb/KGRk2lvRtV5uKXjYtmlBtFCOl0idxhe5OGEWmww0pHdjgQsJ5ZdbkTy0CF
FAFXePRkh62KqZXjvKwBP+dNHpyo3AMwnGGSIHKBwvQqPMbiu+9wiyGkJTpnEL0y
TBGI2sgCw24VBvB9xNgcxeb2ocde9UBew1AfNRajKT7IhwxsPdth59BYynqTwk9z
tqJ5NnDCkZDRG0xANbSXY6yP1mE/78s9Jv08ZTr74OvmIj98v6Ny8TiPxtNGGbAq
knlclXy6jBGsB2eEpupQJJrsavZ7MaOubrXmkbu/kecmPiLwdJAxUSHDqRua0QCK
yFlMY9qQXCCYEQcXSvjEmRQqjCQ+LRhAFkGHZZrDj88AzDwuEnoYTun7DhU62cKR
TnBsyyy6O1AlUP4GgwO7+EhpzjibuIaYGXgzTjowi68V66TTu9JoMQnggapNQa6o
7gE3clx/T8DB06dsrzhKjEvplEoIonHH/Z/AnmGDetnjDRXDUbzeIbdQOcyORx06
034vVtn8PRaRVu3zpGm0Rc8pRjWzpCASZw4Ey47jRluda0vN5ffUajEocCEl4pyA
NX1+oLS8zYZrtWMuv710Px++oJQoTWJJXoX15AA703DL6VjecqmyeYo4Yd2zGDHC
80Jrrqwm4GgZf9wiRGzr1oHf0Qn0W3F6T6w0fRjYimWS8wPq364ZxWHFRcI0qISR
dEMF9b/rWkCOT2GHM2GbqSVtBlVJgwBjmF4Yeb0/UCXBnGGWWVcz14wNTebpFKl8
yp55jhn93ehnAtjcZM9LRPtcKJh93b+AniTvYbnKERplUijZ5QOsUglMaILx/tBk
jHFyC1Amcigqinb+py0bWom4FpoJSrNDFSpsw5Nn5/ERJ6IeC1fkWVPfLHuEHlLB
u3RVQiaNqNXmrIjqturyPQp+MI+F7gJ9Oe6WVAYMnobfqyYFQ+nzScUWEtFOCY6V
8cUPrvkvLPv8p9nIhAHIJQ==
`protect END_PROTECTED