-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
8h3mRGCg/7HYIxOHdDvZK5Wg7O2XjA9oaSiTmFoqBYooDim0z3ztQSsUk5HQKfcY
D8+4YyO6ntNaGHQnmZQAEBoj24fuGSiM60VsK8dVkiZp2wfEylBhDukohlXrYI7T
SNO99K+GC/mJsOA0hoptnFYdYNTZvHLoounSQp5G5b93Pcy758ymKQ==
--pragma protect end_key_block
--pragma protect digest_block
O42wNT4aZkf3rh/J6f0xyCLl3ak=
--pragma protect end_digest_block
--pragma protect data_block
7Uzb49xZw0kl4eKDl0onjXDl7yl6yqlFW1sUReORVEsLRitiAA4fu0o9b6WPpX3d
rObIjNsBvnNgVLDY+mT8OVVrNGfh6YbB5zyDF0RqKmlo1YgzmX9Ux0oaQ4MZ84Cg
GcR/Om/6LIbplxGCb0iIBsNAr6wQR3jck42T2z07LNdegLDhcIZTTDVZ4Hz0zvEm
MfzUhdY5S5/zdiiove3wjy3roM+k+zasm29TD1JGAiC+xq17MF0B6KRoejprG3+B
fEfB2oxCt8bQKb02TT3x+9AouEHEVZ5ttHTv3qwDA8QLuJKm8snYV462YdcCHY9Y
ch7xqCXnRNDP19qrCtnsbn1QLSVEOTw7sk/0XapF42kIhF9Vm9XouaFKTjU6CyOQ
U/kUqMps+e1mViiO8fErvf3bPPIwh8CbHWtU2KOOwCl2mAlR0BhGbBKYBslBkORt
dMxvqSjyM0ST97PczHmVYQn4odL39Gj/PA6dgducxlE0yaKHWkvqbnZGnpujt2rn
XC/jA7qAGPG1+9PqGdNxJ/Sn7tFIh64NTr1JDxrNwBxbN4bdbnuWLEjsONDAji6Q
Up6ackFdPE7uv5Surqf6DPfoCeFoM+VP4Kd0fYqTs4UJh+rT2Ds0ygcSA40pmI0l
DqJmsPPgEus5x6xu9tIkwGIk5yQQfm8dIRJWjAGRNPscj9QHAtlqtGGHzFnxZKd/
LRXPUuRmFVzsodmnVofdBBswPImq83KiiVWF8si2LV1wtCqY9Huxu4zQee8GRbIE
GcI88fmW93pJJ2Yfir4ok0mrFh79JK5+xS+x4hq8ZBNAUBch33yNgJmk6HBDf9hN
gp+WuWx1G/puNqH6p3LJq987q8V5sTm8egy/ebJJLHp4XPrYmC8WGaxTpxPnKelz
KXhL3yQuTG3d/wkGup9Xd7B5j0WwKcaYUjwtzRXbTyTyD49GlhVUPZxTfszSsY3r
GMb/3fO3uqPYwq/ncpsq7BGm0MIpf+4eF9mHsyqWAazh2rVBW0M0Y8JdCG5tbqBL
4i074lwvxgmsL8NSUF2hpPyPr/8Rgo3gRBoC1iXpoyLR/UPdXsWzcC7nA135y3+0
t/5FRudbGRoXxJZEW11YL6/DaLvtzxvXAOCktKSzU4s4qi0PUgebwDDTQsww9u7M
QI8AJSFb0DFf+CpkX8m6WmG2WY68lC20rT3T/8tM+xGSV521uMYt/Clk1GGvvh5B
2HFOainPacKWO8XUOV426arxC8EhytZRxQlrXBNaDvAzxTWCLYmHU5vwvl5tQQlq
XOAP00gRcRuSbLgfaTHt5rZnjoC60ashfrgPa+M0M4tOEsiNu3v7LxNJkfRUo8f9
++BCJZ4zW79Bxib23IF2TX0vapNBoiNhJIq2YXWCkBqohBgECh6OkTzg1ZYXQvGq
nPskh/ubt6r+W4SDqMkyQOsNC7kgiL78WyiXN2BsHJJGDbUAoa3l/4P2lU36EroA
YupmCmA0cxip4Gzl9ht0KD9/gLpLEkKXczDKSWoDZSf5n9CazFoCMkruyc/Do8zA
XBeMbwib6k6Z1UMGc5ypxGllLxI/ii+yAK7lflH0KjjNHHQXuWCeuqQKZCZG6LiM
Mw9+EmXF2EwzbDwOwccuauwvYhriuhiZ7RJubAQA1G1dmoJIpzmLQxwXZix6ubme
DbZ+rq5h380+PlZ54fDGzGrDKIN0Gugt2/JlD4YojyY/4BSTY98KZDCVqCbveSqW
YRrffDm07sYH27fEz30c/amGR0+r/1wrP9++8LOhYIC/Xr7gfzVo2REs1me8EWov
LUwc8df0Cp3rQld07ZKVrRSl/4SxW1m2njBnWirnXgN4mD5W5RyFCbJxfl2ssqz8
qSvpdKrvaFXba5lel2JuW/FibKcZ5GEi0gy2BOuwvbQHU6H7N4xi+0Y7CU44Duj0
MEubsRgF2lucDPOt6pLsl6dYmEf7XeFg+aHEhsYvQXQmjhynuCJwm5dY1PMb9wvq
ZUi3kWk+U112zTH3umXFOp1n3lU493wUa+MIlBUjpsYRfpGhwUJGG9F2S5YMCScJ
C5B6H2aBth2RhGAGmHryTPeVOni1tvIFeYEeyYokg6VZmdJpkHkkZguNBGmkObhG
bPLXDnbSRh9LLR6aKt4MtOx9VxkE/i4YdIfrcJmCoQmRaflfuX8IZtDs4SPnrVk7
SvbG1ahGZlJBc2qLjanmA3W38f+i7K+UMPh91yC9Q6SjAjbPoOXG5u64DVvJzrvE
kXZe9PASb0P3SUCr354yqwvXFQmdl8YTdmPQdU0r2CMWWqy+8G46mffDJFcpKcJY
Rsg0DxGYjFp1C+CEMvmpl6+bfV6pjtN6nmu6oIM575dciU4xB4OCtiWJNxGwVrmm
yfFietQCVLhVW79oWIR4iSQgFM4sf1qWintOGerfiINFYh/94FgijqHbNvZknB/E
wlCsXt4YMXzJRrjc8i6cgpstPKtU+p35/MJw/QmFsuRMuhNhmLU0rjqKCdjYh8Qr
E7p/q2Ei8/EzjLUepIOyE+4oy+w3cGzgN+08k8xfXgvi/V89IvLoRoBz1VP3BfEB
Ph63g+Fqr0ieIwnkFP7n6TicTBbgU2RPOgnR5uvb+EViXMzg6B+b9bgvDuWPepVK
U6qeAuiaZoRii2Z494HUaZei0uAsnqBYlKFkmh0E99sdBmpkLeewDOVfzoTisCv5
/XItbOMj282bGtT3j9jlT6DMG4SR9pVjci12UHNGq3wXR4/DDSE3GE10fIGptXDA
J52JovyhAq78YncPegYbmOx3LIy0J1mMPorr79ri9Zsf0OjHuJxHcKcRa+ud3Yyx
/f4ALv00IppHpHAdEsXUftKVgbesgZE5yV+eSnayi8OzTt7+74qWhi8bBGiIj3K9
JoRnmP/PejSWLptWWL+4vM4WLGlV9Q23kGvejXreOJWnpJ5xZxgm/W/S/2w9rM5C
cagXIPny+JfL1MRtX1spr8ma3adSrXFbhGeDGYH9OsvK5BqJyAvTGg3K+ImSvWdP
LpyA53v2I6SWLHuJhdIygz8IV+ZkTkYP0rKTV+Zz9O7z9+9ibJM+cPKZWRbwH8HM
XbwMwL3qmLo2hcLOSBK6rZWq6yebZa6WCr+3WKgjdC9sYD7jIQZl8qkCslhzLdQq
xKSll4RdjmQGcNAohCuo+nO8l/Fa87TibUUkStazoFfOxhAq2Zsqr8tudk0afkaA
CU8l8ymaUKJ8pHQQbIh86e1X8D3MYjDvk6c87JJOGx+8BcFUUFP4B/oxkq5eDiNq
IgaSLgHjUdcuVww70+2isb4yDblUFbpA07k5OoQwOr7yD1MqL6+/OATSs45dyitS
jBC82mb8enaqQc1wpzRqdPsMCXM516CtzNwWPPQxoVZ+sRPmCDf/SGwNt9UcW7Yd
k4eSd6NeOQob/eXghf2qcsMYWxMGrA6lbENwaO732hGDwC9/QWtaXJCXXW6UAQZU
xWq/iI+SzwDSGBn+ZAgc9zDKjbJs1CSiX2M7B4kA52HB15IihynC5e7tmy30855c
Ff4Fm5xBBiwzaJPxvUsCOick+vrA9LpU7NEAWEopxJOL23phXWdfKdDI9H104eKA
pIC3V/+NGbi2N8sNzei7pdEq49eIIOT4ZL8nvh4wjtw3Quanis0E1e3aQHW+FzVn
jvIygxCAONrFhGYGk13j1fDnl1KNha9zDPH7AWXwwkkePIhbMI+MW0E5UVOD2fRs
w+a9JOkS2emeehWCpI+tCnyNi1Y1nmQjiAvbON3pHZQ8dhWs9A4Ad1x8iLOEkibS
U2EY4G1zhu4CMGtQGlwcHsvTXFppaoi7xK6ynRGiUJtbKtSfer/g2/X83PofIlIN
CMpOc6i7JYj3iWmxSugPfWeA71MFp2bYqN4QIZM0Sh3GB4OFfCfEFO9u7GCrTIDa
csHuCLldAiLIoEwsZKmvtvhb8VmZ+Vimy1l5HGwfILNmRsTs+EmMemxKY91Gvckv
Zym02N/pPJMwztOA88UP1WvNuLjT8qcWOHYaFAzl51/VL03DZXjLBosu1xSMRn2J
fbAbXLbgnq656gmrwinPbXsdVA58fkemL7+oKJk5m0MaPo8RpP9RIyGkh78aVrxV
cRu+GvIxHEshut4gweiyvZihFjUgq4DqNvNE3FQ+hc1brrWa4ifTQ4CnxVLKQG/O
ChuxwIMDAQSGF7WIh5kBjSXMOdks0/tQcZreceduoo+Z6wp0kVru6Ql/pcBjFTEv
Ne7bAE2yl2HY+b1/gQ3LsL3ZfKV0o1W1RXrfpIP78PfzquGsx0wzoF0GX46JnESG
WvmBJckVN43pnPelu6Z403h6GP+9gSNCpjDrNpo6ZIuJpApcTj524FV/j3Vp26QS
sr9R3PAOfBmGCgTr6gfLTRUnkePosMVus/PosHwFp1J6Bn0Ug7ai6fXiZrXjeTrL
mLApyfn99XCyu03l2XsTe+4XjnS3tRR2yqiQ6+j8h2PM7zHsZLmKuAjCDzXz+iWA
yY9Dd3DCVLVZh2t03cqwO0NeZlpnw/a4TqV7bysviqNGLjeAPHKeKan1bMlJDixw
D4MFqU/pk9mut+wl9ZXBtwY7vK0mCJPaQyu1+AerzqZImMw91LTyP0M2Cfyuz2ws
dsJW3wSx4SnSJimSNbYsmxgy/oQ6MohkO/GjTo8u021aPAUMioa/iO/LxcS0oKup
tuB8bBq30pcwuWYJ/ckWHr6/fwsM2fa7ZIkM+ZJotxRwRKzthjxmeMmMXpQ92TqD
mWjQtY2jIvLrPz2OodOArG9NWSXqdVKueZKIaGSjYdXsL+hzeis0VmCHZLWsIizw
slDw1k3QXBpXGIARpfNqtVYFfeBUN410VW1DB0JVO3GFiyvWYHjDAJpH5LGUqunA
W0ePwsntL7oWAC/yLWs663MfaANqBpQpEblGS3YErDKWWnxebbSKJ23EraQirQk1
KA9R4ixKzDqV3IgUf14pGcOOan4nvFIQ8998qXc5g3fSvUfuQE0rHDH/5b3H9U8M
ic2NPoOGg4bF6hpEHkRYWWRNVo2mxeoF6Xh4JADGdDKo4189sxrT/TjwcznT4SB8
+rgPJ/s8MKumpHkmPEPqdBLG2rRPBFANGlhYx9Qvk1a1zbOt878MTC6ktcQsqbA0
Uevr4DPBpLbtkxTFe3vvTtda3Fohgxlz0YuRxR1qxUnPCzgi3rypOPXF02lb/8Ye
0KuBAF03xDiaMA/BuO2/J9WuMRjp6afYDyVTLzuSlKTY8L4CRERlkE+TAZWAIQcz
WfqHqPlxGwyaLytSUp1LuKfLJq5CVnVFWkdiO7A7WkfCwH/b+JEbz4roRYZ0rA5S
z9SqkH2PRsIjs92O3MiNbdfNVt8B/NEWuHS6I59bGzObwRymqiZXRkFyy7Eliedx
Y32iw2AkDrFi4KkOywnmaDW2BZ1vjlEwQlS96Coy30kMVSYqhZyAZyMonOLZENwB
5wSlPZbxLLZCNUq3I9amVWD5ge+7pDXiF73o5V0p4OCvY4HIHELyGU+4CqVnDOg8
ah7sDp+bVT44ebWG0GdcL5mhX95b/0PPpruIhyNuKIMVzLsWIwUcSb3Jn7Ue4S1B
OI8G2PF0fJSWE6OPZMNrCANoDUHgJNgfXTpvZwJ+z3mXywQCYmsBenz8dBpAKWMW
hg39UI3ZGLk+c8BxqiEqtp6oaSJdsxTPlgXJCM138B3617Cc8cgDZatcP0u6XSHL
L7tA5H9+9HdNXlqw6lgvMz/xZQ0oLvCfzCKW9C9cM8gRakY5ccXCoadby2F4+dpI
aImKelQ9crYOlGu4LAQS/slJTtSSpun4Xb7JPS3ljArZfEkRN00a5eQh/9x5c+7O
dJUKVbqmTuo90RRo9150Hf4Z+xtUZSeL0cXAfMvAbKM9UavHumZeYEx1f0q/QMgU
QW4BowU7rFy3MP5vnXhasdL6+gq0O1rLHJo3MxxEaJvYWybZ70sPrbaFXY7qsPOt
8vMfAsUJAnW9vBQmEH/3eHcCIN5S1YX2gz399ZDE/Sh+b1T1unV5l5qAhG1GDSk6
DOY2CRs8q7/EJJQ6BBYEM7E1zbdG7sH3JIwFJFoTVWsIwKQQobLrgKF6yiF/k6Pn
2IlD63uKcWO3PiptiFfWSHp2kZxXx3JUE2Tfjzo5ph7SjkHNPj6HJ4BlgAjGYuTX
K+foOnM2AD+Tdyu66cPuAq7qYABuOWSYvuoBsRR58PCBpwFrAX1fbP5sw8JRdj0e
oHtwc3buSkSwl+fBeDIqf1U79yqhkJkt3LVMVAhg00hYf3MHwB4/LPm7qTeitdtX
FxAtQObjKWszbfeKm9/I1ir5vHztL4wsOej1mvaZAxEFB0xt8H6yPUSkuXsmws1v
agnwwF7mipQa92CnpBFMMgWhUTrXv4g5OIEw27+PPpk8lPkN4czLVQRyPJ701LWw
CNNdBC5ZerOG/CqYGN52SUFlhigL93sjOdKljrO7NpX+aXYfUkBkch68+jiEv/yT
Hvc6leS6RekDkLsqxPBXcmCFnSwOVV7RlwdSIk/6kuXrLRyHBCnFEEFPVSHDFxfY
oncSu8MJEK0BFqv44HsiQCkwUije+qZB4F+wnLWH5y2k9gnsOVxuryCmq9085JTw
bLPhMt+jtVN83T7TiOjtqNusTNnJiOOgvCFzz88hDvsLdYo/faKuk/wMLO0865Ur
OACl1CtFblkTPikCHmaqkTAC1yJG/7PyUmwQY9PdIUMq2J90Nt/Ck9bp+WPo+34G
eLitLMKR7Rzm5CL38xaX3E4SExfzavP1dQlbNDatI7pMTSSYkYabusMchCPXD3Mj
PD9On5bt05z2PSb2xuyvLo00r4XwrMcIYqF2HuGaywCJecx//pwB32BRss/m1Mti
cfBUipykOKGRZKvEss9eG/XgVbOmm2i6WsuLRAS120fPu/CRyOBWCRuLy6kkOi2D
qouNKC60lHcLpy8ZoWi5btO8ICVppjlDb3Jj9Fm43+bZAYfOqV/ib72jE51+EFxf
ObeeXQH7D+JYNex6FKwLxwtHCEgszD9+Mml/7MYxSDoa/jZj4Gd5RjU4S1mZrO3C
oOXWY/5yXhc0Fri2clHeKbeR6qOQs6/hrKYyoYTlm3ETVUEgUCbESZpuZbiRCwf6
CY1MpvvOi5ZslZFE7pTw3ivIGWAXqmGHo22dXscrBDuEa4Qf2X2IQo/I4XWwKPCt
cei11cA6nPjjlsz9XKYGa7CUNqONPU+yg5bUdUNzQ+N5wXNSr0+GN2e50S49AZpu
umA0VpmF0whkM4IIxojBDa5hfzydT+4IaeCmhJF0WEhyFnS/y/ItaE0r4hF3QFXU
svDC7M8qzloEp5s8C/4KXDV5szVLBSdwlsi8Xoh87IfR5pi/zmSVqq2AaihTfzJG
r9J/KfVUxzuj2rHH95NVii5w3ZJKkVpjVrIcSprALISdG9R6ZAT/rnG/gKhP16v5
3/sqcYxomGUoqJFpWOqzpJF/u5Jr5Cs59oxDF/JPCi9T6L3wEKZYCUkyAyuzrk6/
Jupc2TuGpe9Utno600NUsaxfXP+SI/wQO96dkqWy6jsYg/yyo50mY7JVkoAXXzDc
MiDNnDU0BnoW040VUnfghx3oq9nkJE3eFNDgz3sOkNsIsHaaTIJVGIlAxcfIHSWt
d6Xv2PvXstkm3rELpAQIk1zWf5GOAAPjpC1c32VuhaCZmvLcYs7TZNEJc7i4eepI
vUtI9Ql/jJrDbR5ODLXsRMqVwFqetFFJr6/P4gDwTioYRSi6dQDN53dAyBEP2a7+
cxSNekPPttmKJrg4K0h9RqCREiO6BXHtPmrsMhLejooYKE+/e63RNljTMCElFBvQ
rdSPlUXRdHobZDDc7o9KkVna9s3lt16zsSP9nDZ8bXLMhXLiahlUUYytd16+2B/g
l5TLIgAPiV4UarpSkqCznM3pdrxg+FCUchnuOae7wDnZp5NNT6vQuGZSA+lgwElr
53wtH0vjuQ/25kQQ4qZKYuRrrLxwR7h7tpuP3aq3OALN6XZ5hIdkJcT+cXmGB81Y
zTYTp56QIpLN+kh8NZG6SpAva3b2n2a8gWOZW2pVnwMOJSUGtLo/VnfqNpB3LoNk
NwzHTitGm4cxG5ZR8tMsflWvt1Hgj7hvNwDq8BXEFBKroMxmuyl2TKqO4K2mbEht
VORrBuQdvfqZfMjoMkRXWelJcTjdjn4l3H4t82Gyad8UuVZHbmlktsIOczSnAq5y
AKnghqRQcDJb78f/3NCc4/kjcpKK2nw/2nLJ+jvrcl39D8MFf8GRbk/td4Slvmnl
9m+Vwsm1wfZb2dzDJD5Lz2ZyzlfuZi5WKKS3IcPq271RiAT0U8yf9rydo4uRWl+U
xUeNe3kYO6v9hw52/h5UIKZv0l5ujQLy20nll4BsPTNwhiadsexHkDysyzpiTDDJ
NS/yva0kghx7AxumG0hjqD19bZQnDtgTEdDG7FS48H0w7PkuSf/3rsVCmI/SIBDQ
mOyJXzC1BfJHZrQ732W17Mi5hbYnA7gduFLrTbPa25IwIF1HcQLBxtj1EaspUZm3
ODJJiQ3E9tA0OJyOghq1Sm1h5OexQiho5/mharchEPwi9vi/ny03aQx7VqOf3cQ7
NQx9MScjm26H2ogLXGLdjO+ypkStDPVGj36G8R70CO6EfSYZLQ/UPySfAK5NgtJ6
2WwFf6GR1XrP2B5hSw0HIZgyUoOriKyIxIUpgyxPWU+5JFvyt41vzuWePzo9LHFk
AA9e8on1KVi2vEmVqCB2rBHNLWd56Hdn1q3W9k633tvakSWCnEP7MFFAEAIkdO1t
sbdH3TZPk9PARr0MdqyTbgmOSJ/QxFenJx9G0B8nNMDb7EYCWLRGvMFeunw1fN/C
zYMZVOqwGvh1xV35TWHnVhw4KkK7sPq8ScuJ0EhAD+M0qej4lLPc87HstcRxvfkg
y959Ng5eBVb3y9gw3cueal62a7kYfNOTABilfnTNO6oK2mf6h5vdIUxjZt1fsufT
8endGzT0jojo2HG94xiLX44nkncNZPM4yo1ywr6GDv2AHkUQX2c5fpF2s/6SjpcJ
TfXpOi9EQGt5wZgk8sO2UpyMqty6trWmo2QdQZ5QKXIPcPkCWttGWMeVvNpHDPiT
KhGEf4ohZ8WOhPswnaBnRj18TC65jNqnZX5cjMpnoVxCheIgS0T+v02PtKqlCq2Y
KVsQAf9+pYxNclWVYn8nunVEBmK8y6HRClkPnWWQu8sjSLBf34g93YKCXB8hO+Ew
BU/cXLXL/+pNjBYVD2TwSEa8sTQm2e2I3vOYe6rMIRVFMTT595DNBYbPTGrVmps3
TWSrYVP310yKK1+OlOX3HoYzpeXeFX/w72X6G7IWfc248JmVlNqJzZ77rt7WNYxH
AvK2e0OD8zxAjc+JnHTbO9Txs6QwnOZgI9eLJRarePQ1lCmZCpeLNbybamCjRvkM
Bgvn1cBPLYY/z98w7QlsSR9Nw6eI49Gf6UwFl3ldSBv2/Nk1G1jNDWCQ6L1uatuR
6/8saPGXNOq1I8mCxBKyryt1gJjqeCpKwyet1WP/LnNkByUgDoM8rYm0B2gBuzH+
MHS1QjPf5EeHtlboJiEeQcqxCL2gaaEsdHvmIGoupZXdvlQfpR8ROi7oU72SlLR5
CpC900qZRxRSWzo+FfJnageg0WGYiQywyDt+lRMgH2GPw4VDSf1oQ1SOeg4bLMpL
KQXQcfNVdr22zXvunQ1NmEmlsFE53LgPxnSnRVBs4HZBblwWLDXVtTfB2xX4xh1K
nm7zfMSjYqRUr6SlhLLgP7quAbS64rGz0UhdXFomKQw/U2vku2Kk70b61x84XcQQ
hq/+iFEtS4VqwFs5uOR7K5qS9hiT3l1MGcTO4jO2FFU+pjZgu5sKDtMXlv0Ambqx
EFpD/UmYeS1xT6G66UQ9rHHToJX69lll1/6+Wwise6/pnnf7uO10C7URlnJo6CJB
9xWfeUW8XhmGSMX+PKW/8GR2CvIufWrfCAPTWZf8YRh+V2IOCjJQ2qlPCtZftyHr
9e/k3FW8DnLAZyAI0yq0Vsszi+GzoFOkEwQaraq2rYfa+kF/akkFhLBaZkvzP6DT
G633fNU5OPm44B4HV6uxqmKOsLGF+LhBhPyjf9TwzNNR9H2Tc85E+Ug7YBzYsdbd
gOsty7aQnypoftms6eHkJ5dMKZjuaxyKVZjrbDHY1hsn9AYxSoGcBWJXZaYFJ0uo
2jHxThYYCrKuaxvkLJwVXDvaoiCE6vZKJ0wZFGQe4ekM6X/OKS6ug5ZCM7NjGP5i
Do1sn3ZLcQd/2i5QmUgvE4v8Brcp5DX6M0esWFcSQycCarKq1SuY15VpFHvtxsn3
NiJLb9Wk8eTDAyE+wRiqHSbW+KRIMXZhk42wRGR2IhahnYVgTUH4NXrjlCaRFry/
8AuvRDv3e9UIC9WnMNSqvYw7TPZi75AVRNsitrDtsdygvpSUmSGbSU9zsOIjUp+b
kD+oLsz8JvpbvCSxBaPOVNA3vcgvH/DYrtQ0euWd+utMC4eiU/gttfijH6eKK/Qy
Mostcj8NNmi0xcanM97w/eqseBeKyXzWGFpeULeeI0/KXHttG7OKiiLug7RAI1Go
jqTNeVa9Fp/ZqQ2fLQP58sGTYm8YfEAbk0vuP6zIajjiyt7Nlj67f8GEvR3XbLMk
6bO/U2QAvkgVVgKZMQ3haFjulSLwJP65vp9UvLWJK7N2Y7oKYdRnhvJk+oDor/rc
gCz+nADVV3/qyz314i/s7Bf7u8du8mMC105JIqDzg0DNdSrMdoUg6oDRln9V0p85
cwI3rNzaSt6mu2tUQl3/A7OYJTbBnRzwUo3fy3oAoAI5YIyQlEFm7LTbbtxs+6OV
5rCogqC/lpUr37LAgDjXnjBxVxWnO9y22BDa7H+CJLdGvZ50Puw3OT8i5FtIDKlu
3MVvayBEsM2Q2L+ItXJwZOwS/HBzmMOX885P8+xBnkE50Gaso2CygnYa49j/mX+n
ZyfM829wuduz1o8iw69+TaO6KOb0VG9RSutZ8uNgxavD9Z3Bmsho36Cs0QNaQ6o6
5SqtZAovP6qHrAXLJ5JUl0GWY9SmigEexXW8+/8dM7Fo4f+G0R60FG8eyhHlO6Eg
TXlUGcR8w7YRlGbB0AU+CYS/33VrYnX7w1nMMoT8F79TpciVOl5ngWJqvHAUaWCk
rad+CS5/RXZmutrnkJqx7SpZzqzJpSgHFee/LQ946YH+aItqK50M29gWleFVftI/
AGWXVkrG2YOaDUKzbmhJeTeO6atIW5rmE5zbG3YSBUo9+1Y9x4rYNkil9ZUUAVJs
l0Q7+czqqtvfQvXVTdYb80oHzYoLMPagT5cYCgkUTtRdQ40h8bvr6IUinbqq2M4f
muDfIR/EbFl59vDYoq625O7UbNhqYROYppOzetGZ1KSnpKUzPzxEUBspbkgTPnkz
FGUDdP/mP/UqUl3y3vOmryJw7kcb+E/RRmdUc8XeIRNd7KBOIb58HmnyOmERXZJQ
ygiEha1iU5WFs4SvkeMEbZPP+H09M6HPk48mfP3ExGctWsTv5iFHW18wsc9FhAMk
lbA69dPAmlFGajBvNCRl+Wtcbt7Kv/e+7+Bo7+5eV4rc4T/xb6FVyUFJfAG4T2E1
eQhadp2eOXYz8GretFX+dLgB+tBtmexl059VMVJPjKzOZoMskDBp7uyAhml1M2yh
nti//D2R2+w7Y0JAfiEQlVTLdzKqwajVIWs8spA2wgge0IIAHUmSTlm+pZ3GtQe7
tfabci2FI1N+v90ZDoNt0nqaiM5VSOYL78j92JG8d0r9vEyhtGJzpA1OYB6E6WbN
VFGmh1/fTu03xpzUa4zXVcLLRLosQVMb6n4RfZG1vw/gl/aU9lK82HWNdVzCTuhw
7qksDDmsesVRaC46NVql870qrDZ76m1Jer/dD25biTgFiYxYI9PqJAlHjhRE4M5M
AOqRZ+CPzfVxfmQySnP98uK4IqoB5I3Rb16RMKe5gh08tWAiXKbF4v3T9lAm6lcC
Hwp5BDUa5yQ4IwEVbpSSfYQIzoZP4sGXASa5g/mGBiFFiwtNi2PBZWKUj5Ldh0fV
SC5GyRJOTCNyJQnW50of+lQjTxItKYcGFdPQO+DgmB3CsmEFJq7IwrvyFIpsmL3/
9WcPMFIeiqi+JKv4Lsw0cBIZNjXVhgO0Os+MsK7Y8YGw76sEChLirUIQWZgUG58H
rwzxi0XLTjX0/xNmec6tqQ57M5N38DBkWkus9CzX6bTbzLL0ORGIsV4zq9e0IKtq
hQOX7btPhBRSeXTNE3w8L3HuQEzUisJvrWit6HZ65VyZQqcEkuTRRu+SkbacMToO
gmjZSBlxmxCpNwFN+EKrxv/8WbTyT60s2+rn254aVuIeA+2kJFhMOd+Fhjj0th8D
rRMo2Z3H3ZjrONl6WZzQJmpf1PcWNXf2bATealJzvhrWGI5XHh8xVT/ite6Btg+h
d8PD32xhV+jnkHs4u1kcnvssUlIgap+vQjZRPXJqIw3+pg72qqmrc77FEHGeq3KE
G38EZqG8KF9IvaGzxu/l7knYJ6vy1G44TVltz2wm8P0vsZwdTyb9pwqZlOMrM19l
wcmH5tiGrhQYxNEXxNTK1Zjx+v+Vt0e4uhYGwU9jWN67Eu1Lniqu6r8DRhaT4TVg
4eKhuOsA1e7o6a2HxnXCqHiBgY2CFP1ls/5nNmB6IwmgH29SWYFZtp9tGLoQD32A
frg9BJ5DuT3YqkPyX/xgv2AG/OnEb3CqBztE7yWgF7ieaLijlpZVfjSoJWiOZ9o1
4xOHu4xgPLcDtcEx+ririkzicj8zMF3rrXYw4erRwYSAKqnxg6TvkKnvKzLei9Nk
Rrn7kEzt+iBI5KUyr5e+UcpnQUyq4WPJH1jl4uINEkw9M4MTGxIuTfJ8IPEl53Ba
wOeMVwvo4Rk7M/XHGEN+GO/ABA1T3GOLIRNu2oWmgIH2qw/DhafsunDneFEhRsPT
4N4LLH1G9dkc58p2h01w2FaKhDqD+6rYwTCj6BCMukl04HBkt48G4DLk/aV/e4Rq
AoUxuI2cDpb/soy6D1HvCbX2ZpQb+8asru6XfUK1I8/xMvEDEaNvTgIAEfF6adkX
E4W1A4eSbDLN3Nd4EUz+LhQlaVuS3Gq83x99t4lAw4POyn3STjdEisxvIKdAneHB
VmPOh0BBUQokPU4LGmtR+qCxrL2LxdZXyp7OxAZqCP09bw20K0CICkNL9XvBmVxT
qgDCi4g9a5Rih5SNsOzFoAxW4gxVkGjhSfLG7FJv29AFcQQOZXKFF2xDaWhYPh3Q
kV6zwWQrmK6Clk9RPqwkZk8Y7E8YNZbj5lqPWSp2CLOIwgFcwWR4Mo7Tx4QkHYA2
QYA+Cy5QTq5RJdmwuD1k067aHuQKRFv0+TYN+KFgYWCpjYMZaAYAxlCWkwbx/PPJ
JWx+TDPt4FLJ2QI0kuzS6Uq11Sl8iVM/yJdUs9DBsETHPx3ehU7FL8HNTbgBfDnC
JOTRhr28jKCPpSqhvf/VfLtutgtcGazFcBTirust7S69tPoF5UtfqVjM5JVGb6Zt
DJRImElOZsmR/ENOIWaLT3+p1ir2yr2aD5Cvf8z95We4vpMzkKnGAElfdsdBTaru
59jDu+K4Lqc+H3JX6BWYRhmlWYd5iTbauzeZJ7MeYKFlwn2qwNF5O3jDR0vo0ihT
lj/cH7GGSJLSqoXa5IwWJ0YZIb5UJDsq8HpcmFaf8vilkHQBvh1j9AgmFWLHIrV6
dI12/N5l6B5vqET0O3TaMKt+sgbwhACfrjnzGq1XpyWtWO3C8LYgo7tPSS+oddHS
5Sm45UxBO2zBb2CCAIpU2Fa1eA5HzgeMbRWfA+DJy8j4M4WNpGpPxYtQUXWTspHN
6EgcOQaIiWO5JA6zb4oHfk4eFC0/NRlLx9qhvjVlMZjZQcpmG+R5+yth9Hg4lykR
v++PvrnVsX4pt7EYGDmRMWmMkjWN5tz1jD4deZ8ozB+OYU2DLMP+eo3xb10aFbkZ
vQms7CqgYDszWfCp3MGvfJjPPuPHkLiUsM/SafqCwyspRRc31KvWvecFX+/Ulaf4
g3lI2CbFB4zxMalJbWRUWErgtiHhxfNwwaTaPLCAdvHlN42TcuNT/fjgVd+gy4Ti
suOzyscfscyWEWCi9AAPqdniNNiV/9SsccPA0mZ1DwDbu4mDtLsW9+cnduIWMagk
m3uCuzE0cphxFk4V1bkgLn9vAiGT22d3/AK0IHi3HbKUvPPcMahUXl+PKZPyb4ED
eZfMTcDDeT4FUmStSgNAN72hYloQGBKWcAQIYM26OApySp9YdGsl1a3Dc63rOqt3
SPMNqp3qmR1+wpLIEvnTIBgXUb6OW/BO9eH3sT4TdnDkFr8wFSxiADHTCjv2WQXR
xnyCV4I2jY2GIrVacFv7GDujke50E18BfVNZr7I70OPyzSgfVm9wBsWLF2CWQCDx
furhmJavByeCts/fjS0HrSrtGDIrNcqPgvso+snKO8dTmLcB9nJiBB98opSR6ydc
fEeE0vGALFy954QYGtSv04nibTcpZPLZna9n1JGl9uZWa7hEcM9i16csjQ1StJ8K
tY4jsOp5vYUf0s25r/+yba9lRTECZrmk83D+S/8eu1cg5dtf34KqeALLzA03TSd8
cyxe8g51R6hiW+1knKPbs0+lHOt5MstoQJ4A6wGzdB2E060mLyh+PWOWWHFVVX9k
/5YwY6SzSieuZo2giVYsIoA++HXb6PWB20fv6gEScXcImyAXDgFsvC7Zg4TBPlEl
tnSG9dGf303px26oJEJ4uTrQEJeNPsAiiSAM0fj2S+KdQAbqmkthpvyibmfRd8gM
ULPej/VXxFhp4xDoS+qDBNku7wLNTnf4+RM0oSD4Fi8Qmsd8F5c8P8bPhKGqNh4R
KY80uRG6XjQb6p62V+DrJ9/qdns9AINvLJK9JkPpULEalhzkCzjMdFN1drxi4hw2
lP7qKPr543l9m6a+xWL/JxXrdjN4N4/UVLP3euDD2sBQYs+jAdsglrU3tD5im8pE
CZudEzhaNox+/+z2e4ryJ4/SYrTBTL9pVi52cD9ZDPZfsBE+n6sCDA1lprMFLpUk
u7L+9Nhbv1S0MRx3zcsYa5atM/FvuZVGtSlzMBbVGQidAgMaoiLLbx9sVjzH9HiO
6p1zvRDWk5sdqMjHRRJWaCuds1XqDj0J9oT3jgSUtzLdBAz+DGiRScKEsznLPUEt
RJpO21ouANelLOeOZmkX7+8cGQfjEmV67tThfZ81AmdjxX/4v08PciFZhseHsPkO
tCalCemxXDgglplQsyzB8Gf8F87lAPgECUSL6yWNEFZwJO5sv3PILb8VGHJFGAUt
J/OZ0gp5A6fcE+5r/j7V6UTIfPeGb+MHwZUts2fi8oJX0JRpbHBEDIffiAENROSt
BS+7CdZls9T9j07p8X3zc/RRB74iwu1uH0DBsbh239NjKTbpRlSSowjOHn2WOfxA
1JfPQ5SRQLi+fBgUQhdpT7wX0LWz/8DC7ygpriyGhC52qaoW22ZgBWiAls46BFnJ
GMfyQW1yapA+PeI7Emrui4W1y9yhspfDQcqyOCLBM0GrFaInKfnFg4VkDK4x3S7P
jm/aVI0XjJDEVusPlhH4bT1PPVkk8HFBrk/lM6IvTzRVshP8I/+7W23bQledwYZY
vLA6Gtz9KvQ2DjtnrK/btgEXJfugVLOmf4fEon58m4MHH1Z/4u8KkJOMP+KCmk+y
7tuW6rvAo9OoNbDEzzWQDidiAUPH4FPQ7AcJ+anBqxs16g9+hi4l5/FGLagRaTsq
h9mmdVCNMWslb+78W/rIIu5JL+SoBUgdmAGdPhHr840LB2WQ61kzDWVQTb1yfFsD
BIspy0ZidsEDzcKiDyZoNCNbF3sFoK5egsIWMmj+TtymOuxceb8rViEpG+SQ3Ef9
pzVo//r6mMyaZgyaS4GDbUT4wz61WIa8yhy1SVam5XnQzdkFe78qbGwvlykZWSCW
wyJ+BQKhjkJwHfedb6e5vMY7zXo4LjfZhOq5G5WF5dcUbEbdttK1eH0le1wBQZdk
tClgHG661++bjKPpre70g2f8TsmSuJNprruQZ9gZj6RWFNDHMs6dMK23X9e71BX0
bHIsKPHTih87LlzC5WKQkbGxDVZtZiXDPE9N9GePi46tIxCdkx6tXH+SFFo3Orul
6j4LqTqL/IVQ8mBzHBG/DK0437x6AkkN59ZEHKYKnrTSk2utCr12/vbU5j11/g93
xKzMtsMyQj6aKCU7UEkv4/HTO1ybYy3LosDG5IF0O2vODms6A+IhR1BK0ImahpPa
QCAV4+rY+PyYVFQPukPF4H6M6Y8Aatsg0go2/5hpB4x9NMQ2kiok/h41e9cMyGLW
UkDulTldPYb8/oC/WpX34dK9NbrObasdilhfcWA0TL2fJ634K8ULJyIYcoNSFDw2
dVxG71G8AC81qGmxo4Y9CKu3DNTMNSdqz10wT/YmatvaB0+CfsmYkFvtFcVd92Cc
T9DQfGLASSVzOQg0wmTOMpPUFZG+IdLn1c9u2PULyIplGibBbFltA7UZ3lhxAr9b
D9LoorqunBzZn4jrtBKLkixyXz4p7MDbgVpWaWLx8v+b14yOl6+/ZtH3Q5Y2pxyE
cStoNusi0NtGFSblx/VK/yx0m4FD21QNLhmoKCM01OvfZIFd5gT4KTkiy046s9qa
DA9H3r0iiLTrcNooBLvIm7TNb6N3cqw/AeVCeCCVQmTLZcWL2eZVjMHi52eBMRqc
50yzJr96hPF5oFVhXTuPySoID8oeozZLHKEE65X9Na4ZWJW3uVCnP15PAnberI5m
wYqWjoKLAZNLiP0a1yebVRTa2+IUI+W3QVWi/YeCDWm4HQE4OD4oEfIHvkXf9ecP
+XdOEewXdtP+bvAoXaFlBujE0Tmah1jn8VbsAAz1QGjlWz0KJEHrpft/9/jjI9oB
zhuYFmWe0zetf8w+pYQDPrRvojDvj9EIVZisoYDlujHhnKRckdWB8ElGsPmFNOe9
BJ5gR1dZ0MPAIRyucMw0e/KU5HYhK+43I3KgMQ1hVXDYZvz76knwxuEW1h35hQab
FNaJRQ+rFnNqCRbdrKEH7vlviqrPlHwhzImRjdYZ6gbQJUujZslKY1l2mbXxZv0l
nFFFG97cNzdVNNuV3odMujf3cwCKwaCS3WS+bFIucrVpxz+IUCjJtY9/Pr/bs8uX
XOhfSI0hvEDvllGm0VLXhfHDOOOw++DVksRonZpD70PCVyajSnzo3di7/H0jja82
ELYnNmLHx5XgRf0bz64cCAD5ZWWdBbRYsxCkFxOUINTQ8CnGR0Az3BZ3FI2x9c9X
2udYQK/XAfr3bF4MfZ71jLKl9Yyfla3pE0xhGVqQUoD9CaPvuYkBg1o82UMFDAGR
6iSPSrk+yTS9GC8Q06BWxivXJufpikMH0rYkKCr4sLnFezpqbmfJiBtDD5sZHlQ9
XteYUx9+jaMfpzaEtDygCjGfrS0q1pGpEsEt9s2bKFzh/HPblFn2TdY121uX9S4u
Jbbd57/7pNsvBViOA5k1yAfwG7N5JT4KpSXVzs5JVVAJQMARstiGjjalm2az2SQb
jtfC+vYh3MVwsQYhHltpLCImRAYmTTvzAlx87fWxbewd5v4Ar8cvUlZQdNzkJQc1
FyepoMfbR5Y+UtxePchkSx9ug8c3bUPblgYLAUuHRkf0HbZQgWt9ajMY+V3NxLCN
+xUNKEMaUtVVd0JxL+9YEEgVr8EjXo+VTf6h7BCMIlukLcQZvQ81hVslBrRevgAT
N8f0PuJDhNdS/LtBlgaeyqOYBtLJ4XsNLX7na6e9P0BUnzct2vrS8ZaUWGzq346X
ZfJSN6lDzHTqyxUU2wvqzqzl/v2T8IhqEPFeibI0YZaGNo/xI81SJxdRqBFQjLc4
gGWrVHVZ9DqGSGDe50wHAGuZeO4XtmdRLIAgBD9LJlnN7cXVOJFh8bZGAWslDAEB
nh5QQbBA3B5ygO8BqyFftGxv9+M5uCN316WFP8DADCQV52zW3OClArcp7o+R63O5
q+A3uYnvSQAL3Ypq13Ko4NMPjqjvMSR23ddtBUa+c4UaJscXC8aGUwtLsDx+qGG7
ioI0yuGSpipzvT1nU6b9FjI90uP/zAPgHxIwuJvI8+Rs6eNy4TVTbVzOD03sH0jY
yBSoS4HYNQoD1rRb8JjIek1a/Twy55ds0j9PL+OAaPp3wH3d9fYgTDjTyVo1rVdf
jcPTopCYJMG/rx1Zb24Uh8MselYBB04e6arPzhk7pT0+gyEkpf7TZD0hvTEfqDst
Zf559WyrnAse5nsT7OvZuCVohCZ5PdZM4iUEUVe+0KtN3RWd91nWZDHIqmSnkpxf
W0Tf7fLvppHgownGYWWMutJ3FWtPLdiV64nbGjk9F8+sW1jiQD5+6M3ITvW07v93
64f6eNWBP4/ptVeMDTAQUAaGwPI8XJtLcCiiKBUJJYXmMUaH0mQGJjZPtK+SbAY6
3O+bAPwRSfMIoyeRgdpuLHJQ92QH1F1V0sMKdrcT+BjWeAM9XukiaKFSe8D8pRFb
05yDZIy8pAdk6IuzwyyipM3p8ZsYgv0TkFG9x9jTNNBuhzAtBafN++QuR3atDY+l
pOBN+GD/Y9YYI1Yw8eXQ/fCXtzqiWhHD0Lm/c3jqCwBaJnC2+J2oMjPKiAg2ZJPO
ZrwWY0HHT/V3v0AyLvDp4H1aMpbELrijCQ2fZYJkjcoBUyqm5mxAKJ2yN9UFn8vM
YU32zR65LRy16aFbnqI1RxxmPyXP1GExPQQU3k0q+SSgwbFBHusV8bBSKYkLcMt1
5PKb8+X825wXgWGRUFERJ1PAJZ06/iJezmCkM/C+Aqn0G5ml+kbFzMIwII4OnGQn
yTtyHo/ejx7iEU3b0M9ohO6Bp6ml026jFtlPIhdn64AN4w7+8ez8lF6quZ+7fusz
YuJXjYpaAqs+SkFT8/v+yFIFlXd5GxoEOlKHm8FCHiaU9ZqoLk2CZf5JCDvoi6CM
Rqz3elAXReJpjLTKlDnil/kFumJBPVJ5pjqSnIjHj00oUW0i0Qh7ZXoScQ7U44Io
vPfvoUJiYra3frWzvjWzMrw+GvolLs16KCxUna9dz2NWWC9kWh8T+5PXmm2EESPB
+nCENcjU6OlG3awdgn5JxQ6sgcGRZ0Z67VzNIPfDhVemzR159yDdVvIiApqePzbL
Tzh2MQ4MyrA6g2GxsrP3oUV6wewbMgTHoxBsl4Y+tt1v9Ul09nFNTTbtzapIwHth
WYKrCkg2VzuyDdTIX6sYJz487AHf8H6pEjZ8OsotYJdXqkGBmhQ+cAHb5n6EBZZC
BcUkupUfi+h816FJux3dOeiTOZWi+7z6eThoTKckt/CyOeMVNCTsETzG/oRcRp0h
jFkGx4IZ4mJWe4pN/fbarU+BCjTIwiD6B9j4pYGv9gCtJmojgg6qnZJd88JyJdsn
8Ry8DlNUrWilXHs8MvikKdu065G8HIbxkHBXYvJIIWZJ3kDrlGQohcJ+1imsy5d3
PgCUayYx5J/mgKVgn5J3jX7uZy5ymCyL2e8wkZp7TqVAxH27VKJH9+ZibXB3Dq5c
8GtGy4zj/Z2TqbaP88rv+aeQGf0oMthzFL9TCETL9CnalXK4HyypPu433DPSOLcy
wTBmxpcsBQDS/gDlnCPP8fZclU9WshiBp/SO9Smk0/fmMKJljLe3bzwhBeLBbdpg
C3kXr8YOjRFNIWuG3mftUxYBfU58gkxMhgaIERJZwvNVNMhODZXcgOXHSw9KMlHt
fiPD1hSoFM/zFlMFz5He6yDRunY4Wwj9hmaXzc/47Ee5O53IaHbQE+M8r8TVU6nc
EC/2vnxM3OKf3qiAupAND3MjEP1uHgNDRrwZ5kzyqHJ47bC1s5t0VqSKKatr54c8
6nFghagHlsi8fvK9gyS8htS9reCjv2M2ZMzUyl1wqqysDxJ8DvmzGeCAP3x8Mk5O
PcW5LmxaJiFBLt+uA59bBWOYuafusKfsqEQ4nrr9D/si4aiVwYSKwLC3GkUgRwRf
sl7vDQ1XhNN9aq40G7rb+UWGgWtlM5eH6L98D9o/6AD+JXSvxfnzNCs9OIZdxWOR
28VbxMKSXLJJ9NOH0+I4IivMiVpE2khGjTm9ZMLNA3o2u4bD2nnDvC/vISnI8TqW
2BgAgVKm/6V+wlpFLnHk6Xh94wH8n+VPTkPSGetGelU1mq5O7IPQD9tDLO5jxjnw
HqRzO6S4TzK8dp2K0J2UEIjjADSso3lsN9wVkhcksNuC5StQ11vb6qPTaEkgYUUe
uUcrmBWa9cCmXMvamcewdU2s6VZSZEOd0+YDV2wT9cqaRvUogqO+5YqW+7A9YVT8
vSG6eXYgD9h66hAPLRQvAw9vLMbeM3CbGWjJ92YoQnNzMteFL8cuTV7F/9/znMFp
m51UU5eh4Fdd/qdCtfQRZWB+rHdPCKf+65EJAtUb3Rkf0Uwf55/nhzV/I9BvuxSC
YLxvA3ELGybUuRB1X/UuW74JbmooICy0WzjYqvbLYtGVw/H71tnn3twLl+Fcl4oQ
5PD4LQUTMaAf79LvQ+pdpD2uMkjhw9SW7B1A6ecdpE7xZ4MQgsUgzH4S71u0OCy1
JFdpmj9sWQy/CX5sTED+d8xNFdoaSbdRuRHyRErrsiXT44n+649wAeSJIflXE6CZ
U579yCigAntSCd8GxGSWktr57223iPV6Js/M1g9zf+Wqp1u6LeTRMsz1ch6C+3Hu
/n63T/LqymFMasHbRoqUD6czRYAdCeCI4fVEjgFhZNjL5tZee50u54pV6uTD4Ern
LHXhFpNr8kf9Ofl3kqQpadjJdX7nX/0fCMH1orV3lTGe/h1/S0LBaHxaXmwGQONa
pTmoN6066Cz1vf0wIH0r6eVOu28EiRDZVLB3FHiPyPCRRp8b8rkemOl3pMQwLhkX
uexbcQwq2bBy623fyHQ9UqMSArg9dWoFbLYS1sFNZ+GjDqbOCbJzXtoig6j8dq8x
yJsKeaCKD6GOqgbhZNfJfBLlCO5g0pl0EpVeZ2tDMYHtwfNO+FP0IBwTG5qbATTH
yZU4pxz3NCPMmP0uaICxyc5M/2xCW5TLPQVEv3TJTtDDuOAZsX/Jw6VQlNzbG9MG
REePq0o2lzB6nl4gRBP63RS/49LT5LxtZVAeSpNz0dkOub9XF9GE41B8LqOlICV0
ZGcbRJ/0+hkU6nUPs3FnKScnupTzwwaZ1jIDVfelqVH5AJP6WJN4JjHZ3IWjUHOb
L4jtstd9Px8Ciwt8N8A+/ZESRnfoo3eUanB2pxxoRB1/06z4EstBtlMLCH+aGugX
8E+317wZuiBH+6JCIJCJK0mLVz0sYtNmXf03zTBAczLfMgotOBCo+ClrVTCiGmaX
hkzEc5inORmIN14zI6WGkvmjgyfJO9pSFqcaUBF32Bd6KYwUZONtJ7wIoEj4A6Ed
+hBqnYSeXCe3bBjKo9iGMeVDF36rY5KpISqoQtxetQdUy2qyzWcN7fqpsfSS2zv9
iwdD34HTrp3XAX1A4tZDtRiqrxXxG2Of04i+jHLtECK4l23cXqyvwuyQCSS5fz0p
l/ymnFJVbh8i+HyXIma9F5lMO8ZSG/9R9As4uyH6/2t1v+GFiQHsPI+I6jf3ddCe
LOerQk7byjG69m10RIqJL3XdEnzA8G+EETU1/FX2acpyuIpPYABXbQBc/GUXTiYr
8nz6PnDBwc4woHF+Nysh/TZLNiT5UDe1baaptb77cL0UwOf31Gl7JnCkEy+8XBdU
EjKgC64XQ+sM50LpDF+TLmzJzIM6T+C+icRADx3GKCj5EQc4y3x2yhZjXxOuYicL
lq8/y8k99O05UDHG0RsYBZh3EHR3FlGWzOnTACa1/9dONvgb3sU+Ykg/yOlP+5Tm
63GtZz/Cv6/QzL0G7z3ODhCEsr/G2jeKHGI4gyHQlPp37/fQATHwU8ffz8dIjxxf
bRE+pOoc4L2Ciui6Zfo5a8EBZ2otWJfnRAYBrFmvulaERdKsfyVxj5EJPV6VMniA
LpnyDgeZS9sMqplyq7yEP5wha2ZI9ISpZxt4oyWRxuQPM3gzgXCjAHN4mO6O5Nkf
kkh1D/Hf8PJ02orm0XMEEWkf0NUsFLNeAVeGpc9nWQQAjGmbUKe3bNR7BtTx0ROZ
wHzRHIvAmSRY/ox0CFRetJsBWfXy9rRpaweQsSeIjt33EJAVinMW9oZQgJunvgu0
dECbPOsxbDi71Uu10IscXxUyvLnni7/7TV7nw5URW3l7wRmMP5n6goEH6e37hnDI
vI35PecUn9iHYpwnaMGMEK9qsn60NqjLFwUxVfAubW4WiISI7qCSq8liqIpjKjIf
IithYxB3Dj1fYedfJ8LM1hyA7iYoR09Rzc3taZKXlCYR7g1N3S0C8q8wzEpIos/h
MGT2bmD4K4wx+IFHpM646wDLmIjXEUyIM23Xt1bf/pXjCWqyKfCVTmr2MI4Dkg85
K/QSJ85WUvwMRcbtp2dLgqy4F5mnbxTcFMLpw6o3VZHsgyGO2Acj84WQx9mTQTSE
4e6HIQCk41R9VXbEENx2g8+uMxmqZARbnd8eHzXIm6ksLgqbWzXF0D0EWudOak+z
VlKaJkaNNnOvtgwQIbNEPf2x1OX4ylzWF1XIgOnYc5/sLcFGAAFOamQwlHepYlvH
Yj4fi1K7MQHCVLL/4ojc++XMDgIXJtKNRquH5/kKYbJ9RudLIDc5ZAOkDbqCGV9G
d709bjbXnLDE1Sw1k5T831AZcmHFc0loDtzFhn1EKR/QvZqpu2MFKRKkAGpMKtf7
fe/OVc5Z81hGSBq1wZz3/THnn0sllsH/GaiYHcWTHtg/D4IduyHS1CvRC3/bxKv1
n7/dWWn16v/uQRAx3JsPPl4DULOUFvKuP4VdO0bGPfnTSDd6N5/vw8YsH3gsFeIm
mJiEhQLWQu3nYmn9JlNx20PTFEjfiPAPAuwJl/k/3UZg/YvRz9QJt106bY/lS7gu
+gMk2xhMtj5l/qo2jR+s74qmwLLL3hqXB2NOP3Hw4g/rxlOEfcKkE8bGs7PjrDbU
aTmUEzXvXWu9aug28OljA0+TfcsdhCxvFpLkZM0mVOtvScjMWaD6EQQQXdyfXCzY
6yly2HFHHDq8Pt68iVJ0Gk1c4NgfTlTZELcxkfyDkVCz7C1W2eGkVN0Ur1vsuJtn
oDfyaZ7SLYBv4lufIe7CtgyBq1FUlr8+ghKUuLpy8GjXZYXe7c8BFo2w9BRvQW1a
xXggDz21tPUvSTgEXTv/j4thnHM5tBOWGNVTUe/YQ5LKcug6uye0hAl26JI7ZVgh
FTzgwsKPxZcvgUtyRWmDX6fxx7mFIgnazWeIvRT8QUB9CyMeBbJ4HOEWZo/wn0Gk
Ym+iK+2JHvVYb3b8lD4wpdH7b06kCbxu+QizbNhwOYCp29mkQR7eVD65weTQfHo0
miLonTEIDsqh2K6k0BBITW5XMDSGnTAi+xIgZBSV2twWCvrXir9c0rkd6XsTJR7y
G/Za0zyH/JuZpRu0CkrGHtSerSesCk3cPPUIQetyysF9LkYhLHCjf96c2Pcl5IwC
i/0CvOi+S5+6ZGZXpSDMFTd6BeIGRNKXL9lxpXoKIW4MgsrkflCmUhrD0JUJw75A
3zajav2CcMG2xVGk6xlW3SemzGNpSKz3NWtY3Ndf/yOlrt1S0RM8x1msG5nivlFd
cmGFj9kA7ff21vQa3FFN5NSSVsRAQ9VA+jiaFACxWJsc2j67GLb+iRGDl91zD6S1
JiDjhngt4B+UCdRuqj9UdD2T9izsurgGdLhdjKbML0PH/XVJ7YER4Naq8UrqOyw3
tQpwapsYkraysEt2kiSRP/tYUCO/r6NIVhHsEhld8hn7uTQ2rQMUVhR6C7AjorIp
eWPQVRpJMU+lnGzzHprNxo/pvZ3QGtQsKfGN/GkBB57d9qqDABnKvKhn/Wq+XtnG
73goSClVElqj/g01vQ+SjgzCF1hmiEQ5k3pKZWhZRfHRA4LW7PcyHMuQ0yOkMN+C
xreTA7O/lYUkVKqgA9kGVtbUUI+YyArOj0N3GCpMaPOyya6jw0yJTsGc6ZT/ZL4h
4MsH4aRRBOhXL44rt1LdZNAgZJZQzMvAMtP4hQGpDzdoOUn7g1bsfbDQIINVC9Il
sYWv0SLTuQX+M/bY2VSI/IMuNPnfb+4/61r522wgrd2JWj7dcMjoRjxkWuUH65IK
eKnZx7Vq92G+ytDmQlDwqss1Hvf/XFUaq5goLjEhlDo2C7T8BRqcLSzI15KCkfyk
jZyCO6vPjUcSbBnIgrpvKEXt0mzFsZEuqbxhgOOZvMyiBZthgcoVkubC4RBdQiKZ
K0YnJkmnaSN3rZ/RN8KIi3z8HB15nJSMcoqB+uawn8GgXWcXmCtc3vy0hT/UR6yP
quv81kkeyvr2bMEVamEGW2KflXfzzMfRVBWZVf8dA+AeDTHT9yKem/3Hk74x3Pcy
HKW3nnNaYKu7a8QMv1cwEqB5Ma6zI0tpiXThA2rs6L+r67RzniltKsBZLf58hY+X
d1TK6PObAbs5e9MZ+3nz4gBk9BgOp8uHtA61uulRrhS0vPPfNWBoCgB73kBH0p9J
KQArC12Fwc0yOgY9sVOBB3/UQ0sQ2AE/o9apDl+IxogqOyKtCAlHV/SjPQqto5RB
tK4ODJHnxenoTHtU9aiMQLHfTgjEEXnio0vhpR5H6YlFzYlf7Hwvo9NA4jTaAw8m
3WCBg4/ku2fkpA728zxtaRomJHyFYtFq4jA7rBTLq8lDvzUWLLekqwOClEzji50z
SyboLpzD8jNFECMbFsYUV9e0EJGZS2QIlqWRTz86GWvXE/HoDBgsEVPTTjrUeVNB
LY9QM4l3BOsEJmDwcW2gn/O/K5go7aZnSi6K+6wm6+T7Qx+i4cBIwLlGgFXoTKDv
Gm1KTT9QhWXlQnk/xG9PDeV7VT3G/dtmT9qTaokeTMqgTuYgJEd+lstyx6/UZVoG
hGjDlqRepw/RLRO2uGT88i5xT++DD/g4QEHyc9P1ktL3IVlMICCYiYGvhAmJ5Tft
O9j3vcckimnOvXemVJLrUdD3kq6n6pwh+vWcUWFuBhCi58fNj5AiVu15y8H5KOuo
TUe/qFWS9oqdkDIurkr2bwDbAhENCnZAEUF9tuCkPiUWTBm4N/ibQWBHjMrchaY3
utAzoGHnmK9Kvzg5dje2uTeaODGohZoZC4YZYhulJ2538mk61BKbC1KK/XpyHM5V
5ufumLFWRRLNiwqTXxHBwKXm50eJGZWQC0sE31jk2S/JHf+KmS3zmlBnlNcMxK5c
3tdGoO5V8XWGHcrcKOJ3cGeW9Uo+By61p2p2yKJ52v7op3P8DzrmEot/UGDYrdqk
hZJoUQKdSZPBnN1gf10yWSArlQgMXfcUbzCfcto+36YUZh/cJG8zDYzFqUI6Z3T+
x9plt6/nzpyJ8FzCyrnp32Tv/E48xUl0mTqji9paPN8N4wpXb7N90Ob6uEfK2ZM5
p/FmUFNx9owGHGFvKIDyLN5McjNF9dwfMc71b+C8wRZMoMHxF59AQJqu3KvSsU7L
4ifuaALjKmsneEDLLyjBzSh8VV0jBmy1bxmgOfOatUiWwczF80kNZyv1+IzzGjs6
BUxLOKuH3R3xQgFGwDHWSA58br8orNePmGushoRfopoYXnbwjvHJxXUpTcC/V/eN
ijlJ/piRLPXK0oQDT86x1ciaeY9a852dg0j61Mq7f+RicYeUpbQzlnyZ+xTP4oYy
bjw+RhgOgZeTUq8Rj72MojDLhPMF9movNZFACyikUDuh23kdE88M/vTZyyFA45Kv
Tc6XRD6UBOynNZEzK94kgtYIP96KzhLYBx+bkBNDD3ezHeJ6nK8n1n6RK4LiG/aC
Yq2Fll2knxyJD/jfv+855U1QtPnA7Kh7+mB6EQMS94LtLkpg2DSkTnt4QvIGaVFu
itCjXcM9T8Cidpk07ODGHgsiOP+FpTvTashzp6WzYItYb3nX0tEGmWGsXoL1RcPU
mcMxFDaUn28sRGR7aUEHs+AVI7PQr1mDAbrKkRSN0dm9U527fRy6QU6PJOKzzTeo
LypoXqDfcqVsMdwFk7dhom/bK1bTnIepJjylUqyUz9s4tx/I/xAxOLyEnmDg8oO4
AEvrGeMkBlA2ctChu2/tl2gDoIvgldc0jN2ugErA095kn8gkwwY6NkT9ngGCXRBS
J3541XXqGAIhv78RkS+sDp5CMokvHJtPe5C+AxPdGSxj9enkxNwW+44+THtijWrr
32cHhCEKN4wJU9v38r87Hp1oBaFW0ea38W3+A9Eta+bDJKn0WOq0ICH7xNff3ukN
e3zOfwHK38hKZZVIYcEcMhfEouvwLgCdbErvZTrWZSQ5US3IMKkfUD5dGgmMmUky
+yXtk1xWBTSBCkbPUaRNzg4P/h+RJJrRs2Vk9zEOl6WS4hdcuV9YyLI2TucX7isO
CZvaNGalqKlHtgf53892gZzNMVnVADTSOW0pwm2ePvl5fhV3jq7vlkBpQCCpoKdn
SV1u4SD8b3dhI8TPM6fH+z4ytizejFGddPe2L3fdAO9C08vt1T1gWfQGOsjaPLv1
4IdgDBWHdYQnkSWD8g92QRcIP5LV7KeZDVt6G+H9e1V9OvrprRfHY+OGXvvpoX6H
B+ymCsSGLk8MZnebOcT/QuBWP+E781V/5y+e2mYRO+i13M1IbENRY+nXkv5/jbks
XGpighcG0vaHUxAdPjnycTmGxG8Z/7EwdnT3JqcA8SJluksRY905s9B09jY07e3q
Ku8sRBJd2i+EX+N8Pu3PIt7UtGZp8GqaUWg+jI4TBRZZpKGmhzVzs3qDtkwQFrCr
t7B5ic3L2NJP2dfHLR386hrth+Y52ZUMzAOZF62ScMuNpgWTcLvB1Go8BykDrj+w
zhrEb85v52G20Fri+VILcLsdJs218D4F65/mpVY0mYdg3c9HjF7if8EiSMLzzpzw
3ssS30sYhHOFz75sCjPOQ0lnxEZp+sRe46mcEMucVvYlWN5advLsRkfnl8TUL42F
h93dBobAr5jYoowvwfgsAt+4rF0hpqwepoJkgEwkjScezX3rH1lBghyWc+2SPZ+e
y8urLg0Y6Yya9afP2w9eo4R69Hbq2pivmIrbMr3ODI6bHucqGvDPxCiYGiE6/W+3
ypOfWU0qILIwW4D8rJLlTDv45IaEl5xwhTQyBzQiJHeBikQyTeUmybV8MCtqEgN2
E5jodm7rnNI8DCCgC/0QZbMYXOq2UzSsYZpqM6HltUU6N5BeazdgyWuKr7UW+TnG
zddYFPksV80NhX9GNw7pmfgIVThmaKWZhRPDr/yxvSGGbhNMaPD4FIT/eQl+rkPC
MQZHyHkFnbpfZ92LYGlW9k6RVHM5lLcl/rAaCIjSF3aYdhFW0jgX9h9fxBUGKnjU
/gbAtjxAlJcu1Zt8M3puwINpw08w6D9B2F7p+aLacXL/06ak0SsSSTMvAbk4Zqug
GE6MD8DP63Ta/l6lWFhWyMldQ7VttGSIwiEwgarOAWGV3utIo2/+IfiJyP59PAQi
mccC10Kl1sgqX7YUFw771xx15bpcfoKAIxlEM/XDpqa8xrHTTU+nqRDyuxVdbehc
+StOEkDq2YN8CDiz82a3IQ5D2c43SrWh19y2aiO4JuOA7sdQTolesGIgZs12jhNS
xIS2e49++cRxJtnwT1cTVpIQqrT6D6j0F+MaWwerPMIjC0OvN0vxkgZ4j1HitQ9M
XBZXVFQE6rurAaRnUubcL8swwkZwqFCuYQ3lMTXlzqZS314Y5o+eJrFbICWcx2ot
+qmfoqDvSUQWsuv1qAsTRbGWu3R/A0r5eSZSySKC27SzjvvTwceDAH8lOviNOb5r
2TmM6mzLW732B4aGrjSVWfVvpeQBmRxVt0Rp6D5TDON6HWBeZMGNIm9f1UFazp0H
sbj/MaObZudFiF5EnHHiIt6M2NFrbyQlnOnLqua7xmofAeT+RrgFsweMj5NO3XrW
R/GhP0nSlqg9sIMoi7BpMUUJr4aizDGN9SHc6cAwDo8A508aNEQsvbflBy+Y8OaJ
HcHkpxvULcqt2veJjNymsutllXqzNvWxYvqthvC/roECHzvr1SUg6TiZzoyPj2om
vcMa3cNXpqvFTNC/2ynPcgan4oetxnqcLRKLo0nKDRMqHTvX9SkEdJaorQ8AG8Ls
/rw4aJUQSWBW+7sIw4EfY92RQdND7xI5Rfa3FTYw+hOv5up4XVDAGb6tMLlcCgZ2
WgVoTvi4TF5IZXQuTFlEoEZqmEK725cbdkx8gsqA8+/hAzUkGVO/2kDhX8IUdcCm
HgNkhzsX0j9+uqNpQK/MYHiUHaiLkBebEQtCnBR8kCxRcnb+bqGbasiJQuqPf7kg
nXJap9kYZNwQBZAx9QH6rESPqR593b+6tIyA8QY+G/GpXzHdWZutFxjWuHlnx5VS
zz+Zk693/VRKBuQPaoezLfn+vTa6xqzQl/r2eNpMxpxjjFz4vcXtxtig27znZmBU
qCnm7r1H/vgngRj/SBlXNdKW9oSc59REcELHtB6QooZGsBb+eOoNjtrF4x69GbZl
Ol//eALtgFK9JSmYNXm+GgBr5wLWAdcCRaxuepYC30ONmnTEN4QiTZ0VtsDgVsls
+M1j6nYzNlNdgtAv/hWP7SwPTgc5jfSmIMKdvv3EiyISzGXLGL+u5mTBX9CXm12H
ho2N16uQrlSQd8Ltsttm1i4L/a4FRrbLcjzYEmdRFGoScaXdXMeaADsAoUXUoPNs
yo13YpKMtNO1nqw2ksIMeBhpt9Qezv7q5ML+qzNnKQgJCe+WjJZLzkuQjGOcRAEk
hhZlIp5l49mJEJkt5BM3PDswRoI3hOasMuYYBf+Yotn87Gn1XSThlKUg2uqZ+Um6
yuAZoguXL6fU5wk8QQqHVkWYDuHSSVkoKY8lDiDcS4NmBca62oAXiqBvF9Z8mcUk
sVPirEG6UPKnWItUZUM4lM/VasYabj8HEo61MNbP3E2lXThzGVv+NaOvki/2KVTn
YAB1hCFebN7TjzhigR/wqWthKK8F5W3pbsvM9Eyr8HGSeQkLoezxGNwb0xA/KeLs
WD5m43f0kdYVYw4gNiksLub6zdptpvtY/vHkBd18UTLC25y/K9mihESyLpIsMBq2
KnolmvYk+mde87uvydB5ANA+/GYlZndcvktNJMIueZNdVTCM4Uy1aQarzPW5aoEY
So+a+RZOLh1yfbbZy/kWFsoANACMadpffNlIf1EiNOhVlKLO+VtjWNmz1nWlsYu/
DGquJfdY8toB0ZZzAdO6+sy6XTwDMmxsHWuWCjvrYMMXnwPLEjGt21HE+E6e7IYn
Quwz1BzmIH6JnjawhxQ0w5k9ooxH2YgV6JMDkB8RGGWIzIbPvxePf4kQa1bcruEw
OYG1l8loJTfOuri57D4gBY6NPvMPMeWJWSB0jnUe+urev3VFAxb0RC0Ge4CDIjo3
NNEfOiO5x7/4DhFnKPoA5a0OBTqMb7ziVEk7YyurDTpNTFPS/CRkXbwxXdilfJrD
vFRXBsIr9ekVKaZ+zfPtLFgPKZOcccXhJy3T4wJ7IkncmVlzrx+wONXqE//AkulD
vj2DrUQhzPUyI+8RmYYO0NwZBGTGggesq4kjSI8ZlFkcvZPhAECJ6qIJC6ieZktm
m79WWLqIfSSgGyp7LT4AZDT31yNbMza53mhwAxam3JG18ICt1OOzZ3m9WYLmiV+h
yG3AcWQc1AT7ZBPmGJpx78NZc61ryqYI9CUtgeUi2BTJcZTkQiyqNnzjgJkqJhN+
Gt8Ai4ajyvwp1DeU95OMcGniVn8mg5zJTUcu4rfVRdbY4QIUMuwdO/mnysLGFVsA
LawS9zPOgAe8bqmW965khO7w3AciyQ08zYncJ2EkYZR+RUNd6of1YsPwU8hdm6+8
N6Efi4T2oAQbRqPjqfz4xRzVur5PUSEywesOtZLdWLvPnUmbCnrMoMxUGVug4Tcj
DmgAo8tLsNYpE9/hIdZZldb67DU3CrRhCksM0ecJYUkTKA59HxBu+stotwQXQ7m1
rcb3SSpOuOMG6aS+qwaoxZvsppG1MncnalT/adzWSEf0Nuz9WV6KXVa2lUlix8Cg
G737B4lxybf10/uhdTMZTQBINI7wFF1tyug/e7zE2uwnPhmhU049bpm4HVcfSamb
/lZCgLWq/A7kt5mIAO36ZZXuVbbt0WJkC4TJUM56qS7jydiV5+b6He6WpekAjlLm
oZgUq1O1A+3S+8EFky1c3ehXVi4ycxSCsXspttVQRlwdSIgtVElsFFPOdxRNNfme
4sVOk/hDiKM+C/LeBsp/Nc5dOIg+Ypr2F+kpNIf+Fq0ttXeWbGahS124P703WCht
XAJX/HfQy+pIpyCn87G7Bj6Bd2ouq+6j54zCA9WoVxtnaQ1XYxUWVNuG0h4wUX9l
I9w2JCm365mzxFUcfBMxHHUAgOMxOs331pc9zRAyZLkDiXmD4iAdBFZBwt087qHZ
pmwN/tb32UnM5StNs9s5AXcNZ5ZL+DcS5HazwxCLrusuvEV5X2EFSPew0u3kKoqj
Pk3cu9+0RJlwXWE2nffPXBxrOiti4dZ75SxNeqRUIGs9c9ySfh+d2iIrj4DZkiNW
UVx1DCuuGfATzlhVYP1Nx3bkhOA8ZvQYh1A9RyDbIly4Ce3ziMn2oZxDKF/iKpp/
IoTOU0GsxUmnvh9jr5voDdxFW8ssRku3jYndSWc22p/xtFl81JJw34mN33hEIPY8
xt8ylS3s2wv75Jpk7IPsCBI2K4YWlsed9wEc3pY1xM6zr/ppt3Qmt8R1UArjNejo
SefzW4NiX8KZM9tr4/wdz0oePY2kmjBYuxgVbbXbAd/hQozi2ZRM4ZFc2lCa5EdE
588ly4pwf/EH4eukRLWLQk/9RkS8kEpS3LNiXhsIhnDdlJyFEDM4Y7bPxOvYYYv+
/+xJHemyejH/1XUa+aoqpGL9R80YGHPZJ61J/RLYqLn5SBYq3qM7VrOHNnw9Bpea
MWR2rGpmUTow1sMLCUQz48q2CkhNxb4xoPzDrNGA8X6G8b9eMAZsgaaCtdG5h/x0
NSFpQKhtrEG16wPhqCwWjsdwcj5awdRxut032ZwvBdb5qIbTFIZkqdH5eM0scPsO
U9nZqhAQ9xdfnMA6ehK5G7hKXroEJXpLajBJEgzxeaEZmF9Vjv/vW8zNKLfK0KKB
voPMI4vMKxaglnGkFzKA15VnE31beLhGM/Us+7+YmQHkY+ZGsr4Pu9X5Sii1Lsgl
c/3zS0Xy63oDWg4qBY5wMCQLRZFZFi3LKHMLzUBSaCzWD7AZSPG7pmQrXqbdK3kv
t14b+Ht+UB3DH0Q2oshRTKDCt+2zuRgiqyWnJyw73qAjfZMX0jVXVmCamlSODvsO
J5+g2XDbM/oAJhaaOraFD/VaSu4u+uhYTZBF3e9MRAcG4mWVuUrLM/twpjc70oow
54i0wQPvJRHo2nHrwNWjWa3yL1thQNJ4t7THJcMJZMZPO50gycBTWV0ykZiIUP4V
+LrjH5/2M6R68v3PIz5TtqodwtdT0fYaBDVVw6woZ8k9Lju5IMIFgreVIVRKkxHr
Bn2Y0rVcDI+X4He4fmo0XDRRC4SLWSmyM4tmKYeiwvrjlRzpWMHA+EdPpAj3UYHp
7poLhvuy0Vam4fI60HeHYL6R4q9ac2i6P5vtQ9SchdYPrQmUSwxavEYSXantZDMd
UDr37VARbqubh2CyAXjr8Y5M0DRfQJHGV4KV/h+wY22wxiCew5qq8/XSroTMoMuE
jGh48pWLV08bfvFgBFCxJv8m1FUKKNZLOVFQh4bGftWbgb17d9QqSWYZv6F34M9H
a3xilTGvQX2AIxPn8mT8Pr6BeqJAY97GSwba+Wl7D9hEdE5tTHLzo1RoJH486lk6
kE1JFFrPxfA+H2SbeLofxg7JjrMmQLaIQ4NClF0juv4N8x20c22hE9dqS8awt3zf
t4nCGvFJ9zkhF3ukljNqLBLXSj/ehsGIUiG+/0VDj6mLFJGoO23io8HHTN9vbmOG
8Yx6/WxtKU/VVY2UoNBTrUrVZTeb83sOuISaXOMcHxtFiQYhs8EnU7TKLGsyMDo1
VzNvldVeEHjP7SeqKO29sRLJZ4ksy4qiSh2c3Aem1B7REcV1Z2vIunAOEcLBRBNu
tNJ8bI1YbVOUUKCpmQTn5QDuhuhjGaHX8Bien50JL5JMsGPfUO3rTBLe+BdfcmsB
h47uBUVKVrfW6HmoWQGf1I3PGRe/L5Kpm2S4rlcP+28PPGOmBEJVa874g6YsXZU8
Kqj/zpJ/u4r+8ukzIavBLBUvOanKi/0h2kUnLYUDN+LmN7a2pQaz3IhrkKD5d+fn
+DVSOv/Vs+bPs+SNnW27/q2C4yFVHCwJC8FoO0yQYyWooMXUS/5E6fnlgeQ14eDh
PNJD8GJHaeUvarUkWfvEW6BFGGjqx9IZ02Ds3LIQXsoPsBTH0ju2fh+/oov7Zc+k
ue8lo3fU6YAnOTXsflxG/6YAYbPNEGLuyu1yQkHbtn9WBYdEHuhhQqFEuLcUSk/U
F3QtXbVm8+aD3Yphkn41oPwNa3PeTp5PYE/wcdvTTXsw4dg4gDhfjfUZtqwsONj/
aWDiqe0Zgtw01uloESKndV1lldRzPKDO0e+aDdXwcuWW+dwc7siPO+GBADJfd41w
Z4Bt/rjYuD1iS8eBTAWkkU0SI8JCugyzytIj1BCH2z95S2/NwTzI2sh4hHLHEzlN
v945mcWiZPHSLz8sxtXv5AEHfSRHOHkgjtdF9tpbgxSgCb9SFTxYFmuZvr+AXkHk
C32jePOIBV6ygTg+yM/drE01IOIaxdbFGN+Vq8S7zETAyYtB1z8O3QdL/OezGa2N
56c6WdVDw9MWBlrQjOpoKpa64KgJyoqPw5yzX6H7X4lrcdZZke3mkQGjMhEfYvdP
PDBCRJtEP2Y/3SUnSlS1W9CkwNdWURBxCsOm5yTbEgKzdIh7HlxeJ/A6eW9oXpiM
Jn3XxS/02HGsROGjWLxxnpxLvcZLnQfUbYw2zk4SYIneMPb7KKyV/nMnD83VLxjW
zH10BlUwL3kXu2avt64WpvkEO66ecG/zXeD9VTOxWmwEUaM285GIv3pbqdPDwuCM
+GPN5Z2ytI3/0poNRvPIrmFJvw1CVyca+zY6s0aMcBYpsR+WdqYDkP2OACIe/0O/
ywzBzpyGD5avx1H/ntmlCBeej7dWd+/U72rygmZrDZpeS6NcdcmmIw6w5RXaMJng
uUzN/Wid8trxU+uGWkJee2cbg3GF0p2kdFtuYRDOn1AMQSb1Cb3nXtmisM2Im5ar
A7amhAu0mnN3HuwOx1rgbHfY1cE6C9F3iomsrH1ZxqiDVGv3+WkbRqB6yrhxB57w
3wrMegPfke5Jjv/U2bAtnqm5MPkbmgiB4DPb14S6hnMb3F2hzkyecn5yFGrsXnzj
70/69xly9ydAqUu9ESsvPt+TdxNKSG8BjG2wyyNNvPPZa7rOnw0BskNQXejN12H9
ZZ63Gr+PtW1e3NdVKckqCGJXjVqmOODL4C2OzpQmZ6fse/ToIkuyN7jbKZZLbMgn
XyUoqsG3uXmN68DV4IKXE/KRTkO0ug3fCmiAyWpTvNK5XwsBpuyitm9Fmo+HD09U
q1JuI1Lir4OTgfeB7TvOVv6sMbeV/S2f7N0bdiyeJQX1hKe7l7bS5eLlMkx69jso
wCpynajfKpwu64yRa5HoAu4DAazqRrU0iwQSjBBBMQ4LnAeVaYnkJF5cftKGepeN
/F3nykbjmIsegnZVt/YRFl+R9au8kvjymTCjmhgQ0r9YAkM1W++RHa9ndrMwij4N
UbDz393tVUKU3RhrcFjx1+fRega0/7+cgf9hu5EybeZIKXP79kfNh422JbysUl4g
2SMAEeYBoFaTLo0uHCENA2FZoNQ+Zc3LuDqm3o3UgQI180FopbW63nY/6BPz7gcI
zxSPk8QwRYOYmeIRo4yEg46u/UMevEzY2sHXBghK64r+CFcrVN4PpHkw9BEdknFj
YeH4nP83c5Y1UwTgb/7U+B3+HfZ4h1Ijw0SQoi2AaCsmsxTnOICkF0plpUb3Sk9n
TYJQmtOE1UZcLomOFgakMUDTYSDbrgW9NvTGk59tmfxL4I6KiSHW/pQFxVZFq5Li
465a9eoUQP+xzw1WMZhfuscVINTZyRq8EMXzCxhI8xeQ2cH148BVf4ojSJ09cJIm
Qqm+3i5h7IttAIn9k0iXKC6OOeQDfKMEKVDp6GLRDE/OKGjFU9kWUKiRqifXDDay
sCYDIwG7ZR/+tsEQ7NFF4XI9b5Ykaghf60bx02O75pYhqt2HQKBlPvV4mDyE+phB
ufHj/eacLCkZKEXgDO0RxvvyAAVCsNZFdDPLPyO3xBRzUtbQ+s8180LjPnJTAGYZ
rQJNVUxCPSaNs8eUvY8TsPRW8w3/PV7Uu1d6gt88DLpyfjDmMtBXwnNgx3fWU56m
7KQtGjR5WGKCi+nrNnKX47srAQpkN0FB1TR6YS67eBNhxBEzltuW+owBWT0qAJ7H
WYDXsMTLZbKFDQD9itQ7bVjTYnHI7gDLDc3mQdcWEVlL70Z+p/QB/ST/BfQ4HU+S
gcE1QZB+XQPyeUAFcLOaKlMjbt0iwe7K2LaS8Ou3bR9YZAQhAlarUKIQMK6Uo06m
5WMtFXhZAZQvmUhvKzjJ0mvJVKBmfOuVBj3LQOx2TlvIJeEvYHWIfZAvjPabSOd4
/iWGQw2tALqFAyk4H7nSZz2+lnmA6rSouMIj/z+2Acyi60TID8+D1DjtjAO75HPU
J3NMz/JeDK4JB7byA+PzxUEC3wcYfNLPtZBF/TSiAGY4ziKtKJllFtk+waEOWBKc
LP4vWavYOP5qIvowxOBgU5PEgFs3h+hqOMPfj+Vgd/uvJKCOra7iFHmFqQ4bOXmn
OCvIa6AN+PcpyhvsnHIW7XP+ip4w6ucrfmiupFsEymXBZ56GfQT3LPHJCuAv2C0J
+ls6PZeJJ2knSylhvd8s+4BAspxe0FKp+ECWXGZUg1Fb0e73wYSxjgknyxOzpOq7
pTmtbimXHNH3YPLnd/K/s2n1xISTsPVBTFhn5ztX7Y4hnoDTSduDrnN9Nyj1Lx6U
+vKx0CGgitgXSz82qfnb+SN0wvLLANDHF4/9MhzLNPeI6qeL3gV7BOeeN8zaCkWp
W4SaKEDEy5rzsLqy5oN/hd/kpdx76NsrNbRn8DpTJzdQO8w8+UGhXkhZRLS6DAvr
n4cWMAbxQCcPFolNuoFYmQRCHLsWhAUWc2036xiikRVh6yYUQqiQgY2v4e5etb92
ztx0gbxB4YJBQdNtsCc0eiCaQT9shJbCFiGZuin7doyghcgGsO24N7xiqAzPwjo6
ltoutM7O+VcrpCvzW1X0CDqAhCrNG5T1jfkNCHgkbeOgzcFIHdJBn8exCSjdm94H
st3FdyKAEEaCaU5O/tvxn2mC1wqMxIUtTPMlp0QHyTa45Iyes9OefE+lf+LRPcNY
XEGbJji7oAOEnNq0ieJKQSsQLRowsZWZMVJxyk5auZ6kX/r3vJS2IooY6xIX+uss
WB0UyKGAqXOvH0PbdAg9fGQEmrBzpbOuI/imHU64yV5c7Cm4ndbJQ3VKHiqIOW+4
LDUZvMGI2NDail4rwmTB3FSAO/oKYtkArDVR9LrqlYv5rRjvtWAsjYT20knYJ+ab
7IrwK9o1K4aItJG6kjPn91IzvPedWbI2g3LR1eI1FkpHKe6fqeV6M4C7s6j9mITq
sBipBju8UFjTDyNeFzpGcZUsO/grY3TMjvDHthBS1mYEH8reuwocxt8yrTCvo+8d
8Z//JIKdRyzWEZ3yeLgj/OgokVp0Xc1LxFPq4+NJYQFubX72V6G0w1EL7pX91ZOi
BaTMkclVBux6kpKSz7OQv7JIaIIOT2y1FUQHmb8N9s/+YujNn4kMNkRWGhjMgbun
//mBmYmUdKgRCZdcJqfXtCdHOsvl8vEUoA1uRmX7NC/zccLkawbrB7tPe8SG+cTR
HwoDQb1Z2q56XZLvseiPWFc+J0g3fAKZ6B2ID3pSZEOwxBsG+QB0zefNXce/47uQ
05PxAF6d8S42uV0PHdVUZgbTjYzQbiXTczP64yOoKqQAclzql9zS86Y/zSfws/80
k2kP3AYFWkx+wsAcLhLrHUo84RfQrj2E0pA1nLc+QMrRVib0fRInebN4HELZKpTo
llJlnOfx3fYF0j3hwHkeN3DPkJBC4SrypIzFFqPTWdXiBXvnp8Iep2GPs7bvFv/a
mQpfenm3ptejhlV6RRDMH2bmfoNwAg8IczLaAvdyd6BHfch26BivYUfJUrEaVjz1
joRH8Qo6Yn0YFjyyg0PUrWFKNBKjHtVMrQB22O4o+tQB4jYHtI6daw4J8OKwXzLq
hXcFcsLZWzZ/nCCnmf+PhzRZYO5c1D1joUgtf0dUTiLxEqqS/mXUKraQ5tO/KGGX
Bj6bJwOn91pBFvWdigKmvhYtejyib0wOPXuJTL20+fNKjJpS3BftJl2l5jMkhOz1
P+2VLWXfyYOeQoCJyLgmpHujpPmlysFccYUtU0swgs4JJbsA5LIwowKVHUSL/bSS
oRGwWzqad5xBOeBQ+lz4O7hmeHuwNGwDBM7PygGyZF8TuKtdrXd8RVD8vh7jimjf
SokHNi2XXvRFV4vceXCazJBRoxC6hRJQaVvCA73FvAwSSQ2v+30NsOEXuqhzYvE1
y1t6dstBBUte5/KjEDhFK7qiF0mDl8AhxCGoVMYDcINiPQ95bM+xmCJcPEeGoEbN
/Uw+Fsg/GtDwsmfOQEzOkbDEhnx37d4FS4NRKKh4rDemsWpeQIvRnrtHfKzHy3K9
cHQcnMhsxr19zJMhcm2+pvryYQ/LyBh5PesvrmWVDYoUC550ZuWkDPOJKke+LHzJ
apqGTRc56VK7d0D9iZNYphVVn22UHaWtNjclWgYSmyyz52p/qMFWfYuwZDnovkxi
aSwBGhLD4mJKKz0M889dMdGNEH4JAMNBF2jz58iwOmncMRXi6NP4jnr4a6nZsxrp
Ax96WxMBdARUmTOJ2mKGfZ0ro2u/cGbUHUDXQBny/pmDv4Zc/sDVnMfchdouxyDR
5BMfc2CcBaQjiiFjFtPNN/9OIew0NULfvxTaVSAvt76XX+EWamTK0dlI3rzs/J1d
RNUCOl8otiBNqCL0J2S/v+lRqZ9XAm6RjUqzihQ8JNwCOJIhHzeWWE42av9u8t6M
dbpHKiQmf8h3MOKYLEEfVGcy8DODF5624DI+j5AD3gkLmci69DLG3bkCIVSKsq+2
lkUWI8xIdKwLbUlsATRBOaw4GqKE8N0RM4wVEr8REFWYnlGnUPz5QfuyMJjp08yr
9eyc7k+iRqlI4Rcr8zH4MHeeyy1aeXosvdzw0k2g75JAuCmR/YcdndgZhYkbQZpD
cxmH3WpaAlDFX2Eo7BxQ7rBDQrqiAOnOeoFnaNTZStOrEPjToGnl1kiUNMLke99g
3dTuE+r7F73ERBLWNIgQi5bPKf1PeY5HZhjMa+QRx1Mp73dPsMzsNCd7xSKuITWc
gOAXOc7yxUAfstFy/6C+JdWEg9gTL6cEIXHbK0eXHL+Gu7DtIXUl0Vu7ag9P9ytv
BF88+lPW0i4tOappjErc67eSmtZ5lJJuvbpMP9YxqPopZd4qCRT6k7DY29iXoBRy
msHHyR27nYlwXttuf29Neo7PwA0+siw4ZD/PCcw6+8IYZroMM4NOww4RsBjgGhoL
iD5G02KzV5PgYWIoxt48BbeB9YCIleFiiY3wpsJr9jnIVQx9308a9C43jZPupRdv
7f9hcwosNhR92eTqNs3nZVL+izTUx0qtwzng/ZtGHJSN4AhV5mf/+cOB2KF7BNqp
G1svRO4U1qRqSAy/Msns1/NTOYWLrKrWWkFky64atcibNaC8ROSehjlm+FK86EXy
7bucZfO/36wHag7NHFGn16sHopey7W3QwmCytdgPYP0XbB1T56C3JhzhzwDLztIT
STHWIuEm6glLkEzb73jookMKbUBRBlhZEV1QiSrz1Ddimb9U6SZgmiHCTsTdTrDz
tXppbXG8ZhI232D4NY6LO7Onuy33hxub6O5HN0NLBMmN/XRH2/hZ3NSH5mZQAqB0
wBjhzjqBFthlrt/YJ/79+22lq3TdrS89K0L4/zlA9tcd3GWjn8Gp6IflLerselHA
FUor6KssBpShe+uAGnmoZhQ3Z7/nibCl5Sz86e60X1OLXUFQx6g62WxcbzzyI/Z0
zmQiGqq1Kh3ExVm4zz55qTFUup2KSyEM5LaUr2luzFziCyFfPqlNACGjhlRxO29A
sSOV+PafUhSJb5B0Xuz8Ob3jLYq6Z/qvfyxwb/s7s+5pp1Scz1HColiPr/ZSKKOG
t5YoMRx1mBO617xQQ2CTXQZbhng2V1zNXrMWFVkhI/0CFJtu7yrByxfGKQyAZaJp
TDC7FAOofDQS4KT02mHTtzOH/NsBPtbOkdJot8uTxbGNtOP+unWtMjMF/UORirAn
kLoo5JfYlC5I6ZOYmymYpZOJRk8QvlTXMPzrtvqFF93uDdeMcoD0HsswQqrPNiWl
9xktNc8Moy/Mv2C5h79hbvlqr0Bdc3cw9iOxxiRpzhK/7TB7tRGhL/dph15iVWuG
NuQdKY29xFfbT0nWzlkSKIqlfrnncPNfVZftcsNHtjL1+E8gVu0M3qPifD1Ke1nx
Mm/AM4ch6GYdc+kNuhAg8mtymvXHZfA7AfZdCt8IB8GBbBHaS1du6t4VjUp4p/iL
yJJxTnCWmlwG5/zEZUu37gxWFCtvimIBeoIZM8Tqa3kw2p90A0BS0HVuzX8oyIAU
/1ARJ4n+SP6KrfWvHSgIgvcKrvQisl+gFrkhe3CMrdGeatZPXg116k6m3uFNbdLQ
21pd+jUNvCq6AMaUDPjeqrQy/EX+9z9iIALE57jpVJVwty6+TWHliUncJ/zuXj0P
260/8x21fqYMY6nW+Wn7qUfqHNP873nQwwZH+zkuYWWKSG3ZpffySapVOKCBjHR/
HO2CX7OI+16YhJVqwNDG5h1Luhe569hJBnOJegtWoBj6ni2on1ECqXUQW28w6OLv
nU1DCIPuhTEirm1k79oJNzYvh8SI/JDiIA5qXPbjRZwIVtRujuHQdx/Glnq3/75T
m8CzVkPMfMeF7PPP7l/X1YyJLtM50Bf/zv6iRmDR/5fn9eAt1PT3mq8VHO1ITo4i
Erib00o/8XVoafilulXYZerRFeXPaykjCJpOoRUEAIzXItapI2Uox7QgPgUp+fN6
wSR/EZXxK3YN3+ohTVQcdi+roZoGd6HaO+cRD1OT9E1+bYi5D95B1r/lGqatSoxi
OoUe5hGnVnzX0blQc2HpT59BMmZCnVrH5A2fk7mqhx3oHEYDd3v+GL/9w0R4Vr9F
HxZX+ApfyNQeaY38eINhqErHsYZowUK+oUmqgj8QyJRjvjSRaZ0bXTU+E2JzOXAh
8DJJUp+HEBSYMm8u808LlYwEvFCOuI+snD9RWNo/AnE6Fm1kI0W3SdI543QSJURh
G1K4srdtAwOzHZsQwQPZRtcyB5N3DIAI5+32nImxLY28aNvaFUMjAiTtM75XPt5h
JLNL7wkmbFs8i1XWxW32gnBxezVJeOITODtWQA6tmrFPmkqFZKk5RF0qeA36uz9O
Znbb5kI2OHE60nJPjgZn0qD0ji+JN3rn9QTlymMe5KHcxVO3otlyqrsb4bHOwyWD
SEoNHbRkitSHttkI9IFOjamwYdeiK8acCXxBNpBY3Pv3oUlW2K5GomxkuKP9Z6NQ
i5TEtJ3qSqo5hG5RFv1n+P4ehJNQLkYizYywugx393ABHCPd6/hg6zhaCNWLdKeK
fegN77ZqETY6I7++0uWvagoXizDgV5kpYFL54KEi3zV0neC31zrdjsuLYc8x/22a
DioFXPaYWZtQhJTAtgU8oTDSSFO8WwGrpeBjvi1B9baDwuQpPyaBRlqbABC1zl3U
hTbdaXI5KjciJ5fNHAomhSglnlHRuUMTIMao52z/ZmB3FE4BIJ/pp4DuwABbh9jc
mrSxGeyaV9JVMQZpcXuGkuXlVHpV+h63le7z7aliWgTGi6tcn2HKx1TGmKtDYNa3
48jvq6NZaLxC8G5ZKC0VbGQLLkR2COPYSGn9xK3UekdrGQxZLvmVKad0gxS4MLhh
0tDlY20+uhcNQKgWCGqbK7TWlwWinPtPrkze+YGkoMKWUwPHF7aoiJZyz7CnSQ1y
mXLS9kOdv5fKHGzzr1uvf5NvKpFP46yMoBHCx7auivwfz3IbpVQlyLB/+2M6h3/C
nyAzDtTWbcqC0ox06MK/NKhl6ooW8Y93I318VhBxhikYMdZfVY6y7nMyGUWPDZdO
xv3gWGDZASs1954ndZTgFUMchRqrztc1G/kTgXARECQU+4QM0WiYrMon5hNxZxGj
TDIiintnhXKgnfq0L3BcC9llgH/ZrkX5cEb5ZskoVBHAoKJUmE/Eh8f/eqnkRGyU
vvm/T1Kizy+RDkmmPJwE81EISS8VbLAQ/e5Y4u8OdBs0mCE+Z4izKLk3/mOe3fY9
GqxFNDQ3ChR7Yp7zbdg6H3NaC+KwYO7MEnxjtz8eXjuPOEDP6HxX2cELqrsVcqQh
IwOU1WSOpfYIA4RWeJwbyV7/Jw64hS2mbjDdhZ284/z5D24/oNJeOokvbDuB/iPn
qyg0TeP8Q79KAI0978KTQ9oGexTQYRDJa1oVC6Vt4wwUxGqo3TMW5DcOowIJQ+vX
C75HGh6+ae1v+fn/HdDtqmdtNopFEcVVwnosKJbc24c8Hd/Rp29Q3RfpmB4m4BFy
y2eEIwYw4LIL4gEvFB6JvGRZwD5hAWWhlUvBQCsHXwsWvy1jseSO2BuXfiQgbvoy
l2oSxigj2RR+jqt5f1F4sex2xwDFOcNrPEhDGfBEzBR207nGt8npEHjVvjAuyi14
e5bIetJWIx0JXvrNok4HeUqjhmy+obpVNieu9LEe6Gej9AjqXhP0jkWygqamBVqf
JeLWmg3Wzhq0d0ZSINQvveF+EJwpMfa4heDBJdlHhVtLCGP0P0UyJ/BYAliREyGu
UkczH18CiOS1x+PGT2IXlf97i8gF/DZNr5XWwaoxSsRDquH3J7AvSPQijT90xni+
gWFpj3g5k1x5Zcelu5GwjklI6Fzw9GeDaqD8tB2STGhmxvi/3PM51wCNfgP2xeie
BtO6DP28p95SXlsBnpdhQd68ccocYXo8ABw+tBrcsfLi6nOjz2e3olDr9wyR2kpz
UIHCF0y0mjP/V4psP7+LZXSLo+M1YRWQbAaYglFeEaBBV6fI+3zgpha/puwSCUlb
EK176Nn804DVoSQHGQn+X2rMqIbhG1vaKn2psDGHVMpKhKI9V+a1O8WUtrWOcWJD
jtaGDb8ViA/5FFR6Rhdx8qavWiiUNY8bxd+zpdh163oj2tNwEMKEHJ3OEtxRCu0K
HulojPu6cQq3NBBKIFHSmniosmNXnfc0Gyrtz8Srp9PvfVNmhTfOf6shFWwuESX9
9FPjKT3tmItP+h9UDB0fvBTotMjyZ4D24pxyQb957jUFQReWDfW5Y5y26NRuKdAp
jf2PH7HkBkW1lX0Gv+eHpN5nfQRYpcoEVzPXUKJfCDWRTpLlmIcuHQsiauVGoXNH
bl5PqyK2TWSaqMtDSZabpUOBkbn+0A7L9f0/UlPDzOggaLveh/DS7ymendoS1o15
89K/ZXuML8Y1K1j/j8WxxJ1tjz5TuSUoxOpBDWG/3jPH4/g9C350r/lN7qJzl9Z6
yhq9LmCMSp/YSjia+TFPl5xS46KFPSdhHBv+vXYiUCQJKUJ3/kJ0AxmDfpLdNWOS
sJF3F+vxytqb476qyRzyvYycNPEIUGzMg8TSyY366OC8qEL0aGf1vnOZGVL6F3mL
v8o4eOL08yXVITGj3+3DtpRpx03szOqzru9/7Qv3uY25vfZLrPZqeKlPAw2UtEsJ
IUzs8AXNg+Xb2h39aJ+OWfOvcW1XUb2Z0wNGguYQy7LbIbPv6dl/IT98xhvmp24a
JjEXfj545zi0AJlEDuC1FHGFKghYd2WCJF6MEyZZJOAXIlvvHszH8BNHLf5dHi2D
7C38p/isjUI7R7yzTENTiXYkHww3GAk8IZ7TNTQkfqmj1GQYPcAMweWj5Ej5y6Ig
b/7WoG4rbIlfJdxxwn5MM4LMECK49zaup2tih+eWmoXstzXfliqilzxByBRmdXiw
FV5eSTnT8i9pIqpZJTHlM8gXKH+K9q8JG6Y2BsY86WoJHy00k+siyLmhaXWj8w+W
Dp4TdikU9wAt0ZeccNwCXO0MtYS/I1Z+2oDXMDIkqrYhenZfpbMb7JGP5GRRrvpd
tTKFdtE+UOe2sbaggaECxitTZ63AIwqtx6cjz08Zzf+aV85SHymvakPPJU3Jr0SD
uW7oo1vSHRyC/Px+WRSbJt80P6JV+AS3MbbWqHfBH77MAxAtZ3JstclXVSHR8BKI
Tlx3EUxN29GGvF8yCK95NglR0Y9YYksme6eWPvcCgr/kuXl1zP5YMBqohyTasFmV
WACvWSkYDVJb7cwHH8eDNzreh9aYc8L1EFn6rlQF2PhEQwPd+0HK1Q4Wjh1+kYjm
5t8yZAKU4ondsolZmGcHIdisJOFwlpLRPLQcnUyQHQHMtCWZ656/eZ83vVJVN2s8
IRUPnItP2z9sLKhXCZi2MdpJfhqcNQiwk+MfJ2q8S0dn/OO/fH1a1qHmqdsP65ag
X75r4ytKPGVXh0pmGcyPYxS81B6TqDph+52CyhQFQiMwT6gM5PZ3Z1mZRUxy3lUY
9Is1H08VM5hcarPGZCt9gfN+L9t/g1cc/hWWYZMopVWXooaMiARPBhbiwbV+qI1p
sHNJbNU+Wda+HHQoi1qmTMMka9gk1wNa00MJWYtA0Bz6AZPj8kmYfPhyKcl7rMLQ
VGwbDgxFKAYHgugBmrZfaCOOm5Xtxii7NjuePaAhZ6E3BmV1s9dG9hy41dp2XTci
LBIPAAMJXATOCLifmRVIXRV4HaALBPb2fFVp3wJ3BFP+pe9U7zLi0fSflFMrexla
A903kLja602LuK6uN8H/tBi3pz4V6ubQgoVOa+mp+Ok/fOTr183wjwhGhJrg/mZx
PY6GME6WSS84+YiPx1WQEf0SmhyfZPR2OgiRfnXnlrMzPe8gx0iKmsDPy7KKNIz5
nN2gOevUtOc4tx9Bs0JvkWMvPrJyrWcmzY7UIpFjxnWPOUYV0cCyyqzRcefDnuLm
CAJ82vVd+hZI3YAO2XDtczjO7Qf34bITG4oRcploVUE2kf7tn0Psq0PQAmBF7GRL
Ce+ZBD+40PlV018uduUzAPqGjNql0FFA/193KexC7zVIklXFPPI0iKZTkSidW4mp
km3A6SoWuIDzxviUAc+ScO6J79PN9PM/7m+pRDte6K0ue+IEW9rhvw0dwxuHrBT4
wEdgNBg2j/H+Mhsmie78Vbor2W6LQLx9fTyAnu8gvncGdkLMaa1AP4z+2EMBNEKe
L698q9BE3QTVlonK9C8saJ6Qf/PCLtizVJN8Vpo/SHSan+O4X8WFRFrun6Zd6GXY
vIFsjx0UGLRpfQizxe7q/orPu0X76MjZEvfQKyRTFSS1VoNeaQeUwrATYrQ9k6B9
ADF2rZdYPeX8rUevzPg67Xmsj1FbfhyzKDd7z+nHT6p1Kofi8s+nlWWAlCG58Id1
iraP/YfJWG1Y6fiqOrV13zCiC32pPNZ6jd7yuYpqjzDNvJzc+Qo0UdF3+RESPPp2
n2MQx3UarzjKyedg2Ht0OsbZZM73t03ddLxOZyfmD5rhDgG0yVfDYRCv3e3S37CH
JBE7D5oai2QqBM6o/0ModvAhJb0fx5jYt/WNmfCFT393vIBlCyGWmF8Up1wrD50V
lXZVdpbxkJ/THpsyrV0hIikq9QDfbalw61agTbqHAdbiiAG2JF5xcYQNgOs2VuML
8YTLtSG1vmw7U0sTS4IlAwe15QWucrTFsMtkuNihUjsSw5w5QD/6gxLh0J7VIend
vX+APk9nbJjyg+62FaOD+cJmpS/AdkwhYHDvtEjvdFiBisZ0Sz8gU9n82rPpobKR
pVOdIZ549ChgZaQy+sa0hqLFd7GjfYhRzPsv+jRW2KvOQHOIkBbZYLV+biQhOaAO
07QZuIg9hTOGfWTIqWDDNGNYkBX5eyN6o6teSuqXMSna8eSZVBUQibabiSIAhnlm
lJrHCCeXN31vijhuSvA8Jt1m8xC835k1vCV11WjXt9oZ3x/TfrU6s957TMhSnbS4
hU+PhcPj/GeKE3VewG0wb6n8sbfKZvgilYWf9oQtEakUrUD0jL5pdrIeZHIr4QgN
VHZC8hBjhsBMjLUsnTjqT4+I2wNALUYIhigh4hZOjObXxH1MIbmI01lQnhE3gRVV
EJf+lecx8LLs+YDvEDCbrhTy1RSIYSVlb2Qj+YC9qT3VceG/gQkZigoGiv7l0vbX
br1qxHKFu28IO1yaP/JpMFCBPNMtICzh6gE/LWrRnFa1vpm8cskbgQVPiwSHtAHf
J4dqzVNV94deFEXJw3DoNeN9PLJmia4QW3JEv/NNhQgc0Cx+hVBke/X7sbaDFsj9
W3B3KdZAaZ+b4c3KHff2yLVzAXEtEDW+ttXR9N9e01L1V7r8y7nR+T1hbZv/ksCJ
GOd6Cf3hwsO+K/TkWgb4BFBTZ2hDqgg+DDOFlIGsHZbiTGfQcIowfKkF0wAokXlt
sSY7vPK8AiFd+zwPGNJEFHepUCvVddRPLxzwAainyoSWJg4naQNYVhw4vBIRIJSF
ZJdIgIIQew405jFAs0Qx74wWMQ2yrgW6mwF7kh9RsZgHF4aHNg1NXBAU3tgj05ny
bFHMEZcePYw/u8x64F2P8Jna7nyOwaZBUQQOJ9Yy/tb9wgRVIFuahExeSdGKHrWH
ExauU1nXdGr1iaovoxJLVHEsTFOxLmlJ8edfDGJPn56IIx+7x4TvwrsX2/8go7nn
sDnW79297Wb/enYDrOt+qxW7dhaPepXgqMxNcX8ZMM6HzZ47Jzi/XysXk/xk8tpE
VLuNQNvMfJDZBTIzC125VoX/0BsmwR+vFVFW4MLb9BNxCMZE8ob/opcUVfKL5Zvt
bBSCWPihJ+3WQ1jqB1i/8I46PlLPoD3RhFckbgwgyJoo+3oL8vJfs19z0aJgTS81
uSVExndKsmvhJM08lOe+9kA6fisP9zNMMMn8jwj8w+AtP7OEzix44d9/2eydNM3U
hPK80vwjX9xYPOAkj9HR+ObbKtwqYqOYMnOCT8G/GCpUwU4gj/o03uWxYQRnSBY1
K9gneC/KHwIS0syWtEBoLbi16AbLxjgVq1ag3jXdyg7OPdVm+RrzyyJYJC+LrfdZ
MsMMu6cu72mKYqpOY/zMyo6H++2AzLQSsnSzRxu+HD3bw+D9R8+H/QIE4LSgc28/
liG/Wb7XBCQ6BBOcYrTMrFUvwMYTDOOED5lYz99qoWrLmGgDumRT8Dvzthqk51vL
p1R6u/51TkF2zEoNzNFn5nVDkoK++u/sOQuiURSC5kWYNnhDqIiwgn85oT5KHLLC
WCFOUODtl53yQrBK4S0yceudovd+urrWRceLHiJLhpcaigVs5HK+Ikbq4ce2Zpj8
oJU0ZLx147SHYGWeWfU186zo2kWhvC9t8ivYTAtAiaFd1/pwA4hFcaWYpIj7SYPn
A9W1G1WHxOeT4wUw/RGzhOI0Fz12+EqM5AmpU2GCsXEAOxZltazZRsPA1ozg/N9q
mh2uugEW1cm82CzIwdEr+YPdY+ezygPR73kvkjDtniJSCY+4czJP/drUqtqSNq5L
9XSblvvtxjhA6yGqgxFElWjXLhG/UFaNviVFEKn0/6MbbTbq38DuNd6cfb3Xk3fR
gFNprcP3Fisd1HUUHBtPezDgb569YEzQZsNpf6fYRh32vx3Kf4/0BDmXjKpEn9E8
xFpV0NdOFkxaj1iS7lHXXNpGmtZpj7S8ona8Cm2oN5Z2CiHVYPXHpiQETH7+NDaj
3lAvl65I4WpFYwLD4shr3286fypqFSXW9H9TCMGx/E6zi0p68m52dhSHMxsLn0C7
WFyxac8tjW7/m87xiOO9LFaKTaqalGndHYsowEDzkQdmM8iTjZJHqXLanqqnurAg
P1xXW2mu+uXPXZUAdXZ8CKEw654GCrxM541/+9dK4I+BOB8wckRL8bx3TQcI1tUq
TafEc6/pFlMhE7DVWNiwFOa++cYbLPQVXwqkYMoNhhuGiyL9IcIr3JI0T7H5+ug3
vZhSgOBDoaT/TAzDsDqmQP2rDePWgux+dgfWB54kDzWxBilpYQMc6B+USebcqwm1
tvM/qQeg53g66lPQuq5ESKZPKmJbqtcfE84F+w/70nmSiMnkOBbulm83e/Hnher+
vkmL3eOcP2g9SuhrvHyWuWjIh1N5d3Yp/qNxB7JR2C0bHu8L5/dq7J2Lu6MGZShK
gMM6cdellkBQSwE/TotUtro9D1eX697S63hj1cy5BayeRTWM5MqRHs03mJ0sj9s0
RKpQfRadM/Knl6pQAS/VkLGO6DR7ft8Tt1hggndGWy7xu5Xgi0vyIrwAniPT6vTR
SjESmCNxaU7aHEDZB3PkJA+OW4iL2v0cCsbjJ5w1rgQbC6SNnkSt07TaZy5OwDFX
kFYTfRL/MXXa9LxY5uTyccAP3m8bOMjb0dwmTZQPu7zzzHa42Uade1MoPKP9hfVB

--pragma protect end_data_block
--pragma protect digest_block
SKPP63eqPgFj53RUW08+BAjFYzY=
--pragma protect end_digest_block
--pragma protect end_protected
