-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
VnUMchMJYz+wPK2lenTORkRvdq3Lph2exOl5QqwT+bTLn1a3I5eJIsXLCK5aEVo4
cOjzroZcVBGUx+H0RDfDAg+DYqkhCXlsRFL5X/BF73cjn8RDD+lXHnuA1pOyJvDc
TOG7484K7dc00aTZcUHs6ZiiWzz6sLVCuS5kUwuHXAhDrbgeRK6Qhg==
--pragma protect end_key_block
--pragma protect digest_block
qfzoz1jC47rRTNfxwsdYhwvXWDc=
--pragma protect end_digest_block
--pragma protect data_block
ct3WnGLJO5sD1W/6MJzN73XTnt++IB08fj2BWSmrvZr8L8Hqa29qCiDykMQcBa6g
MsBN9xNHZg1qSVfpXK+Yd4qxhJCWB7fdRoo+TxZYp4xi0gBEO8xIuQVoihog/XxL
SSsgO7A6Gwl3m3T+e9MOLokqvB7JjQM6+PGZ8dyPQVEvrcJ1CNy0o93ZC2rDk3yS
14+GaPI2sHGi7B1AODCKkXiBYJJwZAupbqqrVcl3xv3lWlndEFUchA9i+nahA0jX
v4MTIq9Fyey4vX+0npWRPfv63onz0DaT8EO+B1IfzQWS0pD/NYUp2gEZgG+S/wv2
hu+w5E20MdL0VngCSiZFru6X7cPF4KasPb2Ouarz72wx5InEhOugNPgHMvRRfceQ
UV9cYeKMAB/b0zItDXmRVR8HQWwJrU/8kPSf1u+YIwyHsWO1JB4Kok2mIOgnPIqs
4uagVlYlcR1s3Oj4Rm9D4t7u5VgixNOTVP24iYRvWqYO29T5EDkGj0rHJ5oV/xJg
kh5R/Sd0Rc2vqJup1e2AiWIDn6KVADrkA+ikBiS5G0Ae5/tTiOBO+1Mo58bDUsBq
9xXO7FmyOSM9sMzZcluc++mcN8p7AmvzrWd/yf5mBPUhgS9m1aDcyVkG2yMEAcmD
hVKQQp5dsYKy/C6Tv57+PKMmmWLNF3bwMMSwlu4IMJEGuafiSUFo0tCfN9kWEvFO
HSDOBV5QkoflIih/pP/zoH7RGUwQjvPpohKl6iTqOFG4jjgMMoH378ZvLKrPUdMz
ULAYs4bODNVlTCgDkCB0TZiIFRd3VsSowv4oLKJxnE2e0uI/1KPVV4fkHGpScD8+
bDDdSukk+hniyQAezMk5YyAlQ6TF0Bw7T0R3ChVzkWSD4LfLzKd8URGziP3w5ERC
yYoEHQ++jtA8I2Vy2YtPgouNyLwyJCW2cLhMABYsc4LVgP/j4vWanY5XB+jVqofM
35IJ7rkCYx0tjGfabLCRFS/4FuCTvykMAjnSKQ6e6yq4rQmn8ylheDgszdea4m7h
fLKSKDQf0BTDg8lQsHCZpnkYHvRg0O78IvMwp5K8g+zc43GNPb6uOFjKOc/nCqW0
xx3PO/njCd1lvfBfx4n4h3qTyUQzJNad3T6iUU9XpfOefYtvdoi4TVjhlOsZZeqA
yzUbXlwLu6dpK6NOaB4kE5b36S+xWoo3KiqDiidYC7nzt4sdDv8hbaLhtcFfiX5H
8H+tIb22UY5S/1HLfdW11TOjrUqPJ+y1b3m0jCAAY0M7PQIRaZL1wVvLR8J0fnur
TbYoM9ch+e0VIMMVu7sVJSfaQieIskDDJ4m0qQYLCBzE1Znp2P3ED4DsvOFNL9Ua
FrybOhiOZ1rHEOlacant5zHPQAUd17f6RhO+EBMr1xfPiDUBnHAp0Ah+JdjVWVQ0
9cRFn+CN7OYSITsCVEQKpGLfbcZ63f9EIPjIk13tdUG9YhZhEtlxz2SE1hc7E0Bk
y3zqNll0qGFFKG9woqOp/YA3EDZcd5kop9WmaMjKJwAgqzmyyL/hMgH7ImFZVwC7
zo20A26Mq0iTXEZREeFoIVnVdt9Ld1+u0L3FljtXinkO8zDU1TqTez3OR7/F3/ku
844/fQbilSMENvc2Eoi5CRevb73DeTJNXeg/lhWkDWEkitnrocQorDMAeNAU7+Xi
Tl1r/vxX2hx+1DiOKeJZuC/LqUVT5R4fwXZhV0L9jMHoQlzAUetornCvnKmj+00i
p7Ik62P5aHIFG8Z5wYIbHhmCk+yLv+9vQ774vtZKo0SqHv8rJhVHeU+QJb3vp4de
77Pj92Fe4FbBqq+q9EWy37JevLW3HDnvlw469e2o8tJ23p+554RPPL27E6NL0yu4
yobGOWxBu3MwfThJ6LlA34VyjY/TTP4vZ5SBCVBaa467AOj+Jm0J9JNQDwNRGp5u
IPbte3Tl/htJb0pGhL9NgbdpDUQTSBilqAvzUkpq4Bwo8ipnubkBLIlmqeoo4R9T
uD0z8CfYUAwab0oBtRNI8AZOdQtZNulEIaBExit+8oqpLBihWArhzNOeYThsabWE
iBz1PTGtMoeTF2OmX2I+ewLhyIlHJfi+ZPOfr7qukd7KTHyEqLFrY3XmSlJs6So8
SWl8GIy+Bv7QTjoq6HKARpu2F8uv5rm4yOhjGElBBYTutO9QYZOL3hobexV+W4Or
OEA0zTuaXpGcCIzqVFxHlL/mzE0bVsTcmN5hNnh9ZYtlXIOxyLyG2kP8goTMv4Ki
b1DSRpJnmAa0fmJqWOt6im65L+nvXZ3efSDp+GAC1zwQLuNPHp21wqKh4B+JvE5a
b3QWt7yEGdpA1WmbqobOzyn9BVcKTQ8PQekgMfLOo9PYGiq1fPhtSmMgye4uxJP/
RFTwQWoL5ChgC8NaTxy6pJA1b1BZvXCEnrUbZd0kl/PSwf4IPhOY6mlv2Jfc9hoM
zrnmuVsQeokgsG+Ixukksrbi9QA4nTb87balPRxB/3gWkFJoeufyIEPdjHPsgPmk
yZf0vVL1LkNcWwFvwC3qW7mJjLC5DTjKTL5Rs28fYFh7/skh/Di/HHWpZ8Z6P5Q6
ZJ6vy1/ej13AKTegAMgK3GUGmxhzbxlu2P8t7ObUTvG6qZXxniIzXnOaxMgZ2U5o
ZU13z71pvwo5VUcNH8LLXv9RChRVS8qbig/1E37MhnwOsjxNNM42KWAGKyMH3vub
P6Ngu1BqTgjLAPckol6SBkdDXsKdAVNn3oaPGwUbTGKK50D/Fz87siFQ5vAAC8qA
xpK1FrA3Br3k0WFmzJA77Q4dy/vzD3ZCen+mbozWI3gYiyGU1tF9ibK/Mw6m9hsW
R0OLpHSda5iKpg76wpk30xEPCRSe+cTZjsya0HyvHGfodynhjA+gK9gyNeq6d880
wBOP8j8wbdDQR4kW5ZK0cQ+GDKITjso77LNvB8FctU+p2CymNmgVuuYjWEv52Njj
gVeVnx5XAkcQmn5ZJdiGUfwhyWFwjshMeBMg/djg8V7WPRW4+LKNXltAsgE6X8Go
pR5qJ+MDb3djz4+YgVUdNpsCB3sEMmZ41mW9tazupn/+1UnVeB84/f8jkgZFJk9o
gZ5P5mMvWDwwyE4fOZMXMwaRuKf1BEGeIFXsV3bNLn0kUjE1n7wuIxKIQV9KXBlU
dmta4nyvtDE4SbkC7Jb09BE8HdhP82fgqFhoZ6juS0+c2qmIZOQUQgK0lWVDY3cj
+RcTwRyeJasEGSNhPbUQjQ7yhJLjPSEH2xHlyuA8rkNG8rb9YPXF/50uqWnStZ4m
vmwRj2pR6Nyc/+oP+hy9R5vWwH0XX1/2rYkiMEEyziINOBlgqr/i/6bJJGfiwtfZ
iZ7BlNM01rtutRIbiulOQ/z7WeASOxakUGhor19BjdLYwo+T2lrxT4eBINdw2k6w
afw0hEEQv2l+3FrxkFqfgH6355MyE55yzYK0Ju9Z2wjkF1SwCpwR+JBb0J9sJytw
0YRMwrkCymNJYqK9dEgNajIr6xhrhLBege3qjBWWTMfCe9usPlpSvAJn2iai9xWA
tvqaqAgLOsyuh8ftv/kpY1hRZGmHUWbzsLldqZZL/agmO8V8uYAkd96r1AwLAhda
/c6Z0VXtKGBUj6goyIwFJpmbPz09iDl9PyGQQWBO3K7sdMhDy/76yLHdSNBlkPaZ
3Em2T2KmXPLYSnE79iBKGmbgsIiajNxWphcVk/TvGSN6oNew5WvBts9qvcY7ilDi
w6TN2ICwaG9yqjimoE3Sj9E7D05UgnZoBO6ZCFCcT6KXS8EYPVOkNl1MRGNObIZE
7XcGAItX9mGhF53He6CZQyuwLBH7JkrLDFAZqRF6hn84yCA3MfyOGZnYoGUyinEZ
dqPuT/N1PQXGx9RmaoHBSw6NE4aEUjpwJZI+JhbUrN8KM4mI3WY3ghY38AgJJBvg
wzmrT6HtiSC67OOdwCbxtZdXa1c7FKVnwmkfrDo7yIkJJUlaeyKIknEjYO81IkwK
trZlg1d+l92G6f7s8J8JCn/PgZTn+52cxuJaQvgsS+LD70rBePaLJ6rQe0ob5gse
l6qgm3+iCnpH46G3MsOcQ8fjrcX+iNMsZrIKAfyTgC5WdHm+axbkVw06K1IfEjL3
fLW61D+1VTkldhiWASGoM1xygjy9cAWK8uBZHgJcEMbY2vwRd6k0RohDwtfNw4oF
BkMN/AQiWHRrDB4d7zZ7R2PV/H5o8fXdIn2Xe1BDNxEVjYKnLVDRVO+j+bzueAfZ
tOjJb4gMnqV3PQhRoVRdnVsu8aq7cQJgMKv61r86WyG8jmAUsKmszp7bw1eYZ8i4
VtXR+eUgwMyDmPvbqmahbNdiO8zIa4CuT1rTK5U5y8QO2FNkSNSAtwdXNInIMLgn
UgCPs3RDmQSGI0b/3nbnX7AZWva8tzzS0AIA0ggrkf/9xxxpZ/9lka22/IFyU9BR
SiVdo3VjyvLAkYBWI24yc33/yGPVZrJoD2kLhNhazbcgiq/Al0Uc7cBfA3Hc/XJM
/6gfa3gpPpB/uRZ9lYQd4KIkv1rfABlK9txAKyRgRfHK2rfqwwgAI0KPmHwVpp+8
hMid4tP1srSuyLm3M5jrX4aw9U6zk+MKut+Np+5q4olSNSOn1G7grMz+wsnO9K3b
Ny6jqWVaWwvvfKc/j71WfVdoRxzCFhCLHCE0h1bDQSjjJC5UrVVU6+wFbiEngQtb
AGLEY6bPlHPgIWPcLV2bdr+eqF4jFLcYyr5VqdmwvCjiV/iA5ycAm72A9julacig
fK2PJeaf4LOESVEEuWNIX54Cbg9xp1khLX4gQpEwBwPrDoSIeLjo9LErXIIkCQ7G
j9rDl2vSj8U3QCZr+u1A2bfrtH8n4oXOwDq53lkY+eozWZgt8wKsHRbJZk+Z9gzb
i+0zfjNppejmxCHKsVXrPVVhakqbiP5ibSHxAD9bMb5k1QWoRS+nS3eORtVkuHA+
DVRf+kk5S0vdwzxr2HEiE5HZLE1RuuZsYtHPPGTPMX1JI+00bcG9h5vsHh96pBBl
PrAkIR3MV7aqAhv1A9Ods9R23trnZL5lunfrIEJ0UdDcP7T341QwnCrrhX7Re/uQ
bClp3zAac9B3HrqoH9nhd9T+UaS3KfVHZ5LU92acqF4OIwIpMwCEpriY3S5UjxG/
KDw/ma7g+OBKb04fL0e1FPTUeZi8M5TXF/aPAWvJFUhKlHjzG1jZc/XvGQcsB1Ws
J6fRUmAnxW5JyPejaEwk23eBAcFIfZ7cRpz06XP54OSzTQTscxORdzA1HmMaHTez
iatdR4DOwKGwre7CFoDzNlbRpX3GwwwyWIHlH0mfqYhg3qpWyyGogBvL55DLeDVk
f1J2PRfju0bBe+Ory4v7J980IeuJQdP8/vU0xJl575zu9OT1xOIExub4qTA0clYB
aGcqCFUwvLYiCp90n9wpURhMAQRr/plLxJlp4LDRyPb6tazG8fn4FCdiuSIIhX78
jIgBx+ueGqttoer9wSdrx0tx85kr4+de95WPUnEfDOhcPAghgSbXWfRb9J1Y625l
HCIq/qQCosqPubr52xnhrFDjtzgez4AsWhRCrxa9kbeoW8lqB6hgf7UFgmcTUijw
VwE4OPAes1K7du/33N+cakpWkrKsMYzq0bw2dtiJJbSQSSloTUW05SdrxArw5cHz
C3M9b6Ayu1OmHqaGhhWt80idxnsKCaR2hSJmiob97T40MwkYG50ok/PdPfnF4CLZ
HDnmIoAxv3sq18ncV2Q91/OGTWfyRdOwYw1VuAZoQu3LQTaWeq0Lc+zhm4fsZaMJ
7oJNCFNZw4A0iMf8UWNnmWp8RfCUR8i1Ihh9rMjB65R4gZAPRBsil+obRy+dKAlm
u/s6Z+HT0xk+fPpa32ZcB4rjMhcQHJkOwOK9Wt8qrKItwMu+0oadIkUr8le667sS
O0NA54Aa1xBotY6K8dUVupGNEyGQYLgPBeatw45LTthFgOufDCpi5qrX6F8X40v+
ZbzZGwgbjBGmSSExuP3L4TGDNtAU2+ZSQDPpLHuRAhrTI+LD8my6SqGMpv2uXmDk
cFFe0Sy5IgNHq5R7i8NDBVEWiYPEbe11x0A9xA7HcONA3e4ykdyzvNDWnqbVXQ11
e67nw1e/KOp1X73siaSrA4XQueGBqVRdlKue0118E443coLNnPGb9RFQRREwup7R
O4l4JalsBGNfBZgcuZkemrdmUTlbmvV7Is6JE52q4iKdtpkCGbZyv2rsq8Rv8/z/
L8b/wijEEg+BqXq88UbbJ1inC3RpfEzordf8Oba5uNQLdU/x7eocQgYGlZWcqTtv
lHfkmP4uhC1iMlOUvg/y3vl0/X5vtP+26kcvXlyX3bUVFiNr5Q8wozOntKB/kwwG
8XsPiLqd8JrHEraqyKnoP7tCapMkqrKtFE+uT5YPVbId4/XA84YUqJlQRgOYDQpv
7MfEnpPO8BSiMeXD5hp6m7d6IDsaftQALyPNmGQjWI9Z+JmK6DFf2acrTRKS5Ijz
niEzgNh4WvN98dpIAiGpFuOkuFEHMBepfVxzdT4zxOAHwp+LytB/tGNSqgsnsUSV
4V7t9Y0D6c6H4amA/YZ+89fMSzIXnq0UaCxEj+257HNOrhatp1G3rCHpVBoP0QFI
kCzEkiNhYeW92H8UdP7FzBkPRErj4OEP/ok6Cw5FB4up5/2JwU6vQAwjML3VKmYV
kMvSGUI4jsL9OPVZlP6Cs0hfdJ88RF/ARLn0T2IO1W1S3K1u5t/s1bL5wWf1PTL5
ObFGVXCjmx/ZV7ZARFezEsXk2Ge0ymkX4ANiKfu6NsWJZ5Te14b+Wowd9VSFe5lE
Im8vCbYyHcLeKrT6olQO+qcL5VaOQXm3ZDaJE6saIeS3eRJP9LHd8Swb8UqRttf3
Xt/TIJI6ttwLhtFH3MZD7eW9ODe/JykNDbvIsa1cC28TwgLyYEcXB8rYSUMUZciO
g3xuXrn8htEZ8fptKWA5LFcSSPSi8ZQwwYszfyf4RqZhJjsc4ddY3bnHDWbYcygp
9mOyXZqKwIcGu9xfqVQS7tmImBLMaPpy2RnXQilFt7eARSO2bq7yxorvjF2+BKym
74urclnLtpZ2MvukEonbWiqCIb2+D5gsFoXThpnw5MICkAkjK3Uhn11nmYfM9Eon
Q9ovBR2kF65O2q5j/aWivhkkQOqxm6/d1et7nOP3ZNtWQAgwHcEW7HdemiFoilu5
YR8yf/NzOF80xhuYxVY8SX1gQE8IA4Y2eZVaB9H6NJ2VRlGZXja+JtAnELxywMhL
DxBi0vAWfZ/QQ5a83EOUgUbnXoXGX+r955vXZyJuS3fXKq9UBKeThR49vikrYPEf
PFVmKrdldhVieTpJ0HGrBYcUAisHPVvI1CAkGzyqMqiRnfehfXbbMFRwOTLFOtdC
bJH03IVbhOj/9hv93C5Wt8Q3CYviB7/uTTG021Fv0E7Au1dTPesW4lCQjGz1/BJ/
kYnps/l/nlFzI94XRXYi+zMiRq66lBNCAeWq3VgXGK7OFNQBq7g3KWvEvZ56xEa3
NcL6SR+qXcM/3iwMfSUO18RiC+d+mHjjlwOkNBctHik5FbJMWuRu+ZNFOvBGbqCT
kFEt7VcLDCtykL6eYHPG2VBqXJdatNQgz2eeaOYeNDKRmmHWywTRRUtLwaib1fOO
RCDBr9QA7hXpGDvwc4W1RO7A3oSeHYLZQFa7BkjOkSlyE+KJdcMbq+A5P9RgMh19
fyt0KEFMJOdBQb67oMAougDpvXhyl0iJBQSQr7B25WBZyHE1AOLWvo6D0A7PjIJp
tMUEDpwky95MlZCzb35GL0uCnKaraUkfsVuk8gU12O05NLEMW+UaLSb587zQ6Fjc
nrn8K6AYgEd1BDAKItrKMMqqrQLnC4Bu/1Wkftg/4Ymjl01/MgByLFnizG3AE/eW
98t6s73Dp5NzmD82Q7ip8DKKFv6H+vRoW3LSdIhbZboX6dRB9JEKmkYEy9CEG9c5
mIXv3GSHogrVn1SklL7WHCYDb3iHF/zjXq+fyCWQz1IbpT+oqY011GgdtbCNgrc3
7/DOVX7qrBrg4HHFY0yXBXfKx89AfANfc58ADVrYUJ25AQoDmdBbtFX+1m35j3le
kq8Per/9rqMtiDaR4d/34KdXXsBEyuamxW8NQJjys7GuJZu6C96Ewfco6Dfu/hlP
ZHpB1SglrlUqapi+cv4rxCIiW0gX9odUX0jV3tuy6mMUdSqGNPMHqLtYi2pjTm6a
bak4R4vNsq+NkUulPrYJyfyLsXe40/wdPRFA+REf0wHq0ktV2y3pfBhquTJTA0Ui
mpfRNIYajvX0TRIEuKOmOxmykpLPYhm+PvKTLjr+mqsSUwTtULF3/PNeKh4FgdAN
4J76f/kHMcBkfgc/elNJQF9WAtDpP0a49Dmp1s34pczRVSuFPu0xI3WeK9+reGLy
h4C5c3joqNWrqPrIJLTGQ9kzCLelsuLiMN25jqmymTEYuaozPnhE1SQe4clPSGUP
hHEdwVa8rYcYWr2IcuIY+gVNzcgYKI32MMlIEDPd7pQKNPN6jUs1e6axQE7g5Ain
sdH4xHLyCEHpDMsPLUWNDGZjV4TithLaYh36PhnVaAXjIas+Zmrl1nfdTFbzwZ8y
oR17NDLTe02uW5OMPRiklVSELq/SrFiqZ/PzB7axwIH1++jwhpxLaIZp8+XDBXvL
edNL9+URJN5F8a2GIZYfCpOm1J/kGITR7OvOVgNsYFRSYoHy090/QO5aBwagCwrD
7fmDWjYPym1yz3c4DMeK3odA9GDNH5/VLXDqVLCZGbVbsLKSEjix29dycyx4KbWw
/AVyKDXifxaHNKi33ar9WNPGBdXsMT55nStwtQdehYuwxQCOH36IFa18UOvLCpRh
+z3rXER9Eq/D8pK2peuHqZXY3vRmj6vToUSvALiHB8D+vUAYULhvmAX+/CsZ79gt
9W8F/fAyGy8VkszY7YEFYvRLWxInciEgK6ocatLJaSYE9mAxUTIV4/duSCA9ogz8
9StMsHS2cKYjUkLuiA1mlxFVQpwDm2Lf5kqFgC6hIHXldTL3NjFioEsSWf6txgnS
dawNz+4jGUIBnMShjfejMchv+YFkaq4m69VbM8c8uQW7xUkCTJw55uhzfKmtFZY2
DyuSmJk9IaSaZXYOsI8ualAnvkiubfK3iDv21cIOroUco6wb/U6LSZ02AvUfJmfP
LDIubMvtJ3oAysidZyiegsXd44EcKvfdG1AMXe59nktQJawykvvaIphjKQV8T4zP
SVtiosTZRGEggDKAuhgtDacIeifxiHy36hGicTBmzTrPxfQGyI7E34bE2c0fmMAq
KbumzgJmtjMMPK/MVfceC7NZNRwLzJhRuvfUpHJeSl+tUmCfMTr7Sd0WEv5JaWVs
iNGSsQfADLSQEJOka2P5vIpbfxixI2SBQ7DrougJE9/DQcgxF0S8AS5ST5xeQxzJ
vDDxgzTl1LECjOwHrgj/Z3r+CyneZYZOg/qE1X6J/KWMYhnZZ0MaRjvPkVP9QyFY
J1EaU+u0E9RUVqBxigpxSIfZQhiNmy+5/24YBxixPr6vE9uYXZui59OFDmikxtw/
d0hsODYlk605eetjsWKDcY5eNULIIr5EGqtz52kw3g1R0P9AEfMWDLdSUrP/r1pw
+de4at6IgU3AIXy8jyfmiZ58Z5gz7qFcIXVwaA5vKlmkdvtjSXGgyFHjst4lXsXi
FurwLg4QFU7AA7ofd7Sp0DCFbOd3qLDhugtlgGzE8YXgEqdFCFZGsU8bPkB3cnwx
umCbxz65i0mF86/nQFHg/27TBfTtfyw10ZoyupM7jjFOKfNWOd7/Htk0iStDUKOc
CPCil3dFyW5lyaDihc6IUQF7ns/sLrJ9Ame///99aSOaZVwFJCZYthg0hkaOaCc0
yca3zcNLzvZbkWWAAaNBDsRQ/0j6A06qVaXjd0KL3RpiyAWubHKDaTCIcAPAVZL5
sfQHPKGwHE0ee3FwgJBCdOCyvC4C6oZ0AccRUuBmwjvu5jSFaDP1XckXJC5dIco5
4v59vcSEeUMcyj2i8NQ5JTFY7uNsj/7pNRSfqp8A0e2syy4HYXywvZ2v023RhbjL
v88WVJSS4UbxFnq5pFUFz/uMS5Tt/9utSgcIIKJKWOXCqkk7NFjU2cWy/sOiDvNn
y9+T5EzsT8A6nm0M+7qlCQEYgYUJIhgIcmZt3IY+W4Ms6cfTzJZVRUIFYyiI8kom
ZvGvcgGqL3HbDf53Xi6hoxYgm5XqCe35nY2pkrFyqBK8/vuaS9NvsTTd9IiX/6M6
MuvtD+KmvSoDCbEVLzR9jcRpIxzXp37FuxAeCEu/NMeDaAnED+EEapNYhxYX4Ytw
4w42uKNcqQ5WqapUhgljUhSQ0IVIWzKBiGO0Nl8RJ0Vr0gde18/XOl+6b+BYoV6T
R1trlEghV9VzmAeDtV9y2SwwB3K4QKcUTtv7H3w2JhGGR4zzcksKg8sk/y0X/I9c
Ytc8ETagPhp9loFH5reBx0+FmijVUixQBK0KU7rlZ7ZW3keyWSV1/6OL2jc3mHNx
Ihvsc0AGj/DkggTpQpZRxMdDjVLIVtYiG12OmRjGNpDwrPycAHuRiNbPtVps/B07
XAEgnTp1OIxSSDCg7FhBCRofBKzHRF+lGr+iZyxryGfWRSp0HXRnaFOOAIpIxq+H
vnJCGrQeIMc7kxEtIYLgx92gb7sfWcYQr84vwbLnV2sasSdJPocONdc2nQzHL7bL
y+bhJ6SCvsn3/9T2TkgxrYL9y6LZOQEE52ZsZr1eO4QHS8wqe1OpKn9O5MwSoyhd
yGrxpTupjR31VIdxVlWdH4rCR1Yk1Bh9KulpKo/zP/ojH1cjcW5rOhzNcA58+gGG
6N7xjIukT6LbEwy52K71oDby3yHzKzqLKjQJohVcKCOlid7IbsaHiPpd7vlDlFnr
69yXF2Vsn+NaVMVvd3zRT2xU7Uq8Wyl1yM88jkSyy0o76V5rdClTK0qHoqAkJ1Hc
LfEcgCoU0+tZdBO9AmaAZG592tOMHUnLB8Hutruddal4b63neD+L//HwIvy+zFAK
jZjDqSUg4cJe9IMMDVt9lkMsBuCgtRZV+nbB6F52h4V0QYHmqSOutww2L2k0CZVp
noMcgdqVCN/mFGYLmZuMcC+qTlubPuw7Alugqb2hDa8b1OUeBPZ78DxjsdgIh+p3
rngm8elvudntfsY8c2+UmPj26e1bWVSe3Z/2zwQNk72exXeNkdGsD9jjNWSNNuMd
+MGjXtMKQ3mQjOhaq40HmeM++NxgqoU/vSTXA0Kycf7sulGNqiM0tAYzci4T8A85
Akw1KER4ZgwscF5JwcpqywWZ9T/5g824ePY0quFtHOB9QJyRdGBpaG/LjcVqS6de
TufAnd5TtCkVhWkKOnSj1J+a2ElvNECBRLr9FSnz32P4avvOFFHG5rTv02RzQXLL
MfSJNL9CJeuUCu3fzSyK+RBOaJAQU9PtbY03It1SLFiSqBsp4RawUWaSX1D1VN0P
1kD8xZHgH7F9hVLtqTH2RZfRYZRU4MUs307CDKA7nDz1M28yACiquTh//CZCvil5
fxbv24fx0mbg73hdj6szO5HtHn4wxDPGGJKFzCofV2IBK1/cPOMjqFOMbt0iKn9T
II60z8XAmoSW5f36xVMzO2MS8pJH+ViRhDZ6LMUd5PRrQvd3tH6tO+vwnTlfc8dU
ba0qeaNPSJwxMp7BkdSXWL+oxecP53T10u58f7xsNrFC46PghucpwBi1VArEHiR1
eo6feJvbAM1epb04RHEJXFmCvPhckrFwsdd2rQfuVlhDLVQ4iKADDCeTuRwPS8wn
xZijQsWoJ6pK5ploHywAZoA5f6EZBC+srdyQoAyLiQNZPOkCWMoUdtgBG/UTQL1Q
iyYBJGr1sWfH4G3/69yroJsUwBAWIS1bq14khS9HG//bpDYIFIvouqX0kOopgTeT
6c85Up0Ney/4TihjPCOTtT3MZ0LwdbJCay8T4kBP0r6NVybcKEmXNoNa5i+Zq5zp
YX/r3xo2zenHcqekCJj3DwTb0repOzZUVRuGbr1si6d3c28/o0xaeXJzxhj+WNEO
wXM4EYf41OFFCquH7FSuIdv6Jpzsr8vxrnCpiTwlhQVJObrL7W0q5RXqSrJvvA8o
V/jZkgXgdIVFQ/kF37Qef7qfh3QJ816ZJWbF+fmCMTvu1nzJgm1MTrnkEFzXLGow
20iBBMB3ySQD5ugm4R5pmvMNFe+slokgsdfK8GT0Oh32ovtQWjMbc76p/99jHtfJ
LW/ygzV5IfygsI2En/1E/AyFZlnMbuz7ntIzqenyv3utf8p/UbIex/w0H6F7v1eE
OWT2dZsh3vI+wBezhhXBapMGtCUg68IIbdWim5AOLyNgUjYAFOyxUoZeWoGzUC5W
1skZVlkOZEawuynTA8jLx4Q+ftcQH1R7N7emWBzZH3t83+W2BoAE8B+mImQcXoRR
JMIdHQDMRb8AO9iX//RytXDFEx6UjxqlhRT6nJau6eOuKz4kWjk4idKAhCNCyAQp
Q8MP5iBRwxg9cVy0XjHaeCSy99jBKZ5H/+azdKFgsFm0oBp/Jb9U6SK1Le9/EcfK
I3PHe/eOU0iX7jnTBrglt7+Z4A7LdVHJFYlleZMWoQ2008HzXesiddagjAocwCwI
uvdiHodYE42sf7UdsWtqaxyCvAayYT1KGXfcAGWM3s3fWRWVRE/7aNQtCWd8VL24
i8OWPR++WKeriqxG1DmNGwMqnQR1RiX5Le90RLyum7FRw4z7P1qzjfsoF1GRu74/
dPNiwlo3mqF8zUZzVvDbBfhNYk0wpNv3vRjK0zZ7ilHsQaokRfyO1cAjn8vSfEqi
XqypcNknNgGSrVAqSLTzENifLFakFVNw73uH4ofOTAl/9BAxAXQSUl2eUsMQO5Yw
hFblWnZgwXUKVszD65wRvZVnLNS5hAHnKq8uiJ/jcwDCVH9rKcUjbD0racZKytLN
jR975DyfgSCZrXqPAYaCfqAxfPE/vl84PcSTdCjBB/+68wpn+j2huV9mHOgU5bby
G2VrURazwr+3wnvkavrYU4VxAe267gO3/f7JrTDZ3NZGECvlbJb2MwtZq2kZ/qTZ
vVvXSFL0XEBQbWwlVLZqMHMfyn8dFuqErs/P57oul+4aYAr1ktF2/EsIPSk2Roc7
7q2UtvI8hmZqqc1vTd4QC5AkIzTa2P9FHJ0vj6te2k8rNI+jYU/CEo+YGXlls+9H
3QdpEr5naTVaRqDkaidXPz9QyJ4etoIOgSJIXsw3XeBdwjRsZM6S7qSiqSRQnLlp
zeI2IpJnl09WztTxBFhzgi+VNlXFYBIK5WMMz7ksKqTm3oDEFsRPHnmf/inOYKlB
hynA7AkGKsBoqRbdgBRuAhU5LhxgrvE/nItggA/dGl+b/LOEQ9Ftmk/w6TOQs0gJ
GIy6kwKvPXoEKPQGHLlGACJfLyif+VlItSzMUbTpWc5aW2eur2XR3xZN3XM+Qlfy
tztDdZ81yqIZHjGIWXlR17O6yNhk0NSCfZBgwBpP+Q6Q7QNvXyW5WRENJZ0D1ZYj
coWCUCi7vRffGmUbtE82avlw2LYEN1eA415dxKKnVcoZNkijYjnJwNZ1kH4W2l9U
wSZJCFmyVx1zIFIvbL0/J8s55mnsjFujM8WAwzIlPYr7N79PehOex548VVStzxzB
/IM9xiiDePT2bZhg89X2xRDIeRqzhBCpmgbKUFgk44I5VZdjbs7z3CfRbw4nm97Q
nMdZsrkNwNtnUq092imLUUSnRyjw8D90msMge7pR8B0h4bzBsonNe+PmfR8eQYjQ
Gz3SGMl1ISeGTmb/FxUMzBg79Dmah+jSorQj7UZ1l7CnJ+KhAEnVgnJ90SvhE9Cy
7QOUdqm3EbgBN3l9wZcCZC6zs3k/oY/q7dIixeZmsvkfdGiXZta145fgnQyzBlYv
xjKBhdyZsSkxvTgNbIoyPVpj+uiGfz+wONFuPukwKXfpO2b9rkVywdcCu8umRtMi
irdjvUKP9UIsGW+jLKpElc8Nge9G1dwSKWXOYg1/hvo77Jp9YpQWXygxWasyh/02
WikvxsCMofFqrTOu7R4Fsee8FI3xktekQhfPwDDYt0/LaNSevKTKvZQ6Y28GV41J
hvNK+0Zo8zLEGRQwp4haSviE/3qfwf8LmPCnVxKYYBeEaJpZ6RXFJjE9BOgT6Xcr
twCuN46XYdxfgpIsdztymIdyNG0g01HzFo6VQdfX0WXPtMqHW2BbsbRKU1cyG86n
CuhAUZ4KGVs/jcZlOZ80FbKizwipXVjc512BkeKf2n3Qp2teecoumu0nGiVPlRBA
IJIp67h0KYw0nMLB7nl4HET/2D3x4r8aD7mW4lxg7PsL+hRCRo3BADajtT6b1MuV
ASNiksKwT269aNeOW3CwzwY7NtyHdkxpBTqmTcmXOFSGJVuM9QM3z4vikmoG9iZA
u+LohSpqrSnvU4ERGyWzqp7j5hZiBPdPVkJK/YalAJHAgZMeuji+gqiLefQ6tVIo
fCrdLdEMn6Q2ONIvgd6Sua7fPo4cF/wXEjbezSHUoboPueq8q39aEngqhi1vk/yW
Zu7jGjLtlcEnfil5OhG6e9NOfZppG8RKrFFHoXj5abjWuPiR/r18wmdUcT/623q4
9uAXyobUXf5R8KMNsKCnkdifxqKjZlCLhubS0WVfWc//SHENBB7U6k0moI2kEfa3
vMA7QgVksT7YuilQ3n+5CS89BC9C7zDnF3IGIfJ3NDKl4rBwjnIq5BC1mFKXA2Rr
gWgk7xCipyAqY6hAU02iOFvLIN6rZydvEvd3z1y6dntfN3scikBgaqm5rT2YRNqI
mJEMLA1kZFd7YE45AN917nwNaxGRL/IKZHeYyhHyqvCNw5CfWHJ1jJ4JN1avBJRo
mpObDyLRHnvZUUrmhL0ESjSpqXUNiVBU26J38Wsr4toN/AxL2gzI0XLOaIAzfDEK
Ztv29DqAJk94JQEZa16MHoU83/7U4Kmxcgvt4G78+x858RFEhH2eJ7+LfTFVeykj
gHGZl1/RLIoY+pjVauQ7gt8diTlX+n/rmidzjOdowKeWEMqmo1jn0P2Xq5eF+Hjh
Iwy+IWacrXarahX207zUNDvi6S3D/QOGZsSNAtrfuJKjwWJ3sdlEe7YJGqexD0u7
SR0PqbT8t4VfwDMKv1Xl7+Eg1KwgTJRLYpOz5E9xCd3JFxgOSZz1EeYl5nkv9fci
9XYNHHjpUlhzIT7iskleWkriNEj+WnHydxFe5XLn6t9DnKiBO3TDv78PTuHfudgp
Gy4NSNGJ5JIS70D0Bkxk/nTtfvhbE867GVfbNMP6kgZ/oSZBPNjQBLxWxC9PqJaa
L0nhX4VFCUSN7oapiRqYjdGGKPmcVB8aZfbvWytquMSTTPq8pnY9wjH2+FoXGz+u
J3Nx9enbvuLgULIli3atKHy0YYVsAEoCjNIZl8sP4hBp5iOh3wM5e8G9cvQVxWyx
k01fyKWsEpe+aI6NmmvwfTZzot6gKx6ESdaOK3n67vIfHktzDUVd6Clqi7pX9xir
lgvf45KAgUtFicJ8+MfOQfh7F7TwxDRvjFd2MdXZPXL9X7JB1xKzbdfzmVHSVwWD
3Z2xXFzjHIWV5jQ99essvTYtmXOAFq5pIDk+CLa+oPynXiuI55VQq+idOU/0IzcG
l/gtPI99Whr5mzHa9i59lKqheb2HVbO/g2SgIP97eUACVatq+ysXNw2/QW+nikvk
2weVpdNKBUN9WSIJKIzf39CBs7sg6lPMnlz2vqwU/9xOtWDDCK5YnrXOIk+AexN2
uRnNpAH68GIRFLOaBLXt1FrvFAtWfqynj5Xy1XltZC3g+cSOnPEjGaTPl5bgLoWl
ukfgMA46B2A4strsRYR3gZv+CDxKprc54+MHTEg5rlGXAFYevqjZbCOHiaFki/Y5
o4jhEF1bHevQYxU5GpAG6FhDR6udT730rAr0vFfBchzfjUvqtrkB3uCdRiBDaQ1c
LftrGKSXaPW2IDnU8B8zJl5u1wJUgJX4eQeNQZHnBarKManoZMFwHklPowHjBoc/
St1k3quf3GITzFmZi/pKKqFC+SeRYXK/ljPE1rjFCceGdLvm8SErNB00x1QUhEjz
FDA68lMBP03nr3KhJ1MEFEknghF8bm6L2YATm2jlgk+A+siGb5epExgVgelEkcbh
GqmFDWgDFc4lj9x1gZV9SyeKAWeaqu9AZ4rrunXo8Ihuv3pDhn7v/c6yi+FcQ2vD
VncWaUR7WQHGf1E87Zfgp5Q7cb/v06MzczCeK7gcYPYHRJ3kSxHNB2+4LEgVAGF6
FnjL5NaKOccYuiGrdSofDtRRAnsMFR/0C15BMbgvoJTzG/vHkb2lP+XmSibf4FXZ
3XW71QJBNEBxXOfSwhSR4R+THhJjqOMujc+xMZ5Oxwak+mdCI7+1NweAMbyltUPH
gCbO9Kab9IxDIFwpZ4TqqfLubkf+Ew/SRsMGxe48DQ01Qsditx8rASdfNafEdVSc
9Ld6RljnxugOxE2/UGC3HuQ4q5waxobufmeGjr59vWFeyw5H4c5shlvrEIIIKKLM
8SSTJ1NjEGKy8XwAZNjLsrysKXsX2e5Z9K8ueW6/fW1ot/pMzk5CBBu69fUYsdlw
z0PHf6rblObOzdTMJeZXUZEfqEW03gefgD0oP7ST6NGan+wqY1d6IO99CIPCFXd+
J7OxQqRKrkb2jssjyWFcrlIS6i1GX0wZ4Cey4vkYJryWFeY1Ykzg+Ta3Ri5fDa3o
zjDKXXJd2ri9odt9XLVTZQv+hTgfFkrcE8Oqn+DUefS2ebjDS90pcB+YAGkXG1+U
glaiPbqRuijtr9j0pxag6KN5ohd3zULZ5eed9fExKfncoy7DqFAem85EYfLt6D5q
iHG7IrBlzaMD1uTW1okt6Z1kHlDeEW+ow7aMD2vrDT8DqUKL2fyMiEQL1TplRz2V
Uy4gtCu9/HzZlGeuZfyJES7X9YdZN9WE6fwAQPFqvaFKTQ/bbsNHRjDDl4EyygXW
NG5lSlVhrFp1ipZNn/pkXzpvuuTfW8zX+gye/2C2kpfqfYaWUf1Ry3h4WoCzKCQt
b3yRszDk+2ZqZQUW/gpPqJGnHweUZ1uBqAKL20P1L/28wyeWkOLLptMK9vZqtljf
b6Kj38aqO9uHOtliQkxkKPXFj37STqEzrhTCaGInbOti+/oh3q0hVoP4iv3C84LZ
MrgJflreeQ9F841LM9yKaqeq4QG4slznjhBlBLJZXPnNde8N2y6E6L67t4ueXn30
AUSptPA08MNTBt9qa4IFdr5Otl7h3rfyDSHDUexSN/5pE5Wv8+fp77HdVOgTVNI/
X62v4HW3/CGV0tefx0K1uzlk+KnUiTKNhnjUZ26U3CQOf4VBiZb4k/rJOdnBPcZE
WjORqvltMrwwt8jd6trw18PmmjDXs6z6ZUsEFdHCw95Mp7Ljk2rWTj1dP4IGfvap
KObtDITkeQZE3Lq+mktfpjvG7JP4jvtvTuIMPv1/iY8adq+Eyp4PO+090mSd71TA
gIHzQkNsCsCTvwpAMiLfdzbMvaPB63tk/ScYMSuaymU9dskXiJS90ugNvBfu2Q6R
As22tGzmPuTKZ1a8U5CsJXWf9pQ30plaPJVi9Fyf0pvfipOAGY90hRpdBmPPPGXo
ILDaUbATjJ3Oa5j3/sRxNe1ZCveJKDcqTnV0SqCVcPrE4Ongmb3ZjXhEbBYuTWIL
OwunX7lm7Txl68xSxhTS4iJ1WmMnPgcwkZo0DKziiy4rK9FgwDv/pVVadHOR8NMD
+IoaRPYecWMIc/X0dt3TwnODcrGM/QuybVjJSmReBVxjxdIDxg5q+nB2Sft0xgDu
9fzIEpTNz5PKW7FBIy76L0UdyUewuhNgLrbEKiqLnXEmInlw2KM+PIwkCloBP+Es
Ja7GjbpP1Iuk4SmMlPc2OWeZffmCI4pfpnsmDIJweGl75Tk/Bsa2l5Pr9IRQejlt
ywtVVAh6Oi83Q6uESazGaADLylNtYR8t7ME7v+TmEFWm449tLeGbh6318u8WjenZ
xkv2jEXYNpdKYhcN7tFtKjHQ7zkss0cfVnSi1dEE9ax+WD9Hjgjx/v4foJoZIFKn
Z9e+gvn4Oji/plNgUnaslvwwaL64hZH+ZTSFwBl0sfBa/3a+6jSgoSj0iUMDfvnj
2j3zUpcLYLtY/Cv4Ef72WMG6TWKTANJeoYk6raTNg5erncYEx5tNsBwqz4UY4qrB
j7ejfAnzadC3wqiwwenF7j/nq61W7ZmEsN7Q87q8snzTpQrQy3hxtqQu55gc8VY8
cL5EYUYiHTTLEpm+wxwBBznA0cwesLwrV2Lu9ZDrCWcvOK5WY5ZnTDZYcafNYLKp
5QKekAuDInhtRtSJy0kwDFE+cKl/QVuZ9kHrNUVcjiDkxAyVpJjIuic2+tBu3i9P
tYoQHeTgjl64Wq5ZyvuCeK052/6EMNiQvx81oj1E1CmXvThpQcUHnQd4i2XIGuVf
xeSfRj2KKs0QBQj+SNVcwPlm0aQrMveURK2hFAgb5SBa9TrjA5QUoiwmGzQq4FNs
MPF6IFqfhWfWyG/9hRCRD623IhXWeUOjGd1oDfFdKeU2YemwSwr2fb7gHtK+O8Oz
7RGOErdE0uigsCYR/uMxjHsLUagWKcgi5i2h4NExYkf8DX8ne1mNnig6HL1ww4H3
OakRsUNepOyKbd9lPgiAFORy0bVJzURvNSzVfKz44oLaLq18hqWXnrJ5Ungx+R+6
Eu9fUFqzGABHOrAxKVG/TG09yv9+sFIs624BepE370kiOzMT2dJrfmhn532t2dHr
gtM98D9dkDRHEKh4J+MH0XrZx+FD0sQ8ssQ8/YBIBiYe8qqAh0amdRwb1NLyKMJ0
eaGracB3r9XEw9g1hhMPR3T3w4+HONfVWCLlYbTsA9vephNi3JsOhbygncvo6FbC
lWpEJoO8BZfWTze4Zc8uvMUXwjaI7Sdzl92cVq2hSMy6vSr5uHMB5PG8cjk/+6z3
fTGHUaUgeU2kUGh3HXt+1mCe41ktvfeeRMLq5c8GEpD3qZODkwlp44O5TMeeXnJQ
1lNe8dJUhheWdkwwO3bjzGJjzWgAJZ7/YuH4FzyoPp5NvvJpStWzjE/FxMCQW3yf
DaPm9aWMQz44mQhEq01cgH/9cP+eVHrSovf2VzbgY5LWgVa27gJ/tCl2E2n610FY
K/oo+udl+/kS4os3eSxQHfLqXgLBHYicaojpyADgW9dDghg1bIKrUsK4OjUNSr6i
u/hhfAx1VfKNQaUlRBTOFSlUPj2RDBIOmuWJl9dFFr8TE8euyR5GSV+WT5lbEF+l
kJlH9BPv7UvXPJU3j+HAtm8rapj8LUawrL/Aqec1OXJMjIPy6APt8kHoNhrMkriW
Kswoa05gMFTqILujNilLouveL9jWdk5ZXeRROfsxxUq8zUSFsOzPZSCQCMuJMz/G
gD9QrXBflbb69H4Abt3S+m0w3GO7cYGSEz1ISZL2rxZ/GnLawz9ekhdqLp6Ddmtv
33snMZg05+8mlFuyWN2609tuX1subB2VchHqBScKdZx0gulyU1NDxRKvqaX1/x6U
xjr6noRwLDIFVuKDq3yAM/bSpENp8Y/MwiYjhpQ+BtnIgCYHVQJI0V6xe2gpVqYV
BSyaXYbt22hCGrBQWnBVkWjimKCsLexsUnB4n0rF/hcdFKiMSy2xAEZKpnQV1GFs
IUJvFw9NAGFGQVQdECnuycGK95jdVbJArHBJLzT83/u81VM+xYJbdfCrFXtf5clK
idy+vvnhxvfoyqC0Rnz19m3ybJvbLdX3VlW/AMG/T399i7GGQg2EgnIrelc7/SQu
lRcj8EcyNggyz/5cDrEDxyppUS/TVRlJeApP5m0N5C1ocW1FrI/Y/r2Qyau90Tup
hoVgHoRGW2FFl1KC6ekQDfNCjtmCfCpK69aY7GmXan6HoIHNKAvNBVzRLyZC3E9x
+KxaogBjpYZ7mfHzZhQ1dTXp+PvIXn4GBdWpJgMrgjKPL93+61KA2mtXOyloFPRZ
5cdVQFR/XdzaJ7LI4LhRhrK2L7kYySJLnxttHweLfS0QxrJ51tUIs6R+o1z1Xe8r
fln7I4BBTGqTt3l4Ii7Z0ea4CfWx3a19hDBtsgAyP/wz+JE81eqvwyvasfIkFOD2
UJNXvLH8Pp/2FxCKcpO1OoISJL89YpTqGVWEb04FgRo8NLfvccpzCgBvbH4BPQQf
bWFG5Rv84gfhE61VOVDYqojmrX3OH41/XRjB8zZkEq+I3YbeiTRxfQBC7kzCP2Ri
setP+hxDuvCiZNSY5b8PuFm4XmuPrZko2D1a+rGi63FtJCLsDemhFcKb8BWf9vJH
HaSgvk1Kk9UIJrwZTh/AflG6/I30163XGL43c3LP+OMwoTf/dxYnZMVYvPS/uNfZ
1sGaVa6EizcfPP9L20q17SsH8KhjGDxn7evJafJqnjHYYnuy4Ezfv++BHi4jr/9F
LniCrx1Pg/QZvCP/N0xiUZrWXXOP2EW5jpb1kQglv4QTXNZK70uH7q76oN+kbD7u
vlx5ZTwHnkKm8sJfmOAljy6ODSgBXqjf3cocbdKcGeaapwPeePr8amJ8T5zqw2TB
lq9WfSweL0LiDMAIUgac4y8CGdMZaGnCgGASTgvtKJgGSC+DfvfhgspaB6F70RSA
flWn8d7YgToI9tLSpwL90Ns5J/YUgw9imMn9MZBscbAAtiE0FOjbg4CTdM+mR2ex
VpnpBO/7aAukgrkZUFotabcFzsG2uJwUJYxisiOWGD0zzpIuQnCDZGfXpE+Efepg
Bpb8V/tWdU2IzqfdjT/MVEiyb/adFGNt4ECOJJO0h6o/jDalwHHCejjkzUtt8QBH
zi/9s6SqXgt2At1yc5rTe96UfwztKuCPR0FQAhq0DkQQyMVGZuw+2VnI/5SPRrPg
HxvQ75tEtyH5ajb5fm2n7Tc91V1TisaQ/ROEY8Ow9xxZk1A4wJ2ZpTPxnfCzEEu6
/6wmCCxlXwna1z7fIlTyB8NFajVzpzONycbPkYLz15CINc+t4UYWFMMqDy4La5Km
TxlWcNbsXiM3vtbSPsAtpUV5OV7yZRNYNxEpHnAF974+V1/cOKf7fv7i19kUVwmJ
K9BUM9/Ee8k1T55FWFqv/THN52VuWYWiV6XRN0ZKcZ1alTiuGLAV10DsDCFFU+a/
Eh9YdMC24/0Id46dGNcRhxqA3s5xmhgSgS7guu/oXhI8hllEOMkhj40fhsYvtGkE
PxVyukFk7qcSAfAvPeKbci8gz2Bzp5Eyl+NEcWuDOp+nHfPKuKFbxebdNwINco0K
hGBhEgImnB8cErv5wbfrUvf496TEYl60c7UBNWHyWw+i1PEP/+JVyzbxnH7bgQNN
xCpNE/WPUM3C6AeN4uqC1RXN6F/bERoc3DYXYhGFYLLQ0nw/S4LKBPtL0DXFsl47
VH6+SERgUVuE+soKa3mZToAzg+o3ZNIt4AP9V4hC4znSiM6GuIeJFJ1LXg1KFsW9
U8oTqS/U1GkYOhS4KO3PS3XdpweDUhjGj1ONUuxwuwU2OQUa2kkr2ndkR/iTxrlw
iDqnT9J7t5Va21jnM3O6RqYvceoAy+y3A9oSj/LhH5+hffvodxiEr+4pTf2N4WSl
1lndSYuwShXjMuGIdpvQwUdVvd6lDsa97Q5uqZantYjBDvOBNRjdswFqzDhO1DRD
2iawtdHM01xvUeaf+2Roix5pj/0NOK3xF9twLWc1oJPWrPb+asNSOc8DugrfvVJA
QL/gQ3L3gY19SHu4iMeb0xgNMrS6/jkbyYHpK2m5hCTQKdmzK+WAiix3EntvjVyU
uTyQInglmx3xW9UTR42NEgv0cOccEgNk46o2lg6ovpKD+vwWyjtqeJaNoNRnrw0a
UgEdF1UuXAe3iXCRHJ8UqciCYHSCJCofqX4Ynvf4+tzndpJChm8bqZkvaqX64MTk
DroGZNllSMTV+PqLHuTxZdSgFG4eR8beiz5v2wF7DL8jfWGzk+ND1UqToae1IzmW
QxRbS36bMjTHkb+VY/9C0MDAJsT9zdgcvFCNl7bRhcuLWo0dkfXBRN6VUTj0eBDQ
U3HBfrFuNoSskJF6D+K0bBKtYMHlgG992VfICodxGj6jptXjcqVt5b4p3wxGm4bU
ryLnRrrDajr1ThDpPxQ4HSQD28Kz3X+n/iGf5rXuAb4WzyKw3K1dnenTjPGiJrnq
GIfPnvaVXeZBSZ0VcL6wJ5arZqGXomQzADrvAqGMrdGTcpItFVIKKGesqQ42W7p5
S0ZPsrRf+E3dJQlJ9zqzS5gKYjn11LqFgCCgTa6HF+8YITswGb0ZcdZO4wawxETj
M0qvRukaezo8uRcTldMJ4zJtgTDAJIVEzrNxpScL9suWmSOUHVwFKqyqr/bDM33y
C63SXrhm3RHi8NKh1Hfl8VXWy9lL/Emkl6+dZiDX8XZo7FMxjUQK61O1HRdyR96u
bIEx/sWwAtxVUmXqRLQoDcnvlqR+uSkxxE7YBLaCtrqUhEJRfYdCi7x38JHG4et1
APl3oAjJo/hW2zBRr2iOWsyB5my7CZakk3EA4e+xQ18c19pkslbNjpkFyYp20OZf
I+v+UVMXjTC9Rn9F0jjUXnsqtF+RdDb3cNVOAQn8nnuT+ntgZgOSiMyG+20g7Amy
vrlD90u8bjS+mQ9JQzo1IWSOdBh2o3QQuePEluR65gyRPQBi5IiN+0Er208SntLF
yn1t6o94sdwUulGuxOTkSXVfEO32El4Q2XFaL3wX4QDGoB6eijXo0EJYLcgHOx6M
nUm6ynby7zkP4Ap2NiuG0oYS/h24IAUom/WqoUagqXOrbl/tRE8PlGvZ/MB5eBF+
0yHGiQVy+KL77IUZ7S7pN8abL1ybUUp3Aq2k+c1Oo+jgROi9jmFKReWZNSQRxyPW
ZhVtBS1586vyJkeH0Dcmc+q1H4hGl3Bsbi7NjXxLQlS8B5hy+fz3b7dLmFKRCdDS
GbwNU7iJL37vSivcKNDMQjvNUbm4K0SZ+0N0WCfnx/qjjp5TX+VlDwBDiTUthixb
AsPobKC2LEPxE32i18oe45a53HgYy7plJ/QJx3EkqfWpLihCbOJ6BW6D6MW503Yc
dGeqQIdhr1NAIBGPvOa9+r4tovbeySZlpGgHs7271uMFvTuk1odgzeYgf8ORuT2g
GCoS98kPgaFRhKoGPuGP3QgwQXcj4SWBZ+HRUFYGV2vgy/wj0ohB1AOZcOm4YHmH
7sX5bbrJOb3v7OI3O+BjX3WbA2S1LZxHy9cfS2FhftSfQDnPDh3uxHKPUzCgv+y7
mhx8tHmC+wJ3+ObJx0dGQJqRfom9Q4DiL999nYw5CF8tZChv/6/LNO3HkGTHi0Vv
lU3rp4jfcGKBFQa+SH2jdFkgSZvhazwHUh7SdzpzVAwghtbtzhIMYWsqHRpW1lqm
Pz7eZd+EdNCcvARz0hcaN5eKYzkmizCYsydhXi+J2FEmnDniQ8nazj/sjeezOB79
0U2F+c8V7Mi4Frd7ajjsME4XVe9jqpZFUA1Mfnq/KMzAlstX0brBPehOwoeSc4rb
+0EKVVw6WqIWm0IlyMfuhPkwP+6RKwzdadZryjRqUxwRjMzRFkTdS2jujF4tsGH3
oM4x7pXXG7YotAKm3Nu8iPeJoT3//3jF2ZjyxsVwm1d/aeRkFYPClRtIl9XWNdCS
L7xhxiBcaZSAF46IU/j672ZGo8RVPDS4U+pRjNy3Ko77YdbkKnfx3YpQjNQAX0Pd
ie9b4MLJjqj4MoEGzLkqw8cUZzuXYLdkSq/TzIvDqYUnVCU/HDaERx0ROvTWI5KD
UUPKEerC8teR4drEcDmAMQC/SDPdi2yrTOsCf6m8Cm4nEVubw26jUszFP+rAGEjW
FApNuxx7HiTQYjBd3B6VtadKdjhQR34Oahn24wr0CSavAtGXAsScn49NYH2sSp//
2azui2zXictsxM5jbGej0OAZOOgAlCL6NjrAJiEQdRauu8lFzEBiBUcM0KanKaVR
CTjWsag7hq4/tQrKmngMqpxM9f5fuWfrs5jqfoUGthAipqTwS70Tdr64Pnk2Heyn
JYMTkkDJWc9zH7ItcK+ViEHrqrRpDLwGquBQujK3fPUO2XuDkjZqYwHWL2fXq6Cf
jVKoSOILYrJbUfU5ePn8cwsB0X/zW55XBuYBqJpvWM3aOdV1abVJWJZQjEJuN1yN
rsoS2yvKnotaBwyG9SeCbuZeeiEwwgzEWhbeURvRZUqzRrK0Buw+NZ6gd9nfZxoT
t7EuELrS8YDTODSyuh4CmZT6p4O7HDLXzaSRzE4CGL0DLIqzQaTnYfZwULZUYLR2
R51zzwyd9+usj09KpWc4EDh3XEovw9Dund8DZVZsV06kIAoYvsqUBc7yQgwvRWQQ
Qgu5iGGoOh2cYkSh5geGcuQ5jH/TrEiXCIu9fDw0kLDzg2fz4fOGJX563ZESjizA
mIjIghCLk+LZ0nXt6IGhMTtXBxkCnqqsq6cSfb4VpeCr4iFKCRNT/Han0Jk0EV14
LhfAwvzqpaxROg0a7FuWDHaTMx9ipO7VROhvJiIY8RectrKl7RkWlgKiDKJ7Z3Qg
78uXKCDA65cMxZdRrGm26IGHrUS8RcCSPPCWI9l2Mj1w4qi18nU67YpFAmCSds3x
k4Qhv7z6vM1inOrV0B0uHtLYooWLmaBp+PICkTTllA+MnIf87mCh24f2nlxqLHGc
F0hvz9UdplQCZng/QVThszcNuPwJgTC3efBfx7LmizxJJdKYlMCkWskWq7dR6KM2
iybvwiFWOUP+LLjo6Y/nqg==
--pragma protect end_data_block
--pragma protect digest_block
Bh79GerW7eiehR5PXDsb7jq/RiA=
--pragma protect end_digest_block
--pragma protect end_protected
