-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
TgyYYWhwaQhtOBXbnRrMZZHLLPHw22SnB/ILEhHn8YCeCgMXFO5ZkwxylW/Q2l0e
TNb5t6bSHNDaImA+3goVt0fTWW6DFOfswFTdJbYVo/oKRqM3NGR+Jx+KN8ZtbxjK
GO6k+lWiLK43q/61E8QQHPpBDiyAZWx6kiy7tME5dGWNcDRFs3OG8w==
--pragma protect end_key_block
--pragma protect digest_block
PLeOSZvm3lrNGVgP6EedRWgFEH0=
--pragma protect end_digest_block
--pragma protect data_block
cRl4aSWiufILm7VL6WAIZ7TVEIWgH8A7axlS5nk2k0PGh8c/7kjISpHSCLP/KO7j
pwQRYEezYpK7PqYlbc30TE6OynEEKy5yTGC92ZrVzc0PdcT7XbWgMygU8bdHfj0F
3hGDtz8gFdUhrkloANNys+ExRpTwhD01/5i+3yvQO4mpO2Wvnyo1fSAWkzqaqITF
r4FFJF6ndjxejIO2+bxmle9xI5jm0ULlhs6l+T4KnYED8UEwaORUXtmXLD+2oEup
gGt5GWcGo5nLEgiClUTc1tlmXX/RlrEY43SpWijeJmk1NeOQuvS7q6249T90KFp4
1ObDVN5DrvIOXT080bLVIygC8qAdel/bCX+6Uy7ibzRfCM030Gfyf0hHe00NPFZP
oJ97dTBaAz4smqAw4pIu3wELAJzKXaEPDg+D7GkGA6/heSyZajpxVH0NJqMhpUKb
zHRxqMXJQRLqUqdVqAi/C7Xv4rtigy8fwvLISGsBoI/aFHSc3k5XeBxzLxZGcloV
EzRLlex4wJs5Wxvwhaderb7mSmghbsfmtdUrvWkJpK16F2wNueOurdHY426ZX+db
XVp6c7yerIl9nRZuOxAwUnKu8DY3keMBc4HvlNU7k+GutK2C8qFS0uG4KlXgtDTu
PBQ5PPVtfMe+2ES62Z8I1gwVGebKux+bQE1fF+uHD3e7taj1VzE8cvXSK6InlnhO
d9GkwdNQ5LjeAiB+fGEZvtNDd1o0TLuKiliQWszgBZtcgJGAbzFZJSaXWrN9A9FD
rnsnFpWnyPOx1SuszOYjihHGNBxVmgsph/ODQWI4OG91BP0n/1A2ZwuwQRqlqmkL
AhCfG3YeQGh/PLjLT4Y7utiSxXEKZmHDQwpwh2jZHl5/HdyOCiiz+8GfzMRbxox3
/LFvkfIVlfegiOZO4NJQ4htgULycJ2gC2OBPF24KtAiGzKx4wPrYqsTKbAwYUi7U
Wy1Nl+NouB/S0/gyum6RHPZ37d9PcX0ImQcN1GGRzKVSz4jMix9mpnuBEcPLOAZw
OUhoUHjFEEGxTaZscCWaNWFjYnlcssxfmCFURmH9HqoPP+gy2cktLGFGVdUtTrvq
g1ZEt4WWAxzQp9iOXln+MIM0cx9jVjRqHMn1r9ZRPtTfaSOsKRRHVDyW7pc+YA1Y
Uv9ki/nYhqCKxxs+z2vf20lVsm8zgbmPjbPTdMbCO/M5Suo2dbChN2SfJP3I/Gqm
VMOvzQMvvH+XH38tH72sASnHNSiJZi66IZ495b6SrA20G9V6s7V2lSRC2aLGxm+z
0kkDeG3bDLBrB1nJn7eSgkH44Ze0pG5X7Xw42pbQBs3BgcCEtfqE2aaU1hw/FnyV
ZqUN2IsXKmJHHdzC6l9Y3hpiuYofX2Y6rUzFLgTQsQj0uiQe8mdxMHLGIp5sfsAa
KWVUQ2aywwAo0np79Wf8jOyRelVsBQbwJSqTMflFJmtWZvRzXGwPuHxIBje+Ops4
w8iUv5ytdvUZ54HAZh5UCLH5wPCDGYbDUVY4oAdQH4Y6A6q+kYtOtwuin9JMGc9s
e0BYK+zgMx1R+/NCjrglu2aZkbM2mZqMhkw9YssisIM7mImJP1TFRqdO7v25GCZ+
ZtkXsf3TSDLxc5ATuyASmFGynfTsQtIbHbXKO6GsJwAf4urwy4lMFMzlfiTIG+Kw
lLBNVPiyZpLFbhdWASdMEx1spsiZIRo56tC3EqdITbELDt7AwqAgDis03jswb/zy
WRB1yx+04FK9vz4mW49i+FArvRrPovlC0Jt66kr3cjkMxaMfaxJF6juBIQA9F/5f
Pc4afW2rUlrD7tS8CXmhdAm95i0NzNdnATNJtQRagQVMdrBZLZOPt4iLak0Ezi47
AgwG3T7l5dgbgc/aN6q8XjdpjYkO/rPXL+I/m+T+YDMWteflVo2WMpx3Cq9XaH7Y
kq4fdJ5lJ15//XXwccrbTu/yf2TU0md6UDiE9T4ggfryZHWc3SZPfLCrvHBijN1Q
wQF0X6H1Tp0zv66kL3I3qRVEuRrFEI9L2RG56fSVn65SctRTFmQS9iCQkWhQo91P
Vq+GjDKLammsN6sh/A9fyAV4yiyx73fvUA3vndADc4IufwCnSE7KRrGxhJC2VJr1
gxkbi4kZ5Oa2IzurbQwRmZf2QqktZ1tC6nuefbv9RNZi1hcJIE+teWttdoI13bCd
1In5SqjLtmsw0Czmhj6dDubPH58lPk7SNt4yEKp8j2//nvJ9g9X2FmyZggTPNHbD
sAAKesaIAjCccrnGR6qV0WB42bFb7+7p9LMw4ezA7ecYmHlQvWDOZrnDPWVL1h3W
NS/F3NbN3ocaNQtfhRikxwur09U3dS0xEiidRVX6YQD0jrXBtetfUM/iSwdtGjnS
qK4FMh6Z4KTaeDX+W6lIOquq6JBCrqUDTBwATuNxpd22H2/EBnOssxxuSGcTLzsW
yQ/ONCx5a6W4sVJp0OFmLazvg54pdsE8Ip+1YJ1vG1C7lDwgwhlx9UObC78mJAy1
C/bRoZJGYwf7F4Ze3RiA5OHlBXY70+2sKeKKnNJAcEpc/AnKak2so43pB0LDyVjc
me3+caADcQ8oblAK1ANsU7QMlDj7SjFDWuqmKKTWbnG85oHAqOKLgj8Mln7MGS+b
mqGr2iOVCDiIXgTuqeIi4r/ndn0vvJ+7ub6fHZVg0TAbaBFIhOk6URV3U/6qqdtR
0BxV+PofIWTS5vUluigKGn7lCfpc9a6b0ruiklVNDOjWNftIRaN3PavZex61T1LK
/vFHHyeD8j1bCpMAVHKEEABguQhEsVCVmxyPUgmOYHGC4VJnUWxEyAdEBpNbCBOP
SJ7WCkXdMWfAAkNT0xlGnWVaGe4QUuJbwgRSLcm3UnVTDJfl79VgrgRlrbq36TYK
8HMFVHsBzl9D76cpvB8N7KFb9UsIHkbA1XV1ycXHf/PPuajNJ4fkHDBBeffTIu+n
D7JZijIFT0GfKYYy0/HXukt6UFBvmWIPvv838ZSm4CyfQhlZOiEn5psjZepSyZ6d
1xd2ECtx9YZvxpUS0Hhi5onfI6g7Xd3y51ONQhvW6kKZz+wzds672KNPOiT1qqtO
gToTEp2RuuCAlN5nrBJ0GVKGeVm9LeD6xd+sgD5MPi9mu/ecbtPyckINS2EtFZKH
wo1kO1HnoUQ6N8HizBAbUe5MSnIxXH252YhfsviddzEdQrtV8GNGABZLA3bOTOXN
z1vBcTZAzj1kV6lBEtoBJqIqO4pW6EZFfdGHSMdUNFC8r17FJQcgfWdsC77nYQPq
uixFLGD6igwC0AEwgoUxqCvJ3140R+ySzdv1BLp++5K0qYZ15LfcJO/o6fwtTNr3
RFuJJ+aWsdPmC/EQxZwdP3crF/XLM3VJCnj1da48ZzrFmtuRH5AdL+HdRuxOZPft
B6D2Ag2/6FISeOdHc6enU801qWg823eo9RRx0Ye+rDcOcqRFwO98c4qomG7Le9iu
mfCfZlSsNCAFwQ+aZWqX+sUeftxXh4hqG/RkY8Lh4gZ1NCjwxY4rBZ4+4l2lZB5w
MoXpy7eE+qA4mpIflOnhrLt0VBiwHerwCfVB9RzuSCIYNqrkSa2EX4gvsA1YUGev
UKgLMkFoK1M7PrNC9MfPUKB7+0M2QsmdSq1SbF6DyVmtm3ViTcyYhrFuTtQpwLw1
EOFOSX6rGh0c1x8wAZPsfGDXvQ1TynkuiC71x2ZMVKohYpb4RggKjFeTKmWZHdK9
MVdn7JBhR+sL9QMJpBzfZ0R1hYvZ5nOQ1sGGpyG9B4uRPSc0tFGj/WkK3cF00Rr5
48WhVD93XBK69gC4bT3CIcvPGEIVrkj0CdqqJcQM5Kg5yneMRpRQaUAMc62WkBn2
+4DvTLQi06pqIbpZ7NcMnMfmK8mp09ZwGiOwDdc/k/vIRQRtJw3IrR4a5jZAqyT0
CASutxJ8W6yGvrHHU0qAlveWoI/DPNJq4kJic5ZeYNahPLM8Za3e5UYlzWoKAuOi
zXcK7JeR4SnXy4opTqzvFiGVov0l/aPB5ST3+Ba0hooyK06+FWbDr/STIp9CwRkB
Hjn+YhcMfdAgKWtUoxfQkcIimMp40SEl/vdeSxI232Ora5LS3MDrqS8URwx8ElQx
c7MqNz+Wyf+D4n9s5QgTGXVJWbgr+wKSXFQoV13YddkRMpU5tC1EuuqGNy5edpLn
2gDyp8q+SvhUUlAWR4RD/W4qZWGLIOC/F6FIvZzA5NjIJc4nM8vFEgL8ojjsq/eo
ibGNokCi//pLb7xnaD/e8BiX315tYNkTZN5k3MGlYIo9ha0EFhcMa3Bh2HTdJu0w
EsKMwsT7KnKBmVlGLS8XA6KS/5+0CYqdmh0fZMyXaDP+xyFFiaqsypqBN0RxSo/k
QJUXEYWtoi1X7PhorgcEOJVPnJLbFdKYkFQzBsKrH2sqytuoTkhTC4AQs9QdbFD0
bcHk78KUkYIwGmH9O0dUAq1KZ1Sc9TzY2wJPzVmox5xQ43mrJa/8FwQ406H38/BS
mKDRrOUs0ZN5RtKAp/UufA6Bc51f6GCzIJW82e+K2eQtMeWVY1wR52t4bp+h4nsP
+qQE4SXm3FBoU53sF6WGNwtdj2r1U20df21vJmfucQYRhVyv+MjrSjvKTIvXxVnM
xfaLiGPqeHO3Q4PVJDwCd2n7867AtseDuUMINyumvPtUBdLMwmzrxEhOCs9b7g/1
AvUfowd4Shw6pmt+PFHBMZtGwHkxX57HwkWi4gACt1QyJtOdTjKtLAjs83kC7ELA
WTAFcJHWmE9xhOPiK8t1xZ9nQmrzu+7kqHPYDHTD+ftVA8X0oqEmQyiQ81ZTzN5K
EWyfWCa6F0CQQCF5GnnbhTWxnqhxGh+EkaiPb1h5IOO9KTVXF9M9KYpjC9Q5wphz
tXdXzX/gnMYhARngizFNVGe7drv1np68QxG5a2oj4AYaxL7i4tBVxNGKiOHMm13g
rgLFDoIWOeyLJc/oRCBHd/2voqIuH21608ZH4BKYS1i8dqWRxGXsM2NpJYJ8cX0o
IJSpaL2RlmD0nfnxv8rzdFsB+BsNIDX47k5/XmrT6C6xkNaIl4iqcSiOIAjSwnUp
I9EPn8DPVHFiwtQqVSUnnq1RVfFONkJGiXIPQGouy4nYtlxiT4AGaTRHXwGHc5Uk
D8czNr3BHiFFBs6pJCJ2IAqk20lqmkz5KtNOooCVLsyER9vvZR81DUyHTMtWQXWf
FLuxhOFNmBk45A5stLFLGlbVNGwDsyPC1/FUF2PsJOm32h6lGntZJGI+p3WqVI3/
Ku39Rjvv1pnpzbXC1t0nfehoMGjvitBEQTNz5G56zkuRJbjNAU7ayJzqjakE89ni
Hqr6kJiSUgv5bsVEL6yOaPYb6Sc3ItlVazIqxL77FLTsvahtgswMoHkRtQQBthFv
gqY6xJ+hGKFhCDAv2OT0mcONcPhw8d4L10wXgDX/Ya6G2Dh6888qeP94faiZX7nR
GSdY54F2kuUYefKInsaq/Fomb0mAGraeCAoXeYUvvRaVxiKpclR4zctjFwipddxX
ZeUiVbphrM85D1tKVUt2jcoG1TTvV8BNkNlMCYJqvBc3RCsi3mIcatMOl8wYDIa0
Abpy24LDfnQQADhmDoKA0tawNNdQhAnbyJlGQmcvT+ZRjqI7fDabRlKcUuHo60VF
ROzdVvr97SDQuARXLebFS/8l0T2Gtpcco7W2sSa4Gyp+6fnL374HfxXm7FhnBDRa
cy3JvuD/AllYDjz3axp0GIOdnMCxqET6wfvDTYWHWblo4fLODbgNOYvseAHx+0lR
k0e1hCIn7JXUbOY/jZuMghwj50Tc9NlQVAsF9X9VKOkOXB2405FEnaNuJCwIJMVZ
TIFGfHBH0GcoqRnxUqYpWc4UbCp3j+lljYmLwY+seShmafyMDzF4hjpVvS2e9f9k

--pragma protect end_data_block
--pragma protect digest_block
Re5rw7Hc9iMJCHtteCnPYXNHwsM=
--pragma protect end_digest_block
--pragma protect end_protected
