-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
v8rP5O3fQyFzyuEpXuaiLiizV7HwPJ5wIXi8NaPwbI5gfd19xF1G9syg5TEbDtta
pujSap5LxoIvx2yv8+weaJccDL1VojC7wYbSGEk4+/q68xjOPoi4NBAy08lpL8xu
5G46TbkoLZXFtxZrLhVW8RWSkemLOAN0BL/iv6nSZW9UNHCqTcdTJQ==
--pragma protect end_key_block
--pragma protect digest_block
jXCFyMXJZ5wo3Bzv9epxJmq8HGs=
--pragma protect end_digest_block
--pragma protect data_block
DAqYFSy1VbOCAZg9YAa8F3m7y23Ts4y3FugMPNLiApAHMOS5KvVekPzQXdxcPdfi
mtgk5gX5PBA79UuV545FUVLelkd/sJkcfXAhZTEUlqoHg4lFZ8aPUfJOnFZy4D/s
9tjEoX3nWNZ8gioavxgErBPQYXPkYU0DF08K6UmhBJnpz9ZA7WiaRfoZtObeecI/
Htm4SQLEBKkt0s3DW8GNFGwBzaapS7S9Xm3xN6yfqgkhO0BSWvYVuJNAQBJJkYQe
SLjzYnj2IJJi8dz56r200wDyluWVjd6t0SKVawbiUoBWXt7uOidsjNQtiNaQt8ZF
plTmu4mAg6YevfxdcGF9XoGM/Sl6YzjZWVKkPRrpWrygIlMM1qVzubm++wGOZVgB
6rMPBHYXum525/3fPLac186z//atzHwGQqYl9854NWapqpXiXIn15VvS/b6/2Vwy
44JLVpERcr2ysnqNBrLX68hEPoDJWnLR2VRXCpRl6bNRNj7/UAxQA3TKdyAoX/gX
KzYNBh51xeKBEd902AnP4/P2pOghoKlag93mq8aEZxNgAJKlpxCR4ssbAe49yGKj
28+KoDZomR7wsOZieeJF8LXwBQz8I3aMqi3CpzamAY3XRDDPq//jPGBMjmIXrniL
/ee4o+9uyHOuxZn2vglZ1i+kBzJwyFqkjxsoy5sW4oDl26iJq6YHclzPBeDMUKYk
BugZyaCQwI4mPspooExG7nQN4A5EsWrdIxx4bPRjHVKlYOsYw/HtZ3q6T+ObrosA
5NrY1rB2JWV23uIrwetwrvY+GCNXa+Fh9YjTIJ4mFotYg2Cy4SihI1Ztv32acB3x
Qd9hiJSW3JDpNsenH9+V737SgdZS4G0amJaMyHn3gePbBAZF16vISypqusYeOkwF
tJa8AAEbYCVqp1hM9x/hO1Uj7GJlrD+1csQEsf7awmgwt2kWXw2mN04RCC6ccx5U
JCoUmb59rCm4RXnDroewEPb/LJUDOajCDORFDfnCWeWMyMxnnnR1WCgFuVEFAXnG
mNjKSXJs9ohCsaon8dzXI+NS1wFJhqG4UT1iL8CYuzZ1JUGEWwaVIRTPX5qu/GsC
EUnBBAw/nKv14vNosUuj3z5ysnCwIu5pj8AKqxLsTZoSwhzIIo6n7RSNB+gZdNxT
JRWyqArvnm09CHFChTerg98Yo4WN017d7GCyl9lqomkRiJnRk4DBl/ivPYOkOqCt
QOHqkzLor60n8+jHzPgSyh1wVA1pLQcLnUy962EXnKOezCYdhSh3klnMZb4DXRtA
VgfOKPMZ6o6HVJ21KBisTzh17h0UNiGIXE4WyXdvGQmuzaj/9Bvn81aVqTYusWaT
fvkd7auPHUMnm+SiwqZcAompwz7qjEEmYDd+1VJpe7xmilrUoFKEqS5T36oV28V3
2LInVZ17Pry4n3CXfeSZbP8uO9ReSsSimQhipWh7+8TQpPNegjj0phAp4BlyWOfG
lg2l6BKeOBb2k+jdCSPl2LfpionpvpL5UmhyPMPiffGNo7iljqGFBy3P+wzob6ts
ruJus+0KCrD0ohhsJDPvEDBRBcbspWwfdVZnocssUqY7lJocEOJnvTdVtm31Pyn0
reA292yRZ4LP0LUWyOAppyVQdPqDgNlDdmTkthnZB3EYggOdATugN8iUaAE3ZM5H
AY++yKsSj4pUcyOVwcc8hAAlup/PcuISuVxjglQIcWJj6sg3z0Zn8sioDn6Z6HQm
DTQzBl9KK8RIl985klq217sIqvbO1PWB58uY1XwXged6YtYkO2tqVnEsBv7p/+G6
xlcptLtkTSzsNxEFRy8Cog3als2Tjd34YEfEsX5vp/AuHxUFgN3/QLKC8wH+5R2m
oVHHhak0W3YgtHYB2h9t+A5awqdL546eIK/2SFd/5ChA7xWKlsyb3xK3t14BhSQe
D5lTTNsGwqhQKwiaQFld8HmxknJTi4iAr7/TM1g1jilHv3AuPWHnBGVC31nxPdxZ
cGSg8PZDA6bbkWCfzw2BjAhHFIsZAl5FEsuQqy1W+dqLH/D7gzbCzJhQckO7caDC
W7ImYQYHAWd4kV+CRdfvgajQ4SM1pliPLpF5GfUo1udwYqZqV5rtKLrm/Jom3CPk
CgshhHEF21FNQtgNkLr5k+szhxxvoetxMA16gQ8N5d0EZsFDAAvPku0xt6wNL4ln
6ApeNyjSu14SkDjLNRoSvdU6H9tDQGXyMgLrAoiwkuyES5Ja14K0jXrjyMMfZ3Su
wWbtTCTLzsrgMaldDFBOL7InoycTWyu38/xa6BvAy5JFJNA2lMI1URBEM8a0gtKC
S7dS8EoDfoQ7KUXQL6d7yxXoa7+pmnR7zSgx1HKWx/cflBq2PJTqbKpkhvJ1d20D
X1zT3cOpluBOQvqJQpevgT9CGk3E8awi4xfaiG64Hq7BOVmAsMIjSIBapSsmRznv
fF27OsvZ3h5jWcdeAv/govMw6OWBvxbsZnBMb5yTxW/mdakbRCTOCa36z/6WA5Nn

--pragma protect end_data_block
--pragma protect digest_block
lsICeESYHdRTiVhpeWlTS5AiZcc=
--pragma protect end_digest_block
--pragma protect end_protected
