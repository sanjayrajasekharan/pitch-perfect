-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0uZ3lJRi/rB+GWK4dJrTMrVIexLASq9NnuyKlNBf3P2MRGqh014hObHF5LxTbb3lkNNWZ2aNoIQL
i/JmNoWG2DgPYPBaHc77Mhka7TC6nHWmMqQyaSddlhwz8yBMMfhnRp6aYxekh5Ia9cvEfkPfDIgV
9AVF0D4bfO6f9KH5RCIwH8JcNtFQ95Zlz6jfjuaOQwqw2WZIYhWWb2SOuPRnC1Z1SzKrVloeAyGR
H90NlqhOEynxkn8tCgQm90h7F/SS+fRnGFzM3WRIMwUgzg6KHFNscE14yNW2GOmcrYWzblY0EX/S
rs292mGmiacM4uVd5Zo8WviKUN7tjF9LdkUQjQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8032)
`protect data_block
6wbZZtP5Wki1jskYtaFCjvlKoPKYSy+dc1OvJ2jahDxLz8IiHZBe8WzE69V2RiChoSLFczEuoG8B
v4tWOXzGRXtPjmc4qtKQWLUnn8SIKeHzOjeNvH9KE4c6qmaXU4Dm4TuhCV0gLN2BzX6RbUPOlBib
JYZ89edRx8tY/jvS//PgIzWcHQnhq6NKz7MCAFBMpucxO+1pkcQ/NovRQHnlq1R8WZYGCHOce4AT
LCTRHkDOp85wvv+CkfaqkKvlbzKmT4essEIzsN51pe7meJu9TKvzyV2gFZGQE9RAn+A5xgs2O/Um
2vKl6yxk86s8TZSh+RC82e+kRI9xM2Y1aU95p9TdpKh+H9OKeJuGlYnZzZttDDGXSJmx3vT/Subp
Ib65qtQZaeZ5JGeitXY5qsueTD3ZL50JwTzsieLaoZMaDdjbEPG7pZWsW/HNGfWgH2u+K2Hf6MaW
qqcbaeWi4nauxkQRnfTCyk8omYQ6bleuEtDQE0b3QH95NzzNvnz5DRN6wsPp+KclWA2rsogebHAg
POmwiVKHvKkv1gNw9WHmhdPMKt7yQJXI43ADjhDu73Bx0Ky/OgLE4lu/LE08Tis8+TU2vnV06/Ph
tTa3St0Fu2Do0Oc3FPQC6ylB7Nv1CkfMlsnlTrWaYo4Yi4Cn1ogAOfdrKIxGz2VOF6UbskLuafKp
9rCU245bqUFL9OatOt5Ks2qLpDGyl/84E5OTyqhfbSPNYfP/9adr1fGB9ORHuN2+GuqZRnLWoJNk
LQ540oIcy+rlxqp2rwgp+/+obJdJVqQ4cqKegfYsleh3G6sabnMJPNM4wu39kO52qB3fZd/NySJO
XLAxAw3EQWho5Gdi4V3Q8zrNLFBVSFmYuCAJZwCpuPxMJPYWYw9iJ77tAa95YloVL5CbjMy52Lui
D1KLSrqf4EvQ704HzrG5qghrHiwufup4rqLKDYt2jgBnsP6F9LaZkIl2Z6N1OMzjfE8aWIpSbdQj
WNf6TTJ7931tCsn6+x0FjzFV5z4ewijw+X0xPBTXggIglxrdsaU6tvUkZqSekR50IRuE6CkCT/WK
fygEBdC9C1hhC3kfh1DThwthQwinF0CN0dVQ+e3Wq/6G6ca9SzmBzOLqKTti/HjATrHLNvNuIX6P
L7kNGWTTz+ZmCCYE+uRaEu42zeLiyTMhE0uTkq+IJpoZai5Ux+GznEYrnPe/PlzCRVJ+E0Bjyo2e
irwD03Ji8KRFB8IPH1i9sxshdO9seu3G5P2atdd7xivRnf7hRr5FN+qQXYtwechBDapXZ2jCqND7
g+IjQHJ4bq59pNYkPMluEeEjvRGCekvkMDbZ7d6ylnzzLeVvuwkGoNGCscO7r0pqUiTW5UCwTGdJ
feaU50KjnZsbYOAk2SY5KQgAriMGT0oT6GwMo3bZmGqrenb1fvodcg2iGy04Nviqp7gWoGeD8OU9
eKfB6xt0kD4K/EaH4dEbuapa9y7MIa7BNtdXzWKFfccPn98AIEM7WOJsd7etQzxkdDcI382WnE1p
mQi6TY5haklf5tPSI5yWioxLv3UpS67pM2at5RVDZ1HiAKYgRiSpezTMiax1GmjekZQ7U9bKkkrt
1Gxjr54bMWfPBGsU89Oyxr3ilqtcw0Z4uXaftkx5uTQSoVKrhDqFuAhOcqrU5HTWVIPM+5PjJ11Q
GlfiWE/hO10/jZVxHqOKIJkMQgre+zHRpuATykj88zkKXvc3VBnZBN2ofr1rRUBzAGwASV6dJJbh
V4RijdjzKH1xZel/vTp71jmjCSse8a4HTSgoyrJwqeXOVV8hnUE5CBcQ50DfOy2gvr0bzIyQW89a
yoKZ37RWKo3QmnwHhtzxb/nEwqKfgPm/UdCBvDtNbWvDfQLshHHBgWDdnvM7uaeWGMKHSeSLc8k1
ci+y3G+xht+ssV4wyeU2q5JDs+4S+Td2d+aEWGRp+FjJJuqbJErLMAjmY5sjshXzlXe7gcW6MwtE
Mf7wfTVALA0suiUK6Srm1WErThsdFmdefmZvITTXq1gOct05+aik+VbbMX68NowHH4mF9EBIEda5
sT9utmYMdQh+n6goXD27+aB6uROhDL1D2+0Lwq9dYZuK7tNhK7m8vwrm2uN47p5i6GFUzhqASzCz
kEd/GX4moo/ZqqbszLoYDGnMNkI92j1AY/Ee7bIzazDxZP2+M1lqC7ukpZW81f3sSoLgN7XfE+PW
zrxZUmmS0dZ2ZrhqzkSIv2axuSr0uWDJp0o6jLCBQfXTVDdO/plowocl9d6tXHJnYLfE3X+7oPtL
FatlUvcZ2+lnbOUJYIwlxnijJQK21g6hJKVP0Y361R4yInWXjwBYC3hbEz9g3bXQb7p/xJxwtM5n
GVRw1Fa8OeRBS5f9zPEkgSuPuJFXBAoBUaA9gc8vtLrlWZw9Vw7JtpiWgrpXwKs9PFa4sB4QPybk
hcsxFXIgb/0lMr/JTec8q1kJVqXbYQCdJnA793FNAuYNOiWvYjfkRNcv3NKdvPpM3GQrUVG7S1oI
MWqaI/1LCx/8Y/JiEZDddzwDcJuopWBsCj/34tNFHPI/4kpkEWwmgkscCLjJj0Tr7rUnH2oh0Qj+
2UbjZ/MKJIRMxUUfhw1XTes6m7hv7pc6vbDgq3aUoBGdPcdeRNOOwXd+kZwkvhxctJ6x1xSbKMPa
mf4FU3oqSEbtF773cgrFy0CfaDtaYKgB22R2UacU208yN5FQTKgJ+Xs8Jx5I4gsCfsHXNPLdJ73A
q2V5/uCLiB9X2FUJEDTQrZ0n/CP7t+B+BsElTDExIYxsDDYu6cCgzFIwb9QAXI2v/tPlnzcePe/Y
mw4WzCc+RbGvtgxbgoQWZiYAyVx3n2YDvyAcgCaX3bjvGiQhQnEyRorWHfcwB9IQS9Epd3QRpRQQ
qiKmJ8y4IYolSzopIX0YqjbdLqLJNMQnt0q85L5a2VyTxPxknMRSBMmQ6Do2rhhRaYYLbYtd5Y3y
3wrDZyxccxRaPZbE3/X5LaJYwTafQ+0t+4/QBcK4VyJL5Wu10qWEl3hFtuFAcG/KQD5G+tSLUVjx
Hhsd3po/pw/QWg/EDAbAIyj9PyBnmj/OLHSRXZb3vn3W2x+A18kvW98kVdoHf3JtxncoNdPqiW13
VI5fZeUYNzY+lDSyXZo+4/cJkBkMk+BMpX5s0Vj7L6XELdLMfvhAuCnq57sf9Y/Ri1Y/GNDPyVJj
3Huz/a8UAgelUkKNk33asn/KW8/z430t0yoa4L4N/+sdgW4IbjKa8yEr00jqoDbQSDlDWQWtoii5
TlO08irIKZf7lu2IgyUi8aVUyO+gn13RQHoVumwjTMranvhFLvYtLA93PQQAE9rwMsMiDyiMCYNm
91Kdq/iTAiArw4IcGsRXU1nYWF3R52ljvrdah2lLmTmqGtMAxSwVM9qEVNbWdwZuNq0+3rq9iGV/
Y0UgusXgTFy1Hjycs/Tfj5YI35mm26F7S3TS6FI8+Wqn+8BtW/dEIAuwwahT3g9oRg9KVrtFRAPp
mXtznEctP1uwl23QFtRhxuLFrSvnTKjEunZoF9aPkb72cFKkIYZb9iQQasuD5vF2a/6pvjfOtU8U
4pwnO1F+qBgnkxr1E4OT/rslHDoEYrYQ9FzSO8MVm/992a60YJDIb+QAEqAgSQ+aQTAA/dmhv10V
hcr3U0vKxg6kt6gbaMm66rvUAgsqX4LeLf5vnIZBjWWX2UnpwGzKgRqPA4ZGz9YQM9ZGCiFCzzHm
QTERMXyDf1kB0FurrNDpSi87ROEZgdSS7s9M1tbMuzXeirNQ0ybU9ziiMPg+LSU5y6u/g+z3suio
1xcr9cZZ8196SZd5YjntM0YoHsbhKRWrHPCMF8+uJ5SahEqf7/VZ72NbcS3f7BBZjCBExfa7Xctf
X2GY9oVfdvGKXOUIK/9TlbEQUu2GhKZXOS8V+M6TVwGh1/wSg7A/c/T387dYhQv4I1+Up9/4OFst
Vyu+1WEb/DFs7/EItWdy1yRvdOmm8YT6oKo7S6ye/zgBVyxryPbboLNK/4dJAddyMjXv307of7Md
KB9x1WJ0CjFrRwEnu0rXZiqVMxtmcCuV4Kd3yB9IwvwMIpU/BgB6awOd+2wRsxmoxWeprbYz8PpC
1NwYpIlrtraOBGXGZTsIdipTJ/+/DZh/fEdF+Z5sh8buSvGKwjw/xUFkhPpKKjjFTgFUX7aDN+eT
wyw1yocN4O5KJd6xERXHYf2D1Vz654t+tFj8TlEjA4dfW+NRz1UDh/v+lM0XAcagXLVGmIGh06Fa
1ApaB9vcqWqlpl6D+FcsuaEu0iHBXJKKX7E0XVbyUBLTkB6c5wOIpz740mPF6UgRXFIPsM86ARs9
xNd8e43j9WjY4lqz0ASxcX7Fr4FWV+WX7P7yuYkOGUoxKfy8xBeh077G9Z176z8/sc9sl6W8WsIO
XLPxW7TcD3j3//Mc7QBJmCxPHCZC8rK4bB/CHOg71Yp8V10fZZopQSUwTyDQqkg+aWEV6UDMpC0y
WCVNJYG/p8taSYrdmFVUOgVDDJ6Fl8YS/4FqWV78XpULCo9DpQy5TwUrgcW/eXSMPxxiMB2yPjEO
515TW8Sxy3VbTwgt7JwpG9Qm7gr2cHqCqQcm7iR/QE4pe83WBILXuff9g/xcWxgCOi5zFrWh065D
GcG/MDeU74ris7N5hJcVoBxqKT+8augoqHpT6wxOAsHlFkhrOMmB9Z6xGWrN6iaMr8YU3VXbddMM
QAFPDF5eiuh3YEio2nM6lMSmT6SbqtY7VSkm9pcxpWS2kE52wUN5XlDn+vE93s8H3D/jkbsh1CZQ
Ak5bKkgktbYrgcyB5T2q6jNf/cE8y11cVllmkWVwGqe+nI3PejMVK12qiC1tX0bv9sVtGHel7/dw
nCftFUovfwmUZY0GLN9l9tU+U+DLmrqAgWUGv1hu+9mMf+72Nshh3OO7REa38yPWbTzekuKPD/Yj
uiH7L4OqQ2/S1Lc1JgNE3aAqWKDxWD1zoF5p2kxjFUMG/2jfQfz3F6ztXx0VTaz6dWkBZf6Ua2O6
YyzG/8YG/X090776+mLcQVK9Q9qqlXZUo97U4JDiez0KUJrxEUpWJS7t/4nQft9BK7jDrbRBqTBw
A+tJL2OPNO53465dUbhQxyonoq37j7ztTd779vUmo2Diny7INqUIJvklaTyNIFep86w2RlpVmauO
wv8jUhMPwTK4WhYc1vdce8AVErsTWkuh0ihYY3q4P0fX1LGmZimUgngTgjukyeJG+vl3/e2NALqv
boGtYLJDwj0Cd/TAt/DcsDckuFiU2rMbP7B6FodnNFP5DNaHvStSmnTWzoHKT2/QYcn+j90gNKim
Fi3ffyYclZvLRe0w6868BhLcA9ncKYh7/+2633shP15AF16VCOnaI/RHENGlDS8eyjD7yQQm92PS
qbHGmfR5Rg9s/wbcn72N4AgnOYrP44LOCgNaKr5X8Y/hUhelnmeh25iBZmJbH4TQi7//pjox6+wc
6ZDZrLCGY7N2K+bfyEQ5CYgeKThUhQ8g8jS0XZW9HIh5L99IBmXKSbdJwtR8+w3Qmm70NBfsbV86
RAXLSAQ7z2L9F7Z5DqxkA5SC8n93gO+MCn5RBPjKPpdui2LTTWTBDw08SEKwmzh5YT4EmPLYgbic
+cieQNtxpWzKccehvK7NZkBcMOLugpPJzJ+PrtRfNi4zbJsg1qXSd0vR3aQMFnKMVki6KbxTfRRa
QdfOD5dqalWwBrla7eF14RHGxgkBD71g78nJUwfa6Mji7Bc4sVVpz6ZnPrPXLXY2/mEEuCqc49JI
AgGmHrbQaY0BDKY8lM9RAhrfakINAjsDpCpQaEHCLwQZISiLoFKDVRfZ/4U+MJYczAR23EEdY3Md
Se/N8RXxiKAtXUrHmig0RJbnGU30iv3brMMCwAxexY6MiPz+PSDoZYi6ZJ78TquuY5FdVrTRF1hR
nQWzDK0swb4Mf5HRupl3ZM919ipKy34aU9n4k9Gu5E8kHkCjrTx8TKlHGXiIIr93DarPWD5UMvK/
s22Jy8MdYlMVbhOYJsk8hENrvn8YQGTVpqPMh9gz/oNjStqOb4Y/CIWhYYxzEYCnVIihtbWKRwnp
j8tu3muenIXKAOML2fIQBF0Q/iJ2syOTFvz/FNl+l3urEFYL+exR4A6izbghkBehFMYIcDGlJHqp
t8ShC28HpWTymBn0Ck/UToLDdgJHn+JgkdRIArpC3c2UNg+SneWz2dtczA8OcDkgDkOZmBE4y5AV
Qhz9rkI2Dow8cx0fPDAFkh3MJq4SG8XPjQi7ohIYMpLSktYScJcXqWAx2NYSI7UUeDM4m9GF7lZC
1Hf/hRWySm35xh8LIC8hZDIExGB8IZAp+nGSW8lmWntNKCjaL7K6GHlx7OaR649/IVU7FFDSKPUZ
6Zp3Yx5l67cDOak9fAVQJue7hFy25/w7Bct12VEXW5kjIXPW14EblPz/cFPjXtDCjXWW9NC7P01r
n7vzj/q3+BJ3lnNMC+/7l94EuzZz4pK4BU3CWDBYyol6s7nD0HpjcF9NJI/nlnU5RPkH4rtx5bMM
qYPe85rhupoz1VG8CAjjrMroM+bh+1M/IzOY32gRP5LSPkFUU9ElVHTwZkpNgqXS22vrqA9pAG/E
6chR9hgvv02ouLryL4wCvv1k6juMXPsIwfZqynLugT1NFChM+dlzkdrK0IemNsdoRzRvOJptRupJ
yGHDhMxRB0U3xrf0oucYtNXPCmnz1+GnTG2+vB80y1EDzyrYmc5dMNAGPHNCABBRn0X8hMEhRA4w
AxcXjF9Z/3auxCN/q+ZOIPSNlR7pNZ8Pok2b53kTCrjohF0Fmzg3BY54Sj+1eKKq7e33o0UvxdV5
+2gkcL7BtXqmGwAIfu7LXsBePnGCfCycUQy3CdJIAwLdT8QV/qF7iq/lSeM/x2fXgO39ZnFQri6Q
sr0z8K0/fqRu403FjeU331fIYnH/U9fZraL5fZ1nc9LH5r8I2cIt49oQnEVH6XTD0k3Z43VohQnN
R0wb/PJQXc6f4w67BPC3YOX8s+F2DLuIRieYz/X032k9avXR/H+dtcE39Tec4AO/M9SNNYwo1hVb
tDBDBs6+oh1JwOLCG3/sm299sIOLE/keDPLaYUCjnPTysb4iC0tgwCO0B5qSInUY+5XmngIwaIhT
3Rk1LwMe0uVWrR3O6xBwbGdJ9vwXm4IguMCBHsw5OMrLigbb6WtYqnVTockVot8qOKtl6NTSTvaV
ut8/ReFDXZFJJ3OvLYLGURODxkmsLrMq0o5th2Txsy9AuQQlqwlBMEHeDAkCGD0mUYnl7nxsNj3D
Cd0E5pXrlN1K8BHHnALwzieLI0tpOAvSdMrkgWxLQ2siPY5p4Lf33lelfVvEHMfl1819kyzXbWlC
zI1Y1F1OkJUXInBiiKXcCMl9OeYJnD7p1bDN86ibIj/uemHmFIQ6iAWjEUtfzG6LInAksvc4IWYT
JyLh/gKv4/SFphkkc6oobVtPrPUVd2jRuK/k3twzI6VVtJJovtwLP1HrozHHYv0aaxO4RyTTceBw
8hPxB1rv+B0F8pw4INREiziLEjAAZuIw3v6ZGEanQzHC88xKUyis2IbPWsBRtujK/LHJgiXmZC3P
WHyfT59witf2QFpEF0VWBUqFkkJD1DXxkoOtZZzd2oAYpTBppV45act29wi3n39EZe4TehLS6cPL
BGks0oAL7xE4n69wPWnZl9WA2TGnxmxQUYYoYCC2c+P5+RVFG30zwdgrx2CbxYDsrWnY2tohGzyV
WK64KYw61UKFlMRobyWv0dmVr3lU/UdUeXYnYz8qTO0DTUwR8kPYD6MG/rF2GmGQMUhi0U8dzdwk
WoHc5PYBHSbDTjgemm4439ScipXScyxVW2JSmo469++E4xDmmPpGgoJoesYs8ZCpB75KzkKitMvi
3I8iGJK511H2BtTzdZNvnpMw735d3zZ6u7qngPpwaKhw/VlzNdRb55NglEzBvvcr8mo/N05R+IJ4
aEYZCKnrwnnhV7ddwzlC7m6fszdKUnbqHwFJjLD9WT6f9LYzNNbK9Jhjh3kSPqHvA+g/XtUzhjA6
C6nqJZEMpLyg6Qos7Jrbfv7D40xeZjfobjzMSMIoNy90OzcjgSYep3L3bpktHLst0yoV6r2Qt+Zx
tmKBzXFe49Ze5UG61WUMlnRUYsNPGmUcPXhm21B3STevXNU3xP8WDnSkfcT9XaznlIkmkDutZQhh
Qy3QX/HJ5Rf4MqS4+0f3dY02m8c7jj0Ekb/KAPrZ/HZdXj6RlcISmdf84Xuk/tNypmbQcvsQprqj
gUQuVIC7BuPBQ4oGpB4SUW5CF6VhJ2w5vWdmKJK6fNntIzcLLCIyaMs2Ky7RvBfWnJtTefh1CUzY
CG4/jhMJwk6KuX9E1FdnyCWfVZGi823DxB5sXiHktTLoK+IyUrryHWgOuimEZAioRGrBrnjReG0g
GNGhhAbVFo3IDAYjJWkb0+KXO6OZXOZ/EwMUEf0mYjlzRaMXa0epsyLhdAB7zaf9YnXwefslwCDX
tHKYqH7R7Md8oXZ4oix+5eLv/3Qxbv2d7418v9T1egVwP8ka1IhxwHDVm5jLkjA64eRck4nFygH8
eQTLgaeJnewBKHjLcKNiX7bqbF0euT0W5RCpFVrG/XoHLnRxeGEVvt0MU/lyhQKVNM3ds1fPbSUN
Zi3noz6i2HawNqGvPLP5jEZL7W1hOYakJAS4gAP3GXbu6cf9U39TUq2nssDtgPDQzEqW43WyCbh6
EOtGGkWh90wbSv6fU6OZV1PEixr2D/CNo2qCF7TTlX9CJEpibq69TofTUZauuAfRxwivVVvG71je
yHrzUzP7JaqOGFc4ldeDKsa/bdadczlppkrqPJ7YpSuM0Nlcyt7h5kSzZajqWsri0h1wsXce/Chu
ye7bPRGdxeoWRNc9RqKXJG+sXmqPwkP0TW8H2OikRKrdUcliE8l/TtGv4oFpg0KzC8tMXL1agXjO
PIW+HC6jCvevnqqSuJ1o3FAC0mtRKTjGGyH39V143uzwGNhH7BFM9Me2qVvTSODaR1PuYD+AER9k
ufMBpWvbSvsJ5kUB5KlXWn2GNOY+hugCPRh45b0c1OIR0PcIEOOpDaCPKsq1zvru7TXUKo1Z2U/t
BnNQ0EKT9PFCO86l/H5BN4GILbmdBn8UCvVEFYIMowh+qyXkqVS6JeME8BJ91vtlPkpUd95K8wJU
XRb0/QKVRxaGVNl+iHk7ooYVx/2lFW4NN28Jm9zphWXFUDjesJ9t20z0RJzt+IWeqK3uEgxijZlR
YOg8fZnS4QPKw6PP4JzyPZmH2TrQ/98kxpB5N3C23g/q+WsvatxjElxUm6ZmL42W/ShELihb93uo
B6Tc/c5swTePWVaykv+jM4pm/DHYJOrAwJP+NB5WBiNNwVjn/jHEF16vyQcpz8tif0ifDT7nHd0g
Wz0Peotr6Brt4G0avZOHWYLchH8MN+E0vq7+bVKSf33dGf9DX3/n1a+Hrh5AYpSuUpG9tQxV7EFR
v55ktHsiCFQKnSEkUDqxa0O2awDbSfE9PEg9pq+XMzvDLsyw4oQTPXMn9CRmxm0cjY3QlzIQkCtQ
J6E6ArlG2XFTqgQx9pRK7J593dKvH0cAAfDXZhfWndbEeZidDvTklOoeHbnWVbzo8fSggLMWY2oB
F+KL1CXf4PtFRFwcj51JiIBACnvuX5onm8te65nsmHoQawrAUsxOiKaOShtX/sfgqWsD+GpM6XIt
cKFEgItY0Y1kDuBF0QXqZB3F/PnlJ0QqwXUGLbxqCRWyqqfMj8xqffVEvwLOnE69MZkjOqeRMXF9
4XqiNcms4lcc2pwuAvCuzSYYbFSdwzwRPbTMgckMdB2HQgbwncYYEJlnJqpy/vtdab6qq4CGAQRi
dvv74VxXfqQqLmzE0PYt9T93Y05ooKmmFhv29CQKzOss5uWTba7e1XuJgxVw7LSO2k35jMYne/G8
rAQxYHrlB9AG4EDUgg5WQ2DfGzJcZcufXd2DNOf323KVFBoQYeiGFNAWSPKfu1KuMKmp5nZAeMWu
C/7j5xLAPX/pwH40Lh7+Lqgc84mP4jbikJ0RasvsI1L4s0YQGdjxZXMdAGiLxZ9SUep+rXWyx14B
+EFfH5n60Oe60LU0VNZL9ppNx0DOY3D1pp3jRqZYqAFomLncQcSpVMUhhV5t9pStAgq7bjnwGvpx
+02qo1hjQZ9odY+o94ypLJga1tqo6LWip4Gx3zAbaSLIirM/z0Qnug2eveZig6ntZODQPVs5bITV
UESJtqVxUdTqgcGZVkT0e/lN/NJpYuiK+RzGiX7in+uDCM5WMfav66yx/2Y2hkJnLP101XGaSu8K
YAT3nS3We25Ve2gKeYR8BQNPeB9GuPgh7mi0GPOM6HrkuDyjEYirE0KM+Ut/YpKal+9s0JPDp2es
tmrl8Oy7SpZziKwDVatAdgvEEciJUgaMQeNEFW/v6Uyvt4mk2pXSTIuqv4fp84tFrrl397xt74qP
YstAf3aVFmhWV02bghiL0a52K91nAS1ZxN1ZvLb3sK/lZ0ON87Eu/m4KT4sfYc2mqyy7dxpH/y+k
NXdH912hh1Q6HlrEGEsJUMspfvpmmlHEg85Rnp5UopeuKPrDZOKxmOcAtBdlmShksFmbZ0P7FCtN
I3VXGW7TJUSZ7GLwNiTu6Lg0J9FczHH7bL4IjZOHFJSeTq82QqpDDyBIr/tvAcMoZBjX7A==
`protect end_protected
