-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
T3lj5XMBcNEPrRXQruz5FVJZwlwZv6lH8UCVVGEtvlicwrzSC7BY04PS6QRWReKZcwsavypZFpm9
ZokH8Edl1omXak2wfDueBmkk8JZVIhlUfBn+WMUzZubKIX9GZJGjQZ7ZLpRMIBj03w92uDMmx53q
Y8ChHR0G4lAbgHx+v2QTfnlyyvVJME243Bbdt2I4Pql12vfgnScPtpQ3d10faSHNQqc4hZDh9ceE
gUdSuDFIhV7QxKUMDtYGB+EKRLxU8ynoNJjTuuFfYokJrOSPOxSQ+pNtlG1kF04EqKHwKW3rwJ1p
MMoKaqqe32yQOkuFCJwpu66lQnXEWrmdgC2Neg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12096)
`protect data_block
7556Jbtx9+B2p67c5etDYoJrqcwCKkoFfx9TSbTm9Lx4pT/PdGqaqzpWgGTbYPs+vAv6qLlNqjq6
le8TnlbYazjBpbSmfiwkfY1kCaOBI8jDWeawktR9lHSb4hYPNnVdGwdUsT0WkdAewiP8zyl217nz
iIA4DPC8sjN1iYIrQ/p26Hi4dNUPaUKB2YV3gnUQGORPni6+gVXKyQSx5dWpKbXtJhiKc/YsKD3s
fI6IQt/RdzKw9Npyp/LgbvXUQXeYR6EwZDAok2x5HOHY+br5yJ+iXOfsXWPsPlN2ye7PQCYTwWmb
QDY6j1VfM49zm8sLOFF/OhnCump+yKaWbxzHSOqSNOeJjykCHrHBVNX13UDS6g/rmBaUtN6yn0Zv
dP/GxlcBgFktj7XIw0zzxoz6rBlSYytTUYkJii7i4sZnookI2RzXpWvh6RAgTycnaKAsd0P2e9KS
qNTJaINvRA8V/vU5K/Ucfk3P7PTZB6S1Mza15t4qDknOtLaZQYAa6BRpetX6X9nLDM0d0/QK1Ize
Deu8OhjDY7UyckhJ+7tgsIBwLpulzYaaFRJPoI3gDzfVLah5MWERf8ZTSZ7o06YP2Gun4bYE7nj3
S3Z9hwzS2pUr1LHX0GvdoVu26CAH65VZldieMPWU/BO7sYTpMk2tG09EwJsyKBiyk5cBMLPS9k/5
SBRyJ7BD4lhGTzGLYgOI8vahHOQqT69slHyBx4DuUn8MwiyvOmp3J0Uvwoi3wAIYh1wWmdyA3pgQ
cnzNPWZNZrRS+/hVsR9D+D9obw3abAif7u8V3UHKctfHseh/VxvuCAPyuyocMDk+ZcVD6P5YqpPo
pCQsqmaqy09+BW/qPQo+BRE/D5WRMKlUdS860iZ+ZEjAwGyIir2tzKIgs09nim6JEAumSL9aeNQV
ZWlBPpUgk7E2mCnVoCz7gZRM21eYxUAa+alNWV7AXElqmNdSR3g88uS+Cz1vBJgr1zSYrDP83ggh
Gr9i5n85nTS47/aKu+XKe4C0xwSwYSq6NMQNPYs3whaGpc1Hem7znQjJ+w6b5cCd3OUaqtcq3VNb
s4v056gdLoAzoYkrLjp3B9WmnPLEAYcIF1fluy2KXs512Mo0kQ0OTqolFC2NYWD7NzhZ8FXAfFdW
LR3ywOkcnTfUGF1WtFvfjpP3yPtAUtUC++uqOEqQde8fLFrt4yj0KhVniobC8QEcseeM1RFsiAry
wXSMsyaeRTaU45TAYfo5UfLTOov0WrHKEyNEwXAvPhg6Fz+BhSpsyeLlnJk9Tw1sK2Be7+AKgjDM
byeVDlYqQVCsnRYgdy9FYBODY9UAgYIo4+dsAQT2JZsSO8vrWXgzOIzVcTYt4wBKnDtoXq4vlwSL
kGVcDPQjHU5K2xHlrFhYfaEgsquyvYoM07GsmXoecwmY4YibqEPXz6YACXuz/75bXW+twN6hEdzQ
Kbslwl+B9RZGENAz+G1eDxjsjtwsYsoomak9Ry7AB7ORS38b74CkXWNSjO6VHNwwABkHVLhjKkpg
u0HVNuWtNviRRlF2dExE45bVXl7Q9wxvPpbS3+WjSx9RaKbKGDAwL/uJRAP1sYeou9ia1BG+cePa
TbxST6nCHcL/KPakldMLB0KqqdCE6YCbaCLeiU9ioZz2X8DlZ4bdHVyvf7knmV1HLNRiMWEL0yJa
e8DjMnhhNOGspAyq8zJbhqJTbwRRgXRXvSggFqlvLbEyYh3JjShiwBuQGCou71ILK3xFUhBh1rhO
JyyEmixwpap5ux94dVncFi1zdxuFZWvUr+0mEAs2fuL/TAMASUQ7MT+d7RiRWWc6Zk26zo9s+OTL
1+K+Z7mMhsdbZINVz8+6pnP8BDr0vLU8ksZmfBUMg2R9If+shNeMeP/i2Qnb13oMW5bRwlO2DJ6b
g7zqN0PwNPcFPTGXj4l0x3i9wSmAqQdz7jl9lmNDJ7ePCpOgKKyTf3Q7gylqWdDiSLV2dZu/GNPT
zcXDg++0umYMu/OGo28IvPJtSuCceHD0kcDDwHIy6alMlqNHOYxocQxYUBr2JnO+C4KmRPulW8Xd
u+2tQxd+k4BlB5fgxFafs3GDUEA4YNa8pcW74cLS5ssG2gnfGY+ioauFivVN2Y6pbViD7XE+k7Qk
HvJwMgH1GrPwPd3eZ14pJ4dIcxW17uibIH8IJjOEy9gwDujJi42KW99G06a8P3T4WO0kpCsP36n8
/2He2COheq11guyRl6KjVuUFUm06vX0XM7h90S7HVN+FWXGj5DIjQOMM1zcRCwGmqmmb3D92JuM0
H54nC+pkKi9/5m69yf83N4aP9ekHocY7VBLktm5RQ6YE5YC2YVl/zjrwAXiw/vWzWUAtebqyNIyv
EDA45BHgOByG5DD8GA49Ah1GAbnqUSO8q9HRa9IIzCIz0aYfnKBxmDidiRgXbdM475cKcRPjYEH1
ZYjtxmTfqpK98hDQU20WocTcEeZJ3b7tDNCF1AmgpQ6tam5mn8NHKPZiaROgiwGzbY+eAS0hyYhV
n+YyaHxVDmDBh1C9F77vU+6A+eItg/ZD9q2bjDpVtBmAMss61FOz29GnOHEQ8+Khwfc7EFHOb/qu
IF1mKdg1RbV+G2efZPSyvSNVPqsdT4OIA1l4GNjfGqps8Cuyy25tA5qas9QaNM/FWuvfsjP6QkHj
xJmJuoF5JQ2OHd7QXQUH5mXyz+7bhR67NNXX6M8F1TiataQ6WaOIMWSz8u0i1HQdthuhZnZAXohQ
lcqCR91HZxG+tB2l9cvgR5pEja17aPKfK5Iiz8bQZ4yYvsdQcLFis4J1FOTOTP/62jwgapWzkVlH
bl8VAMk7weJJHRQZkggRhM5V1nt+253bdcSuLgMa2BlIw6xMC2jHNlATcjcNdR9Adpe+7v5r838S
3HP4p6Tn6yqUUtn9YvAF82Nn1AAUQ5Bf543NgD0Ocp0u8Sok8V0lw4JSPJfIq41dvjeOndprv9tX
I4oXtg2JP2cnhirX7MtS1Z2Jnqx4iWkZFCcRWx+sJMFdlU6gDqyuuwLWeFG6seziIBIxJls+h6D+
MOoMbPyWf2vTozYwmWjQdDJAgXwT8SN/NZgp8gWH4d4GzAK5Tvws8r9X1bPdpaieCvoYb3hanl2R
6LGdJwGLQH8I/cd55SSZOLxCLDmR8OHrogv4fcOd9H9uI8i+C/cbfEt+IiF8FFqO72y/MATUX7lo
/ZXJs1wFUYjXQA+Ksk9AKHPqS69eFWao+VL8Rsp2+2JI487TRcNvG/uwEmubiOhhTxCdhHX4uML0
t0DOnMsCPaQ7zf5r9+DWa2iQdSiKaBwyhl+bXvgg5Q8Sa54m/8aFSp0SI4tIOVNk6HsZnZpji3vj
2dtj3iZYV2Dy4WViP5KycrgUC1c9QZrymW+z6eZ/zjbKfMitaoOSl1qfKJnuo0SOUWTmpHe68NYt
SLyoXm/nOETDuN0gFKk0e0U5M/7ynARHM05SDo+kZ5gOZZ+4FuPFfvtVTQvllpBZKI0w3sPOnNsa
6jhw+gzEN8LGudPOuyLraLpKnwm8GZTuBXP0wNKP63AMhqGU5nM1zW+2kcKhHNk6MHJbTfH3QWRD
yz3F1QrHIYTy4WU/1aqwax3fVM2a2qEhWejqmCMd9q+uD+HPl+ksh2M6r4rP8y/arB9SoYqH9Nnh
jgXASWp0WCoXy+a5L/ZS72g/GZX9jNHcmeILLDFaen/au29+r3JbObyn62+gDURwGN2+5gzaw2cN
z7zu8mL3RoXhQgGTMO4DfUJ8rlojsM8zyP+O9JRpwkAf1FRVMX1IFgZDammEPxAEkLhs6u418wNS
eZAyfBtcMV2xRkhm2I+FQZ3Ou2EPJfq5dZt5FIuYuPSibpczuElDHz6/NNzL2lKBykW2jxJlglcb
Uv5aJayYJ8+SZnLR+naNQO0h7Rf1LM2RRfkwXZF9HsodsJpufFoXoIEzeZ42vtfJAgyCQV+yG0bG
g06WwjTzfjTWFu6R19XiOFa0+0TdY/Mb/UauKkrJffAUB1K1Nm1GlJBYDJ5Zjao89QpLxZca5Xrc
BzR4oc5jVVvN1wqub35W50duK9cKAPudElywsXyOrG3Ak71hnJPLCtaTHTL3mBy3pb43RBIRWF+8
HlRH9tJdgn/LvhkebuLADFSZx9a15RL024mV2M0kzKgIt+kSkHoI6tHcA9pkS+yzW227R3RVGHYt
cfn2ucwvoKtcL6lnQhQndRoe9HgMJ8yLX+7u3Z6eemPezDxsr44d2lUB7OqXglgetDPJaLwWm7YQ
liYkbb1Nlp1QQHxGyUdfimeZND4du6w12+IdnExpgm6qoOEXRDtqJ1r/GVEzncmWEqVo2Ssi1LsQ
LZEOK/jtfDyaOvBF5r9bYiHhbrLmSZpZnk8Cxja2LES4ksdLpakY3DVrvYmyA3YDpLFa/hjxr8rU
Ak7Rx2ZqltGpvZ2nitcUYGZ1LI9C0fjyTVEaaZ01JYyjjWCXy/EEIHyNEd56kSqr5w1xhRAat96o
ruCVHYZtUYFl4+Kwzthw2Lf7C724qGHJBMQqwZkTtSNZNFWjOPzvUp7UR9mAcE+j9QYGKv27VqZ/
3lmdZKgz2X4Kn02PiGGt073r1x/NosmoTI/xPrcwc9dfYdlsRPH7iguKi+JxXuCAmySnSsczlZaq
9wiGRDLpHnjqYgLSjYrXEsr1fRGRs+YwO1q7K15C547H+jNNX6BkB+XYRaSxQgY4SgPtWRPKRbTh
aLSxo2LIy0779vha3XB6pmFXYIH0jKXZgs0clH0FQbj5XPgvXafuTuz05/OGupkZTi6AXO1F6N4p
tG8+Y6nAFZl+8TV34RMmFaJIHQL27OhHU7IXqGUlnW4Ya0iKNsDLASNPuqbfRsLxC5/CViV2gsJO
ig2T1dIblg7WNTr8lO7ZuPBy8vP/+u2TQTREuOZeVQ+d4gLjevDZUb5K1Gh/9Aoi7BJ+/7LSiCXU
9QHAiWSzmCCBNZQbgHGVCws5DHHr9kXNrAnniBiU2WOYnkz+2StAlNgVKjT5+9yX13z2xLdIXmee
6WClgg4+RDrYo/08Yc8x1h9pfj5gfIeoUDcQGRRBAi5RT3sIr78r30GLT/YBygCfc6iB/zOizFvC
T19Sh25s7M3P0XpugP03Hvew15OMVwhAGeS6z/b5F9BmOH3vGKErPSBYAJJo+zQvsMPtAbROHxQx
Xt0n9R6OJfnvSc1wlzN0q53oGXGB+jbgzRSEgn7PNcGxYTLLmR6isQwJVp3nZZcyUvWc2z6Z9XIO
K3BewEYsu58YiHdsdLO7ls5TLO1mWbyY+gHy2njlzycs7j7ZLIb3h0CefewSlhT59mwnoiP1RgCy
8v8GYXpbGhTGlKB0yJVU98HJvxIx2FmboWAjVmjOSfgPKNcP2erM3j38fHkwjvNIr2pjBSlgEi4e
8l1dLh9OA5f+OphIJBhQe+Vj3g4wdzehY3C/AofAVkRjx1xBixcWPByQ8W7MFkQN1X66F0GkOx+B
6sJk6G3mpZKrsosKHj2cbrtX37cdvf+JvmhUzKOjaX3csfAxkGWblCEG4BO2adPLAhs3ELLn9iN3
F/7GZZo59i8Ot99y53Ntg2SugOsgg39GNR6NK7eZ9jswIYc3WLNY8zx9ftX6ZpB0cZTDf5ueOlzC
zHcVnkPEmDk6CkRjL/FtAyeSeku9nWaiC2oKkdMPx5PHmdwNnK7rHT3ncVfb+eKggqM7aQ9ZAwvV
tqB+qtOZls7hTb0r8ivwwaKFyeK76m0CJUJWBD8GcPN/3FI1bevH0b2MBzKDRSZvRRHhrGikmxfq
g19VulMKaHzO/5RKxDcgKQjIvVL93YGq5OAK1ExjwA3P0AOEdB+zVKTKubQOtfKyCv4hjDW3RHCe
09l2PAhbowr1n6cHPCI+nIyZvqSsg/lRzoafOSZ/qfvxVHAARDE9yNifJZv0V0vc/RE5oyuZW9wr
8ZpwTBRdauCWv90GENqN5haeVrGrp++lh/APty7zZVIf5W27wozIkug3EjAZFvx/JKVoKjwCNDa0
/dNmIRnKubJ86BB4O7jTo+N1VvKrjays4ytTrxdi/KLOzzsgAh8oVGyVeZKvU6qmU2Rd6Kq/G89A
L4UnvXT+d/QGskHyLeQWJyaUu8pxyvZ57/8iVr2NJ/MZKhBATWzZJDOEF4HpF6Ut6UgoK7QjcC3Q
N42uQOIg7z9c3xw7p2BYVgv0lC3rXNr1Yc3EIhxZxuTyMC6bSkmnCE6UYGuDTawkNEcIgk/Xz/dU
qfXGK6yx6fCrLVwi3X14o0z1Y2XYS+85ccXdqxylGvrkSyznMrx6l6wQmooZLqLbokQ1LKCRkHPJ
dG0C7BVuFlmffOkrAnNJreFCdTOYEksEktXdxBRDbJ7mgUbQelAPWKv6BxKCes/BOQgfhN9ZfdB/
WJSkuz0KAmTUCYCsWuddqSsodMgj/fzaWrCUKMyHdoBsfSqXG6gJBoSP/AcmX+hnTjWLoBug7QnG
AgPrgFJdGxUE4nxYunG+oVI7vr7/HsarF83I+ed9EPSL/4gZnfCaJQ9qBF8O/PoHlDjL+TK/fDdi
OPC6UmkC2+6hy1swKpsv02qfMnmt3R42FHquckaUBVl2bYn6bJMUjA/CECzQyIgA1B8BjMx8uTyU
k/CVgRvD8fwDXSPmzuTFAP+OUjRyxC2FV7ZdI/n/qpPuGytdJlySXRRFQOzB1FDJaNpcg+rS9M/a
dvRSEM/f3DBsmsXouRqexVg3MdG63qB4rDUtvWeNdUscu4Fofwbq8CmcEQJ0NGQJwjaSSqlgnnkO
t3IVsMgLOQzDFYqNTfuDKaZi2nJnSPpcgp2WStJeDvTLuPnzzR3qsi5coAVlrEeVn6KzsO1XvPrp
RQvgV1GGYSzK+GJfQxQEip8m7b1/dMDUEqUCgStKb0WCIoySpY3eFbBTeNZkaxXPsmc10Ee4ycOo
unoDV4rD02n4nmaCjWmSryNDqrut+QLeVx7793D9UrWslQBSKeOHI4qNeEbIekdRUjIQfyhBlXXy
JUjCYJGXxwZfoB+/PMtypMb+aUZuB4MH2dMeMtyqCD1gQ/UBuFy8FjicnPtXnw6b4oJfYQ8jsB17
8opnFA687VtB2a6YM6YgS0ZhcY3v/Csb+69E39oxqBeRgn6Xp0LR1qCofXOXTx9GZx/T5sqn255K
TmcUzx7Ygefp9klk3qTHugQMi+8dKpyu6bXvmh9ssKFx7NODdA0gwW78LN29EhRT8+fReyIfou6s
donNdsYcyttf3zRpyo57+UOS452SolH7curQ8/UyR/uZf9ZRxpGSA0PvvQk6cTEaG0wPJP3X4tKD
v8G3pXRiGt+RM25xcuAG/mWE6oCcCNA1WKETFoNtTgKqyeBlbuajE9KylbRca6GPQy5ftw9Vmjhj
KIa06AdiyCiOcFdep+OPK+yNHEJ3uhfUixgtG+f6cuO68KTi1onKuYcKpaxXZEWX79F5WJqS3exq
pfPqRuPjCDNs0SAtGbfKyNj6XpZe7eaqTcu16ajg5hNouR4+WF6VrJE2NnqJQwNrqNg877MqMXXI
nhspeFpXQW8BJ3mvPwBpdXrPi03hDL0Hx0VtkrZVoT/oPHSXHHWPfZYqxmEUNgWQ3cI9YzId9a31
lh9L/xrUb2sV1XoZMRpedymovNUNtoPGI1vhMh4jrOUJJue8vRyIio1dRAAYmeWiFI3ICPq9Kzc5
p+3DTeBg5z3ntqV2EI3C66qJGguSIertS2DBCblULSpXLt38kuJFfJstLtS25oVACDSiiXjXArQ8
1GlPFWs3I1/4UnwNuCvOt95XZGa1Aas2NmCtZT+gHpwPJ8AXgBiMCpcuoxKLvRQfqLkpZYvhg+Cz
bJV7reXbf2iN5So3rOGU7jWVY9ZyefFXBtGSfGOBQv1x44p8zXZebiHJ9hldWXMLKKWDc/Tjb8yM
IBoBKtKiA5ROW/rlI2UuHfN0HzYyQq2mG+RVJPNfpCE9b1wzUQIRICKgnmNq9A+iTFUmHf5adxnx
EeTWPBaYKz+gRtInJwPg9hR7KfseE4uveHHpTdLcM9C/GqHA1wqVUEZcI7k8WjTHnaiBjc7rWxP1
LWO8VqMRl5frm70zpsOqVMTLY3zO0Seqk3hKaH0MI7J8izNW7edtjF0j+rSHS2pqG8m8UMTDQoQl
7kM/InHdrsYlvb+C1X6W5C0qn2p6SUaFOJtDHYsQRdVwgZDl9niKqzLGkFQWsI2c+tV/Ki424hbP
HpvU4tYc31cxHbWVtrwxQ04Tw+hNDwZ3o0AjAiZdrZ2etLZ3HAyIh8Y8LssV6tp3eY6z7Of1dqa1
5HV9zMYG/4gBmVPGwdpJrty5aWpIW9LQP1dZFJ/4yt/hJrzWBYozxJ44wK/+cjPmZImLdS4HLI7T
LVGaf0aXVOcoHLRj9dXSeyAuuuX14I3AJvb66BhtaesdFyCk1M1pD+qpnjg4Y9EEcLgOI+wbX5Ib
wjlzB/8wDtCIAaTB3jNYd98WjlvIRWdNQQJH3S3I3zJ2AVZTJZtFhUda+raKuNqXArr/XjqHVaDu
uWKB2VEtsnNjaK5Vr1qqSizQ/H1DEvBYcovuL2jC1bTeuLxdzcra1582KOUsemSpQo3MAGNMtwJo
994wWunuF2r4QkLOWVTzD5ehpD7BKxyfZSYIzCLbWLGKyqOwaaYKcO+/oJtUOciSw2t8bHGkdGcS
WCCbHL9FvpRMh/uFKO9i2R7+QJNjGlNoQiLdCPWg0txIuFgBZ2OXe4SBfI7s3lpf3GVSlgmrhmFm
7Ip9uuDbW3BFSYOc+4tdVpUrlOrWr0MVaYmCHYtcpQbQRnyOLROql++VK1k7Tn/GzvuBWF4Vk6sv
0WoQ1G1i7junlTSmJ0sKrmdQFxHTgz5EefsVFNNnu0wQTg7rMX0vaWMbniMb55MbQDYkxpiMN0zT
5Y4zKSW8VQg9xog0PbTQ7XAxxns5L0ygGeM2o1duzeM3CraB/8hqR8XgirkmgU7bANpzTkZEVsJQ
0Dv90olL8HvVrDzsM4+XcYgp1eo8dGXTlGuUf9SR+xlc67vzmGQuKJ0J6LSoI2JhtoZnE2w6f536
y42Rpx6B38oRedlGblpggvMnKOkA/uXVcbfXhtHbgI95987b0NU8t2/NJygzyEd0kImG8rXfGchB
7exVxsS8KiRxZkiEGxebHZarT6rgIWzmN1GPaRHcOgIwObXBQmU8iqpE16s3/VnAYWD8AOlEheXM
hB9CPIYmHIJRcIRv0kVxbhQ8XfiuQNGLMsx+QWwWz6F4fLEgLIm6Z2lBKXwtitMt9ymjTOWCSiL2
i+Op/nevW4Sx1wXJSay6+uXb0g6NpI9VdrM/qrPrptR0vMPYdQcKp3M6L6F8rzFRmf8CqbrspMKY
GkwxbGBqLBELE2Dj3xlvfXy6jKApD4vIX/AXfzXFFkTtwf3LQCQSuXFJgc3uYzp6uMQN72b0KvBi
9xrl5mAzTrKWV01hR15GOKLV5mkgffBeCrQqrIWoQTNBQf/VPcLhIypaSXdWnFtX1Ypy7SqHLR7x
KcQDP+iBeAEgbzGbLEKFmUA6Ciwcg4dukn2JQeosfW+qD2CMZsB2uy7sDys1R6yU5rBoGl5j/jfb
tOLCL+H3XPhFp2QXFHH/1QMEiThx9rQJyGLMvmCKlqWqkPIArpP9H58ZddqGNYg82fZhvcz8LY/3
w61gZK+CsnRsX6mgjlAGiOSk2wCGp+7j5zJ2rbc4IfaSyUp0fgGEtYeeCOM6nJfLRpr2hg3F4+q2
h67vbEwRpSSgWqAryslnRbqC92SKg2frP5TQFZ7Mgb3HjaCgCFZbusQHPyI7YVIPUB3zB+9rapUf
wIeRiUyQdyocI2sqpsHTtQq80y26EiPqDhQg7tPqrZckRMD8fA+mRIvjpVPizdTg41nnx7CFFsYI
AOvtsyYQ0WttLVXG/N49hypQmHtkQ26SbQm21jHGM997TVG+WcsJPRpBHvEHr0sHF6SpyD8SP+mY
C1/W3VIlb+blhq4P2NxrojAlbgRcUvbxwedqzxF+PU1nsi9FRNw5eWtqujWpSfglyu0nyX96jrdV
vM5FUwJ1iqif/SV3G71QlHR/HGpGJiDzzyl0dVePUe29R+M/Rg/kPzmhi46gwY/JoSubYmgEcKDk
d8A0rFDJnPmL6Kh1FBjHdgBo+YfdQtVsKJyde32vM8VBtn5JDSEphLIEGcQ4oX19XDHaiCaCol/3
DKDzyfYd2uHu5wY/palbZIlFSEO4I/Im0yLSx4ULgT5ecGF6hiueMU13H4m+G9OMQUiavsS0uy9G
qab+B6UFSuJIUGtNiV1drgBJRAJe/Rl6r38UxubzP+jSybx1NzJzND60pLTfpElPutGaSMtwMiNS
tjtePGYLINVN5Py5JvtlX6bWtMx8Ibh2HD1IjbRuNYtDsxKlT/KOEDXgyRW73V5M08hXw5kiCk7L
jVLnfs08RXRPEHJjbl3YsLVFL4wNaFm04jndT4NXEA6bXPgrqhpVsr3u29Ol+BEi7hKocLyJK5uh
CffTXTi4BBqLMnAXkQRIL0qrav3RDiHZq0Gltw0hulsFvEkJM+r2Hf/ERiWiLH+k7mIvOykqvNj2
NALQR+tKACfsZXzxPlhF743LJxkhLGz24tUATKqklRJUZm+D0WQ+c7fmDkE+wKtVzu4nhhSw0jj2
wv4tzE2GmvgTCr0ihcrOUtWkf90KajBCc/BgzsvEgcCuHQn1Ett84gyP/FcxrShhIlvPZcSYWhgF
XF4eFo+EYa8BB0PybkmodjWYR2Go+KVV/j1afW22PjUaTw6ZpwQ0tXBTNmHBYwArql6SdfYdSP1/
Po1UTYBXgAzEIk1L7iGQaBq+44aNDV0keY8huHEYrLAJwxNsCbEAXyw5/Qt6noRE+UgzpIBv55pB
oRPc7yZFt6E4ON7bdjLtYdXOlws+OrTpM4BQW3yyAUfMIUqgFeOnx5P8iErLlP5dWlpSQm4UUTuJ
ebNEs1X94AW+c3xf2U5lOoBVt+NOwJLheJXrCQLaJZMIXD7ast5WX+1evcbL59FbpWVymNz+5uq3
bsxMRHQGYaQc1Zr1tex034qyU+E1AhBJoDRgaER/IFiluWHXU60MlXIrwPRZF9KGm3gOOKORe2vZ
xce1o1SAZ8eIhWXrVI/wbNDfZH/Mdlpsi16KF1Rgp7qkgCsLVroe56BkNPryOrjaUQNL2yRurL4y
YOY5KZ9rNBYJD4uRegyrcCvQ7Nc652jU3csz9b0sVvfyq3CA0EpKCizdzgL7GjztUfKEAqYE3OYf
fHzF142vNlNqo18+psaXSjuOvYbFGnKY+2sof97PTiPEMfjnyWztm2GpFGK6sfiuDARQ3xBBBZQd
/whadzwCm7fetAWIi9CDIXlZcddirdZdQQri1dEk40UNR33CzF3W72iTJywzkeI80WGyygqrvURB
IO4ODUpOkYQEDntb/3ipF9HZT/P1G8Msa/n1JHCX/IpEhAxbiNi0cqK3VGTjrIuTWrZH/TKqut6F
vXoh6toS21MmuI3Ttt7yPruFx+H0tSnSk2XNC5Ee2hIhm9yhVWQOXUzEjcfMcaoGtWbNbCR9xIEJ
LcxPwp26m+xKL2gSylMNdFR/wUxgWJs0p8f/kvlDJGMdb3KH0g+JYpiUtuUB4LQ3ThaimKpqoRQ0
fh+fAoRh9yZK2bvibGPhezuWv9Sq0Gy28sHLm1a/a17HiwnH4hssU/8i749Qr68lgriAZmlmO3II
+7quSJfup4KeKCHmKH8MGEajqQvGLr92p5jizbfbXZvThu1KhkiLcZCgeHhvLo/7DhOPw+aP0qlv
IDotpmMn9PDOXuWuWIXZw/CQ4gXvSjE6rmk9N/CaZFOB1mtmZycLg7hl+AaBHXfzb3CPRrpFDt1e
BqnxhmR2MQhvfSr24yBC3w51rzRAcXF9t44ldSvu1t6/zJKkQb1/g26oPG8q5dOAs2s9DpAmQB77
zgcQByb6/oGW4Nl9NnyQzEitumQjViHSLgJ+/8yxk9NTZDaQy1nvd+rGbbOlW2PqFAy9VsyUG1TG
rTc39/Ig0AM2dI/Mr0Vf0WjKrZuOXNsF7oax7J+qOXzND94jaTG6nxYM1lQwnGbctP5TftKjxIhZ
eol8jXGlCWhptyh1hu5LHqxNjIRow1e5HUtaR+6QjF5QcnMS3I1TsLzqgYEQ2h/mHKSHhIin87TQ
I5orStl1In+UWqUWiFOp4eKT7Nr1W7l1t6kCgLCdc9yTAaG5264mKFMrCV2Tk5CNBfwZW5MGak9g
rF8Id1jdzDogiPIZl7ImKptEqZEmJ1r/5GcKB8Hc18lRB27+mNuH39vwfuQ93MOzx3syFOacvwd8
QBHZ09uS3oMFLmoEKTmvAIdB5X1Xit6K03bWfDiMeJW19zQWTsLAIZ307dP2qWn62itthadLT+7T
LAcLDq/S3rf4A45a09EnjOSzE3aVaDg0oVq2rMu9UI/ECEjteIU+iR4o083G+G7SCf/WFI+cDR34
t0l04Dcq1xfjnp3VWhOlbuKmNZR/mhFDJiYXRntmQZvUhqZfYvgwwyw9jDtDWreiFA5nT5H5JD1m
UDfRszya7aPJgao6+RA8CQL5MlTQr4IKpMlP9SYYlevdw7N4fY93uq4JmZS4uyKZd9bbe2tQebIN
WrEWuGFwHkyEsMvz0+oq2fQaC3svkJZRQqtlucTn08KfGjKAYwjRwTV+Umz7hxsM4jtusz0GQ1t7
9NfcPKuK8TNzPnAPWpcMCrDSLzVOfES4LSE6WaeQLLykGY2f+CUiTqoi18i4NmA8NgF6ZOybLqls
6tO1AUKazgkQ119C7KSj2fs8CDJZd5AVx/OoGkzEDL8Qo17gbD2Rv6Z2h9Xg3MKCBdhHeM1HIg2h
BOsGHGKhoiyw2r5HUGzHK/7Cdp0Zyc7depyX1VpTIulychHGiDgqxkB0unAOBTU5cSd7LcPzBhZL
0Xly/cv7CzvVcY3GQToRffkFaHvkukOVqrDGiABVxBbFyD9bORzxCSGPFMMZduT9DfRs+kDuN9is
DVtWK2IxDLe/ImWDe54plOKu020G0D+YNpEunU9KmtWr9Va7+euLdkj6goqjGT9j9TPdsp1PsZ6m
cZBCqTA3jbHIcmyVwZ95E4hjVTGcfPpcwY6KVndT727RJ96ZwJlqA88t6NNUdHA2dWWLqKS7FmJn
JvJB0eOjzg1hmyeEIITdI3f17qPFDLWuqUkGkUTFY4LqYKSMNEGFzr0jwqZojNKhf9Gc2puhwO0F
TDNhTq24sO8Yrzm7uto5IhW9cxZmwCj8Bn8xVjPgV6/qQwA/JHwBH7nIicD7QgmKS5QvV+g0Uot4
j4DqEgVGDXkGeQgWKc9bHQUVm+l8C240sUX4etPjEq1sZzoMiThdr271Z5mon68rU28xnF18/JwT
/UGPQ1O3zvO1kn+7iY5kIH/z3sP60V7zP9KgNw5w5aSX0HtreMiK8AquoO4ym5G/mZb0/Ttp7gfl
ElWvnlgMDNdKou0mQDA9zZo0XVgyHk8L8gvDqkd0Kdfk/p6Ogyx5tBg2XN0vkSi65uPQZ3W/b6uS
kFBoUbRnbJszW8AyVwEua1o0taxS1SVLyovkTZSDFUzAuP4iLB1BO72FAATJqNk2lqDjaVXjRZQi
j3QohtIQTwg6GSUO+JK1GrrOpCePYaNhKe+uDtYl/tC5+qcsEFbeJjxhEg1GdL4rKZgKyhOQrppq
gbuDNY5gD8uLIW3aBpoIh5f/68H1RI9e0XzcbCbzugDm6fLtja/ir+1o1pwqCyNOwxqwUZkASOyX
cx0TmlQ1Wz+Wtrwq2jgvBBUGXWWttFOssq6fV+peFLqJezsiSY7px79uxYAW0OC5IgPHcWFuZzPc
ouikkjd6WOKdValhzv8FSodU/Wz0zVED8ue+1GJ4beiII5eCPNx4JXw53h9fmr8olsUcNgMrCtSA
feWG6I1zTlAE5OuaLD9Zu8a1TEdMmrqWD75LHW88W1+VGYfP8ofiD8mm7UzRWIM3w+0pedpqT5yt
lNc/aoU6uvavW5VUMETClKQMkLe6PeVWXQq1z9VPZcSBJmO3XeFcH5t4ls9rYc0tGRIJ0C0YDjbr
95OL/AqyBrXW3wLMnsD07ar6f4jc+4w1684E6fYiwn5cmq4aUnEA8C0xjmf8q8NQRCXURlbBn9WO
nleAbhOtE4LDvxRgMzcIMY+/3XDNhe363To35KY3LlJQHDS6XxlfsJdzTfQaa0VfiFxwQ1qoiqZv
ERH9cOb4EJrpkYTCWIT5VXHhJBFZ8CvM62T2mfmV6xuPuDOxs1aq3GL6DbDf2rzqWQMtyMJywwLU
guTqw6lAKOT3xDwJs3APwbByqAHkdQc6HpGwUhGk11+J4kawyGHjhZZ25ZW79jb2ujdLnkrjdpib
09AAfyR8/opEyahHWE2SP6PezgSsjJA6YBZ6ZH4McwaoxsujeYEyN3JGy58taWQJQchOYjtlbrH4
Z9FFZP8lBvjnq0X+0fjnh+6t2A6ewyGOCaCWdQRr6xYvUE3ptOGIU2qqNGpnrbaJhgp9yyvD/ptf
MoJBVHtwIejg7NxCSuyMSUAaEgbjJ+5QcfhZs7MO003tRhGaeF+1VyX29Pau5xXlQwWZV8aEH4LX
brX9UGWYSIS1t7i6G5Pp7RhP682MOB+wHEI+41V1685yw2F3BchisryCCNoYRS4VtKUTHvs0IhIK
ksQIj78efe4Bx31zFenrLG5vCqERAA4yHj7egg3aAaRhFK4dDw0qmMgd+HDMp24cHTImbtwejFSL
qRV/9N4HgdxLeuErZHLFFdvBRwrwQDixRhKIETjYetyTRJZplq2E7fwHNPL4gbcvmp6Halvqa0SJ
rJLUod0uEs8tUDtuS6xp7MhFQ7VO+Sh7nIj+g1I1ud3jCtppCDJ0BzRYgFgRlME1WZ5WwFlewgjM
A3xmVW3AICDpFJrhaUxs0syc3QmhbpLbsBysU1BYuRUJAgIQXdH9cHTwR3jLWfshrgbhaMdbU5mo
l4RHkKYMSbZ4xagtR/2DWPIJwI64FKz0YvMtV8XllGlpfaKTx/2XRT4ujNpYA8oTxPZ3ef65BrCW
BCBGbA8rJ+wGefgjw92B/npvQm/A3uWUrtVvAMI9+mO90QT3TL/6xh0t0nDEGbvxqRII/+BLZ4ct
s/fX1Y21HtY7+8+2Nn2ilVXUCg7eWCDbhWkyFjx3CxcAL3FRUIp4vomHWT7LmJGbVHjmoZeDM9hV
iKS3OGk0lkYlbnhXmClpstwpTcdXBcV/R2m3NBBE0h4NiE62ZN/EnSDqoTqHsRJ/980T999WZkvD
NWnUhBsu3V9a0cvAbljESYdOjLoK1fS8gZpWodYw87PLx7lJUB2R8uCERfHvQjB/Sleyxl93J7gZ
7Hi7+rnG3J4ze98dNA/QzoQoJlK7Jbla33razhqAGCRJQMuORgJ8KKuONycJ04VKyOqOpv7sEodO
vMCYHbT1OciNrHFdw+sbrZwwfkaJVeFKk5bRjCVppNaMLoy549k7ct/4OLPpUMTD40nbTlfCAX8x
JoG8NpcoJ9WJisUS79a8zysvppeEgc1HYApPTQlaX1wiB873SdtivWYjod8dvNqvUlDp1R4Pi582
tCPzN3hZlqSJdzVmRILIQsskCAV9sCr5IcoBEMpzmcY000pPWk6+ByJ6ymPhgU1LYC7qi//jL/aH
PkmBoiGXhTRCzLeBl1VoZe3MY9S3IPx/9y/SPv6UytlTJNXPpcBbgud+JjeNFaPD41FBtrqZ5LTZ
Xar5S4vaY7eEWN6wVMnc9GrJCNfzgTsWkTGj3MDPly1JuxYAZARiYgGh/PCa40ZgpwUQbcLwrmc+
NGM8YkSgZSQZ3KGJ5T7i8gt3T9Lx96HRRaCtBsF5BKGvYqMjPmZp9ecx9KJgiGZhMkWRMujg+RQJ
pVKS0sD9TyA56tI3nBWgsOTmT4A3kd+QqWDZqrIm++K5YfYuA4EpjhKJ7fH7UchlGDUX5vTUbk71
I7nwfydkZ+h3oklvHiLRyjKaktgW91NiUaURR5cii+rCYZ2XGQXxwySSUS+erfU4J53ehstAro17
O1PSXgLvFyyIvnPF4iWLKpLM8vdJjznQtxfG2KQXupKHdwJEYlO7t0RCb/g9qkpP2CpHtO8hCbVm
GkNQj6poUC11NrF8
`protect end_protected
