-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Q0E9VEXto6jhlXgH34mRg8OfXEbEfjVnD92EmAcNVvz0caxfXV2JnMNboNFCGo1x
184y3QVN6qydS4P6YhybL54B67PBKIuy4zsKbE4P96KD5siK+tL3kmJhZuXn0Sl+
WRMvo31guT3oTq/xfSRGgQ20NOmB3d9l6AD8KKM0Was=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9419)

`protect DATA_BLOCK
WIVSDstV1ifrT3y7cbr9o+cFAnVpNHp3ms6XQMB/4pdTuanqtqNzjMEBGMNENB/R
qRv7YKwy/2SkOOVYwRSfGQ0+tM0vJrzwQBgwPbgjWeEfk4YujK+Vmxkyfb0BA0xn
Rllyd4UtChbgoDoymLk9cj42yVDEWJw+qyczeQtSosQnq8zEFOmGq49kOpnecJ+6
hIBLdEamnHKS4x+DxEJF//PjxpaiKm5y9yfMl6sX/6TEqiwjuKpFuziUTXnIWac4
PG6RsscuetHqbZB8rDRubWG6uFh8BF0R9mfKPKMe2gschN4WZu9G795yEP5fCMjO
SKNNOfNht5CQ63iSMf8hcH/PR3Q2rdEKmDlViZt0R4Cy0jO4Mw3hj3YT0prOr9bw
v58y2kI94fiuwC4WtZZtK9E7Oww0Icw32yXeFwyykpuPEEyVwfiowHohI8JPDTd8
L7cii/XtUTT3IizS4YkcmdZIryUvP1wnCN8k5hC9tJ9Qsrp5hyF8V9vKF35yIdbB
TGI3ECIKi7vs0x042Nx2hr23ABndi44LIYV0UTMgA+jqS9vanx3QYBfRckxyAPUG
1vOtpLmsZosuqf0jSw+mcn3w6YA760bE7cXB1h7XVORSL+FPupiWrVh3dKxp0bCZ
bRTKYwEwzNuuvdNO9torR0QONzBtv7pPQG3iK6uWK/p7ztKIRMZK5ykXQCisd07p
Lw96jmFh5KCZ10fFyP73vLwF6FU7Ca7toQ3pbT2FLa6qqXzGhhZdLy36pTObumSP
xniP9JO7Z8/Gof8Jz3omlS6M1QchdkPfOiq7CuzXqUDIl+xw4qD6vi0dGSadEQPt
wTRpbU+TxBgTQnjjOrFDPsOsllIYXQ6WKExFsz3BpvVDj/Ko5F6iTIb0vsk40gff
2rfMnE1sUQudrA2qrMRW7ZwMMSl4limXYtkJRmzpG7cuy0eHW1tx54saX8ah8X4o
s8ZfesVfQq8rrASmwdMIki5HZz5gaiiqQfR8MwiJMh/2AxnzJiU4PMOX9rmqOKva
FrZINTMznTyFi8HO5rP4lTYQSrheeji38nvC7d1QKba6H6wngvR58Y/0SDcFBVhx
2No9z2XmEgZDbfOS6f95gM+bZIDBkB22hLRSKYesSnMZ/1MyyEpkmatEQrpbf/nL
7ZI57wJL+Lg5MZuO5YmB8KedtTK0WZHTOIPkGnDHe9wPyPdyA+10z7X5TC1DXA2R
DagZFU+xx8FLkHIgU2epUuiQSky96otSGuBn1eK9x18HgkffRb7693+eTQnm0OLe
yqYbtPrl0tBJiVl/k0gQ9AlxP33HwG5zj86R6UGljnghr5W+9wPCjcI/V6WBtrrX
O/kyceHPIehBeyC1BbMen1MpS9EW0401a59yz7ZyjQMvM7Gotjtdjas5uy3vHOAQ
Ten4lS1HX1WiTLzEYQRczJJBluO057ySbN5FbdnBg4Qeqg8aBRlnGI9Ytva4kQGS
FWkZcRpmOKUOANZtpBzop65lN7ElkpJvCCMVbBa+RJ8zUXRhnsb3l5X+mDZHYFJB
ZKtcSH1UzkYohvpJtK9oyC2lkqzryRkI7zha4EZQe99zMh94eU7WBCFy9yXE02Yw
VGVIwYY3Pnab65Sy9chFugJUAjpjqbvCYeuYHl1oQd2XCyx4bDTF3U12KTN1rXAp
97ATtzE4lxrJjTUmBTrznaqj903RmUZiGgbIcQ1aCHnv0UtXgZjHx9z3wdrvqSB7
niQD2lCxuSs8xU6lkhsUccphUEGFKrO2Nl+dYhdPezjS7lHzgzSXXPkLx0x4Pqqo
upZEFRyxyySU+BLKonb+gjb2lqdxZHLvubqmiXSVK2JYoUjHD/FE9F3YM6F4vG1/
RGqRCJxPBm71VhmrN0nBmWtMrpfk0r192/twEsv0H9TuNUvjLFVwOEW/LvQ8MO64
aOeX0pCdRgJK0aBRoNfrKhGDSdEM7VYoZfMv8sJDo2Jj4CnCO2uhudX+5IIP4W0l
F2wxFlpjsCXyx/iZDMSra+gvGy40mRV2N+aQg30svcX8X4vHMlZ8LVLjlM7zh6IN
abkYr02wqdkE+eYtPREprOyuqljzN4FPQTHe4FI2dH1ex++YYe+9fTqkx5lJSfir
jaqdnRq9TNOAaRKYUBqtM2994tRO8WNKj1y3w4tOJTqfY3wFfTFdH8pREUvXvqqx
lpUL6IPin119iV1POEWqmvvbkzt/4tTJOrap//RHJNc8rry2eF0HGw9LNoc2oRWU
fvW8HMYlMcyiVKzyj1LNC2dEdTNyPizM3+EwUDgnGr71/lngg2ggxWZubJ2+cTQN
UYaJyqJ6L57rYHRRyNv6D5cGyb3NOjakdjDpRcggTN5fTC5oKOdTk8lj4B2mI7mn
gAnh6mFeWZobnJvDkH/pGO1qFCRk8MHdzpyIBjXkOX1oxvvg46MeCuOVgM1YV5X4
l12hOwLfmqI+oFGGWhKcb2o11ZGoxdhnNEK86k0XmxDW7t5z5Rk7IdAKENyMJdwo
eQV1VdrRXl4pNUdZFSZmVkhheQVeVIuA2D4rPoUiy1jULV9FtdHKsmkXkUWfm6dI
0lMJmVQGPe5utattZkrIrG259+/m2WXNnYg9qsgXN7ZNLhaFQ/oBVX2rAbrRw0jW
6I5JPG3SFmTbzCziPWtiqnre4l4pXwCXteQMvHbuEApfyonUOMRYjzSvmRWsFZ4l
RZOtSChKHTaFRQaKPEJxJh+1gaqSc+YRSIYSMheQZSbwPzMoMCEoBxnyDZmrEIq0
QIUKTRH1NUB4vRl0sIJt3w8PuLxsaP63pX5TetvtSIJ8oe/Vqx4HikLZAyBxTiji
PTv+FTRtIiYoesRCOBkoX15iCXAXX62aH/in8zZDdq3Ty+8s0d1FMGTC53UGsHJt
2zpesY8YTj+CYgIusjM8kJEO6RjEwGCYR+ZMdfOrzwUHY++EOU3n6D3PvjK3B8JS
/qF5DZtI0ZeiOj2nLYHy/hq+773/h8ai0WylC0I8Zn3dmWaqU8a22qS1yD7hF5An
lyTQAb6CXUNQwiO1Aof16VhqBk5GnmV7xVPNfgx47aso5hTcoKiZRrvcLSAgLy0w
mg7mHnhvL2/wr47B8N8zBWJ+jH8EMv+aJGs/kl4V5oKD870CrZS6iFzD78anBw9E
2iiepSoefB06jV/T/UlObYNZ/M+ov8A+SObSclMzMESY8rifLCJc6kSD/4deTyyK
FX3X5CLrwhiG4GuA9oW8FI7whUDkwgad62JYZPJqw6SrYnK2x8QcoG44ZCbSCAPG
f8bA0HcUgdgLWICdSdLn0wOxgZohkFAT/eT3YFZ3+R0vE8t1JCwd9Plh5vLKKdO/
LmoGOYEOYjAHgYRN8dHY2t5p2ByW4M8CjbafzEF413EtbrtSNQehbG+BjVQwsswK
yd5UyJpXubRXInjDeNtGZEUAn5MYNt2W/MoazhM8cFrxx39hJI6VQm6PLGnlN3la
PLMWCPjGIrEqzqbacYOE93KwE5lrzL5xsZExab+7SrM0h2lDcliWH4k797RlQqmh
O3qnTmcJa9EiQ8MP7/aPxb0FaevkuORBMG1H4bvhpuGq96RuerWeDnXar1rAL67F
WvXtqPDjW0mKgCP36SgmA8b8mP0F1zpJu2aONKwz2ZfQC405z4ih8NBw30SXK3Ws
CmyS73VJBaeTDPN+bl1roWhbVz6mYRJ99lV0mDgVkA4euji94+ftU2s2UwHbU4U4
ZomQkRCh6JSs8mITLgL+PKBxlxJhcyeE8W2KTz7Lciuh29pU9e++u4iU9d9MhqvG
fQDkIeCr9DTjL/n+9rqHiSjd8azCPIW3mnFZzaSw3Z17hq/jPeL0uZB/xhlE159+
r0uVABZdpuY15+6+U+1ns/5BMA45tKwLN5pD+OapPHlhWnslVRZniDcCG9s4+Ybg
qCMywoqTrh+vTd1Tauz7zOKGqxDmPYG9GYtXEFK9q08/f6xSSSmGw5RwDz6aZpps
YTYaxH4bSXqHb66L+gytVwSnNm71wkG4eQYpcFGCIv0ZcHZBPVYGg3ou3dB9UuMR
lUEKjGX6BhQHtNTjOVnbCB8UuWpqueBdSnRhl6D08C7Ys0Dl7Il8oW3uLDb5zqUL
Vhc7tVko/mlPpjqa50fAGfDS3JPHZ4MrGvGw5b1fJFiXkWE/3sQEbAFl1/ftox76
Dxo1XHCUkCoNiltcCgCbTy/3MxK3ozLkGGQkXP4Gu+wkakVdgnRxWRdgmSDR2qZF
jheQ+qGtwhO72jpwYcrQZ2uLW8X1ed0uFgGdXz+t+8PIPE3uV9QbNGl3zWcVDWh1
KCQVbnmbQFhd0HYRJqHslW/TPtLqefsmRfKvK2IT3LcUVJ4d04A4xSlFhf9pK8ER
8En0vbpSApBH49Yx8+8AJLv6q70Qj4Hpc8p6582ytFRkT6V7AsaHW/Hhhz9T5QPB
FhRXOBbfVyOpY1VBmQySIW42+UHaPci7EnK3nAklclpLVmJqd02uQaKpg233uME1
AVpCDGOs7w4NyzBcaGT9cKw4VFCl0yvXCh+1l35k1lAYvnJb+yq8uT1puqcBuTIc
rFuDSa6PgmSSV5lSaELiJjvgLSY5yIBCDjsbUQeItY7jlLsfZECezOM5LZOmS4NY
Ma/gTZtWHosw4E/+VvKpmHdqrDlYLlxBSAOyVB5tfWXg25Ubk5v24qn12YE7zVAY
FEiWdZrX8/M4YlyFp35by8HcX4e0BZ9Os6x5UXZD8viUmxU0DY1KsqAheI5zInfV
a6D9EvOx6CKLyJWUmriJlaXPKc34cJfKMFLU/wHSGgPRglQAWu1JYJTTFGFaGDTm
p4sK5E7PmfN/VMu3KDRQ/X6dlOQIvjQi2Nb94iLbTIdTAkDL//bbDHBIVnIBcLls
gAkVPrWGy7gplIoXQbEGxxu1HEjYHe50vnVKKx8khuOKG38UW4lJbMRqhB3PWdfW
NVJITcRExJBHaQB25P78iwlYbpS1Q4QAvxxTGHh1De10uBcWzeAsJqw2e4EqgH9s
k8fw4NcgUou1yY/iy0cFI1NtWmmREb3AvkYVD4FnVCp6Jf9VVY3y2oybqBZessAU
4URWiuOj62qbFddNHMWEDTLVIX7AYZ9K5mdx3QKJeNNnNv3vxji5QATKdDs+FPXq
MLkGIu2lSFqrDMHRaNifvN3JO9CGYsSezhIEnuYiPY0CSqoiLh52cEfHlT4VPirN
aj/JUpaY7r3zjgt9EwA3T06Ivd5fx04lUI5UtD7DD/ea0tYU9YjKQHLi5LS3pUUg
jwUWBBl3EnCzHQqCXqR2cAuNnmhw+ZCliMBp9eLo1OndT1yEli5WM1PqxpFIAT0y
Ab2MSZ9bXI6FsBeFdE8vsc703SdDQRqAonGew4jHpQbSzNXmVzxM+eUL6D0NciVm
MnWNTPYjGMl4kvBPw+xtl7y9CdkCp+uqBJz4EAAHNBx4EGdJjz5Bklp55DuIA1LE
P4xogr5tkP7t3w9nI+woEtfs5Ap68je/PtOd+B842pQ2pOirtUG2rlK9aFL21yA+
7+/tfv+8eSjyCxsi9DQs3Soqi0POEgPolwZB79NcJD2nfXFpIqeq+j0j0UfoAfOP
kF9wE9fBAdbkWW/RpS/7WS9WozCOY/rHOsAlI2OQCSB/Y8bodE8y+Z3bqq8VSMxQ
FukdGVNOn2+ansZ/EVXXMN2u4So8a6OK7aNITmbEce1rTykeQzE8SQZKR/GmHM4R
Tq9TMnafFXmYdfo2mBn3wkCU6IOBcxi9xJT0b39s5TBMR9S3WGjMX2/jk1aMtZM9
tu2SApH5AjzQoUPRKHlRpzHvoNFVDyYc9wwIj9pb1gbA9VqSmgXFFr+FgyxyT8Z5
hbDzqz1bkxlNRoHTrsLu8SbaiX+WOUtGmyPTAt+mwJSiNxQ1qePsUjDHo54LZkK0
GP5h9i5WD2xPM8mNr8eJCEmvDantbI6ZAm6mI2mahaU5HWFGKRzu2bpbLDjKH+0h
UUD4czShLsaWvSACjDk8FvWYJXsNUpMHHbgjbwTu0MwM7MvDeRWxze35UQ20ZDHs
F45CiL3Q8fozlwgcHVd7snB/td2W0JyDxOBDPor5ZEdGi50FowyEdgw3tiGvaLuR
jwJWAqZsWNO2HzRqkkAIWwQ7UQsfjDeE9VOYasj7wgqBlx8T1IDUHR5Pyn+h9lhF
HnnqPUs979htvJWjgHRxgonC0ib9UDWki86NyqYW4sAODAI9AC7ujKYlV/MkeF1w
KPjdTzehYFMvnxcwRzdH2wYUs+0VdA9EKD0oyvxkMJax7GOLs2rG8nP6YQ5Xg9k2
WZCriJGaSETLvviAij2JAXprQ+vl/NCBqzuctzzH/HIzKSJsqPTUrpQEA56xaVKF
6moyVMEfnvEzsZkIDXj0stKCZi4tiFLLwRcJtgWXNWXn+0QuOrB+9mlyVNcVl3J1
gMCIzurd093g037GBRmCMWVlzD8cLF9X83fLC26WUe7ZIWb7w8VOeYrARa1l3u6U
AlzveTiC8OuywsPuxNOkVQUxWqdci7rV0+uTllFj8a84hRRcMuuXtqjbWP9UtFfO
JwDOvnketCw9ZYVSLmjktALiBOimoO38T5G7nRMa/gWt9jS04YNY5hTTaGXdqmEP
/B++OjzuTQlriT5pIQVcOGjn9Ed4pUM3HaQaXG6keeJXs7T3D7bFDpBL5XMU3vAN
1ppzPzN7HdVlxY1WYHI2AF4BvCo+5/X0TqBHups8dxfynWvxBTOyLNxWm3ll85kL
ez4CFOXKBqx5t80rIL5ox9llgN4wXRu75Fw7YdtAboY8HR1LMoVqvF2tEXkucujr
umto5sCE8BvuHwF+RLPFc4dBy5SllEgdL2hZTjVSETZmVnRgYAuSX/GSti6IkD86
u4YQCEMFLelf3uIpayX8fdp67rWehVTTvGu23YMbZMDyiy7pJJQbcXM6O0rlhW1j
LNzKcgrg8NldoN3W+fESyf2e6Y9kSMyDSzbNFq5GuPcSUwIHDfYAIzIkdnonQk7G
Lrw19Qirp4/5qZ5QWSJXH+HxCA7eTjUadxaQdSnycp0rv3KNieyKB7ktmxBlGPC8
uLWRJwwBdk6d2Jkt2f/uyIUN01F/Zh8/ZoFj0pZzluVPdO4sNoBgov6QUmnXxlup
hlj1nwNGQhkld+E9191m4Qy8aG7l/yZe3YgCstOa6Kcv3ERmfKj5929ApWfJ9CQh
QZqducYo5aVUYDr5J2g/p1TJ8tQF097Z6xRc+hTNjh0s4scD0EJjoS4pris56eZ9
u0WbacYQqI2/BG5I3qVcEq9ma8cstb1OXz8HBVaolKqCgsxgV10mBHPFKoHxz0TI
DsatQk8S9rrAD4bgQslwZ8x/chxvU5tbNUFVD1LhEtclCMaPrSqr3zx4XShcyDT7
dQaHilV3TsdAFmhQZd+mbBrY5/6geBlkagI+cTYcOdbXEmIA3PBk67pbCteIzHzv
ydROfDE6Q/k7/Kg3GeDGzYfRhUHaXF0xiLDcFbPYkD1mqPd03sgpMD2hx/zeVMo8
HoDkoyR8Yw4/NPDsnwqmZVA6Z3VMlQYKg8KmM0NCpLcJikMtIYGdHigY9zKhJvdf
wv6VaJTGILv7YzISzY+sb3HPnO0AF1m7pRn3D6VAVug+u7SPCqP6AspA9h6PuSAq
MrwCab+pB+jSKBeBQIrLkMj5FDmeKJ2cC2FerSo1p/96QhABT4pJxjvWJz5gqIvX
HKGnFexnTuanjd/gNpb1wBniS0n7+zhbDVb+/o0lmKm8TmczKN138thXe9xVDYrO
fh//1Edqytx0F3pvtip5zMOko+RyJV7a+SLlmaek8X1Fh3Wqb/F0FNKQICj4tAps
7Um+A6UKcU4xU4KzBZeTBMcvakXna0MdMc/daXV6mfzpEhdw/OJYpk8+1mi8lH6o
/uxJJ+Pgmik4+o4xtwR5jutIogw+BJMSBAErVRNd6kfG5QQ67zFPGHMqxX0JLAc8
pZwlnQ2Ha1P1jK0/njPaAVOjT20Z/WqKb0wFUzucTvkBcd0hkFSQcITi3DPusp8W
NI0NnOYqPCp9nX/hoDC5PAU9rLwIMGEEmIte7eYWyvdruyEQb9Y2iBXN7lGRG2jy
RrAUoXYO+n9kMPteF38X/3Y2Zlpb4WVtP+ngnmD4H/dbBn1bdvvxvhddTGhkaUhz
29xeSpobTUAc8aQU6jMD7a+aYhLzCKq/B0SEqDTCgPqMJhMi6FzqdnLctMAjXdIq
ll6N9OFeOjti2GHoNNu2jmI7pCwXgD/uPnYkDwTHv9P1gVzBbHjrr2yd45pK1e2J
AicgkrGNx4izVZzjMqIQjaX5/kGqQKRmHVStQ5OJAW9yyMrUeQ3aa9l3K6TOseRM
yH1+JDIm4q0yiK7oLxjpHoeJvDtZ0569Fb91jnDRXpSq/g2EZ/HgP76VWJSTNHQg
RUEuNqDpjmG0vNUw8FqaEJlulUtyDtnjl0+zCXFkXz0WXkaTIPTY0m+facHu+0Ep
cGDectvwTUWNkiwqEqPyYdSvvoELhs7IMBdQ11hQIjCpztbCKi3bdbhDjjzHih9V
YuMoRQ2Wu27An+Xyl+Q16XxN31bs3ZggjepqENEy3/AOdU+yVlFFpdVYAKtt84tT
+sKKg+eKHR01ikdmy1GNBWTGBufTb5yf7pJ4oJcKbTrkPdMwVKqRL+WZLzxoqUmW
ZAZ8JF8h1JQE9LpnvTwSDEJIVLfdJpmYx55n4YZfr2O16/YiLOXLRwrdjLISaZ3k
ohBU4juxqFCcQK8Pj0oObQYKxrx6z9g2GVMUBceZBpLbD2yGE4Ior27EWFoT5S1G
NWyCtUYqAm3bh7pguDSRCjAFGY5c+0DFWk85/ShDXkVE241xQvZ2FqQhLzDNKouJ
WAqZZG1GU4vHNbI50lors2RcsyfVTqwv+cAtPACVlRayUn9Hu8+HwxhhfL0lKV1X
xwGcGh5XBuEfd5nmCz/4vKYHe6YaQXxlBTP06KkI3LCbEL7pPLu5fBLM+xfCTASu
5VJYGQ9s+9QkQQqwoLtCUEX48wRbma6aJ/dO0ztfW3Zj+pOTzclp53A5RqgFdsLR
C9ioulALzNIXxU08EVe7ARyr4nvcftH/fpNWY9Kcf54GnMaagc6FZvWfIJ+v2+Ys
IQGJkHyTO4sSTnJX/lEZndxuUjvjN5O6Q+iGsyK0BCoya9Q6IQPTNOYY3ONfj6dw
cmaVbfw2XZOwIEK2nFNmX+zMbBvXYMSWxfputlAuK3gIkP1zdoCAnjDi76E1ZUwC
x9DjDUC1VoCOMNSVcgHB3KeEmBagZUz5YkhPSnV5HMjasNyUWwMbalrQJA/AWOze
KrJxPytwMi6b1J30eUNXcfkZVsPwlhWwsW8IiKikgwKwCe+73WVzidsiKBtMdWhd
Q7kIwD0BMGO+K4qfvsqwysvxqoUjzaNudTxoflGujZzSSp4Qn2Bu5Dpbx+IyPbqX
+9FbBAW/qIy5t47jHXjgj1uExETgbD/KcVppllpkwD6Kb8LoM7xjt+SSJ7/U+Ohl
YFDmrceH/BazuZsPhBgT7QPeskWhHJbk7nCcK3zP9YPctuVWJFnsCqneFuPGfGI4
68SJg5q9M0jnZEiiWudF4OgY+dm0Qc87FPZGRCJvl0xUqySQwJBOGm0AQsmMnYX7
mso+p9yOlFABrl0O0o/Pq7TKRzgsdx0w+6QWC2nUy41whv0yswCI16dZLg0Lf1f2
1Pird2U/key5A0OqJpdjxkUu1FLtCoOPP+9vFMdLbfzflR6KapArsZ+3jtnTCP/Y
bZn5iiaIXZtgWU+GjUqiu7fGh9jESJ1SsiUroP23Y9GtJikjR+rYx2Pcgo4cO9nR
/Zi38ZjGJqUcEQwSZi2dNTJDafsK8A8IMQRgY110sbuhGvp0SBkuFV595lOrJAdN
YlZOBKjOPbnNJQwtLzNG4yApOf4Ot1tbNVANzkCeLs8qZd6jl7tr+toYHxVt/vDL
F9DYmqKwqi7DkG1xq8mEm2Q4Mc1xYFECtmS0BJPQ9V2OhA+M794kZcoq5XFmrIiH
6kWchzYvCg4oI28mR0b/6U/TfLyZTgEBSPqHQzYUtQrufZwIxi3gFz8lF9ziRHYR
vRMkrMuLBf/fwFlfjbftbjtJ+T4sOqZNcZ3wukF/Kcb/O5ITAPuKRIsp752WsJS7
D6BU4NDkk3VpvjXlVO0XCT6XqpIM0rLpVss3wNw5jdFAMPjMmiBuWjh87fr2kP6D
XQFKq7gVPsAAqS4nA0GgAtQijFwRCHR+P53Evz3eZUtLq4lN18o2MPLSNA7aq0oU
mpW7TAzkwMTR0O+XG7iLHf5izNsxIQtH9yaeYMAOReJpnmueaOPo/UtnWU6xetlt
kyRV4TsGKBwtHi676+oKZsyYhjmRy5ChhJvMpcnD4sM4cIjeQx/PAV0WosBhGyry
0YRy/wMx591rwtD9XQKW6rNFWIbOOjFKNbSDuZkgr4Z/2OxB+05LIiHbiYyJO0ok
IL9D/VOjG2LLGSzeCWN4AkmH8vjBI3RXrjFtqbAuOJGBYbDCctjyOxJ2RBWG0tSv
z+xratK9JzSg8cGhsuvzWFMry3epoR41h5Q+B8KmWrY7a6ymLU7E328Xa8QYZAMO
BrqkQWC5kT8Eb/1wnavYo02gGXNAn8LZILCbVbkVRtieGxeHe33y9ts+ebioodOq
RBNqfh2FIlZsPz8KjPstStICx6+m2ZzjYgRFRb6WEUiyOmwdlifDH0zeYyeC+Qkn
9mgy8lvvh99IXG6kGKQczY4q7rT+ValWF/ZnrzoaLminPZ8gbLZfVTWF8ziRnoxm
WyTr9lf/USYo6mPOSa5xQ6WUhZF7NGAZOxY0bd7PEfMlyIOWhs9iegfxNAf1lylo
fnEprLa4IvpEY8tCXrkgnRTBwuzGVXYVIN7J1frBTligx8JN0uzM9iU58zcyWI4x
/Z+dpbqObRu76P8OnSlbUMi7QuFbXKtmce88AT7zSKR9HACKQwlXuI0mM+2orHnY
2Tp2E/+DyVCZ9k/T86sbV0xDEBpxMGyyW9EZK+xhKW810RXPliPEfoKNgp7AIlUs
so5QqXenshn5MagXWsVD/RHdNZl+1SPQmR3gN+n41ncBG9Ct+yro279dVD71qECW
UgZBV/VgpSCwRUuw4GmDt5KGz49C3bfsqxW8Xpbs12Am39YzBEmkHcaDKI12JVVU
n0Cfk5guu0debpbeksJCSxhcl9JD65DbPcB7HrrQtsUPDKwsBKZU44jpbuB2xheo
KHx4w1zSw7H2ElZ16mcyTWcz60L8UYW3pkALhlNaEHXEea3biHORsC2vvIX1QgLb
MEQm3Wwu+j9GCn7DMmxudBUjcNTNL+4ed6qEepn6XziXGIhs4ZHY8qne+sxa0smf
EGwuyI6E6LsbnZH8KBteGRnYSj+t0glxvQ5OEEzY9P1i0LVTw2SoLUgmW2bNQXB6
tYy3oFonMFizrOYrAqg9bagwYfcvqWNdM2IhSaecdvUG/Iy5K1CBVkkp2wn90/3S
lcsYdiS1pyPIbPFLhQok7Sq9hZKHOVNgjS8G4ngXEH8tuIUDOOgk+4QfcgU+jpT9
QvlwLuQdsixo5q3U87B9eLvAlqA4F4VO9+IU47TpJ9evktIafAIWlX00iOcrMDSI
W3nYAkrnqzbJEfmVhhuCl8kwnFLmxq/pHXO3HUhs4ZJW4Y+t7DcqXvXt7nvL8yCm
jHqtdlxcRFWa6Wox79DFT+F/Ju20tjIhEFYQGp4OO+x2392euShQ3dTfVfaeuygU
PjEOnrqHJzl3bFdrNs3M8YXdPUkl92G2zCzOQQA86KI1VX55r+1C+hVSjYhl953u
dLPef0lLIbD38u6XPBr3y9ieWYFhlSk8VspYDnA/o3VfVhQefzJiZHt8fLjDahJQ
4SVuDp+H01YEAkEhHQ66Ygi33wVqD2Jzh85Jl7NGUr20cUkTLfpg7++19/mWZJ7o
jTpHtVJEqgBMPkFJ+sxK+OLyQiRU2HTsOo2QvMIwinW7KpNoo1Di4xqG8B6yMtc+
3LG6wS9gAOdX22LNW4GtH4qFDzfcBAdRFd/L3dqdfETu3+acTMgYc+fIokyYa7AV
8B0GEYSSfD/FlWINl8wHrCv4kUlbS8XlXhMopxuNy4T9RFKJAvyMu3BCDaEn+t0c
p7K6yKSdTwfnkRsoRkRkhN5HZ6FsmReH9AmFy5SfvmFnk2i3QYimjuaOX1+y2aZZ
btnUVJWv4RUtNAeRdoNL+o3fkp1TQ/6ybxl2Y0xGlY6PZQBQtTAcmNsnO7R1dleE
YHbdoeuvmvzKzqGEo740TQaPCjjaVWpNlrQlB+ZiW4IlbTCvGJBF4vig/UjBUF3E
u+qTsxM2++YlpDayf496j+gwBWJgtBESBWUNMoO26v2HFJyQ0pgkcyWkx8zgovZm
LIx5G3E8a8zMSzReTGBH/CtVILW9kUobgLaq/CgP/3RsbQg5uLUxLkWqReg2qIZT
Tdjl7uTqpMNgIg/7t4mupNaIb9fdR47R2eXm6GGCp0qZhZn2P2eahXkBmoJWjxB1
rSsjlCwvaaLKi7OziCikm6z+xKzwgBqbdmYq1fJDPQyxrERntCo0VqmfmQDd3H5h
RLijXV/4uxSNyqpCYS7cDU4UAYW0fziHIFzMMdKLS18=
`protect END_PROTECTED