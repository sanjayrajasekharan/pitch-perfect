-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Jg7r++nmL5epzU4ZfhY6Gwn6GFpuynRyd9i3xF0b9kJ+0UbA+KWQu205XRYF6jRq
vqL+oW4R/Uxs3wH1IsoQd0BqVOQCxP4yKstW65LquKt4RcwNnPtovQfKsDt91/Gs
TBUlcUlQ5U8yBrZMrM1GZ4c6P8p++L2zUR86VTcISkY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 27994)

`protect DATA_BLOCK
2mh+OM7Qz6tLnntxnD+5AtFLjTDJxZQPgq+G4UJZmQ9wjVp3MV4QKirL6t6wxpQA
7L16GWpCoMHORI5EnyJjxCyh4kXx05Ac9lXj8qyHZc2IYnE5hvfbKTG6g/IMsUJ0
dnHc+pOhdbgPJbSSR4Utgc749I2QeJMPSD7hBIcaYVRx/eh7i/NwNVZnSCkZiS6P
kgu81YxHg7NMbqievP4/VffSGhtGnenZOZ6OkFn1rfgNUkCaVm9aWkh0Tu6Flgfi
aWsA49o9A8iEcGEMxHJpiKy5AMnO2fYocYtiEptcAj74udPJiVDqOeVoAewClh8y
592X5lssEjXsHNRjOBIipliYrbPdBLX9zdVx/gFBPhSCxlhP+nU9hT6+oLvH8GMv
6ifLsmE1t86Q5tDd0Nfl6FoRJy0/Z2mnBrl1GO0n68sQIN2r99CoKAHr6DYzaUBf
YrjhcNeiqMlIIL91u2TszXJkw+LLFRoSdnDk+bVSUkwFdncxpTl/jZhsCmy93iRe
t/4Lh+bsMBv8QOgYSEWZlsRLgLaLNnOLjfJebntTeG1btx1twIYZ+9jiMSc0j2ry
Q9r2l24UXWV7rzlTwKMCMl5aTMJH7UWNqH93CYoJp1pqJCo9A5MizfQbKy2kIXbQ
EyM174H0kcIwZwnugU7L7VduH0q/OMuqbq0Jvs+YaiseO/edZNrKp1wuYy1a37yE
/xoE1M6gC7lI9Nk3+XtA+7iRnUgeAzCF1cu7y7QBUAMLjkC9bDZmHpYzJOtuPPTI
uDncewZ3f1JwyZdS7D/g/GeTiX4Khh2dp6SeXQZGJl78zCU4yQPCggC7JHvJ3z4J
KObdY9Q6NCrfqqmHB3KOJzPvVG4yX2rFKYsmgLNjk5HnLtk5TeVIPkT8RYbnce1A
Z7AE2yaWuZvSPNKYJcYF/evmKGO9LZceWxSb47hMkGSvAG2fZNueI4e0PHTqVjdD
KgAPDwQGtQH2PKVcMKCb0eL7dDbQO+0xMESQP1p2R9ydtViAQLUnru4vElM2VPU5
XevBIiUK9r3op2xAZ5CucRd8S4e8uJ1Ykl55vU6TKrGgTZUnvQI0HcyS2TFtGb7m
Y4cdc4cs3cjiOmI7BT4I+yW5O5bC5+xCk7ra3Q2dX7k1Jgkjl/4Vz9oMnTuD6oix
ttjKUucoN3ZB856/SYNLPHE17mWJvFng3VmE3rGk0HTiYq1CI5wYlmnSpk3hOFfo
pWVvNGHwKmp3xsYq/P71UCS1bSi2/QL1su7tr65OBmjYMLYyLv8Q0czX1XZCl9sN
lIV9Db0of5LiO2kfXifxARcu6NvdG/Fto8maLGyd86Otnul47s4jt8n0O2olOatU
QzmIyJ/ToUmHstGR0QYZxAKLV7O95/zth6oiEZpMWHmYJ8f0CQChDVukA7JbXxUZ
8nxjnziLHHK6UDHallElVmGBopw0ErpDg98dEcHtK3whJQ0jgbe45LaJMrgSk+Cz
b8jxetEhXF2atTP+uDj9q1rir4u3yMvpboPqvut1qJnH7lXlS3Qv15B44YJgTr4N
lUzC5tt2HVvUBNvZLkPtGmFYU2ELZjjJCMpJfArOVvafuEWWBC4XVB74HRCAV7K7
2WC13tWfNRuXzlSp/G2o7OdWsMrzEAxID/vgOrLS0l5rq8IFWnHttqAtWwYqFDPG
jjO/9eCjUVI1BjO+dRMWWDhgyhOx8oM99xZ1PT4PW2P2o0Iux4v+QBlBmMxaGXih
97LzWRaZGbqS0elvH97l2r2daihNOgRncRcn0TTmxHQShn/X6sgYVXDdjQzOLXkw
2SGWNPUKiTE584Zen8LguZ8DZ4Svi3J5OTM8splwvw4Qu7EnalEkWMRvmAkCCQFV
6ZOGS+VwkOdYrL37LzK9Z6a0MbV69LA/hjL3VWLGENP2wwIKbZPJGbejvSHVZ44p
CCG8h9jYpSFQULWPk1k/hNvo/NFdy2J05n08pIwWwAlWCgOZqJtXuvH34tmlf92k
3YDE/7RT6+/SWLbNkflD9Cn7braZggtxfN9H65/xdtUR2Zsq405nWPGgMnj0OF89
wYIC8kp/lHPUk5Flna5rb5uP4EyDJ0rpkvwHOc5D255uUJRNy3tEm8EXE7ib+Enc
9QTF7MQNrEtBN2AhVi9dIRkkQsfaGjIqJTod26RPqmYsrHL4Wo8jxSFm3bSXLFBY
zJvOeOEzitTBOJLQiQfn9HDtX09WxXrYxo8wTtPOteMWKESy3PlP2gPMXuwp/zKT
KReDZoAbPiJ/vf2DSiTWDONYDllao1/Y7M1EYRcY+oJvB+qGnFts7TrusbEe1u/G
MslaV4HFwbbOqkNKUpEenAmVqSj6jYQTQgijdCgLnb+YHZnAIwvg9fyOd6ReIIyJ
yYyBJ/PIrIJhPpWwMznbdbcM89yuN0XErSjg5vbSI0bHAmCXDrAq1aKV9N7koh/9
knNcArZHyMHivS++/su1eA4liPUdmb4tIIUPxx8bl3RyBlO2etVXk6KvtE+NQeap
l2J8UKQCPwpmduFHyZ9eldIq55Fy+tNhsrn8jn9WXhcvwA0akRW+Qq0Zu3lGR1Yz
h6s5F/6T+34jFyP9eJHbZaiG9Fhv7EX4M7BMv2uawLb6vs+1Ff4dGA2AUkBZDULU
HTcF7jzf5v0sCkOitJM0sFcVkov8h6ktNQ1C1X5RIaphMBHP0vUqKnlwpV01456c
s+zMtktDCQNcDQ/+p3W020P6heFtFMkJpN9PaZuvKtBymRNaPvpbyVKBr7im3p56
c1vdRjhZsudmNEScSBR+y0FLqpJFigyBnGEkpKbxNXJPklqo3MlP2m1ur9v4t1MR
uCD2c8fpYjH3S9ppCa3kfXD72Eb3SIIISko3iWMn1nJw+X2wEmhiAy5TZpiUy8Ym
ox5rDGKIG1gRgWZbMHLdx0yGhTh2e25BjeCJ71eZm/4so0Tdb+NS8NeKUX0MWo35
HoOquNoczb4zrQkN+QwibpE3Byw6oW9n9yPm5flsGrKdoibUMSIThklnXkG08On6
jSDN8uGBrps8H8i2fuM1PAP/JQ1OtduWERghabBX6JG3MHiM5D4hrv3N8/yO3aAh
zKg8n6hpFszlGux0tQIGRYEcFSLDtSyNp8oTU7Wfs4ZiV+jAFHdbu0i/6XbSMSbm
QHT6apEkwLlOQN6JMxhx9UA80Os53Sm2PjZ7kEvpKYobL8Nx+htUYeLn44wDeF8W
C+sxGvjQTYXdNXfhTiERanOx0yWQfjrBb8pHIu4VZnawKjfWui8ca+leEjR3icjm
DKNdIkZ1sG+KbkFGb9CnENY4XBDRXhGxQWEms5UDEUvZTzvTnBkZRXR5vyiNGULJ
04dncf4Wi3YJqP/6m5TioIlU36MOrABBR/rfFobIztbux0UkY4H1WLFqRjDieYGl
m/iQEk5FZs37kt4cdBaXPiLLN2Ll4U/iReU7cFjImnqD1TRt0zVydE6ACGqwVvfj
McLYLE56T7Woqb6XKQqPXfCV8LkKUS65nPVurMxNGDxa51NuXMMEzaNBCA7yyuw1
evLYlJufKlUKST9DGLd22fS3WMmCos09TwSmn7EQ7wjTgq7hCrUSnU1/eJoVx+kn
YiILFotxYUiKMoqmI7ZwtprKX7nm2H0A8Z9gDlPoqwq2XvAHUP/Cr2h97eZMrE93
qa0pjAUniM3boOGblcKcUb2b7nG87A5oZEKDJW0xafjaPQw9e9TDn1t3IjgAj1an
p4b2UsATrKAawCUIpBRt6/OJZxkZEBRc6C2GorXrTlzNqfS2rccobrOjAUOVhyjB
6YSxy1h3K0Z+QMgAk0WQKkIKFnsV8fZn7P81AIFO2c/qgxYV0yQXKGafbQxf5vOt
Ah44Ifj5RybPY/6WkuSHTkIJV2A+jr59zvocyqlbbjh1AARuHqAZkFNUfQsjD7zc
zhN1fraFsj3WOkm1hCZ8dakdnx+dsv4UewhnGqip1gVqA/q+zVh+WAvS8QjbnZro
IWT0CHKt1Pq6BjSXkrZpbZSsAbmMcP7SWfeYytGLfSpcor07fkmPAPzRZ/4tBvsm
6pR/uhjR3mo2qWuX65RuCssXQM2B/AaxL+n6xrUQk1CLUluUKzylYTDn5Tru6PW+
6P6IZQDTNbqq9PHn0aNPfTV2nzKjH/QArbWR2G6gtRrYDggXRWIuB9eplyIQ5DKG
TOtuxw9nA/ar2dYBdC0cdhD4DQvqlmVZrq1y5Ofbf7G2ihTnwtW5FuMEizkO727Q
aP/PXSgdLMmTo1ssboj2GS/xbCnbBsrv0ewlIcycxlNW3KliYoSNLY/eoqVmzhFh
JO3OzJdJm5lbtG4ksAM3gyMe6FOFDmHNV0f9qavZT/B/mYD+f21R9WmZ4RRmcgyF
vblwAj4I0yWOLqUgCPoc/os7gk8ulPZ3f4qno9xNT2XNAfLMKazoqqWTDfoIpxt1
K56cx6oYp1hALkdLmOSgV5nBPj4SajlMiEL/AJ3etMfYK55/u/vqnCzklFlUWsPW
uFzTH5yP4EwZhUA2TjCtYLB63u147eE9cjSzoldfOD056I5fC1prnnogInBxB1eh
ZXaQGXveG5si/aCmOlG0Y13gjuKvEy6uZS5K1xIfWseSn9niTs9JkXr0DHhtwgDZ
n3QhI7nkJKV4enFxE/l/U9dYkP0dW1orfSgXxfdEeiDCw/RV22NmVya5Z7SkOYZf
3m4tYwf58JguYUqs7e7EBJMNisWUJbnEVzLhPVk3TuICn8hnRoVxwiSaVrq0dGRw
pf1KHf99tQM6IjeVbiIQANnHK2HLwAuPzl7fVkE4nas40Otv4Y3iN/yun3p638aL
EfB3awd/FW27TrQ3cxuBXQIjEK/s/IuvHTNZDckh2RZG9gqD9iKg3AFsQJFbKUIG
m+R9m3YFVPr9dKf5B3HIVnKR6x+HGsJNVOTT/UeJJCUJuIWBhKUsmYiwT2eFb7Av
DC2MHyYK6VKJ45fL9GPzjlOlXfGSD1SYZWM98YkBPniuNWnMlk2eJyY8LT6mR09b
D3SFi3/6mlt7tWi31nBi9fu6vd+1m4vjxu5CkQoeLjQP65TfmjXqDfRRpOVqP7wB
cGAg1eKPYf/sf8laFq2+XO/XDR3KzbEnsP7+BG1QVfaffSol5f+OlOTvvDj286f9
CxCAdewqYc6+9B8PBV3TbvoSo1z3n5D/rVbUf1652ifP/I0hRbHotn998ruKN85g
Fdrh4/QwBfcXqZJ3NvkVfM+9ZWE2m4O7T6oTkE7Vtljf/cBfI7QrzHeHvG/PuJpf
XXcf5IC1YuNuVjQwPnrmEpEXeFUiHogFZVTU/0zeNI4oEjNtvLFI69nadlpWlpEb
h91++rv5ujIQQsVoVNDavMGEcV0Nxi1api0jguq9S6MUGjBMvqEQGHbp5PIFbmaV
U+E6Q8pS9dwTz7eUm5/0Ctfy17pK1P7yVWbVpbaPw2INWXH+JiZkpl5AIxhaVLhX
sBlDXKNlJVRZJB5K7abCjSE72u9S06LweDaCskVXNm4Vhe+Z9XDYCH8CckWel7ID
b132tOeO/T717YgKi5LQWHXGRVTBKufHSZJCl0NYD3Bs2AcISLACwQLm39eIDcPV
Xff2Dhj9O8yXsaHVJYn+MWJQ+f3oH+ujWB2V/uhL/XFJ7Ktxxhmhs55tocOB385u
/TKSfIxOqtQ4NqACOWKNzziY2rZZ35Fkm5DGCz1vF3wa5H/AuSVJkPZ9R81wPRxz
b0PcDT/v/jrpLK7bJde50t/hAZ6Jn+N7wcs1x2vzFXMk6fW+50yqXoX1YzMOh3g6
UPPJUlDam4Vq05ym7jPyzC7lu/UE+yEO3kLZclAO/75cHlONnQAauFmd4lhyC6Ho
tEfBzOZIMkXXIGsx7ZPHS4jOpMfOnY5yf19sSToy7a5QgGNytGb0Y9UYxX9g4Opq
AfeFCQaxI0AIu4XhZyG8Et+meVSEi1K/Zx1VxWk24pjhmJ1MqNd1QZtDbfMN/vm6
LhCatMhFBvReDZyw9M3kUx9OS+5ewIgHQ1JlEShhJShxA7VH4HjcFLJ0r6c3V0QT
TyhlrNid47xHDEMlS6qDOWydvfJQwWO+MdRMTfkkDlhMx6SqYtZFKFKzmeG+QjSk
NFeUaX0OG/5wey9Xr7lJX44K/Q+M0KtnuWNGqV7O28Hx9EtTmP1H4cgtZHf3IfxL
KSuVIRLOdSZYFBEXEfMr2Ff7XNaaObm/gUTEdTEK5F1qDl7g4oFnzSUz5eWzXzzW
dRLBm32l6MRHGvFotTvnNG/10p1PHFf6B56E5Xyoi6DAHO1+lAUQFQ3xd8QbMi4a
JM4A7h+rIVHdOg2esoJrQkf2N00VaVa0yMpO/ofTgWwe2rHLT5mwByffAYf7tUdG
1M0nqSEllAoSsOUEUhlfc3rcHtcHd8sA7OdszJcx4Eq9+BH+Xo0NRGoetj4TmveC
hzze3iMK7WF1z3Ir4NfSoFVlpE4MSoUNd6QqxNuieMA9Oh3DsaXqduXi+wdiDStH
Qf/qStqqyLwrCVZXPuECbjz6e6yv/+kSSUglztL7EmPhM1zdxMZXE20DICx9NF4s
/WqkLkoARastZLdJn+9RGMU7kvwJwi91wz5CISl6CHXjC9EPWSX2sCF9ZHcYErGI
TUKocPkR14nV6xo+utA1tmO77zN8PN7BozzUfmEsGob/LrWjm03nbVbnOmaqtmrx
ZXCsP7qMAzE3SkisybUX0i8FT85csNnPoGQp9A15j9d/lI+eVbB+TzsV+GPbNkOU
4AZH/ElgW2XLnMf+xwO3R7boCmaHFB7doGFMkWQMdP918YjPlznSdvVgNHN5qon8
3unIrpJDJvUqKkWmMwCly4tbV9wUkD3pwHks6O/bkTbRUIGgca50Say+Vpxs3Foj
fuwY+PcTdIZgSfNPgNL99zlm0jy5GV8rCxLaHnseNRUDg1i6Ab3fTKo3taZS2Jl2
qnEkpSIevm5gv5ARPlbLgc6kGtUGE5BUpEBdnWF3hFR49g+oEi+H+sXlaedylJ+h
YVPBxmRKtddXiNPChoqNN49M0FebMnwadRqxQR7QnmgWW8sBpHMkLBgTnJA6KgvN
nO4vzXBhG/QkAvnz0boaDdxsL/MAhNrbbsDIjeDlQA9dznsRRdAADJFgWikDX8Dq
N+HHkuIm73mNmwd+0xYju50m245xd/l3wPB1w2oXoV+16sSZ8fP7vdeVKqAecpW5
ESRWSCTn0R7wpwgcMv+pA3TShR3xWLQmXLGnPIBjGZ4mcZ7U3ljhlqTv3kahaEuH
7pNAgn5VtAZIhi7v84Z4mzfN/9nnmTfp3zikCxTUXUveAfztAwGzwAY5goKPUNPU
Okmc++1UWdladlUuaoRqk3F/jvvdZ/nt0JjcG4CJs30vZ6hhAJZabIVTr10/ZrMz
WQolLs0GgcNwQmd4ThwXRWF0eFfRktFnO3NFFBVyEqh2gNPGzG81sO+XExPWzeV3
CDzFvJCEBGzp6hVjZA3gxe0/uj3BxFzJWRiXDyMSUYxX47bmfQJUxqEi1NPAKW/5
iFaeu9XSEHbG+19A/xmJp7JPx9lj6Hx5UKjIL9Tzgyo+41CE//2rRFT3db9pC/pt
CaZmFoKOL4WBEjgm7LLSJiwcBzjlY4tEDiZGQHc7dJ5BuAXqBbg1Vw6YY9xruhwL
Lz+NQQc8RI9RrosbG93/8IJNWCw8f7ICNzevvMl2tQufF/zS4yYFeSzDxcCWPMV7
dnvc6VGM2UAlzL43JSZ1dWXXji/Tnu0+CaQXIWGi+eFtVNY5y0eQgWmpyKdOxy+B
oXZ0j+16xwMr1uQfCFqG3WrmyY9+0ui0z7yKzSFDfjreDDMVE+sEYSN4V2OVchiq
NuYX0quWp/U++Lg4r7KZPn/7zWdWpNarMu0PeUxj7V/e5zKxB8DMob097q07TAau
TfLvMDxnDIENq5lyadPcGSATUGtlYRwiBMp5IZhEpUzDIWrADicL3Zeb50z7oUBw
A8ZBg3UwiZ8ZupU2xmjnLul2lejygbXwGgrKzVtSZyQDbhwPHyfDnyaI7eBoLYSY
9B3aL6Q/fcZzmFy8cWBpC0nabueda+2yvrqEdMi6Ab2pqhQHtPTl+IOBKnY0Pqby
8OXU0LNQLb4U+e8WWfOy1LEGvjXaiLXRzP2qpf2OH2h5MsqcujHaYGJfqrmtfubc
+f0hTSlkZRigEIKvS/h0Ek/ohzVOBEOT8scyPqWIO2efqAB3Qf7a2IyANbk1ePQs
T4Ftjy928Kmjqt2alC0/dcGyrzbAmVTsL9V5+IGIXpLwhsNclYI64Zk+Vqx6bjcr
xjIy//50uBMCcVhECcRKRXnr/lLQMc5Ez628swsErMmIEngfLAiLVL37FMPzuxct
BdHPEmYLBxnXxfkEy5VAb0oUOF9GpVS9uqhWhCQUeqUAeJJFTo9x7T2ihinSHopO
eA5YmREAG5gFJJeQjD9+ygeQ7R4OkWH7eTFdyREV43ZUUJgqxQvCmKn4/OiPA2Qi
UoVQaoRqN6Hl0ejXfsvFQ1KSGtnYiMhHM1/Ph/nR2yRGQLpESS4ivjLwnUB9PfSy
amVPzNH2w1LpjIXUBaZCIsqKK4GhKA6Ciap6Df9qnwLCaC6GXp9yKNR7xkwkKQzM
8WNniBYPgIofFaXLU4Coy+zwRBpKHgrbP5KvM3h2982Ek6UkussZ3QubqfrCCGHc
QCNE+U1rj51XnAj/FRuil6lQuvSxhyhCxRMEDN3H419tD9UoOoe2aDcnxN0kwq+Z
Jo2sr3SCIeRFz60FT/TfEB6eJWeRxFe0sNnPCHotPc8Z00RVq8k+0/QIOXmbwP4H
/D3h5IjioMKe9vlEO/dIbI9mWwc+7jE+cy7zKw/TVowqypSwn2S3Ve2U6T497/9f
RzeDdJIzwb3Bbby7YiKpEKAHENa8VzAHZ6y//CfVFhbDVB12i+St3rHVLpXeeCPs
ccrL7pYttBGVLHySkVywOzlc0XGBnC3LdLxk55NVe/GKhA+hdfdEMH19C63M1da9
M7bwePz7tz9L8uhVsu49ACriHYeBidHdtP4Z1XAY1/rcuTrQ0uO6XZ/C6Kbye0kq
2OjZnjI746fTzRONzhnbGkqBNGLunxnT/v0pBr8T3+tYH8wMXxACCEGwpwRH2+uU
eFfXwvVWArfqj0socHIJ7E9VpS59uHrQAKA2dGLGbzlrc0tOaZVs8wOwCULc/l1p
Mtm/y6q1eGZJTSXkPhaYz1iwBt9KlFvxSi2QPg/BK7DNas3Ec24ea3WD8obh5oGa
kIsaxGIfDOJrxitcAxzMnMeAWl3bhpBIIoCUjNOQ6ezvyB8GevmtqxKycHlLPQPi
eqBqESX8oM+77BfsysPsV3bBd1LZTE40mtS0cMNMrkRhNgNhFdcUK3opqSyyA4UJ
yb0C/nEwLVLxZfTolZArlMcfOl2QwUVhIDHhUD8l9Hn17sEXHm3YoecinjgEvg1L
VYjB/tHqZq4rRX0V1IRSGqtLgFJC6ziud5JWmorb39Ef9FapJX3n3B55RtY9GhIF
wVvePkgcsPWft7f3yx6eOmOySYhWHwl3dJWJ/JN4VGm3SSWwkLZm8JTWGVpneJa/
dM3yzjbjecZR6uDIjVREYPMWysYLQiITVHUi684RQ2bDDGR4I5a+yD0C2f2j5zAa
BB+Hmm9Nva5q4UfJ1Nc/rrabshmZA9rYPfZJP5wSvXTGUVIDePtERTMR/wQP6zTL
652AQwVfqoxRu7wvNWPZxceAiIpHWKpyOpRYY49+iX/dOg2Ja4hy4DGLGbXvGfhy
Mp2yW6b3h/nK/ZEDG2P3ldW9uY6Pf+evWY0RcpNK1ljaa6ypjqyMfVQx3OWMyxcz
DmIQ7fyjDQrcGhMQiCVwBZMlrMpMYYgNo5V0w2k67ojhRAsJUgHxHG4/7NgzUj3o
bJK0iph3riodAiqC8qGzjnyQVOosVZix2W44dhjTCaePW2h6y7USK0SKMYzj32Ah
7lFiCaHaLhoalxMuWAlU6jyAz8GaFC9/gtc1nKn8bkQfiOcrYS08E4pP/1GQX+4t
oGI1/P+MrgQFMUNoo1C5L9xrQp3lZLqv9LqNqVFZgyjNvOUvaa7Bt39vSjL21Ghw
wITXE0Wn4Izz5+8RtqquXjza4dhuOw5g8ou/AwtOoLcqsMVmOuSHPotA2u4w+1IM
fLz1ZHwaBCBnutpEe387DAa8R4B3LlYCp2YVfgaxPGsnWGOrpG1L9DRrhBbBEgVt
vPXXqfMhZUFd6nB7Mxhck7KyEjX6J9PxKVZ/eNF+WMywg50qAPoh2/3xXace4ggZ
gKF7b5g6rPXLKwv4Yfbqqep8BAVU3ob8n9lAmRU2fM9x18TgZoVSEN6Zv9xSRSk0
DehUwwfLJ8ov1p2BZBKtUj24lPXReg+ijHhLk2SObuNpzmJEnaf5skv4Sl8rW9vt
8D/bEcseIWaaQYa+q98rTjfG/aTiu2rtxaQZ8xsYjuLqCjuQwJWWK9BfDuSsZNCj
AMjDguImmf62MtHep1ziBOvjMQpNOYUVnJ7d7/04V1pS9UN/b7+xJDzOOLy5koID
5kEEIJJ5gApoElsl5BPd7BprGuedK+bNJPgjpbTQGpVGRtx7lWN+NZ3DSpM9d8xe
7A/uVooYg1GYoDmcvNu3k5MF781+7qU+B9wdq6b/CbiZmGg/uJQcjIIjOSGoHLKE
6doJmRoM67OCttLYDmcy6UQZkeZyN5fzWE6XoREBc3fGSAEjpSp3Tib6yzaTvVOQ
jkeyhlX2XoffZIOtUB8Rhfmzl+ndpEZxflQeIxsc6TWWsW4lBTQBtZzU7lFk4HO7
avdHlqP0v2gk/WtWK5EbN2miCLSvpiRzNDfTz0D7CLUzBSJv4h0S5N+XUCAA9Gvw
v4L6fGmbZkbpxZtJRjTHRrZ6CqGdAvmSKI1i24t1IUgONbpGAqrzbpw603+pTA6X
cxNSz6fF/ii0Qe8OyFTUkV57jGhfAIppao37iHckffPQIOPmTvYcQyOpNFWelyYj
uibqybDW2oJ8oSqc3wJvbGTS5hbNCbrIEY0tqglwwELRqoMVpwJZel42Byuffkq0
tSgFkH58NFIvsKrbLV5hnCk860OMNoWlCRrEm11NK7MuvA0wu6Yazt8Tu1u0npo+
XpifP80xGLY+mAT5oJhNDnBHlL9u0jMotX/iyC8abs1Pn7BLyTl7+OwnjHrEaLG8
HqznWofyscHMx6T1ygBBsWOQAx2q/9qIY/sih6jI+e7gu2oWh+GOp8nXWpl6tYi7
4usFNIStEmDgbn8FkGDxUFcJl0nxU1SSy71pxznX9op5StvcyQf74LwsTid/4EGg
PX5cQcKkI8b/rIo6u0Uu/EPjtJHHm0nSvXOi6AamSSS1ODkV+nEl/TJem4ZXhZDA
6+uYDCJgQoff571CHuCF4ceSejl1mFwlUNv72N1jYVu9HqJG5EdZz6oQwJ8u+aHh
hzJnFW9QZpb631/xwKDUEIhkl2DQpoedrNb0K50qc9CoChnRV5O2lFppG8XXku1Q
AZJ5Nntq22fXzeVFtUVQr3069kkHWKknmfLUwQC4mxfM2PSJtel248Uev+1XYdgS
t9/GuNRvse/w1j77yimgP0INpJwndRyyNY6Jivj8Bb61mPoMr6jyPEY8uoAG8oxy
h8u4xImAK7bqqemiXl6HFPzB7zka++pg92M8I734HhQEDGmpC+JtlVsP1o8uVopl
3zZAZ2ptgMPQmFxxnGhJjBZcd9LcFnm2HxlEk5LuUQub+91TSLud/xpohxCMMU0y
QcpP/1+OMfT2gJijgz+R44Y+adZHZHkHQ1iu6bcNigVdq38s5IMc4+CZ3/5gie0q
HB1EP9a9zexA/6UF1Ji4iP6yK6EXwl1MgA+0/YgGQSpH5SPO1rLzAFYWgYo0xbGZ
mR+c1anhQ7kYkY//ZPXSttWEGvXFWyRTW2mkBE6Xc5HCRSQtrYLQthhTAZwd//b5
eyZh0w91qLXqO57U+UCAD52LwCBWR4Ur1QrFz/2pvBsUnPWo0DetXM6/CYeOxzlm
8PeeRZvfk6UUjZUUewXl7+KVnbZJbs4mHLTb75TmEkIE72nI9H0X0pAyyZw43wOP
jZU2E0O5FINctmI9pay4DIqeoyVUtgXSm0HbECWTHV9ncYGyILwN1vSKbxGIR5FY
3n7/d3r5bWPaI8a+1zA/QQy892ZzkF7+JbYs4JU8PamszASUSDPFcsJlAd4GkRGk
X/4UwfUkoWbXwo8mr8C9hhSSPR8M3h9TExKCKbUSIPprJq3X2F+ImVOlsXN8ojzU
cajQvfLGfVq9uFlJMiN/snObD2YpbcCHO7GTsxV1Orcy98iKZWWGFKQZHb5Q3HsR
v8IKVj+/MCbgQGGH9Kwv9lIT9LNfL6DcDbKG6gZrX1uxc9xIanW0SC78Bze9C8XD
Oubxhl1aF0QmzyQy3AnUc9q8pv4UbyCPTk73Br4beQqxqOzPY0xIH3YwL6bVslhd
IAPwc4eJVX4pRBi918aRdRKzto9YQEWg8eBp3LveToKZAB1fYlzvTd4ltBPm6bKd
PzWQpflid7mV7jSIciQEx/Ber119MgVyw5xoKKrtxiwvPBqOm1G6il5CyzFibT6E
tXF1X2jlIBVpwiYG0fMUl9EUmE5muT3RsVDoVc8A4v6aeE1jKYMFykFNYLVo6OSw
96EY7jpnWglhvrhmA7RnbQGsVLrmaCReeQBOXti6u1c+5HPCnM6PyZXB637v5D8O
H+RM6+LJSv8H7nsnPFbG4K/iELYdI8XwwmTFXyOmDtwQWOqWlbhTkFcsjp3ZdZ9t
8ZZwcWdy4NzeB2ITQoN62cKOG41shJBpcukOalDF31N8s6AqRKQ2GS7d3F42+fU6
XgPSWpyhJ8eEJtdnpGQA0CwBsMsbFHnrKf5yMb6/Ycpbprplab/VKr6LfH/cs4ux
DS8Unr1p9CKGcOUKgBYhYbPsN4ocBGqb3ZSMhsfkS4g00ad0tE8VDfQJbwmSuk6O
ChkJqYGI+06gCLHXk1Tz9Co1ashzj+PLhN00m4/vUTJs1v0W4Ot0tLs09k3Z/RhW
+jy30elf0QMZSGxLex9ZzOlpI0Kuhm+Zolwy0M5wd+lISRX+0D/D15fB97NndXAe
gZXigztnD00TULyMPoapFA3EYFGXBcBmZbLjwYheBv2U28vb8oVtl6f4GQ1OkWEr
6Bk5g+fB1cY4rgHVhxIESYTNDShMfaRovHKuWOoNw/oLOjM6aOZeNu8iM6hg9R64
Mr0nKsyjw1G6ygH3xzuPu2x9MY43z7MQ0e77zgr84kPm9PV56VImdWjHJK67YLdP
EoFUfJTfH03MDOhrIWIGDpXpN1/WgMl5W/PsbxHNagqy2qXabxKYwmEcApP6rw5T
sSd2FpD9uYc96cGXKz6P2QkQ87MhcCMi7iw1FPXeUkYWv4VM7Qe7Pzvw66IKICDa
k9JSrJgcoRHDZUmLY1rC/rad4LdL3jzitLBgt1RgmmKvy59k7oZyLK1t+ugmSIZi
/Bd8H0Zl0CRR5+HxT2pjXz9XF9iw9+86GJPsgvCQ8Lww07m4aQYsjs78t2HeHnRX
te6xaoVv9Q1w4asfZHwmLpH+D3vvoXJZ54pVdUAb4hm8E7yI8jYoUaoKgkQ02PTF
O5j4aJYs1hHdg5+L127AikjJhs3GJm7J3bQHsVtIjGbzo5vXCZa8Dhp5i3jd3iFA
hhs66kgkdeao27EsTUptfk0opG+7MGqSpJG+zC0uOMP7bt9/WQHukyoGZ0mmTj96
eWKg4gCFjAVX1pu/BODPUFqUIj+kR6T1oZLHT1/L+lD+GkEVwJH7lJ7nR+rYrbHs
ua2CvoMAGyg3XPK59P8wXgWYfHmbg22ujPGmVwrjHvFLa8OzapJAuConZHJlqcxw
qOL7ivyerXDcmo8rUvaycsIZdG2kBQQqfWSaWGYf4NvLCXRZzDQg2ccqwFH3h6Qy
dzqiYmyr4FQvEQZzbM9ROqBhCt1iHJQfrlYpkBuDzN83cE+usL7eaXoYQTI1VjQj
YoH1+1s7ZsPRyxso531qLh5317VWZL8gZcgWN9hzvcI0IriZ4JsTbjt/ubNfysYW
QMJsHxK+i1vUjiz0nIr0adRXV1HMBpcq8DR0hnxcYw7i9Nyd3lIq8QqIFsFgkDnI
WvkXh++GVXmhECZkk/mTKq8BUsXuczlMX6RgNHB4HBx9vXv1D19jGjX9x6lRoE1F
2dyzCjzil+slsZOrqZIwY8H5ZJP5tKeqhxHA5/kYuh19oz2jBjdKQI6q+0+ZrISI
Vg84Z22eNUn2komatzeiKRYkrB3hoR52uXtTqFaVq8KbASBF+5tMn80t7XG7k1ig
SgzMmznuYrYLIfPk+aC+x4bxc3KcfxSPhWOIqCbdjCdraut5m2VbeAuX6pH7VkOy
EzTUGveAJF4wOQkdijUOrpExCzDnVRS7vv/DAwCcotTCw5RUIk9DjS9Kx/Eylmnt
SmG+koztiXZPdzAVo7QiF0woFntsWSvE9viMY7dpMQQupmrA6/6x1QEgbxiIaXnO
xhHc8O9/Q7oBLy3yaB3oSzyrTuKkVSKVRWpN0/lg01ylJ8ei1ehC4fUFNcT0OT22
lqsTxC+FnnafyTavuXqvwL4RCe0GOIftK5MeAsvtD9HDT2EmxBK9PJukqGHVCMYR
bYt4A6E8jqXYPvjIkTZJy8Gplb6wxQ0/pAgLXvnIgpbRDUF0HfqvOLvDl1smFrnn
VsLszjXOtkNcwm+goU1vqKfSm6d/Lr4fN15RSfOXI+FcdyENSTMCihc8C1mNoWhe
SO9nM2swac7FSWkk9Lf1A9bgkmAxqRblwpePOXNo/xJaQOjJQ0j373OL2UV18clQ
hZ2SLf6bsPL51VLo+cdg/8Wj9H5JLqvLWwKj+hSN9z/3eSOGu1ziuIiQvlOamGuC
P1LqbtkN/Y5TzRLW2igM23DQ931J+nMweQc30in0mvjWJZYtk8n1RVVkWxOEC/GJ
lw7yYxmQmygEmLpKAOf3HGGo5gqWUD9mAqJ93tzqEmhtU++frewynUDvxRbDAzxQ
H2XbV3ov/QC7lQ9sJetM8LFuDZqy9xEfE2aHyMbxv2yFzWLwNVaHja6LJ+Qwm+PR
9w6HIse72MPUQKAvDcDpBu6YfKqXZD5sVTJY7xsMQCNdk3RCHWEOcNH3/2rm0Qgs
ederTM8QCSPih7NCN/aOpvGgB7DmEBHmMxCVl/un8gdT3bPvBlCk1ktJHhgPczE5
UNCKR34e0ftRsOv5AD2wVQlLXIjzclXjvjwYSdsMonIivwQKYZX/m1ABt1v65Nrx
ZhT08PcxrqUALbz5KbcZ5wmQA1RV1kKpjgXHlhRNR3U5eadtq7hH/uYQ+QZ82j/7
8dVioMPvn9iuTpQs0dZY1094xFhozUSTTMH9c3BnIlq84mMa4GNeMmYZZfGLtuML
FI4FC6KiHY/2sB/YzOqmDQUflqi8yeb2vtPY4AwYQss8jVNfx8H90Y5asmNqVUJH
oNPKzXIosXwEFxI3zRWKuZlRH3lZ6XfjFCCeLoCW4B8EglWmtyo6mVbjFnRZQCpS
vDE9nap+/WlOm1yhE3vq2sQWPoIrsogVoypfh/NEHOFjbPcLStGRoUT5QTuUOxe2
b+3ADS8M0m1QRSCepZZsP/2MBE9kpQFAbvNeue5hDAtGxZcKWH4TI1mDV2pZzYzL
WqcaG9HlWbp+yN3AposWZ0xIrQuCfJZyZoJv59u4vZrAZ6zkfT9aINcCPc3AJPxl
AWyGnb+UjgZ8a1jb4rAsZAysCIbZwTnVOKIJmG0gJZllP5q8aokiiFmPffbwtnSq
VWZenvoxvjSoHA4RZqAOw5ydDHrRTg1K/qUw66ZizrMuf4dlqY5UZhHAshDxHsHl
DeW9VYUca4TCXqKmSMX2g+D1JFkc1fHw3J3Mcb83ladnQEmxi874uo7G1iAP3jSb
xp234+BfaReP7IMJP2OI+Max0QxzmKpA/lx0c74/QaXZlXR6d+NHuwfM1Ynq1bGa
+3NXKzS9AZR7yhQO8q9ULiOg5Xj1XlwA642eJjEpEuXsc3JK3TDC8teX8pLBcKfr
khozBNg38rIMBvxaKIDWyj5DjqT0qQRhd7X3VztpV4E/dCYHxIZ/SDta0+8+N75w
pQ0ovv9rBSTR3t97BcDLdEzQpLiAcWE36U+duBCp3j6j9gu9oIqIAZh/p23GxiRp
avoHK4hHaTCQJnvmjIPZa7npg8ZiXZ+Q1/EQiKOje+Un6J0xDBl3LHaRGNwYf+rC
0MXQJcnllUNgQlxy7Yo1wCFY88clWNr8lbEEEYc7+HsFz9+X+8TvFKpqnJVeqGmn
EC6FsIdSBo2t5t08neVoFgcWD/lGH+rHzfGdcBmYzZ3BAWfqMHyHZKuSpALZo2Nn
oHz9P4iZcL55alb/m5DgoLn/rxGAUu5lOSQ/gp9WjaAaZ3mF+6LI5VXES93+Nhzw
ODubqRB863GRNpRAYQEND8NWYqr6aP4CRLuudMDi7waoLvelNem3KDHQYsYaaEkG
GK+hQxgQSTRRbt67381v/saAurdNX3AevWsQNdG14iZ0+DhxvdLyzGM1p3jqGDaY
jzAW44HxIfz542OMq+uWI0PkDvOy1omH+nR6Ca7dm0IlzSx/hzH6s4lun+iTUMz9
wOv/B6IDFXtQqlQ1/U9vwu9EXUFrPm63iYJ91d/qgjA4ymCWo1dSBkpERRHrxkjD
RVAvbjtYhM4ZHpN3w73Katv4h/nOstwCZuVYSiOR4uOUEoRKehIeRK2UDCH6r1Hz
fjc97JsVL3FyiF9S1J6ICkqGpJEFXZl+47paCVmFBMayR3fKPXDJ16+kKprDUE7j
JNzkl2Pte4DlL1OEN6X/7EOVqYbBYeOXE7eD/nJtxjJ3S0UXacnO7h359UDAVKHv
mObrjxWLcR/BwVAw542J/48cOeaVNKX6ww5vN3eucP340SNr9Nw5HyE9lBxqsug0
Gb5Dpx9/c/gtiNwUN8FE6Ce30v17rYS2OX/ZPffrtbMxfQl2gjCR3EKvaXmAMrmm
P+d/hLLV61CxF3epZ/58gk8t8XJyMQ8hWvkPU9V2sEZH5Er8ST/0DsT3Ua95F9cf
LZsOgbwQGnIZfZEeolQCEh4KLStiWRFBwtjMUcEq/DtnavMQMeIG6pmkihzFlmcz
EZya5maczyBDWPwWWuLi8yk3lAcioccTHUxXpx5HDtU5UMLr82wq6qgtBbVQ711I
+Ww90SzVGI15i0SRRIa5ILI2CQsHlB06eWcRktp/H+S9tZOpCJ9GWqOimD6H0jqE
C4a4qYn16R8+YIrq1N5omcnW6rYhBNg3lNdkzqeEVSYe4WME/vmRX2P5bD2iWuS/
3gOYXZUAoYxaB0H4L4wIQ2+AxklqXJivigdHPYf+An7the6/13BDkFrw7d9vSDRY
56sizuFq/FEJZs/2AxcN3sm+YEWMkzM+Ttj7wO+7B5q6uHXhaD0yjVrewosaqnAT
q06VF9UiLC66aagnYgAgxaul4iQtyQY29F0Z97YI8yjtB6gWmzO0Aj4JZGx+ZPCv
S6ZJIDvoj6uEhS0WS4hGNjPKEXFXBTOBD6iN2DHn9dICl4CqldHNl766HjGGd6CV
2e2lWXicZVHebShiK0tabTT/+xl2phhP4IFIJ1F9vaA+mNqvfpzpcp8vT4wqH8KC
Odl2B1k7JDpFLSWtnJLYyD/3t8+9BWgzZrDSgGWJMEzoINnzrgmb6MH8D2FvG5tJ
pDxyJI70zuu5c4jN6JQ2Sfxuu+amCcmcsYGNT4iGidbjkd5RHgY3N7PyZNJXxXHK
btNbsAvlj9JILUYpv6l4mS9FxToS3b6nTCIYcrS4/sQRsiISHX3fzdVKwvGBbvNK
AnDW3CZryxJuV0C2F/AxNjsiyOu0KS9vtPGVi+iNS5gjgqHQBTx94Nn3c6nPAyfi
k0gs2/sMvRAeQkAkCysmccp2bnflKLrKsOp7dS6kQQ2y8aTMkaVwj0lWsRfSk/Az
/e2frwgowHauYa2UtZ3mK/shCUDZ9IsXdBPRcPed0hqhbD47/UzuQZTI/X9BzGLH
4zRrMbusFo60GiWe7MHGCzPuH9F0lbSpPK86vANtdejfp8xFDrWgxBSEcVNiA7QQ
EOCMnRYfNBxpLK33Iq9qKe6aXI6C0o89mCLLrjZJHZjy/+eVNPi5Uh+in5ETDyQJ
h7IQPG7zBtBJMksSKp9xBOmnMaO9guw9YyxqIUymdoTSBjFKR8iW1BhrtchncV7E
VMLg34wsaijUR1xr1vMKIcoKJ9DPG/pQgqpjjmWCqMOZ08d+cmMP91CGROA1blKn
Tdx+dmrlconsdkdlx5hhUW2S1T3TBdIERwE7TIzHqSDdI4NchP6HQ4KS/jxS587S
lB+PdeuX4TrQ6zc+ZTH7sapOCI/7iWPkPZTRN7i9VO3nCqYAJwcqonQaranYnKYg
Y2QICaqNbgyqFaFFdgFpQc4i/rWL9v+VIzIcx10N1bZtwR0NxlgJlPVCk20RarSX
tSBFf37iFnffJZ4/U0DCl3lRCU9x/KPL24qTkDG9YDaYESdRi013yUgiVXmuRHl8
40VjWf2nkUatPr0A6B5onLqElEbuZZ8WyT0bOEwhJjVaYRtvhaxfIRtv+RqDFbbD
lcqJabbDS7fgG5usZqVahHSBEJhj+NhkmL697tr+rXeixMpru+xdpitpUyOey/U0
E8X/rgL9tnk3k0SLiC0uoBgHKYEIY7TC9d3JEyQujzwocP+h0/t2QjIzAkBCwmlG
K5UCSFiov+U6NGt4uBuFEGPLYEpaN+PrizwRMFsALFDl2J/Kf0fpVO/HcMwkoDPg
PuyM1m90vD2gdTOmgM38/S9NhbAR+MmBeNmIVvnZRN+UNwxVRAyQWb7fO9C0orYF
D09jTak/g1Rly+2GGOByhy4BX+om7gG5X4Ja1wrk28w61XBXiWI3QeSgp6RmRrBp
d6I2H/6UXP8b2VlNY6jnjfLfScWzB/0bRmjAXZD3CHGQH1Hn3zO/WNrC2RIchomx
jQkBOKF+5b3Hf60qklFxM8uhc5Q+04r/6xfUt+kU+POc6mTzRtpB0McrnbfiiLr6
aBi0YQ9NbMNRVY6d0ZPzfSjN28oy2Hp4u325TL+zCtUDm5bvOdxUFtsoztLiM48n
O0W4z2DvvJQMGm1TGWmFYUkj4lguHvc1YIxaRzC94gF13oczhZmoLtQ5PDWasj1d
/pCsPPbs1kFQVVomtnnuS8lBKtvG/OlS2R3kWLidVfiOfuj3gD2os6oZa1gT8pDU
roBeqdSvs+6OFG3yO9/i19LLzD09g4871Jr+K6Cjqk/unMNgCkV7qUCv/8kd2+Py
fyD0J1h3sNYeBYOTz14vC2LdaKIL9vjiDZpf5EQniiYqnxvF2m9wAOV3Te3c7DHc
gz3S1SgY0qivzeUCZGnjy84Qhsg5q9ZZriSO181kYfF8nl+aQUzG0plGvJOTFZuG
tVmYzBdg0UiVj1Jldc06RCaiI0pqtBTS7bFvluJxzebE/vwevBpG+mhM2s2PRhQO
5qHV3/hJDXTYTaMQzsHrmSU3k6DO556gIn+I1bXL6Tx++GS/V7j4VyMupLDVF7AT
QRHfZq6oVRTTplh01Z9W6qW2jlfPWvyHER6lrRn1pyJchG21S7vLfGI7M6l35x/J
Q4hdwgS2zZ32ti1aOdRqkCewuQZBS5o8HyfBku/1gl6XlvkT9f97itT7lGXYmxpZ
w0ZKAYz/3lN9McezA3ocemM5dlkXGC5DZRQw18y23ZXetur1tDmwjsXt5lsWZ4mj
O5V1FLEwTR0+WvZhXWBeNMY3Kmo194lXH+drcBkLxnR18NEpN5xfHYb6MiMYLGXx
DVO/PV69C67hHtIYTMxNNvyL1oyEHpEZz8ss2m6Vn1JUbxnkU+vh4UsKACvYARvD
b8hg78zKuvEBUkP/+PQeQI0Esngc3B5blAI4igmxtTbYVER0KeCtXeMjeGfhicWp
3C//THC2OuyJRVoe5Hm+znasU5bb9iUhxmGzdhF2QI5Q7HCSX9+cJQOH7Gg9P3NZ
7kY27tahu0/4IacAdL65ubPC20fiT3SIODaj/htx+t0pmst2kk7qawz5PGlbqcWs
qssgKrN/x8e118fgpN3ojsaoXSVZFhT95nwPwjCSwIPbdErFmOAvUYscQnMLWQbF
KUuPQ39M3XoiFET9lrTZ/OJjdPGLdtcpwrADF8u/4o/SGb4+GqJ8UGGdj4Eneslc
DrdOyY1MRr89xvSTpj0kgB0+fkiA1uEWmeYHoJonWXvVfFRgverbM4Pj4qNJopJr
ANoOf1r3cTbdVif5a3cfYomO6D5rQ3DtvXJTMNcQpIIDkjTl0SXCTqAiW2HO+j44
MT2gvJxMnahZzwuoEdTg4Un2xCyjZ435Un9K3HFHpSF0NjggQ49w5LSQaXv+GUk7
Hq8OuPtZsMyTiPc9v5sAsaWY8YLcM9kxYZJC87p4fvhz+AifeTxL3BldENGYy0X9
URd8sfN7DTmiC0FPr+xHgqDJe9un/jj8piQZ4ns5QLNy6ogxq6qY5WArG3+S93iP
vm1b4AdnEvUFFWXwE7060iNgNOPrWd3W9YKCKQgPjxpiNOC/SAaPkFl8lg3FS7AB
irDXZypOMwHZ9lzL2g3/aP/d9PG2rOmCbR8kg6CseYtSkwQGbyXx7djqFfPAazEr
+sJRzS39abYrv5KtRtCtONULbF2kNSzGOU9O/ZnvFVZ2RHjmHAiZ5nqafOpRNIbv
JJJ39j1uR/WC/OPzX6wWD9H+jw0NLurWhdTemAmrH9/uo2vAjQ1SYE2L6UZ664lZ
NDKUbH0/p+mpzg3xufzUUHwHjIiwUUlsdUNNy9rWezEIWUXvZnAt1sIhiX6nFtDw
2A9PDsU+/Nv27LHBLcRYtmU/Zu3HtSaHwjpb6/FynmLRa8YSeCwDKpR1OvkZzt2F
KWq9/sEyuVUIIcXLDBdmC3tEsSIvnd5XPzV4XccqPWQjVI2vzy+3GAcEcwertJLI
t7D9doyUxW7ypUWGlD6YRtbDOWUldg/Tf9PPTKkpZWvyJlqm/DJDbIg+x1odrjrL
IiJHo76EsfWhPsTAHNrY2H89Ph26bZ28ysajYbfDY/S/3BzgdKn6LSPU3glkcdS0
MRM6zFbTMEKWEfn2/+EV8Xj/XUlSJdydNKfOT4qie0DfaZ49K1nyt1XaYLIs5Ixs
oQxV7wX4aU1ayFWeECe3EmzLBpolFC58jxZiFKmpC8W54Gajf04SLnlaTkGCJseq
fpzwld8YZGO0ZHrO0IRUzdbNQs0QUBVUSosWx5XLtNxGfY8YTHPfminyoISZZsDe
+kwN6c1WbqDJKNE0eg8kTpSFls2y84oC4WJLrZfJu82lBssSL1Dww1mYqhQoLmIp
2ea6hrYSdgpN52R2C9sZrthUYxeHHh1r2n6VwPQ8AnN2Js5E4r+/o+uTqgh24Oeu
/U/x0q0ZXEu0fpnWnx8TDDjUeoF9EY2eAPSOa1W//k9AynAOuEhny8sddc8sN7Rh
h615FaCuljWg+v8CgLo7jVMVrf8kZ12WFxT/MtlQ0kV/+SAEeJI8FcRGa6XBcA7Z
djaBJgA0n3zyrQjhcwmJNTEXCFowKMxOx2Kc+SCpEnmrlf5uvihDDPv7uP4yRPnG
d/Pzts4w6SiyRlWzEnZcLuQsVbwvEYkSoozEKjV+FvBoQh/zdZNrH1/XX9ty9JEf
sxXTHolAiVoC15x5FQrLcbHFEge+m+lN4UADRMV00EU2tPxyAAMn0DpkyAPPumNF
G5b8XP4gfF4ukANwU1rzrPl7mAHSe2j0fTDHez64j7XeTCaNBNKtOro+1LVKUSPH
ic/AFwfhKD3E6zW+PK2usUYM90PNJK8HYiHmjfJoaaM8mz8VoLjl/BRSx8bdiX6g
7JEJ1OAAlAGJsuenpk+iG7KuklqFZpIcSbQd39BkRQ7Xxgu/biSPClFjA9zvyuBT
GYGfkvxkQzsLWrT55f5Lts2PADrz1tP1+w0vboB1ZWEhTuPH1o+7a+ixV3XnSQi3
om/71uEbxwq67jRbZ0SvJE8tfHzPG6bNbnuMSRimyyZXVN155ayHDRcaAnvUs4Up
0qk/VuzVd0sVZant35wuk9pxbzieyzQqR7fKjqFXXqSytGwk/tltn+f9LC/D+cRm
+d5V2tKFf8vaiiKYcxEXZnKjjqS0ipJkdZh44P7PImzxznRlAuWwHOrGhv+hk98B
qrffxjBXCTvfJU+G54hUHgq3utRU3BWMizkQUPEzs0uLwtzp+EhpkEiWzcVUeuNR
q4F7hHFirPLE+Nyu6PL0GSF3tQuN7HuKVjx61Vc+CPxnKttCCetWqhSctJ4esMeC
DTkt8k3dL5Ndqo7tBrh50NnouMHkIetbvHdd/brCLI40pKoExo1ZDp9qYjFCSpht
jvucJZTUYo3WBD7HvkSi5hMyxtBSMRYYaiwV6TDEvzHbiq5MD6bOmELyiWA6MiE6
JAg2luOIzBY5YnfrtZUE8G4tJ0w8lvMANilHy+o8BRpsJPqiTHgMmuSrshagdgGH
c9/JoPp7R4qExFJCH1p0vO+6jhEWxGSff5mePyhy3sGdKjZSYtqge42eNRSB+JDe
LpyYDKUc7MKBeHbGraPT9C1F96YQlpT9GmueKd4lsjt4Tu2DR1Pkaui6dY/SjEym
nWQf2dqrFWL3nfmYHQY26ldA8qV7awt35qGppPvHGuh4aKSdA8gAYPaBbHVcWKJK
W7BHfB5nACCruAZnykBlb2IePAwF4s+JAfD2KoiJQ2thzBsLnRWI8qCjtCHAkLOL
304hpAAIZPgepFp6q82qRxc+f0GGbk5fIoP8iTC6c/EMcIwp3JLk56FOAkMMXuPa
q2xsAyWZMQcuTX7gOrFVreUVdVPIb7RoXjhrih2KAYG2xn2hkAF7ankqVtKZMTV9
Qy8WVEaZjqve7c5RAuWLGEYJlwTwbxiFfYtDrcx88GGzYuiLsHiJql9zskBtRs0x
HtNxA1TwVXVEDddoZCeaJci9AipAZx1c4ofxgnPdpIYTm1ROeyZtqYlcy5Q8JMiJ
fLPZcMzmU5n+uy+nTey62LCbZt3FAPlnMffpBjIn1gPUOU15qXRAPlx+DpL1HX85
Yd7pwwcL/NrMc3IHOziTPSkeVeztEsT5P+VnOl2WPzFf0kqvYnhhaq3cS+c2uDx0
4gQnC/Gd06/xlCaTKqPmSajUcAAo1gHmMa1pbH1VQ5xJ8AJhPuj5lsS3MWHI1VC6
EcD9teUR70aqV5/TjcO8Rjb9qeKaTR1VhEcOU4rSqbugyupJIawObDWnAL61dD7H
tVEBUT8fa2ius8hR94W6fepd8RXJISAnR/r+5LgmCUcp2Rgb2CLipISD8SRPVMNE
rdJM8JgjCBBeez2UhcvHR8ZK21EquT7AKpOzmHYON8RSUEqTBQSoHbwKmvo0isKB
C4ivgK2dejTS1znRGDT/lyaSrNt1WbnRRlKWd9G/wqrGJWVfDsGFjBqaJV2XuI48
+JMJK58BBWGDGkQkR7EbrKO3Q9b7aFrfNjmozNk1AXTV37Mpk+IMQoL2IKMVCXFt
S17KMMJ/q8TzPCtUCPWwemrAWEzXQmSnnSiltzDyWiatMxSxmUfk1RJM0qaiO30a
ocwapmJAl+aXqoCGPRe2FDLVYlxPAhZUu6RogQH8S1q9+879by2ulpeQRPFIHZzm
DU9RtdRa3Rahn19VDYUALUnTkM/+8hQjBkTdGqjwXJkSz5LJA3hOWJhZ5+JGgMgY
JLFg6aanq5QtujB8zINsUWczpf1nzebiNtDV42gTkkvUNv9vSlv96K2IgVMCTRmX
dB/VO/t+YNY3JkCEJSUEeMe+z2RbJAhxOKsysfLDA2oi6NzbaaX7ealFoHfR1tg4
7GLtSkPsYpjQn5MrB2z8qNKCsQZoj/DKIXS7dVk+A88zs38Dlq5xHpG9C+pueOzT
TMxxAqhji/2FyRFz9vpEx6WW7QG1K1buAGW4wCuXW6ojEH8P1Kf4zwVh5rJity2h
Q579vscMeolcqba5+eso7T6TqbxfGCm/NZLyxek9qDW7rAWwASsUEU/5ZNZ0NNEn
2UU1zc/BMQeRscUPUPFg7s8A/0OwUPPlQKfi9YUfWSCZ9h5b9DO22oSkEgYhdmhC
hnIGCgw9/t+DBvccoySDEnqPNrDKNmCShum0VlhyOcTBvXESPf1LhCF6KAzE5Pgj
G9exFkfxVgPO/PsOD41HgRtYF8uBNW9coEkQUdpEFa3hFaMEwn9d/fyCZRKMqwur
YRjkjkWCQtVQHS/mnm1WrY4taoo0zh96a/gK2GD5hnNdmT2cCDNMfpIoDfnEdKqs
H2DWu22AXobrEbniTZV/Fw5SEvJvMcnQb5GMYoXk6zKxHvKMSN8n6MAsNPHbkHTT
SU+/iErzJT6DYZg01eFoTsDFilmAuvcZRn/BHH8jfUUqTuVF12fxPsvsbS9eVFxK
oqJoFyRRtddmQ8RPtUR+nopD5RF9+lGCmlN4w9Sbu9LAO7ISPHcVBGYMPenIcg7u
41A+TXGvuWFVSPIOzk0n/v/N3dFm7PEvIVyyxKaDeDdSssnYOPZ41s0r4RCT99Xp
uFuMPLA1hVbRKyM8+kJz16525Mr0bVWDz0lz5XOtK0zrSiv6AbpRgk/IaKLJNUFT
xn3MIdDFj1yy2gCiyZtRnM9WSzmwOFcGsEBelyV4ApPDzz3fb7pyAx2kaIW5oYcI
jF2h+NnZddVMIF7Zu3lz31hglXiNQs4AskOxD71CYbGgo3kCxtDqU/ZXhOJnIpWz
ak9qwuRmKq9KQfyj7lW7TifJrkfwL3U3m9TglYDj4ufasIRQ0jwkmJE/s49vRNJN
FJPNhHbPPwa76mnX0DamaYRUG98U+7Ko6jBE30oA5WwOSdukJ0FcDf4PemL5KXQX
qj7tdd3CyvjmXJ+5JRz2sUBK7Q+AWot3oYNdL8aATL67DHhlFmFRWNA97YCrhqBr
H8mtHSqKFH3dO0/d4T9IBDfeCtuSrKzaWxN+rGMQlsFBZ7jK5aBJnUmLasSFdXUP
3uoYoSb1DBFnR5lY0T/vZsqxwDagSUt9LxxVDGHWFgnMqTCBZzB6eg7u3/xdMtLR
77p/GsfdZDsk4hDdSNbALppEU42Hic9YM2waeev9YKLVB+RilPGGwxbgjBZupIoE
DnfDO/5TBGCY0iidJiZI99dw4n+vgI+E5/omQeHLrDL29Bbhc2W1qbaAdiOK5wjn
3tIShSsmOK4fpyYLSRuh2zj5TRLumVFLPhI9H5114kBDwVsJFO2/UO1oPVJJk94w
FWXVb53ubiYuEBHMl254B8koI1efYCy+/ibsg0SagO9GkrOLsCydxoy8Qn9KyaBx
amKGQlzgUiq/kwLHkAdrS1Rn4gSq979FzuoWvj+tmIBInd3DNNXBPrM5c0LvaLO6
0afOtzZ/+8pMILLd+tPGwdsK7xbDaxuvhPt2gTCfSnIXRQmRLhIsz5lHGbpofI5z
S9bskt1sZu+aD6uPJaEHQ9h3ZRFovJWPEn4O13iHS0FvegeUidcT+Qr3S748sDwa
iQNNwYgPPWAK/AGKYogGiS67o9O1nL0HvNVzAKplg2fSN6U2FAX4D+LfU0nPuT7W
nCP1lycviOKBxYND4kBruvmcXA7GcYjndfQg/YSjo6fS+r3Ba6dAg3wHJCMg9Spf
xUuNCUVI7sZhMxZ7GgAEq1Q9FOUb99pXQ0cdC2TkQ2tUKryOLwV3HrZAiFNpxDlJ
W7Z1P4Fnh3t29HKOLScP4xH2Er9sq9DwHsOOjiFLvkkeW3ui0fQuhmPGSZMDIsXV
bBkQbQemgRtJgPQ5wNA3m8vAB2k7jTXjFsWQw7EVnYjhdRkEPKijk1oNd44yvSR/
TfzabFJ2xjQ6a0AdQceeIDGpLzXkaH7IR958fpNju3qVHXSb7Q1C1wUUHXQHCn1n
uxv1RL5/hX/y7uB1JIiClGXXXOhHbSiM7hc2etnWf0ZvNWN9kqNPEUSZeqbwATrn
7zHJh6XLLIU6lz6eiZbZ0gHpaTEURjSfJp9+HxZBCVugSO1uPnqh9hVfih9nu0Ed
7MeKJdUaG/iysh7tnexnlQ6kys/BN1LDfn7jLDGRAv+KCHgCTmj5MQBXifsJn3oR
kolENtkhT57u+L1LaLCxcOH9lvH2qm2X5n6LARIymVuUeXT3qE6OKKsnMOJq3kBx
mcdrqkGAoAl6n7RqylDHr2/X/c15kM4YPy+nwdWSHcZp8tXb/1xwalFP6q+q7hIU
C+Pyev5D2pu5lRZDkr6/oxHJ0w87HMqQHOkZKMwzviRszgTkYTOvMi/UGJRhQ1Dp
LH/ZUqPaGv/NrlvHt5RJn80UnaJfD1RN6F8x7E6e29hLdoiEORjJR6tjcHlaT3AT
/7CQVQYCxEaBpucda205GHiSb+3f4e3jsDcc3qSYpzECMX+VJkZW8jkqklN+lRlH
gpSDgRYoCx536DRJX81NFEn9XBZTtH3yj936mlhwLwxzw5jgOQsvQ9vG9PbbCMnM
LQI2AfAisRsWt/5ULcnMKe8dqutx+uhOBOEGln5e4r7kIJBv7iK42gxTjHAxst7w
C7yhs1YmPdGD+lREaBYisZ1EongRra9Kmo3gQgOb6dGXvS12wdOC/V7GyPxnOGSs
FfATWdPelawHiuUcpQe0QkJPGfqmqeW9Nzj/gIkPzOmBg3de01GeEb3KQklAHwi8
sZMFJlGGwAYOCm47uem19SkCWoJKQpVS4qHXkOC/ubdS0ySxS7A9RdHocXK21615
nCr+JV40RvKqHBD4HGVpGwIrQtMx17uxCB8TafWZWnYl3Teuh5E4cy7PED1a5g91
Em0ZKUzHILFOadwxRIzgat3YhUQ/aUUmBSPgTCxZxzkT1yk0N/rKDH/RJOJNbaaq
t39JA9F8kluCAHWxrUttAr2k+4qdA69U8Zg2Cnk4RvjAzyOHJ4SfSX+ekPoeVni0
pPl/HIJSJLIdBxeXZOjN2ydLsZekYj+LIQd3GIHyHEuZM+cCtFE4zIMzK8hviqzT
czcWtLuMPvQKray6ozPK1WKr9gpJipwMDsaq4YWPSmgWZbVvGSakPy1GJrNzy5Jb
mGO9DuI3wAvsVfJ3jMB8JHUCMFBUEaa5Cbo980mUtdCj8vzTO5/NLyPqcllPhImW
Noh33lvyqmjpfiZmn2CGSaH8ut4Bx9fE3d4EMWFAjUjUfzeYCdNjRUrVWwqOiMJb
F8AHbTYNnwbyH4YwFobisv3rGPL8g4vzQxWWFSbd68loeSD5zMV5HPNXIZtwVaf0
JvTvhysAGfQYZnIgw8Bhu6qJWI5xZ0dHllSazAh/Dows1W8pUDX89L5CVAvuKaq5
cOUZBHB6pjg9MORwnrgo7VgOhWwM4ujcHugqwFKVscnwvYR4UT/1fJV4/+Y73Ez4
zc5iEKSqgYwP3iSsxmPkuKw1CHTIZqoaKAVrN19Xv87gezz5bpf0xS1Sj3hRMidC
OIrKDFTyBlQe4ggh45gEbnkj3z/7PUCn4X+2bxGUiZrmpfcU1s6zPbua2mvEHVr8
wQA5IsTuIc7GwKbofLwaqaptmpI1HQR9dVCxlv3igLjH+zNmecbIaK9rEoMMcJ9V
LC2YofY9S9VZaGEr4vlId1GtuIxizmTjrzG3X5/bvsgOP5gkY4jnuBxp1Ntbpcu7
wIXoJnM2bC3HB8JLyS68Iwuyl07/6GK49eGsxTZbykQ0Kors4aGGTK8+aJpeTQH1
gj0ul406UVkU+6q8Okdw9+0l5hcnMaUFKu6OsCTqv3dIpGoDD0HxMOTMW9TQ/Cpx
8REYFT41+RggTU8/GnbpkJ6NFf45gmsWOYKtGKExygDDUjfyXPdChwEe7yt6YiTE
sRKV6/7CZziz8tcQViwGZivZQGvD9QFnCmXoL5KeNrcHfYnAIp5g+JtFyvAArQF1
Cf140Vlzl0XvySxVRWhkoPDr7fIMrzcXa9Pe1T8I6IQw9WfQMMUgln20bFjDDYDJ
fYnrRe6DpNVpPXgQ3Ztp23P/jg7+y+CYIMIACYtC0k1LCEywvY9ejaefFJ1bTdix
WW5GHPE9CtEhussqUSIeq+Y0c4KmL+8M7eKFRt+z0181JpVJmniVZY/rrIxW7pza
99sogyGjEcKdhvfsS/vpZ4Y+1DUQvfjIIGseoD67qr7yKrFGUD/F+HR7XNRuZIza
AQAlPeqvyHNvNS7Ff3HNYj7QjuRKVriRks762dkBiqdHhwTXsqBSTlgyhAp8PLLR
NcM+rhPrjH9f8cu6thP8HjtGgJM9SHmk8kwuDNM3fT1E8gl1SvpymeGzKToyjrga
5bRHclOkEZHHtlS6CXfCibIrLk1WGl9SMAe2EgA47JnNYOUu26dsc0a8Gn0Z8dKM
42xe+5Rq0m75GRxVkXILPfXDSJwvznBMjThZjZnAIxaCp6xUMmmxyBOWrycS4U1f
xlTiorTsjdmovlpNBS3b6ft20qE5jp534mEcDYmfs8FHl/nBSoNLjA2cGZyFey43
T5p/jv/E1khnXq4UcjxKGHqOif7Pz8dRW2auEnLOU1PHgeNzMRuh34jPtr9saojg
+DmniLbfy6s2VwqlxtUsn3+0wlvdJq7AKIEfmaz+6+HpGmv4UeHRb/w4NEhFkA1x
Tpg2EVApYvyM4zS/UMKWNgaIcZgOVK+u1mrAwG1KWq9XF2Dn99+AbKE6P3KuhTqn
ZYwd0rkOHsTbX2vkma8U5mEu4VaCc4Xx/Nzf8vCJbefoFvDtI6iLVXXZZRHH2ZQA
CsmF8hC6RCgVZmvdeFU8CzjxCpo7pCLBBapEKlTqatCUSHN1QQotRq7fkv/Z5a/X
/tOYSWI4nJqL1g+Tql4aND3IB7DJUwBssOaBk8K9oIH89PrZT0FcW6606f0qoXCC
qkYbqiw6sLfA05OTWqo/iWqR2BPQIrApifdqGXWtQVXnLN5m3Slz+QZQoEJkxk3q
uZSXn+u16hTFlG7gGUdH/VILlkkrPOkWN+zFZUnZKTyW/onvXxhIZgMvCf8QAB7a
xeoZbCRmRL4mJKBebdJLvP1+bdbKUUEs+1tDxlMIYghaLWH+7Gi5JTPFd49vgxm+
50DHj6aZ9lY9TAAEkhvdxSpxkeiaZebN5+SFqvdoUT/uC7mW7lBMovh8Weco+BCG
JEaWF5xlRpQkT0QwV8P9403wajFhjlx8ONcFoIoNR0EavfDljD+kiEGISPg1+71E
3DoGSTOdtugE1IzO8RMjruLwEic/YHxBz5NnLflI9sBwAKG4VJpTtB/AfELysSNl
jEr4KweMQiEqiEufeqr2+4BPpMxVvoA0jxsd8zYsO3l81hFdDL1893a7CgukK5l4
NFAsRE17H5YBkSbE/lCUeCCc/d0RDszzqOah0Ecg5g+Fdi1hiD6xDcshT8haKi2L
8nwvC3qYiVtqPIluDXnYFANEXFLOxkDrKBVumktk2zxULjfwRo0A0DNi+wM1tlpS
54sD6WqfxeBm3hsgDLDwA16Not1RzSVhYCg4Y07KAEkt5kB5qsS2ZL2j+UG9kzZ/
W1i/+cYPWr1Di8tXZObPz0FEs5O+jZ75pVJhSIhc0wpTpvMvG5Vevqp170TC81Yp
MSPC8QJxmDXqJVEFmejenpXgAn+ggnacpDPbE0HDxtPWJllKpfm/kOCW6fws10vQ
muMjOpD2j8zUPOA5CyZnuG3n3PLukSxoycbQy50NhjMSGavumharNikO3kyQOvJd
u9vp8QyTNHMIuPoQuqhjmJK1DEYTvGayxEG2v934s4YRvtVa1vg2yIOjREm8uq3A
wVG1rOjNbGkhAq6MiUdbqmGM5qzUX8NR+0T4F5cwfzDprtaGGZ8r7EeGlZq8JYdk
/fsj8bMDu84C81IjO+pFxIbnDdp+1FPSUIVo5UGJqtMiZF9UBQkVyis8JzPaR9Yq
lASTBRLDjfA3ZK4GSy9lI9YzfIQ7vTdg7P1pTGd6WaXYB49jTUWpUWwoYYKhopbe
KlptGw4PLNAEERws4ZRkuzZUhg834qrVFr4LwUN/nXg8BV4OLwIDB+MFR+0LxEUF
LKh3okglpSTyOSmUNUS+DDePmFwNKPI86EEcpS/qwtCiawk2yLsvJwBkd8jhZm4+
yeSS4h4renxl1G7c99Wobtvt8jORTDJI8VdpDbnobZMJsyYsj2nuSxJxHr4BYAfP
ORflHwhjfaiMiray6jgs8X3JdpImgIVFhSyFuMLzcQEGFYrc4J2pjrxG/MBfyPe0
jdswzAIeNDPAT8URH6hFMHjk0bbG3k7bVeeFEJcCDsW7TgirN/YRpllW8bUn3tgf
jwvBbyTlWWz8Z/LGsdaM2Av4bhwabT0hZjBu/6Q15ybeLCPs/bip2dfwGDndWURB
yNitvSc0CgtQVoZ5W9QI9VZXB4Xz47f/KmOM/LiZNmk5YgMuRIkYoPQ8YQ85kdoc
GkE5YQqGdcnoWfevueb5CdnDgNPU3o92KDP7gDvTPUr2T2vNTS3SuBoa1Q5gQi3S
Ccaar2M2rqeDrLrD+03yHscxolrLViQeciZ2hfWmd8EVG6K9ZGiiicYEP/5smyjt
5c+CBaOCjHtbmeGvJtwQWKN3ReSAQZjhiiu+Ylpw4EZwdjWwQyuQvouicacskUte
ZhY8aW73urVsCYplJ74dXy8va/cuniE17/nNWdLu5iRX6fOaKIiWDpmLyBVqp3OQ
4HGfTLQfIXEjS9rh4jTYfRjXpRzJVIyhjup0oCCL+IQb8iVESooT+Vl9IBsly8za
gNslcJ1Zbxf4ECZxykIdR+bWmF2c1sdDQLdk+Rnf4niCV/MVmT5lfTb7QxG7MoYv
7BjK15t517Vb+bTXJ0eB2AgayPib/8WiYCNhwRpnICxn4n0eg05xh2gI94nPZekR
YXEik4dkJ9ZMlBBzEk9yOz0WJuw4IAExffFyou2x6op77dN7TsVWSNOV0qpzWO5m
m+fL+jKruAjB5Xuso8PPmEddHE+84KtUPkWMFKfivr+zfXMnhg2DtWItS+eBD6Ne
lor5okfnVaI2Cl/Mcqdt1M8wNawRhvHncrqnkMLqPAVDnOo++bh4Fdd50lmBKQTA
Z94GpQcusakXV60Fh0BYQomzs7xyNKfyU+FFBbAjRszzklUxGvK8I2sNZDys4b/J
QJ15gy5Bsk1trh7GJ+Ojias++bakTof6WQqQjuYyTiGI3NcaD5BWzRUPnHkzZPiv
n3ab8xANCCNuo5iaehF6mg9/I7x80i0FH+v/cIB3RUEIQjWt3enhp3lXjiMxsQOq
ruyOXx4YF9uUDV2b2RCOMQOGIPo1R6gxjs2dfbs+uTOUJPpVQyuU8alLFV4v6oLg
dow37uESXBJZnHS930g7k3ZROizN7cAECKR9GxqW/OSt5WqBO70peeTy0C5fTeeA
D1tiCh3pAKv6qukZckb+D9modqeOHzUwf3uvVWefxV+TutWPOzC2a384x6bZmrt4
nuIutbNutR/WDpSmfxVm0ku4DFMyi384fTPJBWdG+qILsq4hzikYJ+1UBgZVVjb9
ZxlKyv/mmm8gjXapXTxX1VALi79EB1ZTMW+j/ywM5wmXQvarfwAQeko1LJQ8jL8j
tYy8kSGfqB2055tYZmIFSuy82YY4zGBQRyYTx8XHkpGuXg+3nP7OaqjJo3PaGcin
lr5gSMeEEnrtYhh9nc62AAf4l5kl1ri3On1DaaVrnk3G4ig5xLTftwS3sJFZWQFb
yTgAqqG+S8n2qveY+q5ELYmu54rTG40W24VF4xjcKC5tH6WTZEUrzkhY/g6iIVFb
sOEobJNsxeqlth2wDbKkYHhXo6EVahsnbh+Rs3zgvoOtS4krX5NhhF5SHPy2HfS7
4nqEmuwjfOaki6pjnVzjmwr+EatLCU45oHKTVut17I+TMdIcFOyVJQpfF76Z+A1S
p3fpVRfJwmAAb8SEXrrqxJoiTfvqW0D+sRc9bOcKz1/toCl2C0BL/caCG3TR6ou1
n6qA4AiooIyoTqRZdd5ZGKi9Qq9ouB6yKIK5c7d83Vi4+Zt1G+wpObIX5bP+b8m1
Rr8aMR5KrP8AydmW80zwfBOgdJosulWrTP23yF4fJUV40vuFUcQjkFBCx6sDZPCt
0ihzLi5xdSyrllS8mt3LlTa7Mc542Mupltxh+jpmichezpSQBC4J3Ns39Lc60QDr
TRG8JEbeH9KXz30ncfjwCJTnYuWIWWyEbJzddKt4WZVEM2305fWmvIpXCukBN2ls
q/+lYGOtMhH0wLS9Zuzkj05qcepHL1L31Q4bfk1stt0GC/BJfxhbbGktEjMq123w
thzGWV2YB9+b6vYWIVWwiOc//Sjigqrofhc+rl7Eo0ln4Q810lBOCy8Exm6rqNdu
tCXcsZwTsviBGAUIP+QrmO3tUUiNtxtvAcufNZXnc3vrwgunpw5DfuMA3xDd8XSL
bITLX8saUoPZNuDs7VJmeb/gTDVDRTpRM9fJ8qLV3QoTXpZLj83UBNiu92Hn/tOB
MyuLU153yHzsZwo/AO13V3u3k8HhtWvwTa4wZYX+k58Ekt03oB82VJni6cY6Lrem
/qVC3MBkqECCjb0vCEk1dfezVvrJc7JzN67GMu8P079CTEtO4JU6MmvRwLhvuHTd
yTOqY1aHtPmEzpam5/O8zW9jGNyNE1AEHqaE8QOqXudUV8CNe/0QxeMbppwavjwo
TkOex0fnZK09g8Qf+eJGoR7bl3QuN2rdyS1I8uT+MRvnKYM2F7euzeR7Lg4tMlnu
bDYVlB780NDdcEs7+Briw/73udBAnKlwgWWYkUR8j6VqJDnYxcA3nInHNqIp0F0h
utRSZk1Kz7Esqs8Jm0nEr5EIh5g29VHTXT/aYNs+/YLs3lq0O1zkjAtev+Mn3qGs
xsN6BEZM9ES0atdP54ySCfwVoksmm9yW2dblGz+AJ7KH0oJBnbjBtdr/ziPH9egV
Vgv2hc1sPjMRwfqCmQqQjcytiFvBSrLLujh/v2myBO3MsNRAQ/gBK3w0gPaDTn6/
E3bdiLZQmYVL5ofrvh6TasteAd2zdzC0hHiB+lwZZvS9cl+bRpzSztxqWqspd4H0
05s+n29pJclyg3BqoSLZVtlgsBczpLbtYeTaoLXinYxg6H3HbHe+8pGhdcPqlm3b
CaxZh8vhC3uAAlVOP8FKcJ/sXKjrDUpiLLxPHD97pFhVrVxPAeudB6s4i2stx/LW
HJaK3VQZM7TkaXyD8E5tGQhZJIKWV0/kyqQ5la7cmxjmshBbqHftbHudtzRIedH9
eqZ3iT6MB7HFVkPrXXdkDnCJEmXxXsio9wetY9O1RgeqHwclvaLkE5O/LiOmjARO
nV/HgZWnNochdBj7lQXS5u8f/D9siIUX94dZyyvjGBplnBXxf5LR4d4wjvD7H+ZM
lqYUOgWSbbH93di4y4GUyecFTybFQB0JKTafbk3fPOMwq7zwpxUYmniBj0pt7Co0
gcW0dPv2QY+ku5uIUJu6eFDLhQIb4aHgpZxh5jL9/Wp7eHLxrYGUrkJYzuqFOZK6
MZOfyajv05ytzFWWBgbXQNBybk4lDAmHIgbpPqY6mGdJXvkqcm+5+Csw68qPyumz
pSg1cBONtTqshegjmZ/8+HKe5LEFyhDXF7R0d9MbO8dnNiOH0Z+055a6smQZk/rJ
jjYDUZBlR1Ldq/cb2aVUBXtWNR0xXgC7QIIpBQHUc0RCHjHJ/hf8hxXxKZuVuQGy
d/Y+QSHGGIRxnps3ccK0D1XrH5l1DgVUtGkaJbbYMJATLltX4x7O/vpQeVElAXjG
T7qRcYVMlE0qNM7MSno3uU2F1PicfCHzuOEM7Ip8NonvT6768MI8gJUW+sq+B6XH
SIKXo8jjP17IKFS/m5Pi9/3hMIg7l40FZDMhrSpnzt+m/FmKmFITMQuXmrRSXWrU
t4CGEJ3COtetIj2ksur4Lqau8+3T2w0+0350KYe0HAZafdKk4Wt7ou1nnLhU89JS
vFzKKFzh68hw5YitHuA2Uwx3XbIFpFTS+CypQ6uzAidzPVTy+0gAGnAtmqi2T6Oe
Jtj1hxG6NaYo+CT0dQU/X9Kpzuapnx+EFRO5X2bBqQgeVBsO/E/piAoIlsIo1a5K
se6To92YYWiMMtpnymPLeub6K5lS5K89J1W7JmpwgE+8rBV0AqjGZazs8HEtL6KZ
ThgH78XfIKtC/U6GKUjzISJENksHBcWNwbRcep79a1fmd5UGNDK4/vkahdZq7HDf
NnEsMhk8yLuzglRgsWmeukC2E4JXGg+B7Hf1T5RjdK5Tvii9eH562nqXvB+otD8B
tvgImvMLMBOElW0b4XZT73NSz0m/buQiXyI5ZTpshwMYDyvbHZ2H2TPoi22XizdD
VDYgmPlEBXOb4vG4/Sg8dKD4TTxxMotbq5g1JBNrHUfjmsayenoMBFHQSzgMbgk3
rnbvOaFRknvzx6xPiJfBmmTVUX0ogFU0N2PpBBmilfZLV8FjXehXRoPcwR8SL7Rq
wjdiZ4S8ptZqyxxP6cYkJdoxW6WSOeJbnNYxQ6W+l4KzamRmOg5dARPKI16zo3aT
k8D6dnwbl3YWkmCRwtcgCF08ZF+HAopaozKfh45svy4IqNL23CxFl0iM4bDYMsTz
SzZ4awFLRGi1Q4Pgfc4/zTLmTrEkrS/fAsi/KGFII3QWCXq1/PyWN2GqM0kBhB/E
ih8kGbH9MGKIWrsa5cdLMZnPuMRvKpIFm4ZfOW7wVmr1nIAXM3bDjv2urRzSxIbf
Y1Q4L7GQAz9RUuZzfwCdPZEis9mQByMvoXo3b6fPF0a+M4/EXDaSbvGS//o6jHga
Jsv3RtVUIryGzz5vGJQSfeoMQQokFSeuRomuP65CxibZVQdxcwFzW5i5l8EB+vlJ
LnfVA9ZqC45TxGAdKWouFzpo39sahsXt4u80wVnu6EOlAPUxMy4MQ6P0eGplyrVh
VHah6va9ely0x8XhTCndNIq8Ly3A7c3uIqMwra2BRsisI0cc2Z+XDj7bBI2R/0TM
xYYtLhkpXUiarHbeLXPYrII7bSuJHWQcqM3gNns0XNAPbtATuxYprdgDxMpUfzzP
5R02cpYTCU/Vn9SP0k5fqi2eOpPS5ei2cyaCKWSTRgJ5DzOAU/PKBrcIJUFQlgXh
0HA0iPRsp/RTfw6dza5dw8hm1ZlVBMS1bBbuxlLGlqoHneP7asUXsRp+Lw4hm2Oa
DHN49MDmmJx3L7BWqy1XpiW8MijMRqfc0RLO/E++yZniXJKSf914DD2nUkl5ZqZu
iZ9wP+rQ4URq94fbsYWXaU5ax3HzuB4yShbuiwcI0UuX+Nq7VvxFP3B+yYPSu2jY
6YUX9ZfzjgsCPO0mlBqqRxmfkgcWKUzTg4Lqrkx3ly1veQ+McG7vbx1+hqAE579L
d0bW8uh4r9oWZv14F660F+5HN7G/Z3R/LWRDL8nl1tFRyzMxM4AXjYUrGHbkD8oe
QLClsAtUGJPL8tyWoawR/EPdS5rwvcaKLGZFxSLCdAMdbOAyxMqiaeCPWdDm5ihk
fHmD6WK/nYVDZiHwj782hWalIpUjqPpxXxkJCCypkY9WgUTWJieLiVeaNk38APBG
6sLgPPqwJRiDm9tZ5ekbwajcjkqT+wE6UGxMG4IWUF7JTmnHM/aSIyIXRsEmPiBp
tCLEhbmM0TFXTBT+SLxvTQ2LmI9Hats6dtDfsc9alpzQ8kTsOA0UdZc9rC+A0VoB
PQaY0v/T0MrpR7bRnAXf/48jxnZE79A3G2XsCPQf4xWlbT8IqFUgzfswZcpsjoH9
SKM/lLherBsrtgpWCFAaJ0K0+N4Gsh4W61Ba7eEZs9Y6oTU06u4dhup0oIJyEbrC
lVoS7REOZfJ0NVanJLjFknCrNwQdjlxmSn6EXSmGLTPN97dxjAAk/AsBssW3SRop
HYHInRGb8dmQHZwHJYpPmZnI/wgLTMrVclqNxWJxeYwx9LoDuJxOZquItyDmSKKE
S9MwPRWATIfGRrQcw0z3jEcOy/vs6pU7/nqr8x5umde10yneTHqPZxFartbMq6Ks
6rKFl/y8eJKefO3Zyh2MoRXaTebIbjLKiWE6OBGJNsjRgDnQ7ZSdhWA/KiDJZVhz
R8yWD6ycWJ9Gce93M7PUwn0qpWe6BhArGbRBGLFPUpr0tnEZveEWnGfbDCwlA2qW
E1vHUnCH2465ROJym76oitj4a+kdjnRBgIqa/nb4yzMn3CVgToeAGdv+q4nHWiJj
+MMxXvt/q4r8BDXY4MkmI615kvPesTuRTXz0FNekWxZQKnVq/kwzAOSYWkKbv3Ze
x2i33D3Op+vpHiNKGtyzVbXoaMhZMR4fPEjXqr6vzrLwjv3hhys0xWoJLmRaB4bG
y74t+4/aHmhJg3dRABeyo3TK/G0iLQWSr1HHsNEEpaQ1vajd06nk/ZZwI6rFy8u7
DPkHFQnVfKfKayBNTC0cgsBSPfYIfyKvdNq703KPE/QSKOiWen1O6QGu4rlOWwFT
6IynOn3fLi5Uqs3omj0V+U0KncXuDbNvDX8gi0D3gOwi/aQb8kb8mZrB6RPqeiYv
dBwHdfxZXD2go/qYDPWuRynJn7Mq26zxyGIejS6dbkFztCEqGNrtImecOJMLxgtT
ewOaTQ4PYzeubIduJqh13tsCStJGFlXqc+b2SLzIA8zRVcCU7Vb+HYdagk1Tqpxr
Ze5uDbnTotaej5OnSsn4wDj/X8hCGU8TFVT485gwaH0oKdqIIVEEBwYlrdfNAGpw
3T3+SlaTHPRpVfnQejf+8CXETdOvZpTn2prxdtSWYFTzcSFPA2cRJqprEzPnsaIL
tTBjMYJMHItlZmP/47V0kB/6mfkUKIsoBxE+yFbh9R5+VSuQYdw1o3gUEUcSsUzP
PTAlgzw/ToXKgfiz3rBKUCF7IXgcAm5ytAs2o9U4v963gdbSEU45z82oNN+GgF3+
LlGrafCDOQnSYQF/LiiovR7vOJddDqL5nxBi/ZSiwZ4vRVVcbqT/+QhXEgNE9Uuw
ImUYZeMWw69PmDjBo2S8pT3hLzgTWANjx4fVYvSF2HrPo/3uL90Eac4N4u6wmIzS
Ssqmpre83l9G5Lis8EsxQ62CpgYzrV95iQ5KVjZqnQ3rPxr+ylE7tRG6ZEkQndBP
8d5tQ2J5B98TcuOkhd8PnymGl60l0OiOePfSFkFNpAxi2+CDcojB2ecW2My/zQOV
/28f1c+uF3jRwzHK3xezbS+K0tgPMMom7nWfcH5nOTj4HC5KHXve5Np1RnatvhXE
dvieZ+5hEI6OKC1zsoNys5SJt0GG++HFFfiGFoDr0NBYoruW+Of1OTDCk1VaejDk
gqcrn1sREjL43JNoEQy2FvVhX30t75ADcoKf8g3WK+H1mPA32TO/3+YJ3AbokNmm
LdGTgzR2+4JkJ3XOigWY7vx1FjQMd5dSlHZXs2DPKZBA6uP1LDjINPAay5cNwIHt
IueS8yavLM30Gz9P09aHcEx0XtBtEqQ97hSVY6T9X7I=
`protect END_PROTECTED