-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
vlG8Abnc+/ZehxCKbBpZIdY8VRukOg0Tsizd8MR0rm5j3nXQFZn1ti0F+AUej41j
1YIVAzbcLvc9z/cU3IUuD374rzP8j3WSo3qrKxjLtH0wjwtG1/7wEjHvJPDP6PZv
bbe8McFBXP4Vje6XK/bGndMJEvHiFo0sLi2X6oSluN4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 27776)
`protect data_block
L9ppvykGWFfsf4HafbyQFeOhIi6ntCGUvD6T+iInCiYj975On1rzDZ18w2a4YJ1m
T9l94rhmYzWgKVy0AemglSlkCnjyUg/afiUNhmKvMJVT6mE6zUSLoyb9I+LZKUKk
AOn589Sk8jGzfTDoA70JEyUb5ztK9Wlb/r6Fwxc0jq2Wl6xjrpRWe7GeGQnlQBu2
2hWI7oJYxqgvlDtquMiZBUemrAVq4snYiIz2JHI4ZsSn32SAlAYv5u0cANFAIPV2
rZri+fonxZ+KdgaWYuojdDY+0r9ytrD5nZlv0oJY8ORM6p8pL6/wrwE35rPBAywV
TmeVfUZ/YA/ha4jf2JAWbHasoN4jj6/jaznSpPG7Rbw/86vB2oGFC1So/H3kXK3C
ecUq971oGnYDjHSQhuzFeUTiL98Xh2YA7iFmDlaa2cqyZRt5Ttm931GFtk9deqjt
6YDdFbYVJezWx34ZoQuehegFFVWxElu3s8ndQPxR5cBZKO4SD/CiXN7yByMU2S6Y
wkfa6+GNRpDkmft9gIV6ZFkxnMqFwc/Y0I9ll6LJGtdKDwz1yjobdaQEtssbCCUK
VE62CgiwLhPluAGhwnB6u1UQewFvZ4aDC2geMC+YOC0Haz3LgtASrwIoZEMyF9JM
aIYAUzvmGNM3MW+c6WbaOdEWroTPn2CGVaFNRP3D4Uny24CPon+ApIsPF/pIZYiE
C80/if7gIt54GLGKH03VDUnpUcOY0Upzx7yQRWV1mpk0wHRKdk25sycF/NiyaXkr
Bef/5jkKFpy0P3uyqBFLXN3oE9GifyyvUuXoEAs/jq1Yo6xyJI7eJ1hCyF1cPkDK
1pTWUN6wBTLROFv5/dhxxRarkB9q9Lt5lhSirTppoF7i2zRUpvyOPIUYTTQVc3YW
op3WqqJbqqwfvFSMOkD2q8ywhtbj0C6/rj32KAyZr1uAsfoEAavpa5GvuSeKpF0e
4wJjGrKycD04+LPTj8Jirb/rB+FQzv4w9tK4AzFyT2EpXI679K7x9GOrGaXy8pbG
zLBZQnF96GnYEaV1YrgEyoQLnAvtLvn8Lb1nvNfPP496g+E9xuNJ31yiWU1rhqcE
FZ2G1kpog0PF6JmTRHxAxprpWwigdqZeGXxOPmdR6H0K56MPg6QFA7YpanoIWa+6
LR4hz73SxrFMSwJPmBps/eo47o2rWOpQSX1B0wLjno7/dhdGoQoTp3JHKpc7JgzO
rhSV20DhhCeAi15+sSBaPocNK/PH3YcsTUDIZraI/3j7G77DmmQaPWEUVuWEF4Xo
3zpZ9AfCUV0hyfmCrROdJMhVYKPd1OENfwT9Hv+DfK2vtSl1mgSFWZDNbidl9JKp
4FAwTNCP/eodGz9M+oWTK8Wg+gahZFaXc6vBra/8IE71TODUbEfUUDg/miob5t4+
clgjZalOCi/Z/LnRo7h02YjcZ3/ZcibyTTFF4wEELd7FaoY0VoJGliUTPK2ZJM8Z
5Qlzk+yZnxPzvHgqshtEBdZSVunyY62AR6VxlxZWe+mzt9eOHgKVVeOVZ+NPuFuW
Hk37hSEg2ZK9BW29eodneec6SoDzj06EXRED7uvfQz6pTP2KHh1Cat/2MqBa9Dkc
HWzlVwiUEVNMkW+qu53m8nyYVUCDPTnsf/cRSKM9S6xloK09DavPEd2cZ3m6Wt3O
9s3k9Z0RbfNBxWXoxL7hBjYtcgV8FlF8RvUdKeIa04TsVvR64lyX+hPyqOsnvjVg
E7gifXrn/vIp1MMNlmhKWrUf8tG5B706zuRFqcdBKWbyG8/P2vAvIIoN2NVo1YRV
p4A6sASK/GK1PM6tELe6p5l6APcYLWP6PtQmphXr0A6Fwso4wJ4D/7OuJyc+Z7R0
J8JvsW3RA8E9js0bxq3h2LHoZquCcn1s2U+Bk1dwdXuCcDXRWR6QPjetQSOtX4Il
qSvDtkf6Hx2EAHXQ9OSqZLMxYJhsdqNEPktFj2+ToEI2wStuCf7QmOVwWT/11Il0
nfF+kmDh5/Y08wOxXgNUMDxS7JvFpptjapOkWama9D/gbdyDFSDqCnB9q4kvdLcX
Iw0VHYlKVIFxObE9x5LnPC5QMkPUfF3eEFpRS6hKM8xZzEjeIC6fcm4cdfTQY7ol
nW7qiX5kVIyJauY4qoqiQxrzQf4mfgB71lD26xFSLyDmHi047uaYToUw2PK3/h4e
eFmm2CJw5D/u0hiPqfk9pkmcpaViULtszkEaNatGBF2feN1U8eFP/zyGp1QffK67
uUEhlyyIdCBDgVnb/bAmXWAeKZiqxodigVIrzJ1aM0RKgPFKW7E1raI7s5fOh5tW
SbpORix/JjU2xH4VM9pyPQx8EOyjD1EbrE1LX02YM7kGzWg3ksDrP3x5VmDjGxnL
RKLD2k2isSshb3sVkfHxNXYBY2KZDvgI31EsrQVS447m75ZtYTsqAItRIeQ0rAY0
0qfUTHE2p1FK0zorXSl468xq1lXzGgbc+Koh2pizTlmshhyD5LUtEADMF7hX6Auv
Z/WekIUOemPfmM4E8Ihz65QacPzrGFbRmEEwXlGmtnq92TH+6F/t2uc7XW81QPbX
a38h79cT6ZFBC4+q41fxXRF9Jjd4C4ziOfHeFk/88IROy1OxA47prsf+iwxMATk9
Y/M/CrTRVme2IjUJkN6/QZxAv0ZluxSpAKcZ3AdZ1K7Ruyp/eIFcj9FnxNPiBjdG
jjnEAAwsLNCWJqhCCBPWcQy1uogITV8h+w/79+H/YMTQweRVKKC40bYb91sMUIOH
foSj7R778CsE3BwAlp5z+FfO/rQMuTil/+blRF0Bjk59iVhplERzd1tKr1AtebtR
mzDCY2VsQWyiKAu2ltl2MLYOVxF5yQGCVzfoH57AP2evbH0Zalt+AqhJyH68QWSH
tsb5g5GTNgrOMElgJL/kgzdHobOdDTcWkokYn1R0dbP39uehCQgwM81HH3/462hE
kIs3MQovVE4jLW3rCKcQtqUWjHd5XXq3kyYJEdRPJed0VfdOS2qRpNZpK2z1ZHOV
45GAcET5CJcX4TNUCR7zzLFXVeg10bO53z1DmWcl0h2v2IS8tY7+ec7hea5ehp4c
5BtJwgychZA56JstiNj10fk0OEu2i4hY4utCRgSBOa67tvJz3Yv2kt+DjbxYKPYv
8AQV7f2f5hlGFb+1aOyxeJejyY4noa/Y1Ba8Tkvs3Y7I8T9Iqj9Tw7g86Pvs/7+5
qbLD22Q3ET5ASIh3Umv++83JNLuO/bxomXl12x3RM9ZEEqjFPEEt+EyqejTm0/EQ
O8U6VQ5YQPjzVkaPQczpPcjR/120PCtBLczZyGOV0eBqdiERgjP+oHj7NNf/XEr/
t2bJZCEr/oXvHQ4KAMeKzH6pCP+KAhq3h4n0iW5YYuB6uO8lM+DmGIamiipviQMA
YtDlEPYhayWX99P2ZqYX4ktlVs8JIwwkPCc6JgHSsKQxC0R2rrb1MVTP5uggua/t
pyZVCK1lBV/1uDfBfj5wyjU+BFHqmLHCBl9JelZ9DtAIkPccrSegGPPdZ29mj8kl
Vf359yrPXeRTecLRs4YfpLm5gR9fS09ziIypxxIAiyselNwe7n8UMVUW6Ocylamn
T9yBwRh1GTj7280eXCa5K5acwC9PRYLhoBwCuiceqMPXuZEBAugwA1LSBOfqj0zM
oVVJY+d9ohX74ghG0ZiXydrLxoC+pGKdunsS559HVfGVXQTDURYwDchC+IybD+0n
Uwe/J6fW2qLjI4RqVf5W47uW6Fr96WfdXow2CEjjPBw7NkKe8jyz1sRgidyJ2H/1
HR7hU9SrW+BucVGqLjknJ+a+N/Bo4eqrJyIGJxoPFy2kTw3sYuwbCqFJwloThvYK
XgeE8a80yhNHzpOvmhfDjmeqRFeqBgFz5gj9QUtyzh3jr8v3X6+C0pNRpt5mxCKo
ud43mykYHfH6r8llObJy33uDJlqcJIx2PRes4hQeF0JDbsVEtPJnlX0UyDPXneGM
Sq9tzDcWShXvRIDyQACt3yK4teDtEHXwnKWvVdAN43GFqlzDz2MBMSKfPWiKRXA5
H4oVmo6tvmpETDoI0v6Q/xAyoQrPh1E3LUTOiEiSOYpk1vJZgbOST701owTqf/OS
Ytz0Prc1xlgXyy1MGRbYjsoexYpDNINsV79u3esVQXLeM7h/zpZwu4eOrYP8oMuv
tBUpimSQVd1p/qzNy+8Su8d6l3jaNO+NfP97fRsvSuoo4zZQ05ulLd4xuVkNj6Oy
ayb4mgZwqbh955V7vlrFC8psn/qoM2cAQiBCKsXyuaWIjfBh4UhDByhvOKIgxyW7
Hn/Z0cgA4FQw2Z0IrdVUNDFP/9bNgXBSYrl25m9W6PGhxsKK035zdXAYLfOGAofv
q00WSpBMEYziphR4pN7uBtfYko3ly7P4hQDpE97WjGmFYneQi6cb9uGRtwgNZiPZ
Oe9tJN8KVURCyEY5OeABhOoOrbBW9rqVdlGSopNsS3aI/u1FLRGsyK+6+7CZ6tgG
NpCIgYqfuzOP3miarGs1enVZ78M7Dz/RTUgmbAoTo7JD6g8XWlDl6BN3ZzNQMuzv
TzgVhbP3JJBtRG/9koAwrSJ6A3xrBhFm5db5cxLwQeKnF1Tej2Jkqw6ah7JCqet5
7Yd2Mz5LD+V3/KZA3FrKP7XBifSsPe7efXgq2TBS8ueoz3px9r0mjcdssesppgsT
78dUZan3254Cb4YBR+JUOrWV4xHTRPzLjqlvPdAEv98LtUUzGUebb/LqniSfd6HC
EzCN24FgPrd5wtLn2EoyoChSl1+MWO9j3vj10K7RKRcVg0vCWusbAcyazPW+Ut24
gq8yDTzFJKdr54DGZfVZsX8fzgbz/0QwSwD4SjeLiSyL/+PLC64zeoytMxJxC856
tgTN5Z1w3ptKAdbJWsgFXVcDR2CgljkEP/zMf+8wlAQE2Jh2ASMC/WG3W2JugTTm
6Ipw8aBeeNieA3tTWUMRHzjEkPqK2MbI6RvT4ysG3+GhTc3YzA3cpJyJjyMd4TrQ
ZVvm/P2Rp7fBPWHRS4fyX9eiJjp+Rz1L+fA7FN941/7m8yYJfZ0Qwj13Mk+/jSYI
7BEjNM+Mb3d5kBKtMuGWPA3gNz6LqgM9UZ1aNtSii+JFWUwGvigWpbfYBjXBwgMe
NReFVz62uRljXbe/Kq4OPUk5iF6YApGcghynkyN3UiW08rw6lkW9xz9xaNLJtTBb
aO1FfT4MIfH45IADWKl2KlT9skOwbUgXTf8PdiHqPGLvzrQ2zvPmOSeXy4ne0LeH
pBePFFdnN4n0gExg8FVSYODqoYD3iH8b56Od2xz5yq6RphJISTgIpiLIzJG1z13p
ttggPpMEekkRr0B2M0dVTZfPhQqbudFKJLRQp9Zc3K0Q1eFc6HzxRwFD3z07KoKx
Uf8JSwQV5fzKAPtateW1VfFbzkWcj7eAyQhZn/1g6IE/3W7uy7PpHOyh1Lm+okUI
DP3DCi7z/+Pb1x6xDoP53195rXrBHHMfIUNjnhrkyEB/FdkU7WZL8kCDhUVk6S4Q
QI3qnDj0geE13/5d+QzxFpcsBw4E/vY2JIqVO/IZLbwRcbyEZbClv92DryMOy3yy
dmcx+N4Ad+nIuXxtc5gfHz7IUHlLpr/puLF57wiA/rO2VE9hBg9+9XA/R7GYkv7a
WL1Nan9ANuhREsrNemtuExS7hNqc+NiB2clT+DWuDMjs3cqjkVqVsmiplvrG9T/V
kUb2o3hS0RpzTz5oKxfIt3aByNxZbW7l8gGwzE3Dz+kyfW58LzgSaY6XCYaL8G/i
YD7S0jt4MM+DeIQK48QVZbtGWh0Qn6ClzQyv08g2L0VKMDkPuzRD1MmdoB4xVnrF
LQ+ggqMZ8ITa86Xa3bW/iLy68C41z6EDCNTDBEeC0po/MoRbweOlu6/72jFsjHzc
6lrvenfJ/fIS0P8ttKqjAv3IO6Wc0YA1HG4cr6zNy76THdwwD8Gnpl/F/2kX2ndr
y6skWDjR249vEOmHMud+LDiMc3cGaiwShb91AQv7DPDx+UF1d0bb25yqPm4HpR9B
DyztnRX4vcYT2lBlR4CWfCjZuVO84c6mOXPr17cdmtKaQF7g1xVZubppbYz+6/B9
BWcLADVvmktxNd5N/VWCHvhK093vwc2OSItTPK/BsLrXuHbs9Ai4Ruc3eG1xIghu
aEh5E8GFAxexh7kzDY4ELYjw9EonvAs8SHHwaXX+DIqbeoD7C5NyS+TJ3tJFQkjr
MRrc0FnCK2feLIGpLb/9I4qXroHHDWDy9ieUERN4WWO3rFkXW3SOids4G3P7ce58
Gea/Fr/DA2bEXJ8ZH3mAjfrY5valbWkdO5Jd3QhbSA1/BO1etCFJCDnE1x1yZdyw
XzQarNM7D1+nA5hWhHS6Hn1Y8d0Gc3Bn/LdDH4YvCFbilvcLr/boE8QPHa86hkjq
j6PgIMDQGFfSS60eZjHq+JOCilGYB/wm241W+SR0qSgVwRfdl4M9t7OjdVqLTDJ/
cMdUMIs/YOdhOOio5Lmq3Vth+xHSCY8eXnD4rqxoFmRRPsVMhViYSh9bydqGwVcZ
MBu6Qx/XWEh2h3KK35xla32f/eYG2cZanlRCEAB5ywQ3xnKlX7PIzNqMzGjDwel9
6z/EeACvyBoMuRbC9jyoam4DdZia6FEPHtjYDX4Jj+b/MXbjHxt87d6B7ROAA8zI
ZNXaOASJHoDRF89FFg3hcOOjP0MfKThXKIz3SSMsS/aSWp6fItpNvNr5F4HodyfW
3W5h2gYb/W/TprSJwwVEk0Z4Z27aYUJc/XDN7+YN0J62D0DBMYxRLzN/G8TgmErv
XvhuuNxYwwV5ROmCskUZo7qPFv4hz5aw1pGvT01zFCoNh3rg8PziDfo6Da1oAjHQ
CKiYSbfb4bdtURUtEY+pv/alOw3cAv3Vko+vM/5PsIUG4XD/MdWMPaj9YXXJY717
sPNuVHd20aMxn2mzHac3TbOpj0h8xKivFByHVZsLISCzmruL9sU0QeCXM1NGg8UE
CR1Qtj9Q/MWnEvMhnjE6ftiIwGvWUG+6I4Y09QTqsbTKjgk4bynNZf0qmk2tmwVz
r3ih9cZd7U9ZenOxKiOfXQnCyZBgC4c/HbEsvXwjJBgktYk5jYh2NlxAL+a/DWw/
EiKExyJZN9szuapjQY3FNTws8z91eeOYuZilKFFT+/e6TpnLnTWVohoE/85DwJn0
hq7Yh+RPfr+BCgsHQTgcLry+DNqbkSwdH1Fk3mzgVdhmeUC4at/kMM+VX3ihe90P
qY5QqtUNvlDzENWoZl25ZJ/iIG5l+Y/rkuE+X2irHiHy0rVynDjfDPFUgwgpYvfk
k7HJstLPYG0cZm6QxRVBV8fSrnFNJfeVJ9Yro7SDz3LRe//tHHLloaZwBrX3si2S
Ww+sGPJpwWFshYRvmF+yW9wzWxFW2x3tsOUKxqdq6MuHTNSoqAzcSh1/cW4hRgcr
0pCC5OHD2h+3054y0agxAkgYyoR9EhIDwsEVhfouuYi5E9UAq8Z34QQ8AXM1QeUS
iEmaQQS9mflQ8LQ13aaFTAiNAgYmaypvYUkPW2K3ikNUhOux7T3nx2iQ4FvWE5SW
ALTBtjDvd6R8yZvbbacykDHSudnuH+gFx4J/CmLPPBF+POkRM8et/XdPz6Ug/spE
Qn9wkphqv47NpA1SKIunbJOt4BdMNbA0EJXiOii5KY6nxv1JTJV4V76M6qrHcSvM
voncN04HUrrCUpzfTFWaOQ4Of+Iqk4FhB76zIw1PHT9DHojZsKBQ+cZ46sedQoxx
X0kEIFcbCu9HwB170ducTWwdqM7Avyabja3nB/xAlBUMuN8DR70GVAiz8n67fv+b
s2IupJTpVSN/nxPcm0BG87r+ZuM+RYQ/+ZzDlOZXCfJNc2d5vc8vxR7w8YrFIzXW
j8OtSletmENajXEfIMXoegbBWUMNDaTrPPDNdcJQFXdh/EERb6R2/DSarz4RxkCS
Yno4aOZCF4Jty/1ZKw8UvnSuMIuEKSCgu4LgBqd8UlaWK4imrbVEdslMoqkQdKti
Os99BkibAcVbA8Fe8Fiq8pTpGzEd322ZWnxkK5+ct54w74wAj4VjK8ayebOoYSF/
mZ7pi2vQdMrhrd+P3AzLCM/qLqiDCRDOnlZJ3y4LopRGZFlDC8ElBWtgF/D4HnrP
Oo56BW6cR2dgwhLEzjxp5r+SXlbyVeoFhFFylhg2W2YLLEC7z4Ns1azmhjbL1c2G
7u9Am83oeLlMkqtdKgOQ3ysLb7WPkts2PBpiF0y3Pdu6/llrdPwDsCXLfUvPexLE
4TTf+YI83M6gCYGdrNp0yNMxstFiwysTEwE084K4s+cdG+w2o4bX6Z3RP3SiOBar
5EPWA648yI8E8Z66AJLp38Zep93Ck4O8jXi+ZpX/D2HOVe4KR4ZHYDTUQzyVQJL0
sssvq1LI+CzGvmOQGyl5djcXVW9PLtb4qDJtK9oWxBu9NU/Ma0miPW86Mdnuhhv7
wKHFv5FFaEpnVdU78j+9qc6IgQCmQJ8tYGfkUI0LjA2v5inAfJM8ZC7KUISCG7TP
KLsbNIHfbjbNeM65V0iNbqa6p274P3i2kDTkfOyFVl0UCejB0k1NJHQD/a5+r4m8
qOtgKHJCif5D81elOH+vUqvd+FlqrD/kuaOG3qtMSbr+N0RIAqFB6/YSW/A9Ae8Y
QpM6hAQ2L1MxEtPKaN7i9C3bM/1u4HJEwFdKidAEj8FylN4/i1QxHXbALkPXWout
YAN7x5qG1GzKNnMFQ4+a7NPdxqTF9ASIsYI7lTULNAz/PuCJky4s7IwSSH4S7nt3
ana97BhQDMODyzuiPzXmCYwus8REbVrKORnogcnTNpwhEmXtEa8creP5eAueoBN6
fVW0Io+JVUWojR1Yq/CVzcGEucYVVvC4UX+DiypDh5+KdUtCozmLuiJeo33vdqcF
OAl5Rzr4OLo/Y5YSc9KIGeZXkg04I0biI7X03eSOQBf+kFS8Nzh+jjszDR7UUdyU
hSYkuk6XMS+U2vlmkIYC93RIGqnoGfwZ6zJgVLCthn+fJuFQQKEgYjKVvnJOxfft
xEsKvXgS3tmEc/5xylX2sIMBtltKl3bpymGZRoNluuDc2DJzA8euYy2Ay9areJL2
RYTkHHn07dHO0zShV+yWyZsI5m+qcTxktwDOx4TOAfMGphK2HoaX6Z735sm8TV4g
g0DfS2fMyxmc9dnUttAgE7AiSjtesfkYXj/S3FlO5IomaDNAj4jK96s6wuo5rKrw
w+805CiZ5ou+RIW/hFUq8jApsdkFOP3r/k8nccfGdvfHZY3hMt5SB3GTqCLlF2Fz
8rpzVnUOB8FO1gIsnx10PPm2g0W1AwKj8OyGx5Cxr/ASlLCaN37uebKRam80onvu
Esou9VenvUhxuKXg6WqoPYW8IJZPjn24n+JIYWEOPbdfUN9Hd6LLKzgf7d7DZ2Bk
FBLWKc395AAj8DSCsBXt1bqiMKiRupCJw7jnPzu5fdUyniR1Ka207IjBOxYZQtDP
yAEL9uhpbUfHUYbNz7y6iNZLcc0Zf5hH7Qztg3/SEtHOBjlp8tQ4HGGICB7Vt7vf
R6FOaGFEG0MrBh2Bqsx27Z4O3qr0C5WgQ9CPjexrGoRqyhFjjbGadbVmHaFYjiK/
IYuPAa+ty2RHxmVXBzSUjf+g8tO2eiInmpXLeZqxDvUQCYZiOqdc6wciNtgrwgD3
C/EJnAEgPJgKJWM3333+6l2ZerTW5JOiD86LNm9eL/TSlnfbTzt3YNf0GqynG8uQ
OhraAeeuB13PwRjeUz99p+6JIxXg6zLurthtxZH3s87reIROV7yySPdUEfERejOu
Jwx5hrr+JKKS/9Lsc6GZRut27jBYhJKU3yjt7LHRFStoKYyWSnhW5HPTe6KEi2RO
7KiTYX3MWwlG9fl+228Rohw3oGMxma4dpT78LoXjP+ZGTQpbuEZGIX23fo/iT1TO
ry00swUn/BO4TnRpfu3Nemk3tbBFGLzXwk9yY+TnWAwEjhX4n/duSQQN+2JxBFwN
WfpGWrfd59ZW5j9o04PcEg69xwSYVKYGrLvhpl9Gk7iSoPhMp4Rb95aeSzQ3iM+B
Bqv1vjOU4Avb8tM+25/axJp49f3HedD02lfuoEN7yc6Huu/2D/Rnem7MDc6TtR2k
OlO+GNRz2hvFU3+esh4ro7LNTCJJT34oosGaoT0/qPI/LaG4mec+PMD3MbSkfof/
FtBus0guHjLiCfwAnZIqORKyXumR18ps0tcegh+rnevQXCWG8R/WMzkiLi6rncCd
LmdCe4ptbimUeS1filu0sYiSF/ZK74xaoONvzyCnIeZiwlX7IAU9jjPDwV13neG6
E6TOQJLtFORkhP/KLYoFCGTHYGxFMFCK1QEHSPq6AVLs65q7MprKjt2cGsLpDirh
fiF8MB/BKwahy86tSzw/w0IpMfohADoYxxtnX248i6zm4JiuTKumYYIl8e75cnyw
ysCadXhy4UGW4/YUQjb+1CIb8ttKGW/HPH9TlMiIlLoRLmkPTkUdo/ylD7b0BDpH
OMbWbnjoIN9tz/BtBz6cvY9r7Z9OXEKj1+Q6B5cp120hHMVPkUdrYCYx2jI1XDpd
8/5e9lFH8CqBv5t9Xwzckha0OAGVbDrgotrETu+ObePWl89Fy8Uq3eep193BY4fH
aVRysd0DEaMB680b+JKcaNhIj0XkAJ3MI35gf+wz0vYy2cBZTcqWE06dDaTmE3Qj
adsxmr1JxdNE4LR2n/cZ8/GQVTwPzTtIAPruSiqs1CydX1VsUVqspVGXNGkiYo1K
Yw4e6mzMJmDKHDmnk4A0nt9/uIk2YM+guyGBgyz/XU0CI5yUMoHM1sUovEo9cw8D
ZSFptcgqm3rra4SAGzJoXW52ZlvTUhWWqVp11+JRbMu92/2RX34BXUCxQEBYSoJI
CQOWvE05fF9mJjNv+3ewuuMj6dT+XsxCLiD0huTW3itNSJP/IwmDtNEXog7zedTi
+XO5PiqJs0SeIWBNkbOKiU+6xv/4HTuptMbkq7sa8/vF9WvsmD3dSEMot0+efVve
cm70oOO0P0RE/CpTunxIo5wPQuoHZfGOGLs3iNsNALIrrN1GrycaBc7G+gQkYbYv
7s+rM2lMk6orSrxevWscamgRPgbv0I3Yue6R11gar9ycVYjWMxAatYDfoRHVWNGm
evPeGzFBpyX6aP9xjCjlAP1u2lPBdgTxgeuAX/KsqkcLlLSe2abgwn1YY80cxOlU
wjz3CIX2gmFEVRodtMU4lT4wLPWa58AFvxsg08cJwpJL2KVlSSN0RsQqWCiAPEpZ
hIJVpWTw7spZhVZHpNC93RTwG8MG7FqvtCBJGRigGwCI5U6XNS39VK1K1KyMzLPd
KzuUdI5fGtPnD4Sz5+Ly54rXmNKt6sDQz8/9BaBwtYLykuvxp0LgXC+OmexmAeq0
WGVL2XmCjCEwE8gSC5pmwcjp3N3XAIMpaS8wks60+9d15nvKZw59wHdtHD7eTw1s
FKTX2OtbACWFgCah2TbjdzJBxPMf88/i4Pq+lbJ2a9/JwR+0YeN2jo+7/FgRKAEl
SPS12z12h4oiERlLBzwKAZeCAJRbSJ0x9K0gIoet3gjCDCdSnBCrxG4RjBTtCaS6
OQa4sEQx/W6RQ/a9GU1BQlZZidANuU9oMiDK5C3CUjg0IBPwBObfpgTic7PG7iF4
Yky0bEuMZxaa+bhww/sdLqJVgZmtj6KH7ntePylaG06TA/sfZL+Yry3tZBRN0GzJ
emcDV4NMlVd71DL9XNqBgXPYmYMYoFvwjWk2ouaeTxoH2ZDiJ0qQZkd2gszQEzgG
Fgvco5haIUeHaZI9PhKB4pc6I53b/2ZOEGJlQZmcFzxdxObR44c48npe/PAR0hgW
yXU/3j4zsL0lhvbRMoif09ch8YvYX6EqJr3ZNDeKGjCDhH/57f2JawmjIJxTNAcY
syYeaQ9l+PMDtAAwS9FLFO5DvrHNf7sCBVCtg1kF2b4IesJAtINUGVd2DmMlTdsj
7HcCsEtdWYRS7A4RHYhBTeaxQcyvMH++bxmlviae8OjIMm2g3JTmGTI1eCAFWVWW
XR1UrRIAxAIH+q6fboMaSUVMdqKf0ZFeei1cRR3wLDT6pNAh3nclt4g8NR629WEX
COgri4/v4tX4WVSnZvyk+F/2CraHebksnC7SrsCc8nPbDwmRj8e1JgtoOz8Ytkbg
vUMm5nRLzXIqDt13t6wo3q53u3c8i9+uDYrzQb3Q5tIBrQIfH3RelCUA4u8cqRLB
/Ng3KZyM4hRmvX6oYBn+O5bOR9s5sjTOnQ8nBSTwJ9GKj/Vui6z14kQQUvuAJAp4
vyq27wB4J29rIsxeET8hqzV3YypSmndMtSX5xA5Wy2I2+K78J9yobcleNbloWxTd
qQfKMr/xg7gbagCkAGbSRQzRsQJRH+URCngitWXu+YDvdMk/Nuil2NlomScO1Mlv
JwIcHODHzRjhmFBR5VOAb2SHtQw3huXe4Tlgt5qmUSabAKnKuLheG0EqIMmm8rRl
Twe4hQ4JcnDYeVAUa3dbzMNeyaf0dHmLZlwlIEW4NWfwjxm+uerx8UQrUP988R2w
vbfnIvaW9J6kcXZNeLetKXnsQhCgb2pmOLE5R2fFVpBYuiSQ5N/xUvVZ94IC7bLK
P9fiLMBuHzaE3Cgm8FqFmQDHImpHKXmwJlRawVpzbhrZUxmgQfDOqQgEj2swrfYQ
InSfxYddbtFiUhEREW6Qc3N3clYV4ap2wjS7l2CAU1vqRq9ZHD2oZK7A1xYeM0Rj
3IKHO5/s4zb4HPERO7sSzIB9BT/zqyJcf2wWJRIfCpmz9o0xTmX9f3jPmc98UvQk
YUTfd/pFezsPKvjcDLKMWWBAkhaRQFnfibw9yAU2lqjXMvDTCYziNecemThLIBPv
EI5m3XR9qcACYjBWr4p81bf9S/SYfdIZscAUA4iCskrsCtWCA0NH1wB0iScMRrVQ
uVXa/wdOUx1Su9d6RL+3WqmUq8XnOub2YUY7btdTUE9JJFvR56wfx8P2P0K7Ifx+
a3fRzonjwvgXHVE7/1Ghk83Vrdcp6Nh/4gLvl/C/WbfOIZSZOJ7mk/H63KkWcyKx
IH70UUSmwUELEaf6TnaNYpQb5VRClm2P4/NYXCgtlNlIGSIQupjusdHnI1a0p/zA
8RR+IyLAKevTZqagAJoorxyy/Xv2Sb5WSX1tsyeq+rc03AF+wOeqBHPS/cnkQoM4
DBSdSjZZiK86XwgDRKrdHRFtOMtCMx9ObH1liYEz2V4MCMSMSa7vATeyTKq+OPOg
evNhD5p7md9ic6AIKAt1mlTs5s7zly0tUnAr3G6BWyIBRiuqE6JkQ0LOdxGZa0W8
7S4d2JSs9I5H7JnnLr215fTGJMls2P3bK1HC+QWTcbjs0SsrpCTqZnsADtIgbgtV
3zVsalseLg4r9VTuDUnrZvPNEuFVVNNZ7alwXFUEnTps8zPw44DLMCCMb+38vMQq
ySjlbkk/3QrQxCg+rcXFhBGGPR+bGqsPgXUDkdhlr13j/p2joPJm1/GBSCUYxziF
JdNfLCK3S/jAzpUrZtoDmqwXJdFROMaHz+Rria3Kqtq7UTwSfcd5GSMsCtqd+iub
j26ZfP3Ptd/qaOJ7I5rQ23wvm0ANwhnsypRXXQMofWkhl1J+qz9DdumkfEUIwDnq
m4dY+LvhKFLH/d32q20roGjWjfNVFNAqw1bY2m/GRFnX6ABInuODqdvOHc0KrOGW
12USW8oyZ0TQTdz1HlvWARhG+4Qhwt49em21+8cd4BI75zaz8jQrtoOZMY6bDFVs
sbp57Tze5f8OeV1kbY8gIO7YfvSU2D9Cj1ea28gtQ4md4uwX3mV7NWKkRhumdzkN
XnmQ93cYZVLsmFo/xQmT/ngZUxPCnpiQTculraXFeS4SkknGHMdX9pEASLESsXjB
DLGVG4KquPzxKt1D6cbsvDsO2OIP3WZFFZREbe86mcbV5FAGhV6ALAyn2N+OPrEK
dKUhZcsy/wTgs0hZq+W0+VEE+o6st0taTZDc+muG/Xok9ASLOfs2cJUMknvirEkS
2V8LcL1TZ6Hr2UvB5tGfE5g3+T18NfW/PWQlDhFZvCv/Fo0cnk84Wd/EI4foGm/J
3qbbTLCd4w72rVUoS2vpBKlgo0o1rDLGFTHk3Q//unUxRl3nF3cVE7Q22tvOT8mp
qw9TxEHTEJ2T1KwwP58ahm3cOAJbVb8hYTaUiqGUUSnGEDMS/3UaqY3TLlhPXX43
lNcF/2S+XcQ06agdW2LSTDjHGFXzE0OOo4+JPiR7jD0LaK4mrWWX9p11m6D3ifjJ
2F7eoCxib1V6sb1vrRiuhr5cy7+1MgM3fYU2Hh9w0OhTUWmhuA6xAiGqzWfCMlPA
Q33ETijsdVnq2VbLguIMkCavI7UDULtQlCYBCCPuoOKTXw04Sfej9VQZXQcdCl9B
TjyuYbX2bj+gjH6SjXhy6rKI11Q1ca+MZBCKQvb/K1RNEjrS0FRLG5UQmWoBmU+k
dB3dq3dOjqClPCapYdrbLO0DTrtv6HSUJJdC9thhtlYMHCDHBLEolPpgbKVq7N8u
HSN102oiOwxNHpwLRYiWaD76aMCIwyjOM3y55Q+GeX6lXV/6Epj8uY7Ti9doTh9H
C+FSTkhXxdvXbkO9dp4fPYUSrSG4tcZn19DILoHxyWYffKRnpulBihZn7qDEpVSs
ZdmbIWB2nzXhrM90lLhPWVyEj0yESOjNzo3FGuailWdJITMxrbeS5MAsQryUMYbp
eOObPYHrI1i75wS9hg02b5WZjmQMHTLNOIQ/G+UuLcc3/Se9Jns/oAQbb+RwxWpc
e4wRjOO7jprJ+oOoJfb/0bZBq3b28VphRVgOgP5GwvOsVlg9JJZRAw7H/CLRDnxL
60jsEhTtc9CDKJZjMDO/8QxGvRIvWRFtmAVlQ4CoKfgjmR+QgkTp4CIuxJHjkVUK
AJM6jNP54cygZIIvN4fIk6VUc0PrzEqnV3Gy4biiHEfuSY49WdZ3Mmqmg15ado+f
4bFbaxmZl1WPapQu7wIB1kprhky+NLwwfJ4GA06LA6D6Lyd6raxxsNBZ8yFOlXhc
0g7nBSN2BqOyhHhVt8WgP27Iqosxq1p3pKF1t+yRXPRl3uZHAWmwEjBu4hP9TM48
V7xeAiy8r15By9ILTjctipXhB9+VTT2ba8e8CHqaJd6L01XM4s1Q9fm2lKaEniY0
DuEsUtvt0WqMmMBh+uQJOZ9LCFX9J2xZKoFMvg7mPCu4TkAdUcJU4T9QzQFofys0
yTaLZ7yo/67frwGw6adcVZXFcwmHL/BVMdA1APvGWdjSQ5Q9CJO89FYFVC1kkdxL
/n/eoRocockqfP9N+J6oWm1sIinlbHCTEBnBCS/huD6oKo3WWCBBC+LHAaflauwl
ZLl3bh7r38padCVasqH6u5hEMil8ZiIfmh+ZN5hOzRe97lSwb5i1HjiMEdAplNW6
eFQQXLJdjPV89RNFRUxXuSjzVcUeTBsGxGGW2RUNSbf1bscjKV1HR+9rwS44CxH/
UgOdGp93tmhfe6eaAcmGlRN3ZQjXKnehvD09BRXpP+YxOmwmB4p2L7oY61pnmtFC
cAg9HLKIB5tmcZQ9/TBxp22OCKQwPJUWv5TCIeTm3Q86KRFhRuYVS4EG8Pa0yfSQ
zbJZY1STVH5nn+UOYDGooYKRAwlCOHV/zIOjNS1+IXmTjzXrriybvmcWQuvSXtPY
aO7yM6SOk2/w0ZihK6syJGMesRO2dc1Q1YCTUnbyHb9SL33RM7kn3vo2Cr8z4gJC
GK4PP7Htm1sqOxO0m6anoSiTNmNHIqlIJ8bZKLdPhBKh6kAYZSUWW2APautDcBgr
CU9gH/e5Xk4bmLFanJ3extD8ZOVENDc8l5G3warAx6iNaYRRZu9HhHnuTjcboZHM
nO7k3zgTubSPSb0ze6vA5NlFxBiT0WojYDgQjA/aF/vkx04YwZIzdDgZze9ZA1G1
Y3UosY/8bse41vOSxmIrKCzNZQHp4IafZ4cqlQcysk50tmTsaVqb/8TX+aq40YhW
4NoHZn/3VmrZoBKAQlzNfQnY9ab2M9mCn2/sZnpSGrkn/8If4Q1x594hMqI4okyH
OstPyASFWGN5/8sjv9zXRUGophlWQA9fQy99w6021zMGIZC9yt0ilrvjVrftNVOL
ecyOal59d5c/yKfqe0w1sUsDZL7YzzYIknKl53DKEJnWnJzKN/1aYGt80fNYlHUh
zE1vVhQ1pS5QfRRJeO3LTlSJ+h2RQT54oW1UPiYJziAzN4ICd5cISAUoY5Z11z4i
WvlPHjAxyPQ+tvAjDm1czczSkr0uYvtTOeGz5sVN/8olM3OeizruBwj/9i6Mz7TZ
akiwCASssLG/VVJNUbeJhWt8X06kz8IWmES+dBXmqVjmSyfh52ejhWHp/RDzcTNX
1VjKU3CE2+H4A29xcSb2QQ7iHJQsmzt8IKjCmsJAouIw+d4rsv+MMIXPTn4OlinF
xK7DVAth8z2J8KFKeB3Yk1lstv8z4VEMKMYKrljz7VNlM753SaKVMrhGYQhGLRT1
TTVpQzarR4z30QzZ6OnVQm4wu5S7ZqbH1QfpNAYjikAJVCT/fxtDWnbxQ71Ywywt
toMT/UsbW49/OG9pFio9oc3LUHCRmYAvZKyc2/hPf3c8ujWpKk1pXscejPGH55xS
h/wB3Rnkni/ZUr+WpXD0tGVB3bEYN53WnhZ7QHPH1K8jQRHLuCy0xL0y4LKKtcY7
W6zqmHasHiA0BSx2f5Fx8+zj02gTW0HtohLRP9hOjVxfV6YWHcp0Tw7BLXxCh8nu
f+hNWQRc+pbY0/G0YvM96npuUVgyubxoO1qp5BwP7kBz3WxOuZGkBSvVQW9bRx+t
WmyQ6+XSjTXcWUA6AHIaqEQMQpVlgLZ5F+WzjdHVTCTjgTlueU1hVg1K61oAa/Se
CTV2B8Wu9AZmn5C9NdcZEEX2HjtR0596QypsFxPZDcxqIdK8mWnYA90svjOjlVKl
LoofvW6jtdlQ7ZOrItjGPcEJP/78IMT2JCbMeBs8y+TE5myZhKT6Zbpkl2P9VK6t
USR9dJHz4ON4d/xK2itmvVX1BSvX24GM7Wb55YJXsyN5xcbwTgLCHxrRc4bLZSP0
qU57IOFD/0qxityRS3Bv0e2g+xOQbwysuc8RUneys157JFTLrlhn824/tWDwTXUe
TPLjU+j5hM+sJqvbXCHGdWrpha9hhG6Pg8+b5gykp5Il0TCEMzEszfoTxlX0VKM6
Erw2nqEEr2Mm1JMI+dErqfVNikirpJENQsndtliQP+qd5BKkWIVeuErMqLQByui9
t82FDaX+UtVxDotPrzJAbMY4YaJV5GrzSDA/gmXRbQNZd4L4QhsyURl/5C8cxnrK
5b8r6QYwzFVb/KJJIxJulSOeTZR1sKxbJ7M7khrTm/iT9XlP817k12LRZrvBbPYu
1Tj0Brn3/vKHA4zZijYQ/UabyCHNblCp15xyuWXddccGdL00v/3L9dyHrA8mpGpH
vyuAR0b5kLEGERhNg8njcCvf1dJzx5cqaNTsyXzGEncLD2jhs6MveGj0RSouIm0z
2dWFeiJX82hr+7c4n3KoHlWR8jj2agGgKwLFVZTmu8yYhvSN7WY/U4X9eFpgzIMP
9Vm1gJrgYyEcZGzuGqgqeWmDbXHBWQ6mbPBbJCLD8FDRNdwVnyIlptKY4XC/IRrP
OwJQPG74pe0ByIZ0zR8wTst6z2+ffgcYHTaoSeYZq/ipd5NtUZhANuL188TttrGm
1s6TehD8F6v6sY/Q7u78Omf0ZLxhZ/HnTULjwzJuLGXzq8ev0zv+kMIfntwedyUS
7udfaekBr4cKAA0kkj4xFMQPTs+SBpOFAAAPYPSq+DmjEv9bdSMXFleEHCzzEkjr
BbwCkPAIpLdLgUfZ3pZNiu/qR1xghlS6L3AS+62BD0w77YXrsUvQXHBdujYvgaud
etLzjN/Gdk6UlgbAzrAenUo7XAgnnXnGhdnJn7B7M2ZuqowF/W/rxvRVXcV20sAp
Ysc1FRQc+ekR/17oqLe5lPbHGTVwcm9YU7VTfQ/kB8PqLj5RPLj9qEKf+9b4MQIF
HKlDYdbZ/q2gf83ojiAUClkS0Bo0VrYexHLut/U7DGkSyYgw7TrutwLjnb2EiMUX
W+XyV4HFLZb5IsmqVPzoH0+tkd8s1RkHHc2k53Fn8StKUF4XuCvb8C37WyP3dhDx
BS81kDToh6sFiB4b2pzyMdcWSYpndIAUtjUT1cne/dQoHBSNj+4geNcJdLEbFFwO
QrgVUDFu8rfHZGkuYEABYBSJJpxF4BWXzfx7t2Q89LaeElepr58RKaotSbFszZZV
+UaBWGpOhS1dAcs+A4bNug56HjJSQQShWmdyIQNYuW7FoZ7+vQG9z1g9I/5TWV4T
nCTs3disN2165qeiJL2XRCRAKYOUScS1CE/S83Z3qYZmtO4PN33XNdBSKOgE3sKs
Mh2rNh8ZkBb0aiPkALSt3d6vXJKuhQ37J7VaGyPOxfMEg9T9LHlfgCa44UBuL8bS
RcBaU2q0KCvLJ1vYC01hT7Q42xHFRLmOJ69No7Zxxw+ea53gnqE09BESSNukC8Ql
3ZzdXf3SNsvJd/Ol0+GQNMeCCtrtld/pifefriszNa3KNoa3ZQzqGDqPaOAdKx2X
f0MrSVCZMUdmR9aVnc0SPNbk1jFYiPDNweJboxWTPyx0ocr1BWE91SXkVVmSc0Bl
/rq1zQ3SdlaEP7nVEEnE1p+z98TDTknYX1fq6XuGqYvvKg/bBvAo0vanMvlOxCzO
ORKedsdieBnvD3F77L+ocRNQXldwgC4WCNbO4xvKU8Cbe4yA8zn0M/27kx0mDekd
l6IdszkYKRmdR8EU41yKFZN6cKVc49+QHU7++/PvuIetZ/ZvrBQhgocYDAzCMJG6
/YkSmEoTie0jeul8z+cpb7NgGj84dyuINYcrC01vTaqMP4NpeQghNq6w+9jE3Moj
HtnXf0y4YO9pitqp6Dh9b4/071r6YQB2PxiFbyqn0AvO8ENyTd/w4sVRg0GCgrAh
Csz5DrcZfoJ4riTEPDS2sCFPERFrbQQsmPZRvqk8pJQ9W5qeZEvONoq4J3d630I/
UHADlYEn6gp8BPKeUXxZQNsBPKsGzpXwyizaxNysW785I98KDu0ahEaBLBr62yhH
NUOXmfzW39zejvEuD426HTanincojiSthEf9NTkRD76blSjmeFEOeYeuXaKQ/BHu
MXsecs/N9ubrdLk4T56G/v3HaKAkxO13G/34RCI2IAG/i0Uv1eA+sgiQgkaeDiPG
YHPu/mKeUiLAFYuB0UHFLmkAu5mD4JYLpEh3ISLNwrL0btuo/yITZknh4/J6IHrZ
ksH62UTf4fcONAzQNLbbI+u0VF9i10D4OpB5Y5mf1YX21rlJQIXlcvP8q/fE/1EJ
e8LvHCXNuP56L++KqlysvYgXGDDU8HfAqiw8uvxKSsNT0IfQxuRxYsIdIfFpmuY5
C5oPUYgQ1vDqVsTyIBuzdBVCaN3RCHYrjRitJ7tC3zsVYmbuidheW+pKmzqytB8W
fyBNCf5hGyYI8/bWOSoUmsFKI3z5cYWKX45GWU9Z+OCBQ4alarEkbDeXEZK3OILz
QPKmf1UP59oREmyDneXOs+Ben6FGqm6ACKLQQpgVLC5m74Euxn8FVS8xV1B+Z5/3
QNePueyFlTZwMbMGsW2q3VGW1wRqaxpaxlqc5C13b2Km4YBA5VRQ+YUXuYWRC96+
1RLbyAJBDcoFG/cxsnl7UM2l86OGGyG3x2JMUOoS62xqqWGi7ATJvJwZntrM9Vcm
5Z+aBM8IdfNPVb5jmWDCOQvr19xGR86t5EPMiKMCfb0hrnw8iYYFRpuzsPrWQzi0
zdvS5/+fHmCmzN05BKqBzROVNvRRVZAJm6tYGHw8+mUwNA5QuEfp/r0/QFdqtHz8
K9iZ0aw+LrSwUWQ5Bm1k2qLqjEZJFVMKk6Q4o1Y58Uoz11U/ZJc8aeM/+yQ/Mepx
x0Kx/oYGn5XV0ttbonwJgd83d7pUHbCd4vImw1LrWdTI5gRNzc/EU36N2czUhkdH
mpgTA8ONbWsRGfbkK+CT9FgnueY1dfyDHILN3WWipvGKHR5qqBhovzPY3SG/rKbE
r3jx1gABypA77w+QU5Qt1bJ1Qip9AT6AhorLGUyLE7YcVI2JNliGYO/ZJWOVd0I9
5QkpSQeRjdjyf88leHLeoIfqFgv6iktD8IQAfTVKDEHgH6F9ostVgjFa7DRXkXU2
DU/+KmSIdz1l0q/yjBxKvqbZmSQa9HLIppGE1vNSWqOZWydJNvGbVq3Fm5zF9mAk
5+/wI37iavtMG50CEtEK2X1tSbUd/SRy5abSXhPjXoK+aNowlu+tzF+ALG10EzJW
xV7ckh6pYH3IVInHLH+ACSmRj/m57ACNHXgClu8aCtvD3ELypUFGAsS5hPzQ4f8E
GIxSH1FbB0vnrcQ9IamsvBTUOx/kpAfF4s3sCd+hFVfPcdsxIBnOSoM0bn7JSwpw
Z3Q2juwSDThIyJSgu2apwk0VO9fTc37ufXLzgWhL5r75YNFSeazdAKv16yt6nvqw
BOtfJiXyYjA3h7jiS0d34399yzaL0f6FOYy0AmPGWarlV8rqd0sxem3ucGlayQJ+
QurMjBpxkUI4qIBlqpm0jCLGNGucDSD9VdLY00oA4hQl2ytIgV4deMP/OQzeoZZP
N+1eO71267dlthWMgeM1vXGKG5nV5JkN5mPnS9I73UX+hKm8/NMwIkF09ONmpkSW
5OXgZqSUROC+pqNRFzHI1/kE7n9HqT/0wQLyDH8akeoOb0GJL9ARSGLNxQcIuAFh
RJgvDigVGfMNQF4SEIxFr0aCGaSHGG0rEN5+EipNPC9P+8rMHZZl90EvWKR5DIXB
yvNCsiAb8gpAn/eQbrK74U+BTfdZ/j6aURN3UnhEFe+DS7SYeeCtXEifttar5G25
BnKqjXEzgRHP984xeYN5f2eXfMvB/LJPZcHHCr4wux8nFctPTOFb4KyGsXusOZWa
Y0UVfLrYmQ2cB77yzSuete1yc0PeAbOvYl4jORV68vQg08oLPWSJ47KmR3pM6trI
2LVFdCPtt4KlgMXSQvsjsB+GQ6bkPwYcNrBXL2Mec+fdYZGfkRCiaMY9pvh/ypq1
d+T4mov3V7zGpe0cM7kcWlQLSdH66bGfo5AWfrrqKtmgt7MBcOQ/Nubp4BT4pu3j
kaUIkJ8ehRl8DLel9/f80kFE75KgipcFehYCXpLivGiPv+FS+LnefLBhnRHwaWHc
8sQ7I0meBYQ3Ilq4HZLdlaVFeg8t7Xb6BTOunexfJBSejFP4RTQyBnRE9EIzxLG/
SuwtKSfVuEVfrndIgk6mhi59w9FjZYGKhf0X7QMN5Je7cZuZLsIj76MW5SHuLvvh
Z0iqaDPY6W2UNTuDwWzGdC9wINDMfBzuyVAebjCzNk9mQVXSb6gR/9EPFsr32SYt
4PSc6vjmDx5IQAzLytiAuV7hdSJ0QA1vkaRtQ6mJnuDt4PxGukTRPSUBPx4WxNBP
1nxkbCIko4z+4hQlZF2MoFfIInI+EpnvB+D0U9ep73a3gLl2P3+qMc+foFWz9lja
BuHONDVxmG9+HnG3j5jifbCpdMFADb7w+OiEHGwj8XBcni9pninv3mlcAkxF9n82
422sLEtCPV5vjR7GnUhAsYIULOIf1RJ9n3KRfDrbopk6ILRJ5v7FYWzDUJWtonse
LhweWO4iprQRCtD0FeGSksF2El+nNxmT+cqD8nqjkdf6Z2WQcac1BuEMB7A7/mRJ
0Xg3tXEZIH4oZm4QDR4mgftJDg+xi+mL0YVGjz7a3gkYPmCHw9JJezoyhaVdWzs+
O3zw7gJ7LHUG4nsg55A835CVzh61TDEJcF0zjKpJGpCHQfx44o1VqDsiql7AJS5N
7iZVoIzSTxtY88c3cYne0SoP2myDHc6qJjqVZ8Tc6dNr2TqUJMtFTf146cmqMenj
K01NV6nxtMF3SvX9zf+6peDqFNY9tTC8OWeZ248WM3sfXNEem0mBVS/3CsHhh1Oe
k1VQTyHUFwF/e+rtrjALmcxbn0SkM9ECLMcoqZ62O0Z5DmduCkFRQ5C51fUfgHpx
qvtfqY5rxcCSeaurxKtcrMGRbLvOXS6kNDQV3/6rVH0FSahV7WMwmZpI57WgkQ+I
vz0DpDTKDamVesiIrNXGJ3cjuls3AfC41Ro4kqDP083Zhc8O49RYGVvgWi4X8XOA
1bUjqOpO0W0Cu8QjOtYAYuklK1avtLG+MK4HV9CEck/suz7v1RI01PB0jPXRlAJy
mcPf0Ddn/jHXo7xeImzEEQpOVJJhKbw16YuT+sCRAuptI71RFDwbMvDdsXIFlDaf
PIWU/TlVhISunFpWYXlz+bB3C1whb0iOBAXpyLkqF1QZPOS6ASCkwDQwo2vwKPYf
/+p0V+lNWfkyyohY+60DssC9HAmjSgcwPmJbwVrMXnZadNEh1LV3OJDG9z9tNpbh
aHzliQi/zV0ebSqJtRQFZDer8wSF/7a88v/X31BCY01x+qB7YSa8VXdF1//8UeIP
HamKhNd5FGbrF55CsZ17v8FkBZUWqz+NTKdxVCZElOaPbNVLdLb3lY/7J24td+zp
fSzqPSznhHxDSgCU+H7oG2JkzjQc1/DMnYk+73BbHWrnilP7NZvG/gHI91NwUHUv
mlGuF8x43qLHackLTsvfziBdUTeye47+5BSYIepXMRmKWTTSAIvsyc6hWY4HOogy
Advtb2D24veOnCQeckhQbDGcfcZMBXTXSXC7N3Jdv9EHNsH9i5rNKYabXCjl6yQa
Z3iGxLvYJbJTmtvE+2fT3z9PBGBgALZBwLkzIFncicML6rvk4cKcpF3Lfq70VxhK
55K/znilXuU/+CEdkiTbQKqsbYWI3vLZI869DDTHJg/b5HpGZrm7R157sObYRh7U
9hfN1u0c+S0OpHaEDy+TPMkgXo1gRMZJG8zpjF3MtABx3k9CkIOvLLfnQxKv3iJW
wogEMTOgtbH0i9YL1jifiDV1yO/N91xV2pxb247Vl06NZ4MaMwuxbDb8wDcw3wFM
LV5+UVHOIqzwbtuJRuPJq1s/CI+Bd2GFgLYSPTUuQvtYRWJDlY8nlstTEURZSk7A
3t4QHUXqWXJq2aEH9LC8Mm+gJqPcbLDddkabsu4E1u+gj2/Q04CZxvjDwyAftIIR
+9ubVpenadiTXixvH+uK5aeXRfOjoFtCD3qjtBaNXRX765wYzZwlkiqBiohxcxli
zY2UwIp0jqRclPiMPJM4wy4i7v2ClTHPlG5Fhc191ReakZkvRZliLYW2rul/pp2G
U9qg4JvGmbbKP22ilMJxmHCH6jX1xohIbvxncfnFteWJVrcRzxMkug9QElE5k7wR
sau5vvCOob9FYbCPJ2COobDgiFyGq6nLPdI4dBOqqzJ/VjOifrOMuiYFTsCchBGw
1EFmDVZTGbqW1YojHdCbmWO7rxhC3OImq4RVCrFYIzCIRlHGuz18jHNkfu/4coqk
cULyKdbPPOBtU/JNcyGfn6TL0o1r9MywR2IO3ca+HdNHrYPtREtNaVar6koX9pGr
pzq0VfJQp3UWJJPNRKvJuA8PdwppdB2/Cd6YAuUxrI2Bq424DMsUhVbEgZGAcEim
EQIK96oUFUTNVdyYko589YLPoyEDL9xlH3TpvQQaR6Q7YjAYGzXH1l0eeEJpGCmh
UIcUv8ssDKP1x1emzEsrKaaieMTnTVhq1mGF4x+LhqCljttYYaVAOMW0SWJBvGwM
OtHcTRwZRcSQVz/3OVyCR//HlummJbZfT5M6mtGRLBJfTGQAsrIInWTkO5iuN6vl
dJO6uiW++1QjP0s6rimTf2iP2EpDfftdqN7qeYQNGa8tWI6tVACZlRqQ7fDU2ISt
wBjR3LPAv5gxjVWbfJFSqC2GZEwOpjLtRF17LDgOwoxjCYdGMjVyacdeTiyvlVE7
A3Q1/7oXsGPUhCo1ulxENqi3Znxe6ThUL6oZSuznm3kyOOkjG2SACZhN6+iYNNfL
AQv6VUSJxovGh/WTm++o6AgZWiO4/MqUDrhh12mulnsbcnabP9SA8zaeuwmDYN4K
SlDn/dy53+/6KOrvu3VRKVXOZtQtIM9D0IT9tL7t+rNy9XzAVGrw8CzkCpHoS/VM
g3AoE0xaCIP5nvDRDyfeM+/z6RpGxcJsVDxAHQpp7r8DKZm0MYysbNAtD6QB/gHw
KNBnQh55ssLEGm2uwa5uO7lTu55qFBrcn5lQ7Sz/TeY+65ebSf8Yr9AKr+HgRtoB
gTFJwov6b9sIlRwZ5Iq9spr4waT5w9zKYs/e5/JQg6s38VOaQjZVJjp+xF80yaOh
p6yilysvAUdD/6MDLc6o4jUcqknl1t8ISie3zkTVZ47LfwCcLjBfzURO3eSxYW/M
5NZ0gEDFUObbi9mGRIgS5KBgiagEAYJyQeVEuvcA2Yk2ltsfkbiJqR4l5vNAGPG1
P8Tojsxz2IG/dGWoAu5V/zgOn8M7zFT99XcLEqAcAJNdE9pT8+pt1rQQ6RjolvAE
judORfAKWARo2ZckXGLJ6vCWpk/OrwZX2HWeHyw+jOT24AMBS89W1A9d0GYj9qjn
BLWwEDjk4aeQWjiId6OBsRGbLOluHYmBBiL4lktG02Jq1FLfe5xctKfDcRF3k0EO
xLB53i8iLaG3/69nZjheD6WXq7nZNycST+f4wuonzTRcVRJ9DU+T4blnlGNzWBp8
3o9YG4rKtYu5/2SANu6YFP2iTtfIH80rk65xuWEUhk5RthVuYFA1MjcHzqpX+FJ7
bQAnAtHbaporQUUEEAQ5R77envuYd+7fMyTL7+P4tKSy9WVa1XpzaTegj2Y2vsCU
63Gk//NNlusX+44L0bUkSdFDe1dNOmKeLutjmcaVgHgwkjstxSUefxiMKD0yQvCH
GVEP+1b/b+qHQ8MIaVco8PUb1C/vfldTkDLtJnqyQegD2F13W0vwQ5EONoKPbYWj
su7m8FTjPQpN0e6AOlkKYkKybCdqNgSJIUXrFcF2iJQH9XvN/vR10EEJfgoPoH1H
RCJITAcz7FpYWaxllRjqgZppMOwnDh0tglj6hPUGcbLbuVdZOcslVZ9jaxwEi2sZ
++FzaVztajiFVprE6dHKDGRPhcRAugRA4peGwuvCcb/n1qNFyNvy2yqhIDcUbbhD
xDhX7Rvb9sYnbLs1xE1MCbzJv9J2JvHur3uiFpbO5ifQKq/lsXRoiWVlEPjIov8F
i0MW97j0QGbPIcSt8F65sKKuESdvilQxlvsclDcn7eP8bcJk+MWXhOvViXPAOfcX
bMBvm1CJc8lhc4E3yoY2s6rkaVIMXGFwCayUegOJGbKs7GSLdDq2pordUUTsZC40
K32UQ1sv3UB2p0uvU8BKYPCnyQPdao50J0XNaOkZVtzLbnS085E/pj1F3NDNqNhx
QOnZm8NObhroQb+nwL1rhTek1GMWJQjBskJmcBhfSd9FIB7QrhMdL/onA0xixs1U
2nQK41ia2JnAyWDFigbabx62WxnXdNuhTUEraoJ+w0LdEhnbi8JcPdHvaOfMNEgu
SFr2P+3ZHyvre1ssaHVwQCU0FioRPEVDHTMmHxCZl9JQHs6NB6jih/ytZe4LyY2u
ktZ5L4Gm80euzwiT5qNIPiU9skg3uFTK6WIzryCQ5dKBOyeOTz3JQVD939ODhxcZ
WCgBpqsa/agHwVqIAImUCNh6DEVx/2GkdjNiMkW92kIsEv43dP/CEyxAlhF7e9u5
1lNvF2vWQcfHdiYRKYyhJ/Q0uAmo+oPe/HE7AKj9EuVSpv2b+BvAAQyHOuTiYZf3
u0hvqpeqgJV8qE6b0wWeYL6f6ma7Rw13cywHnVFx4cFhX+0x8gUG3EWFNEJl9Gw+
JPDBQ5FeCOq0RW5R+2ReQ7d8iXQGtJg9aJqzW/dGbWmzxv3GZ6ejrTPTioCJRDJq
KpUux0InDbuZKvN6A+CFguUn0nz9lwEsIqBpV/KjTGvaiFJc8c6c2hmTA9R02bDM
sPUQUTxnv4OFojesvCosPdiiUcjh5EzVN4nLD+Asq8e6OiP8g7BPw7P59lGw+Q5s
D3RG4O2b+u3Mdywbpkn/dnye3ltaCQK3RCfFY9QZXPNDp9KqtnX9LIhoh8ehiViG
uP6Zb6TFYIl3oV3LC0XEwN5/gkeo9ua5JOjqv9Zy1xP3LuiRKypdTs5Osxjf7Fwa
V9SghdAeuFiGyZVxeFeLR9CpwPfAAHkwNrEzzqTObuor+QW4FZdZWBUNvBJMTvGM
uTm77p6YtYkCQwATcezidN3cscY/MyfP4tCD+gSQaszgE+IzumfH2VUnS0tr/5ar
dEtDChuSbs33sPFcscGyI1TGGp2Q1h7RubCxgx+vIFgNdoWJcNEP4BKO/X6ZcKiV
1wL/Z4+PHQPqlx7NZraHBWTRkZZ2cPTzbgVNhtibCS9tOnOpkEVfHzSjATqhp3ux
VqXpMa/ePw+V6UrHanQGrwmzCt+acsQUwGIKmDcKWHYbRoEeyYfyNqdxwUivSLG9
p0Dc/BO/lXE4cBdUwEhnPBsU6kRNQ6wXh5DBwhTjyA6q1IzNlqsK3oc3/MeHyQ3L
HMjU3x61OL27s8oHlxfR1hDYvoKAwVfNJHLBERMfACb/ufE7ima3S8vf1Cvo5qXm
nNgiLdCfecPtnGPguyN9hLfcKN5599lsIbg4KWQ5hNFnsCLn0k8hlUciB1nAkjyz
Dkvse8S0RYVyuDDh9Glk8svIYGKbtzB14Hw8Txdk4DUwzLnX7fdAm3cSDmlMGy+Q
Sy+icGlgFsvy5D76McZmfpYCQ1iaXGuBeYOhEc47O8/vcajj/ftarcUJm2XTDRr5
3SMBJa3/YbKt0APqzIbHYLNkp2ySnOcPsqwdHTlhP+b1vbRHzVoepebPQCyUboHD
IdNX4Yo387jKS6pQIqoDQLSn+IJ/XxjNcz6/5rrLXYQMsIyZWr+NCZA9UHxu5UnK
8isN3XDlfeR+rswagt2UJ3TB5yLjzGeMuPJTAYlVnL0/jXxzwupI0hcg/VvYAboI
6IVw8FjpVSUM4am1IMvQYvLZYFZ6zAXkpvADYetsGcYp7YcD1wQoVocQ1ndfwJ0P
6LpLU6lutDB+WJsCOoa9wp/wbGHFPc1pl/HpNFcDe4/5/uyiPKKksqO7HWL9o+jQ
FKSSTqRPaQcBF9YOdf8j2mZc6udlZRoYIc7/sa4xyVZCk8r2cJWNuk22VqQ7jHQV
bIWCL+L9RRTX42TmWQs0IyU01GPGMc17eWhOM+laVtH1maFRXVfa7cS/A5EshBJL
P3AYm3pJqYqwO+JTb0I2sZOdBY4f+9lpvoN6AAtcidkm5H870MNOyDUOIh0E2CVN
Grk41rhZ2IpWpeOo+0DvvfgGSfpN0IN0uiPy5prRY5RFtWK179KlqzpxfwMduact
Z6PjoJgOwCBNfPbZ8vKKGUap9S/LgBfbjRcYHK3sv4d42HH9zPsR+zZ3oV6nrnUx
x4rnIBrb3RA6FZBURaaydhisKu4rEnezpUdM6B4vT51zDdvMy7KvuU9VfDGzF+/U
xht0JCcIGh3RWgAtjSNq2n7Oofx5qxsB/ga3I17XZbAjDtqDCfkc7oKlLnn2btKu
BjEb3zbG6btaLZrSg9c78p7AwghEi+AmthbcxSp3VtF78Or6wlzcQlJDrUN3QTbH
lyMSzyWQIGlU4wMkUkVbfi5xUqsgAjdD8u08FonouPVgJBAka0ECAPh0iJAF92vv
zAUKK4FwD+fpmuhM/GF2Z/uzxZRCz+00hQ4HdL8JRFRrul8z+8TrsOujSox7AO3m
bZuRm+zYdATKpWiGDrPJCDsx7DfqYJVjYiJ9wO0aE8ZEO8Btuu4LzIpPeIMXt53N
vDVA2mdLS8M69+Hu625JIPxjLQBERjuYRrZ6A1QJRlQ4YZ1yYVkA4nnpDdS58YnN
/uB4k2UjaQ6q+fNf/Z4GoMZf/hRzhYjJOAzixvVvz6XR2LvazZv4wUK/PPBSwN6U
1qcyJZOa3OBbXmqiEsLQo3AxUcTjslg/pe8nc0mulZG7iH9cB/E7WyVDQSM195As
PFla4AmZXE71LXs7m9JngNPpD0iciTmYgDko6+Pyh7EaoXP7taI9L1a7uEbqM+dl
5nOyZB1Pe6ZRR9oSvQTuVyIvht3WQtr4m4ZZqhq5ZoqUReH6Q5dVFEhtQBO6NQzv
tMxwz9lrhGe/c+NULdBjeUNHCw2E3FvqpX+HGxVjv7D/OQ0A4dkrAAlM+x4spOFi
eOp8i/v9ms2Lyov2h3/ImdP607yKHyfmwnOGjoYO4c70eoPKeDGJv5Wie8M/jPs5
aNpYdULpMn24HCDcJgoZxeLP5iEAWxsPv4E8Wo6QqQloa16kHI/uD9AntjelZpUW
0r/YZjmR54MP+oBI1zt54mxBtG0yCNesg7J3lpJlCjgHNIw34cRiW7xm7RRM+N3G
bsYsY2IUpn/l+dXg5B4PHON1DRXziMV80wN8Q4KEuY7V4oUupRem5a49+tbZQubx
5l8+KyctGaUKVvjC/x/0vRqvPfQBYiCRg8xyGRlBEjAe/nym+RqqG2Y/ilsITRlU
8NRnGA4PAyPijfLACLlQNP0Wrl6AfSBrJW/CWGy7IbmuX6qLHLqoyH/dj+urc90I
8lxwLOhv1riz57feYSsNQF41LTssmKP9c0SQ5Frg3KI51DMu9zegWSRk5KfBKE+c
L1wrMLdOcGKGJYYK3qxsI6mb6KvM4Ae9AwoW8OwAb1/RWNjhd0eIsLa1/KJeF3k1
2wgZulhkyYBmGDZ2UGy4Oo1c6Bld/1mBB5RYczigMEjqSJbSh+NLCxSeYVEIbctM
/QLADNS6Fxh8v1DRe4oWfBdixtE9rteFrzCbywB0H6MRI9l+UP2d2Q5uKnbRV0Ib
uiM+5C7u/WMWAUWLWIz7AOFhFNkbOCCnmoDDA3MKGapSkfJRz33k+Txv4bX4kV7K
9udFhnFV/lhOyxBSwpTJ32ogvnBR7wthI3yfsrkRvUqkddseoLv9a3dKduNMVLIN
/uPyk+2u7iE62uAgjHWAgbZ9Gq54Xk1tSspF5Iioy/Rn1mvUyS06/vs2P5h652dP
sLVgDjXa0NpkDEkJS0Lgkmle2VDn6D6hzv/05CHB31XTzmgXtpUzPsdquxJeYMyZ
/Uacw2huCh6lBNVBF50/qCTeszzO91wFISHNcBNGVmPpxBxGvAa+k6HGxJr+didP
IrzTAdQRD2+5WJi3eGB8uvRkHpI9oqOMTXUpfwtur0CTsfU+Y1XiNIfrh2e2D+zU
Qx5PQoqir3M9Xb9/tXbsRAMI1ZSQU9TUTgVkGgwCsFbPdMgtDMLAgmGPKU35eMY6
dFUvMCms3tUsa4+cTXTlePHy/31FT2pWr8c+ZZwSG5dVX7qNuJL+60lGDRHWf0gA
4YoLuPg36zJjx4nlnzeefDjQ+SPWLZSwje46AYnofvQxL9XMW0vcXxIjsSFzpXPE
WcFXYVE9Oell+P64xhZva/6X1Xd9Pq/8jOm3/xiQz/t6cJe1giel/vHtwPzYn9zF
R5g9FziHuHPVlPLNWPuQHrXASDxZ7OE1VKIX8og/fWzFCV4hwNFtxz/bMt4cVb5m
xV5hGk5EUi7HeNeQYhiXIzjKRoR8m2VtLatU02O67e+0Qh/z9PbjjW+LXDD6HAOL
4Buc2kkQd30QV6y+vMoe5TaiG6sTnWjmCDDCs3qmkzE8uvfej/vGuF8J+VbLxB9J
uUs0Muz7ju6pwU9WwC2w7RHmn0Q0K3mYXN4mIkzK7RnTJxU7GV7mzW1hAY0EEelJ
5aE0GCWuCzF3pnDzdwHrOZ0GVvo+fhsTGO0igOeAO4LxvlxAjlE9DxIZ+D4rKo8k
i8hBfBIMBM8oCZuEHKb+lHSZ+0FBSDhj09Jt20mlcnDcTZpwSwubTBBf0qOIktq4
xZowiqxeozwKnFPKCeU9fhGN11n4ZDvjdlH6ZMQvyU//GSu1qoa9NLKICzH0z/Z6
4uiwIQnN+kLfkvCxQk1xuRn5C8D2E60bXXPmSdrO8XaVOZhVfDAAkycqAGn4FNa+
SuWb/zmPWeXi21SmrniytY8cLjYSKuvuHQ82X0W6rnhDwtgA1AcMjKWpKyEKIuqg
30t2CHjPVlyEi7BwrsN4bD+c4JaUYvCQpP1n12LjC06A/FPxSoLB17N16mRdl7sp
uteFqfI633o5zWUvGSIv2yu+9pLzcLHUuCuHI7YLqdZL+iyRCn8twOKJCUI+cAG0
bCSsNhU9Zx9lFQMWfKEvRnz6NObUWUU8dSPJGvZFhFBwHfup55BhnThf7cB5P9OT
4zB6gsgDYZVEpBRLPS27oDrUBsYy8die1nKTAYPEsHkzQMDyh+0SM5J/HyOyPui8
qWdpgnYlqIGE+9vPX7qLTFlQUuNOcS3Y6zGnlYkGtalBTTG9u55zPgyJcznDCd6a
XvNNo+PoDw9861Fi//9UbS/mEI40dstrs5XNQXfy2LDYFxInXP+PrslVwRPLpcjx
t3DqsZMt99MV5ob1ChoaS0MCfg+r/mmE3bg+FHwlBrMIwI7dB6PFrQQYGxoxCs6S
41mQokk0Q38wFGyYQde/n3qJ+mHsGgnMdzWI9w2Gz74jA8mcYrm3SjIbebQ4ml7I
CsgT8kVz01DgDsaWkH4QPVo+yszwO4ba9uQP+vNpNOZU6I2ShtSkHxFnUtUivG4D
ZeJlrwLwic2V+ZxLVGwvqYac2n/v/MzKWEPtvGkOER3LMyaJAuqDJT4Xd2L7wVzj
b2jKOhDh7gjqPzVRHn4yLG37XSKFDVWEgmNGpfMrkItePLYlvsk0hwLZSoS71b5N
ZiWUd/Zt5mAEh9TE5jFl9OHRUYaWavMJ4YBBOsMfEGy8zUdGe0ZSHeMSjY0MORIJ
o3f0PGtf9mVoRCQ/YTYdSv9W+B6wlsv5rcaqvaRudjpGoinjTyaMx/Y3Q90zdgcO
JNiBb9nzBxZodoPd++2wClQcHgA+L2DVuKdItXqToUmJFG+M9N1ch9sPC3usLHK1
1zQEWrl3VqdtlvW7uc7Nw0Ax+UMGvT64Emchu9GV0N+T/5OZZmNu4RAnvwv8IWXC
aNRYeZKjh6bj411cFQ8jb3tvUNx2S8/fc96rxDZy371TMdc2af+1DkgA75RsdhK+
QIxlGWCEBbCiAj3U6ZBnqgalrSC8p1gs6ngrS6hVRCXn8mmMK7j5l10bV0A0ndiH
JQ3dfHU3G5pMUvEuxcoZGoXjApUySmH1uxthE3PmAr4WGDj2JVL1YhGBAOthKVfz
IsqBFMRnLpO3WSXCEDX8qM5C2XGIG40JPLCvdBn+ewkI2kKvTPHyuB7gm2NCvBaD
Zv6QGWHCDOJbRiX7Sz+D1ZKB1nwfv3Ezt7yTYacDc0gmwvJlYny5f16dFRZ4wpDy
fy+ZJCm1/zjx/G5wfrY5t6cih8BgT9FiiLaC9+oibNmc9pquTFW40cMZ5Zl4halR
Vfdo5hQr2q0aAXYTnZM79gi93oO9XbTIvqLjso1KyRwhw8Wjn0hUs77Uy3wP4daO
LmZ1lIYMIOTGnqQXpIGvx4cmZZdhka5OqjLnU5Zk2Z4oNJXWzP+kJFXWE5FG/Np5
LJNkfl3gUkA1Y6H1Kr0cWFNsEzvA8JIVW8o7ucq9d3K4slImGvoy4NDZHlog9TLR
xDqrlo5SykCJKD34yJuZ2WFPLPfHmxzi9r7WYIGc5HcpB8sl/Ez6jznBGxGaRBWQ
xS1ZI50jxeGpulWqYGK/iFoJehT/mkcBm3yO8Tj7Ll3mLQvFvIrLWz9uPRnsKPvw
2LzaqW6AiOhe7KvytyI9ccUGoIUXM/dS2UeyG5hZUf8wZB0/+u9+EpFBK5eqMfAK
QfLda4jbgx2hGknH6F9NEnCwQFEq9KOtS7EsdMd5Jk+ZQWBKsmNjLHqe4oxShpFt
NltHIrqiNzhlwLemthowj6XXwixTEETvPUOvPiZFJUZJKerW8x96h//7hSxsH3db
a/uQhLRmGygdECNicdcbnYSXTuKD5vB2+sa7VaezqWwBpwjBQPzoPRgiVLi5aADR
pbuRh7LTI6Dm7KNa3YB0vtMLjzrTGwcj00UTGqFJQEGVFJ6DwpxU4ib8OdEcKEDT
eYKvXRu+9nraUREJdEnd9jRsjJkZ9QdzWuE4H53UmZq0+J/zqYbMBbmrObmHdnX6
hpMzc+wEkIcxfRwz4cmtO9CgMRn5K9XsmrYbUsnCg614qOJSe/AvokHTfuurgzrl
iMrZT499XjxRP0ByE6j0adfYk4ZNCFS1peVByuKV3g5/z9JXkfwOzz+FyFTVCFTK
nt6xPD9JLaX+Itzy3QJQOPDt5qR+mRPu1QFoBvE4+t82o2MGf4UroMuiWgmPiAtx
l4KlA3QcEXyGRMqmBAGKDxsPJFt1+ErnR07rAEw+dw3OUhRiEp3cyomBz3I1nBEE
QSx4Yzy4jp8onIITRTzOhC2uw2W3pvL8LXkkXShEAOpShCtQmF7rnuEDMaCub0fp
bJ92El9CAbpstuGyXQ4atBoQFZE57wtXSz5tiKENW2RvD9fgwoBqfYFMAXx/798x
v1P8smcZQMm64/trUIqg/u54kysCBU2k2Sawakufuxh9xEXQm4/3Vb1sgErv/I67
AgUw3EGdUFc+FlUM9RCj49VXQ+RAn7AhCMfIUFLa30VBst9z4JAIIQf7l9SWDlk2
i+yKeJ/lL2Apt9v6aYYNjCDnDYsnVQqnSXRlAKeMNpy3xG3ACzJd1omu1kHzTIqi
6fgrTNrirl/8Pet/W59wasVQAz77rJgLdD4S+/wVXHLxuO3x8Xk+TVT+LC1ydMtA
I5cjuWrjnkfmetEZL89QxaSx/WqkPHrOEvXZiaVmY+BK+J2cZgMs+eJ/943T8GTt
2lfkxasDEdGbOhKBytLkDxGzHGp8OEdmrkOenw2/IK2mKdn+i33XOkd1Jceg6pLB
fK6fyAM/FBtWEv64R5noYvfpBRLXyjpvBrsQtBcxnHEP6unzT/WtA0BitTQ4o9I2
5p+eF8k2wuRhsgic8d27kGFUfIzzPpU07FPwMYdCkQRfhOxLtqw51iDxmfaZEKCn
eAO1EpRNkjtUnzgJm1XR2crFRezXKH/lPlT9thK3Jcdeq6h4xYcmP9XZtWHFTfjF
z6RGkdIedkFZVetszOek7uBzTvJXETE82+4yNV4X9mSoUdmYk1RiaLzFaZIB11f9
LnF1LhinRxcc1GCNOgq5S1G6rgjiwpCwind6F68u9yITBIBhvsyZL/6ydsYMFsLp
ei46IinGLMhNWo3OQi20pZfQkHi7NAlI3sfY5pKIPwvyxbcsxEBHNO+Bh1IiqNwX
cw9oBFvaQKz8Hahqykh6mZdnT/lbCMGJGmRIWfhlSXHuSyOTA/Dum0plphpkO350
84fCfV0/Jvb7uiUd/DGJMLDFJFs+qdlonj65RfaYHDOh1nxHvNTmi7wlDCpgrnGK
8q3DKRXwCIP83PgvUDg/SP/nTjiMOvMZcY+Q97Gkqt4f/WXfc5Qt/tbVdnC5T6kl
vWnKXg7ivUTwNXSwQTYIj1ER70vlxQa3B1fEZaFLQOgWawrxYtwXMV7/TQ8LwSsH
z3EN/mKIQ01Uxtp3c7b6TzaWZO0bRiGlHJnAzCv0ReQ1IAX03uS6EnyR+7Zx5loA
WR6ykEolewDK5kLZ7hnrftlsgbKMzzeB3qTy/tgRtvmdnGe9aw4fh0QUt+ZNwvU+
aCJV8pTaBn2UtzF/rJRZTOFgsgxKLIjKRogi61fqmjYCrSMfJxalXTWedNIFpZzO
+J7a4eCCjiwI/MTXL+7pslUJtRUazOchuDMCKsmPoRpWmjwx3efx5YmPLjPC00oq
fk6E+AngGBB9a7ojl2r3R4VLuzWnMlwp3m5EH8Lw/piY1SioOXWGUP2JyXvLwj8f
cAkQSD1GBek+gt4vwt9OGvzVxFMrx0r1kw9ttNwkUs+6LCCSx5URbyCIQVx+EmB3
mmoYxWZH8HJAK6V1HeCnCoveomnbmgmg31CZ97oXWQVtokpOJJdbYRFOzC9zEXfY
jQAwtDkL/dt7eZsADPAOjqOiSAiyW6UM8tqdQh7D8b+flypzLxPYB+K3V1JF4Gij
5uW7VvVpBRgAOWt+vV6gnBmugAnvFlLDDd3VT/vqu/6ZozABCEgTA7x8zJJEEu2U
VXAfPCNvUcYt1K8oSkf7IiWq1JL2nif35vzv/Xr1vvrwU2MYZ6NDySTFBfLvGzOL
dldVfT2AKlXgo1NTl71501DMTlA1KN4QnNmJofE+UX7xUHr5kOKGfy4J685B8umN
Rj7R3MUhGKIzxXPSRJhYMXc/uF4bEAru1pxAiZVgYv94ysY2brPJ5MZHZ6jRqp40
PxwHsoLUMbuYwoPz6zJN29HWr1cvznzwbmkWXZUBQ7KzwCtvc/YbK9YOxZxmoGTr
K/lXwbx1+3lg6g/lORtV2fqfax3WrpfuuYYaotukXaMVo+l7Ldj9/ryPUv/mtY7r
i5/Ja5aCbYC30h2QKTsr0kNEFcNKyCL+XTxPYjTqyo8AZNNactNt5fJACyD4QEcd
+3PGIf70DVccI3pA2scSEdx4lzEbGkELRmBdD9MBhX61GK+Wsdx3z71zp/mbb9jW
eBonxk3VFPAqoT1D1VPfNq0+0N79QAUp6YK5tzodihWdvVDErZpjVxKWkChfq6vb
VnMH9eAztuBILPcjp+zfdu8bkWnJFxEUd2nKFSoROAIZTrFZsbQDEnxBhFP5DEIv
wE47NiCdk/U8DXL0xu3Iswps4In057Jxm6Y5GoNpPbYepsR/W76eNeF984M5nhFy
rKbEnLy0C3oQECPde3Q3rvnGxVQfSpf4Ht3qx5GpCluuKwEgf4OroKiaUMSwqYgf
4VwzmqAS4px7a0WVE3Dg7MBhXba4NMiupMnfdPYR2HPoPg7JQGOTGlhXNpjAEHfu
Q4iJszSa5enTXC4bjVCt287AuWrvjgAV6R4g+NKXOFnnnU1D6Sjumd6HM6COu3Th
suPKgyUSC9pRfs/fezx7MQP10bNpu1orb3kLf1wu/jtlzrwQLNGbtNBKQK6LKiny
H00O9F7ZtivOj5dcgTwY0hRSgE3W1v6K7+ELG8nU+ElI9xHTc5qSogrr4sZDY0bA
o8hnR+PKe/iCjIN48HKGHh2oTvXwRDQ8jOMOpa0s5BBgBgaNz8+sAFO+xld4mrpT
InzDLbmU9sL9K+oPIBGW69OFZ3CAo6kXkanBh/C0SZuRcR7ia6hviduRPl14Xy2N
UGJE7Po3IQUXxsZLXeYtyb85biIRzpc+PGGJ+ZwV4N+BV97j/Ki91euLSSADBljI
xropbYM+eTAX3I/ObicnBd9xBQSjY9dt1SCTMLEuzerlxtUXH/DDcywhBDMoPuMk
Bw/boessXz7HxaHopAmBpZqjkRcu5GNx+UKaTjspMNbqdvLFtQGCWjVnleIMle+c
IJ/RADVd7CUuGzs8YWcJPfr6iQaCAgmY8A5wtv94ZaEm+fs77BFnX0tfrhVf2dwf
/mlXq3q8C4DMC6va+7YZumIV3DC9bRgWwm+nOBcHORCrTNagwBPPizJMC0hFdgK+
rYYyVFXttQnfTOoy26QKyNcHy/m9EkeEw+EE0Oj/xMvHMBRDOg6qjfM5tIc7lPI3
R7XF+/TuXG8z5v1vimaxsVvff6gJTDXS2XoRafQW1k4elcNZq6jkB4gg3WILvHl8
Y1Vyuj+iynyYgLID7eUdj5ClFt/0+u58gdz/G9LD2phwDdAC15MX7Gt1SmMdagH0
MBhEm/Nri5SJPgrd+Ux1dn8C79DoS8gwRV7KGehb0291mTH8qYbUov2wJDtRB1cX
JZz44Pwp0gCK42viPikXW+N2y6BsdPgdKeRjEO5Dk/isfrdnZFtT+tjEk5iGIfBO
o2rmvcIYad9A9PCOGYhCSKQmwZOmC+/RHZ/QNq4tXA/KHhQfyqTiqp2+ggXqhL4o
l+gJNvhYCBVRZkZo+gy3BV+Q+UBF/Ddr858TTyblmKE6J7R5vNfEGS5tpocgjwBM
VzBGjRjimHuf0+eCpELDYq+LW9yXzO1euDdR7773uHfenlgFDQCWcleTYZ1xIWTL
vHKXZP5LPLIjIgq8PH4NkqeLtcNAAHurPL3OhAACt5e2KIPo1yMEdww6TWkpKNmj
IqT18IMXr8HO4s1pMHvYUjF3r2dUZWddqUtufwdwOpT7jNk7wJo+c/s4Spz0W08P
zYYWhAR1ofdHisK78aim3K+CFXqMZlToZZeV5FSIcA3m3yJ+qU/HBAorjKLVl9py
wPPBWxZMwlthGjsuv8S8xaRue3JjgQ3NjVhttD2JuIaQmyYaT42IvGKXkDQQ//0f
ye1qlSrSNFaEXBnYt36pCH5f9qmX9W9CG8yZjl6PiP20iOv7X6TNjtUxZi/IDY4V
G0WJGheLDpcze6f3FBdCdd3juGsP+WJNiluqHXncASffLlKrgub3R6Yeod/ozdf/
4Nq/U34Gd6/DcQVVObJbDTl+HnCI6UkDrxal1w3/pi4AiUAuPT4bGlHydHPTLMto
JpkISFyV8ZDnnImQXLCY+7Whi8scOVTJHwNPuDqq5US+gLqqB4U8QeSAAm06u3Rk
wVPzhrAahrapK9oBFOkSnamjItV3Y8Rie7j3nzscviwF+zZpvRwvMEjXqStLuCdV
kR7Ynrci8vlPIiaLT7Q9M+CrDZzS+mukdbtg1gvp7UuR1j6A2G0YyIAOdc4DAfN6
BgHcCAPjm4dVO0+Dbz4fgwVxXGS4j0i40D2+lDvIG0J3ULZfkwA+wbXlx318q5XC
rU0oOav+jdTRHvWiIkxFkcc4SZTVxYVOCImgVzWcdqqxBsGfp8BxV2T6FDhSJDxz
oWP53S+k0pjUOeI6PCJTbtrJ/EHPalbecO0GuNlDQrQonnVsza96zWBLr9tKvSyx
GAT2Khbg8IawKUiWVOmgJP9IDV8yXRdfvbMdV46gR7zuXKslvjMlNDWiJLT40Htg
nbHiFy7QjNdAwDN4vb7Kz+wQgFqYJ9zBQqB16ej3vpXBnuUOEx1tLHnGrrUGksSm
wyJU+tA1vI6eI2krg5iKxF4tIz5ZnSlMenIhhx5cOtg=
`protect end_protected
