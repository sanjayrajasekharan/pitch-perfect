-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Tfejh5PE7ZAc+y35TUQipI5enbn5qBcVYMjD0PIHoLo+fXflRPLymBYBJs4SlnT/
b9Dd9//0BFva9FH1YtR8d1a2nob1fGkbvjpMxo65fAze5VCTB/CJ6T7Pa2OaTnbC
y4hG2fhnm9MteyDCS0cc4vL/ogsbNOlLBlN1nnZEuB8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6062)

`protect DATA_BLOCK
PZkQgqWzKymu4+Toc3GmU9lHOOedGh456gWnTaU5inBvnqA2bW2Whb/2zDiwLuzv
uReRTFts3a9jgRb8ndnlv8QCN3I8A1di9N91fJpKqwy/1stCfCsAktXluAY+NPvz
X42/doNGE0gE6+Ic+uU+NdMGoE5f68InbWUpbrUPmFrS5yiwWTKxjPyTl8O0+1Fy
X51a1Ff/uEqGlVB24UxeIkBo+9GAZloFHCtY3d9HmRyfDolgD9Fir+UUQu2DId0x
QEP0VYr7NilCuy+UqSUeb1bVhmPZ4vGUMrbGcXoy/svVkHDZlsKE0bqZ/XJLeNlN
ta39fsmDLUqgdOdSm1J9l35TSKUz/2A+6O4x1Rmb83dNzdCOkOa1QLU4VtgEisJO
65IgobmY/3ZTu+jit3F45qkQkGhh5Ot2w3xmY6SfQSUkDItjbVfc+5cm21CjIR70
11HiupMcKrPWoG+/9LU/ejs8JIV5k7ZevhDjgNTaSVkZK78KcP3B2FmC+HA55Sda
y8KvGkopVui+x+31z0kOc4AacV0Z7kNNsuqd5bUK+6CWOBpC9GBA32rG7hSYN7xd
4lzBcbs3vGanPN2aUiOUrdSkngwM2WH6mxGDRiIJj4j3ziddKwH2me1gfgSfZOK+
NfAggvl+B5+cVwzoO6Oq8bw+fLBa2LsIsdfkmQS9njAqpRu8HhLpw3AJkxEfIJgx
dTMmrIsLhgl8f3dxeMAiUmPnUZylRtH2VU6I8IFwADa/tt2bJW08o/mcIxAvhYbD
tqAcUdGWlCLLm2Dwo2J/GenkAGCj03okOiChkVKwYpVVk/ktcSv5blUZkrp9zuLw
jX2WVTqz0FqzaLmHHeytXxs9eSlyz2PgT9B6vESatxsQ5ZGfdxoQHc9umUDmDNXY
8a6NHwUecP/RZs7zT+ZKG7lqV+jE5Nann6E7QCSA1x5zX3mZrB11+dz/SEFt0KWa
sEngbF4tqHTXux/yRyj8jxGwZWT+cfdAhllxJ8P5217IeJOEPpS6Q7BHNbfXvpAZ
DNxZg/FUJfqH/CkRkofSeGa9EGUDyeumzuTcwMa0jESsBFKRC5A5jYPduYkxG2hH
exHBuPinMu/X5KFNmNzKynImB+/VvqQ7bFydu1GWbroneeIl1R2XOJL9HhBPWLck
ygrnT3dWmP/RBsJkBxkN2CoRn4ZilHi3aKH57l0+oopfv8YMK2VZ8H4AuYgXAwaY
l3BIiLJP9Nwx3AGPFQ0bsgNsRdbA2BNNZmmRkF5ETGNDBKTcCx97BEBFuUhgzyuX
UA7OMzV6YLChO/U542U2ErjFxz+7A58IRQ3znwVdzHEXJ0mUW1ext1XrVV4g1gzR
2i/Ejd1iGlzWlSa53XYLrXtBwIodojaC6X4s1q30HdrH+WAqnF4n2VN+EEN3/0l9
7p2Rzms8vNPrQJ/aXlMFqEkRPImvP39sLib6yBQJGbrZWp+oTadga0GI1iMNn/xD
dv5B/6c0OzlIjYEG1K4VpWM+ThbNiHXqvnWxOExM83s1y3fnOx4xrtao8ZLvZNUH
cgEMR8WLNFr7UcmHiwMxcu8S+tTyNS0asAfitow2O2/mal+i1yg9Gn1d9hlTVnHE
Xx/UA37R0sVFx9P16WrGx4zm/IKJC7EnrQpvUf9tyk+9LHIY85MRdCdnq24TKcb2
0DVoZzNc22e0TJ8r99uL1KGNSg44JWuBmIDaLbMZbh2/KS6qSsh4mm3HsJKxGm8G
vUvJsRdNekjr1WBUIEWNk6bBIYeZfzvOjd9Q6zg8cGk/Nl6YqH3QfC27omHEJC5J
33EWWkK+6Yl4ECpJaI0q724lxJMMs/tAlCM7OmRf+zUpIjgA+JUCJ8UwQMklt0v5
iTUqDTFG/Xggh1O2nuYpNODVtoRJtULifwcl5ZvD9FZhela2XmLEDTO3ifnEZPBd
99Mz4Q0Tn6hiVoRKYw83+oQkev/UlCBMh5iKe2dR8/YFt7R7vh6X28z/yL8FnRPm
TzL9i1PHe9M65TCJ5VQB1JD4rkOS57SiJAqnosmhgDebmnM2vqiQqFceT5TlxuIz
pPd9LOZxxiagakCj35tGzIBnyxYyw06b2/7N01CxKP1vHu7ybwehU4TR9MSHOzbG
LRqFZH7bIlG03tRwOPG8qkKAJWFx7Ap7g01FLSVCanXg/FeWBi3VUDRz+q66FYk8
G+w5E5gPzcAe0yyz0tr6ilST5eFBmtGcdavsFx+NL9cbjxZQk77wYBngjFI+xgbX
iYYDn/Mnj5sld8JIpDFgNhH+wOLLK5LBUWpA6KlkFG6qV43ZEPSlCarzn5PppO59
FGVL+1qpr+685PSvfFnKY4ou2SsGrf2+fR4jTNKKE9z498pYIlK+X0AoxIQx39M0
BZgmV32aTUKrZZYUuH/45biTgwQfhVZfmEjJYMIIt8LeptGEoCSzsYZBU3nwgDuj
tTKEDRz3UzPJu8tNDNOIwyBuSaix7/C3MDy5lbe3ElIzHDbX2Q9fA0K3NrJhqYHD
m9aKxlnFmVzEyF3/Y/zlCywsI9jfI1CUvCcA9VXPBSezna5IiokvC8q5FpQnSbJV
iR2F/529QcveFOBM2iv1bZpL7r1bBcg5z/9vd/WM9puYPFSAcwVv9KNWpsThDzbt
tUMSTRBdIM3t/2N57qGVeLgYIHPDSUNUZ4hfizU5Na9Qf/oqQHtHy1pKJujyB71d
zIj9itRklPYQ0qM+o1oTb6gyUC7qHc0vEqhjG3c4s/GRWdDjPzi4ZH+sItFdG7KG
tTq9/z0tnD7OqAJIKVLzYYIsz/SfwSBF+I9/ZUmZC7o7besL7/p2l2NYFh3ojNk6
xRBUF4W9r0XRDoQwdHmFQFz6wUhRubMNsQdDs0BOau9ViuW1tNebw5IeJ2Vpfl6R
8JkiPrqNHXyRT5Ec3cG7FmluF3BxWnjwnJvH7XuFsesL3DmrEHJ12UWHK4bsoedA
RyaKxPsbsmOiAuse5h9wLP2dLgOB/uDj+sy0w8atyyZE5rix9w3cJC2bTRmk56Fb
6DU6d8VXGeoD59NAFKQplsEmQ4y+iWb4ifU+9PBaFUT/lkv+BoMj2zAwXj1c8M7h
O4Ip/gXHmmxGo8sxrPXDpxWLCpAtY49tbO8aT6X+fXvbd8sI80lHej4Ckwd+sGbI
BoW4sAyhCR4IuTnVy1rSTqO16Dfb3V0n30Ntav7akZHljo85+ETquuJhY0fSbz+R
Mr8hJaNyWfu0i39oxTlRXAi6V18ExhLW8m9SmTXvuEdXHz3lHuuQDixh5Umathsp
XrpXxWJx06I+CzxkG2Fzb2xw6Gd9YefAyrnXXTZIlnUmdCzEefyx6F1MdY9oKAGf
V9QdtwKR1DnrETeu9PqT1Hcydm/jPV+zdKRB2his3u0NjZFOh5sf4Zivm3vAZM/D
rKAhvvIvwXOUfnQGsUeaDuSwmPy2LNb2r/vO5wzJfib8iqhWKuIH0w0gNEJOyAcj
e7gwrW/A2mq+R0LzhjU3Yk8f+8W3ccRCbB0VeQaJtgNGS9nG/ejsu49mXebd2LSt
IWJmXupQBgUqh1CAdxXU0cmXHHk85skqQ56VuMJjZlOQrugSg/fyIP92zh+GSiPx
UcCnoW+bhBiF3ud4kMhVPERT1aANaqYjYofcUpKrVnt5EwnkvvQXcdSxQHnZvXjk
l8R0uxp2/kxCCZ6eEQf/z8OZtbzJ7H4DqzTIkWyJg5GHNT3Dq/A0s6c8ITR9ZT3h
CUSU5cJspciiZEq4MJGBb6mGxPsBge5a2qvdT0F8pauyOgS8yApg3rUXvpOiF6oF
S7YeOHBkB48XM2+DUHXGvPcz9s/qDIPgz25wUYrqkgd/BomYENeGlJGeYvM36C1T
SO67bCgMFBpm+whpyAg4wJLt3syGBHnDuj66HO/TMHCQwsiq+BJutVjGzRbsTaSl
Y1Ki1S9XCyaUi/qlRH4oIM0F7QzLJyJELthqbbIiaf/89bKqZDg2PZz5uGt/47jH
pXxChytAuhOOIVp4Io3rNd7Zj2rVe8LYq2G6G3mXfni8Lnzrx/x1IhaH0Ny2gLGt
0PYRGaOSHbRKr+Rgr40SV5ct+mwgSR30Bo5xb0dyTEGMAiGfPYHuC3LRakfRbqSN
0l5p5aXogItVZl1QOa/LLnBZHBXGmZ1Ik+ZSqVdhsiNDdkVTH103qKY+iS4652h9
m44SSMRmfpFwJD3vTOOP/3eCyYJlLC9I5NdTrbUf1Ksuphv/0RYVpR0giYPNsAGG
bApMcdt/xu1nOn6AGbVZi47vcDZmDRSblfOIJZZxMAQK9lW5+fn/dxR7nKf0HOIE
eGeSKLOiNBtXvXlRJ23AxyNlkcSYNzWzD5gWUw4EaKVWphPhF9XZkZPbJNr+PHKK
WKw2lTBCFR7khZP57gky/AlSNBPOTUJ5kfyjmMuvjrqvJfqIDb40JJXfP+mhwSPO
XaBugPiBWmjO3Egb8Ve+Q12chV8eYw86fzgibOs6dieO3eIl1ynGbwxw3mpFSjXg
DA7zi9Mw5ExC9+PSNwpB6Jmt4kMO62jOk0PbsWjQWI2kCF884E+uK1SdUKbaxTiE
/RssVWWF/p2NeeggVFz13kH9RWhgITXGVmkpDrIxX+OCbtlHEA+Bqmm04w1V47Q8
tp86UTMG0KM6iAo2W8xkMn+PcZtEP/15EVPVnVd1t+qSDrYZ/Zrntt1X903Srj2b
quDUXJX7YYO8cHc0ivIATB/+x0q8/JDjIZ0wxNrsTlhF8yZMt+j+HWxyFeEYq3iN
dfAda1HeyDOYmASPnfSYiLCLXlyoENzs6PYxcnisxhucXpgAaGL4q/6dngdtVPYk
Hr1sM29qex7/oiM+VKKx/FrGbdjAJ4bkVVKjFRYnhbgbqoeaXUIDSBacHdAtjU+F
P5gVic+oLMWx0B2stoNggUSXjFL1Nif0OOYaPGTJx4tvZX2wreJEzr17VWyiPU3W
sMVZ86nw/WmozR6amVoFmMEk0bU4mLxyHFEpNWl/34WbvyVdl50vdxQJU9t+sTCV
YL3q5Y3pWBxRrtn1KOLE93izQzJKwGTK9N3Fp8YRLy9iYL4ldEN4n9TIy8p0wgq9
kiEIYXPFKqryegJ0aloI9NY3yA/gD77/BTGJvyiuuKVqc+jjm4nLvkP0YAxkW0as
68Lform6d2dzBLitheO2GiiCexeu+kAqQhCZ17GONxik24rfTQYyy0BV1MJB0j2c
gbBMhpBYx+GtFT8wFBd3H5fJvmgKDrMpByeE4oWRUX2Y9DoRSztDfcZT9MEKdM5z
tdw9hBaE/aXNeW20hkMjRtDtkkiojkve5leYgITavEev5y06oacWPM/4m5zEv52y
HvyT1Aw1kH57rM4KDg8W0desnjnWtMOv5dmMJxMdSp0nCaOKGagNJR7fJj+i0Chk
3UxAOkVJwwgST8hafXcoc/8GLlpOGsnhu6pnb9o3kM6wf9zB/Mtr3a/EC10EmY0+
ueI5js9LTpcWcQFpcZ2TRbON5nwkpitPUXzbCHB7IIp4cw0I5vB9/WAy/yYtYVtJ
wAR3IXXS+Cckob9q6IdE6hUFFNyflsSbzbt01Lw6MLg7XY68Dom+0zfdvPJVFLLv
f+qhLVDGGQmd5rkhcbnGznnIkM1YN8/2YWIAHrwVt+/7r+WBzqtO69MytQe6IV8M
2iJt/uKG7SWNsb18OcWhs1kopq+tzpAXJaBVElgiXKby/peOAjzcj/w6AArYrhDC
cnOsQQdSAylJODXDg4wIEjOsEUQmeV2+WH7yQuBOpPBVT2FHi/BCKMt0z8xH0UJw
0URImHo7b74kvpDepq7gyAuj9J6/wmuOh2MB1TLJU2OB710g76aZCPuN8mirxYkl
/6E4ca/MssPYluGXRLqzVmTY+m2pVSYm+x01zMd8WwoI3xkexg2HLkb+yNDHFiSA
j8tujTZlNP+3lKzzEvg4mlgPmoLJhq2uvOtANi8RPvUFkouk8el/6kbnlqZ4gSkQ
TbMCQ1gPyCbHjTX70XZeTM+diYNE1asnW+SvTJPD9lCpWvYsqzxJDQ62HwJgRiCj
cEJGbVyY3P55tJGQpJTOb23vbCU3OK9TBBfD4sKkS700x5KolperAvbKGAgWzrCg
Z1FrV3sT129afT1QyC7txCqndyEF2LEqOUyVUDxiHx8wI4OnFm03qUWCnb8DqSj9
kgEIApBphAsDUSQvJNrkin4eiphiPe8+wI/vfNh83etTfpuk7peYX6myg+rB1gEf
k2x5fNq+ZA8mXSYGxxPHjjq3qUqbJ4KXU5AJBmr0sdPXC78LmEmSnsN8M1TH6ywF
//4AbjjeGUfUAcrvYMlb530u9I85QYxla8E208ef3U3Bc6/f9RIF42kXHqcUl3LJ
aFIUln2gughSj/UG6FU73EeMpCb+mAB5wZGxg7ecjiAosv4bz2oio+NUdEHJqDKK
fJrUIx+eVRRPOYI2bRkOkjtcebYoKqdJRNsGprsSj1h6cEHYBUoUQCXtxV7V+gVs
tvNrhDxgPfGowglsBKGWHJAmZvJLq/R4lLn23jEQXAQvZjqXZ6EFQpwTKhk7GAuk
/ESQhe8sEZO7c/psRGnhq2MTfa9Lx0yZILImXFVbNhjldgq2N1Bg8oOieC1CAlIq
XwfZ0C4+nmnYEHstjet86mL59U/yCF9mtTfcVcs9YKf0uNINKqLk1ETtyhCLEfVm
+LO4ycmFoGiLMv3XjGqDXEtksUnsFbf7dhnuaPJWzIcqesn8+h8ZFurRKYy4HtYK
6hI5EnIKpaosFO3SjkbD/vpyaDc9RrKlDWCXSEYQTroJ9aYPDKOAzwQAD0NhS9Ub
GY0l0gd8LtYBw1dIGq4LPoQVcg2wddL90Vnu632vh0UxyOgAPulBkYUicl6UzUvA
ONTmfyiUIorFv9NZP9VElu2Zj4ZsOT9F0jRvnSIsH/TthBUQ9+2iGR4urrbNS+Gm
URbSORYg5oaxwaSU+P8NZp6SuQmMDVqamgDduuvv4kvc4+64Sv6aWhvVIhniS93t
VKbJra1ehbc6mXbkp6b41w4PQqSTSjpXu/rd8+9IwzOoWi/dDWanSgfX/5tlsYgy
Rp+0ivX00fPOY/v4ZmTfMYXceaJvl//6+aChoWcVaozZK2yHewqgPJI+9h+PVQBo
TGOFKFqieixzEUSCN2ZKL9MSi3R65or+ro5sfd9Pa45AKLxgye/tJJJG3iKkgzkq
giHbd9eKEpzPVgawG57cKgAMmDuwe5NnR7MES58g03tHjMBTxs4ZD5mAsCylbVqS
zsNhMLxJuOfkx4VFajTfnv6+v23PqcAvbh3GzJdXeg9Ma67pC/ssvdT0QcYNQzwR
usZFM46JzRCk7gNwvfblFEFkgaeqi63GMHZ1+kgnqFa4ckObWo3lEtziU+T3S3zp
NwSBlwXRfzXUJUiqjl9M8QMJ8eHz2SNCZnzdsHznihgNPKcMOvzeuwkSP/ier/TF
ouu6Gefver71mPZEp/RuG+Z7jIChpv270SMcy83qeNOFFkgaGoU4eJKOD5MML+Lx
1Pp2qIiXWP0+vTx+bVWLLLVfL8r+ESyNuq6c3dJtVE8B6ZlR77s83yAJf8+vMLvo
AmRrfHr8LZShkzgDNjcGbCX2vRMG4aBl3S2dO6ufhphMSiIB7dmeJJYZ8R+Rmlzl
NU6l8JXimLgH6w6XhSM6HCUvabDb/zyPt9MZEqxMTwNuwllfAaX51fFC3hwKrSEK
1qhxOCwAzRhGqiObOtREArba+e3NthgzbxW2/OWZpXRfS34OXeqV1r7h6CNMrflD
Xq+h99ZE8GYvkAiv+Oks5U2h8SHHuz3NUxfvUSfyeYP/rHIyYmzutOFUmBh5uw31
iNt2Pjlp3wzFlyg5yKc4rFbd1ECVHijndMjPQXkcBcwqXaWgVeqrR3oymagoqlq4
ZA9/hKYIGuho7l8EYLDwO6ZiaAq/uC5qijuYZTLlSVoNe/Z7sa7WkcufiKnLDl43
r1gZmWJa5d+gsYf8JyfdYx1HI1MRvsZjDZWyUP4uCyNTZKo/V+Npmj9PnAFJ6QWz
thyAcYFyWWukOaGIB5X+H0hch4m4CbOuBSGycTskcWXy9+e/KXartOnlzZlBSpPQ
pP6MyUCa0kd42x0ORwgWUCfs52w2Yb8nvnAYAu7IqqA=
`protect END_PROTECTED