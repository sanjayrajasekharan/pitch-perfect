��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�������B�ބ�y�)��X��ϡ�!遟� e�	�)�){���J�v�l[_&|�vm�P��\r��	A�R�u�4l &�Jx�����G1�[٥lA�W�2܇k�UJ�i7K��%-� �'quO9���)�����qIW<S"���#���GY.���s}�e�@7
@�6e���fY���;୍��
R&Wf��E����=B�H�����8��=�;(���[��������Օ�Xjh������
&���_�����%��xp� �YCF4��/�|`,�z���!���?�u}_H�(x�ޑ}�V���ʬ�mL�N(_A���t2��u�%��4tG�=(�
G<9�����OU�)����6).�rXU��.�dj۾��Ivp�F�]}��#�Se���>�%"叓Ս��짋H8��q�P6�y�i��%��kr�q�pէ㎷�[[�6�g�J�"�͖.[I�S�6O\�>o"/��` �xE�*�r�ӫ��,�w��LW+�}�����[zA�>�*�#��,��(@��i���'���^Z;��è�JL�,��/����>��E�w?��,��
�s_����[����\�b�o]���2C"�2�o�qAv���<��,��w�-WwZB6,���m�����2!��c^�)Z�$ ��b�9��|tF�i_��$�O��A����a6Q/���50�I�}M+��n�Mؠ���d���7�-��V��
&)���,��_
�y�&�����Z!N��O�f{^tJ��La�i���3�(4�֩��LEm�U#���A��� ��-u���-69.�������<H	��;"d�5����o��
:�&,^Wٓg&��1m�M,��G))����tɮF���At��P؝D%�����ֶ��к�;���D�.h-�U�}��e1h�L/��dr<C�*�$�=m�2��ʉI!ٛ��;n-�)�d�4�W�g����i����?ݯ�BE�)��%���oD"S�@�"I�<�\��P��<THNL�B�z�NV�z7|:)�'m��i�n���+���_��	k�蚥���OP�3l��]W�5������6ަ�J=�E8bG���^�O+GT�\��؞��߃u.���_s}_�S�;bªo2#���:�����f�	ڏ@6��������
�3�)ߴ�V�tY��tu�Gs���f�U��?j�⎛og�y!t�Mrp�u�����`�m�JH�BR��0뽨��)�B>�9��}�����T�x�E^�pX7����f�ՙa�������b��W��u1d��fX��9d��\��sU�� =�]�g�����R�����Ps*Q?��U��l�]�����5��ck�c�F!���o���3� �:����M�$K��By�0il&'w�1�ˍq�76��7KH��~`���b��|�R�<'�œem�qOfp$�nx��(�Z���|'�kʱ����D�;|�c1`Y�u�2
����K�e��껄�[�K����\���yh��h���a?��[���o���/�z!<�
���3t�3��Q��%�a�5\�2�G������X]ޗ��܃/�+I|� �>//c��a0އͰ��m������h��=u<w�}	�f/�K�mF��Q��u�[�������=�y�%��zF$TKI�����i�/]����W7$���Nl[��=Êl{�@#8C�d��V!ȓ��F򴝓���g�aِ/�EJ�pu��ԭ�giK���	�e��ق�_�X=�_GN,��ÿ�9����!�D���-F.���l�/�<�e�D.I�D���ᎊ����I�7>HǓB̚A�7AF����4i��D�؎F!�u�e��$��'���]_������8	�ڂ:�39�t�b3��%0��V���k@h[4�d# � U��[S��n*�+��Q��O�i���v��^��04�p�;}�,���za�6vo�������Tc�� $�	��*׸f�=��"
6	9�1aC�{.(,5�V&	sK80b�>�a�u�堄%��bJ�C<��ziŢk�ܕ����~y��`��yL໪�^���l��{pl����貛�W� �Y�� ��=�`��	����2�L���{.(Z�`�g�o��n�iՓ��`�Kc7�QGF��Yr��+�;r�^+�s"�&�a���!�#"�BS[fh��?�o�1k	�>�f1��(jEk"��P+���3�I�>5��4�E�lԫ{{�6�*�
�vt��	g�4������6�I6�gʙj̅��'Y�y���L7���j����Z�*��2nÑ:�P�v��"�}�n1s΋�M��*��QC3�n��H�2���)�l��]C�z[�2/3xt���
�:E��Pfӄ�x!�1����?�cUQ��4�(�8gi���рdd��ڑou9��=uʶj��eM�dl�]��5���k���"J(�hV[<����Y�LS��������8�J=�)� c��S�,�YC���BG�Lc���!�$��߶09���ҚuLT���\$���8����
`�ugC�7���Iw������4*�FWY���*@�$������n�H�\̵}b�ڗ�΁ZY��'ݷ5ckh7�
�X���:�+�~~7��a6@Y�۱f�f;��hr<Vo�����PD��:�[���v�$1��2�	��gc$>P)q��~*hni���]Llq�o�m,���n�Rʴx�<��P��0����rd��V���k���jx�1�:c�OO����M�CG=̑�%R�[}����.� ��8p���4V>�`�5�����j	K+�&+&@�Y�3��(&��Jj��5$`b�ן}'N�@F���T�u��L�.�	=E5�մߎ��6�?��}b~�E��S����7��kE"��-_����z*0�3�I��������II��=��x-�� �v_s�������F� ��;$��k�>�����>V��f�Í0.�=�ת{S</Fk�l=�K�og�J��TWC�"TG�s����Q�^�4�H�c��Q�MתB�q����,ݼ���Ei ��-���`笡DEļ�� ��3������:�%��*Е{����; ��+{'B<nfΘtƓY��7�{vE}�[d���vЃV����Y�ϣ��"�ܴ��X-/��m�(	y��\n�W�����k����̈CV��Xu��rsaT ��Y	�:eX��~��%[<�YQ/�(L���*�Fڶ��բ�w�¯,׺���"��w�`	\�
���-���n�P��U��S Xh��R�-�[XGw�Ԁr�F��۟���t��,�E�^lM�=��B;�ܙU`��gF�rm7.�#@��>����أ@CΠ>���6Y�U���@v���NL�T�	>j3Z��J�O�W-8M�0}��j�y9��b>�U��G����,����*�}^��yha��w��q��.���֛�X���{�
����5n�b�Q|�U�{�M�G !O�G�.H��96�$�7d�^�I���w�q����M;6
I�_���S�����a6��A��<��UDɟ�#��Q�Swkm���mn��"����hkM�j�"�LƮ���mֆ2�B���R�:4�7��I���<����K�� �:��N`�*���7�<�2��K����Q����ͩ�7��λ>��*tFQH���	�i��j���^�W
ܚ�g.H�?P��W@?ԊF��*��u� L�p�dM�*��x�^nѬG����n����_��,�����Ůb��Lx����Ѩs�� vl�+7��J�R������
��;�d�,��H?�0?o�����5�{8c�#^�Qr���4��k�&��Ὦ�r�L*��ʨ$@�H��Da�!��q>�c�V0#���:�L
�S��4�Vwk���l����M���ǔb$[�xA�g�VO��&�"A"c�[JT�86�qU&v��Jٔ���f�����>�=���zb�)��nÙ/�
��rB�َ��r�o��ۍ��&Y�S�����>�i��i���T��	��H""c���Ÿ�S+V-����������\"|G��bsM��`D��C����L��c��p/�7A��;�l����l��üQ��`��F[X��FLT���dn	(�bܤ6��jH�{L	�Q�I�n�����U3
�6c����]���HQ���9�Ԋ��=��<E�#A�>Lf���r�E�s�	۰_N����8g��k���.�
�}9)P��|
�J���dt4���K$s�)a�R�.�C�2v��4�Vz�D9�7pp��N�����и�,f�\Q�f+T�q���CKE �;���u������̬B%��sz��juŘ`����sX��ϸT-.�z��u.��AZh��Y�G�S���!*�}��^X ��೭*ʹ��#G�X{ƚ���]��W��nZ��in~G	�-�ŀ���TIŖ}y�9�|F�̈́cuPc*��v��@��H�{��о����s��˿����ZQ��G��)�ԡ��s:%�˷�A������oQ��_�!vf�p:�7W$Ж�x���4��"ð��8���}�9-2����Q�	Fk����z��L�b�Μ�<,�!n���ˣٵ^�T�=������v�Q��S�N�H�9	R�L�ϯ�:��'�Mv�����C�=��H�u�OMmf�d�'65r�������Ӆ�i����Nb�E�Å���
C�R pP��Y��5�QCoU�?�����)��p�/֑��޴3f�J��ic�"�t�w���+�i�UU��\�J�*A	*�Ϳ/���$ʻO����C�|I�y�����&�����!��DNM��J¥(�t�P�6����9hw�_F��^���ߠ���~��;R�e{K�:�k�A�F�w���"[�<*,��h�����e?��㨱ia��Bi/�4�3w���|!���O���j�|�Q��1�M���0���㺊e�R�5|ɔb����D���	�{��r��h���[=$`�g�`��#�^�t�ANN�q�asq���y�^���T�U6Fa�W�&w�"s�s}�~�.Fj�I3:�3�^D�ݺ	Z*+ApB
w9��>����x`���aJ�q�ز�xȟ/ �$������-o6�ti������!{k>�n�%9�aZ�/a�/#�o�(���x��\(}<���#�sJ<KΨ���*��+́u�ys��رs�<z���j��q�m�la�2F����%VR������\!�6 ��~`�.ԀG�m ����!���w�� �m�����#���J�.�.�Y�b:��0���6�XԶ�>���cX.�I^���́��v�����G��~ĩD��~�RS>����uP�k��Jy�I@GCL�81�߻p?V�13�mscVܞ�D�����|���*Rv\�{�ٺ{h�tu{�>1��G��c�>�RR0�ҷF(e�f���?]�"����;B�]��d�"\rN@Z{S;- ���}�H��%ݯ�����ZHn���j?S��)�w��uw)�w�x��ӟ��4�ga�$0��IQ�5Ø1Q�>��B��\�A���Iɝ6�и_ʡU�\�5{�~y�Os+t��Bn�{�5���k�)�Q�3���Q��-z�2�"�u蓑��~�:�g.q:g��hX皋�/e�5<$v������ߚ�{T
 ����FT_c&�nT����5Z����P�{1�����{�S-�H�� �_*���&�&n�D�J"���6{Ѷ.���������PV��;m�7�/F�|�Fp�_��w���)#�ۑL��/��Бn�9�\��a�����,����.�~�o׬�7jϗ�J'��V=Jm͔#���Ҩ'��t�~kf=\,�F���U��BZ��� I��rs�2/����ɲ�g�� g,ןʪ+4�j�\���]��
�xE�m{��%�ط@�~y����Q��=ߟm�j����|��=\����A���8����.�	���F�C�sD��v�*���������+S�lQ���u���w�	��c�d�P;�z3��������G��:��GI����BQ3A \�t��)�L��Uj.*�(�8h�g�Ks M���h�a��_R���&=MR�&+G*D����߳V�*
$\�<�ط!��*�'�J �ƛ5G6;�lb�~GD�D���of[q�iJN<w��=�B6�0,H���^��O���MM��W�$��-U:�����s��bE�c�J�[��U�t�� �c"ُ,]�$���:�	X��a�{����zV�s�hP��,�|?8"��u��iC(Ce�,C_5���=^��W!�ʌ:����i��*�6�agd�2�|6�P����~��S�>��M.�������X~?<{�3 �E�ހ���:�;��[�Y��/�SI��y4�/���3c8���;�,J�'�ͯ�兀��N��q̏T/R�pR*�����+�8l�������g�����P�o�k캐Q2@�T�MU�h��n��-�F�D���+p8��!N�λ��[�8p=\�6���G���#~˪~�_S�e�����Zhi,��w-�ƆƧ���ʧ؂[B(��z�[���a��â:���%!�Z����\�~N �:�s5{���{��\�B���)�u�`ٗ=�؋1 �V��n\U����&a�rS���bOr��ΰ0���}�>�\����yO�.��T��*]6�6�_�uQ�WuGk��Rm�֜IC]�	��Jod��c��"1sAi�Q�ǹ8d����n�����L��q�Ie6��4H
�&��W;A��)#�bY:8Y�ط! ����[_�����_5ܢ�\M2ɗ��u���R ��H���A�u���������=�"ߘ��6j]�/����������e�d'��D�5���e6�Y��Jg^�;{ou�lI�YR�2�5��W>�O�p�)�3�v�*��Q�dU����"*���!X�P�AM��������Wu;a�.��|"��:q2�^����y����j2<��qwU��T�:�������1ce�ꛆ Ü.�zd6j�}'z?6��l�B�g�M�$�����G�� d�45�/{�S���=L���e�	�Ry��ңD���B0�F�\�Ո���ݪ~���dI��_�C����lzcQu�R�]:B�̩�
oVi�����O�Q�fQ����a�ڏP."�����i���>,�Vk���w�����*2Dp2UJ�vp�V��mX�h�FX�W�"��$�Q����t_��X��])�h=�8:Q[$�"8�J�;��'qy�Յ<�DJd r|pD�p�v9���\?D�5��@~q�� x�̝��3^�\#��������7Ր���F�[��A�eD���f�S_�nS�@��~���H�`�2�.,���D�Օ��c$�l��Y-#��Q��C�j�9}d>Gf�jw���`��*���ˈ�!EQ���p�A	,$�;��{V�ܿ=��)h�b�������h����7l�(����?�%��\'5�)��HA��YLfe�孒������9�7���Xp�G���q��=��jz�C����
R� Ac��/L�c������
l�s����7���Ge�~�E-!�mp�
�{����4�������H�k��쓕1���s润K B�����E����P����}~4�C�Q��G�UNA7S^��qA�i.|XT�w������z')];�T}����!�����
ҹ�u�7�G6�{������kē������W_ �yY/�R1��l-@ߊ���As���>�������4U�NB 8�$��txD�l�
�u�Y9�v`С��Q�$I�(��a����)Vd���n�W��_�iM���ϥܔ�@I̔10=U�)T�T�����ʒ���N�@��>���Ӯs?�,v��{t>��y���(�'��;?�m�+?�ӎ�;1y�%��Ɋf�m�w�8�37�L�u[c���9i
�]+)Xr������Q��d���B���Z�iG��ػ�^�]7vcH��\��[H��k�.Q�����¡��kB�c�0
�u����
4s_6(�LBЂ0�:�PTt�c�ު�9yU}�І���9P�7�x����#z?�1(��m�68���A��.�I�?�X5�L��ld�b߸VlʿF0�Ut~L���|W�w����U"=G�U��} ��8#��f��wFĳo(:!��q	o����u2�
K��>�* ��g�YQ���|�>�Y[��r�؛+��	����H�_J&Kr57P_�f��f���\$u��>���*�QK&6�D4�l�]��Ȇ��uO��q=�C3B�H�+>HIc������[I�D U=�uj�޸d���c� ��:{�"�4[��9&Q����{�1����� v�y';��"�޵b��eS���NZ
*��	W�N��Nڷ���GF���霟�ض��gyo�e��kũ�R��*GkpݴS��Jދ��K��B�f���z��G		w��^�$wx782���l��1��p��2�E�Z��
���W���H�+�/������1��H�*�B9ڨt��^�?��s�6}���������v��g�NkW�2񴊟���b�ݚ�t�_�F�m�Xֺ�Ѯ�M.�SF�}��ZTA!b�P�����hsN�J�l��g)��nM���L����o��ss�,�?�������wq��g�4ȃ�}&��c;�n�*��a� I�Wϯk ��p�|���IS~_�@�p��*�HkЫȨ��& ۍQл��a�Iq� �JXY��5~�qH�����Д���,?�m`�5�VQk]�T����.��W4 _��!�>ѝ�ŷ��U��I	�Iv\+�04�d�� �g�7#��!�χ��0��γ���S<���~<ry��O�~�4RY:'Q8��X�KX,Yp����(D�m�3hW���N5B�H@k�}�yWOixPB
�ku]%+�f4�Uְ�,c[���&�.�æ}Q�\��˳t�����"�'�:236I�����B�C�?��Ib�SK���`���Ur���i�u�D�@�4`]��=!��bFk�{�l�:�(��C�������qyb}�۝~Eg늠�1�đ�sB�����u����R'T4ƒ��Z����|�,��.7����Cb�<7[?��,l'�҆!XI7%;Qp߂����`��O7�L�ud��ӖЭ�=?l1�|&�x���6i�	,�MeK�����o�%.@�\*��`�VXR�E���%�V��1���G!����_-��=�򳤲,&�\4�:;
�a��	��Vu֒�{�U�����rF��P�jLa���rO7����М��o1��5�ػ�\vr�`m�Uӭ���f�X��N 
����[ĕ����P�) ��Bw�����y�:����r�3�<j�N�ޔ��Tj��!���$���¢�R�=�X ��U=.mNʭ)XG�a_a�b����P��o�$���g!��^�(���|N���ʶʶ���������`�@C|VD�����p�3:)\�>���F��_L�"6����O{��H��R�Z.�IW�H	��z���^g�IF���8k"8���!Δ��pH����-��N���և6�ƥ��ױj$��Ghӌ�Yz�V�W��r;���N�/���y�G������� ,�^x�g�������D�_�BM+xe]9�?5����^Pjf�_�L`�t[ˬЁ���_��S3=���BrA�"�2��y��
@/�CEj `�82iS��[�_�-|E��f���[�B�d^���=�X)��)�L���fR�B���e��+��wO�^�dV`=�1�FcPv��l�'9�Z��H��Z,�ʮdh�*�
�Z������Ł�����˫�&��е�O��,�bP� �� ��>dh�"�9�#Y���V��i����0�a���NF�$�~����_�����Mjbx�q��\����I�nbMQ*�7e7�-���g����Oܵ�Mmo����8k�����ց&3�X����Uw�-#��A@$�в37Td��\��vF|�c��bd���g1����29+��r���U�Vg����(��ϕ��ʐHU���.R]0�ؒM$ɐKWSp��%�۩�e믄o�������7D́�c�0K�V�;�=H�����E�&ΰ����|��<��B���;Pg��[%vm>�"���A�J0G��,����V�B"w����}�1�����y�S�+�����z���V��V@� ��d:o8��J�>i��3�����L�(lcV&�9Y�.QЌɲ�o��E+���=�`��ϱ1>⽺0Z�G�
�pȴ@��y�����7�ĭT� "�Vo��,�'Q�1 ��O�-�Ѩ�6��E���Z*�o�z�����G�+�µ�p�Tt������w)�y��߽2�ə0����������6�S��:nM�����BvC6�����9�Ю�3���X�S,�>��>%��R��]5�Oe7| ������k�W�2�f���}kI[��6�~Ha	��0���xGA!�KS�t�!nB���&:o�vk�b��L\TG���O�4�o_������_]�l91����u\�I_T�xb"6���`��eNܜ���k��͆1ǆC<5��6�����((�J���f��M�g���e�v�8���>�#�;��x Ok��S�.{~�	��#��\v-��$���ʫ�mk7k4�+�;���(�mxZ�F�� ?k����:ۿ�@$�k#��|�"����)�Eb�y����頯�/���p8�پ.Ŭ|"^���?Nf�9��ם�+��ZЮ��V�*WG����H�i��5%��i��	��4����?��_�,���$�)S�_w�>���xL]/��m�Z)��?;�C�_xq�i0�L?-�O�WQY}x���'�$�_�������B{?3���j�Ǜ���9�/�C�p@9��^����N�:���md�&�
�#ΙJ���W�C��v3�20�	�� ��` �J$���z���>jl[�]�θ�u��
�@�V<Fid��%\BU�.�w�XV/�B�n��P8���,º�EXʃ�}J��09O�w�V�1�;W�m��n�]*CdCE(F^�QX���z�Lb9t����T��(�m�S}�j�~��H ��ɟ=|׻�T�2,ɗ��cQ�^�(OL����a��Mi��SE���)�b{<�S�׭��Q�M���-��	>٨] ƿ��9CX�����fJ�kW8�|�%6ugo}b�p���7D��X�{�,┢R�J��w��pG��6U�;(�9��P"<)�aWƋ��}O�VX�9��oRH���#y�f_E@�w����&%U%b�Q��t�]�p�W�R4Vx1R��/٢���U.��$������E�Ⱦ���x�S�C�U�u��٭���ǚ��N7uc�����`x��2�����ΓAC퉨b���y���#
?P��Z��׸��*T*�W�%9(bL��'����������Ҫ��'a�{3��B�D��.T3#߈|�+��JǠn��� Ī�d�p�8E�D�X��P�`�0���ϱw\s��3�Fm��-�':�@O��Q [j�W���W��������&/t��_�V���)%��܈�S=a����i|9�����u<���7Yg�1�m\�c�`����ю{�q��,���H��Q�9��d�6YO���/)�� �ob<-K���L������ge�qLH��-���QVѤ�/�3��%k�<Bp�^��6����y­�|�.Z���1��=� j��)3�G�Y�����12s���]y��S�II>�8}3����=P��έٵؓ������+۫g�ڶ�;y�gx8�h��(���8��l��>������ ��Y��r�A�-��u5��J��\#�Ζ{qT`���f�:�.����;E�j��>gZ�����P�tKz<ߵҍM�C����}�.j�0؎j�"�'�F��5Z��EÏ������ _�{�9�M�q��r�Q!���ۣT��6����ޗ�e��5��mT�2P��Gh������ut�O�?h�l��Pu�r����}zt��fI�R��R6,��	Ǻ� hsC�?�X��,������J�TӀ�X�r�]g����M���M�`i��uT[u�ÁB�r|�!�Ŏ�{��?�b@�t;� O�tN:���y������O2i�T�$�M�qd�W����WN�;��h_N��{���u,Bt��3�o��=��y�Ar"�Wش��2��F"�i�d��I��R�	E)���FR��\�J�+��zB��jJ��#�S�W�AZS.�_,Y�
Toh�K��T3�r��_�\~��=O��:�1��'h�)Z�����`�B��P-���O�4�x��N�Y�#�}<��ԵiU=�\��/��VY=�)l������q4F��)B�2+�㖎��kh[�D�2�J�;h��(A�k&G�4J?:l�aG�~��"�=�rٜD�z(����'m�v�Q|���j���)���s(���CS��d�ۋ	��SC�,�$�%��U�����1 6�(ȱ[�Pyגs8xZPÎ�^!sVEϽ�~R}�'ߧ��em�o�tV�����,'3�R�uAm 	0�5W'c*ꨟuS�a	h�+9#C���%/1�OB/�sO��0��\=�����e��V�!�M�%	��W�L�N��I(�TFX��bY�9S)��FH� ���R��ͼ�;G�&��&�ΓkK�%
�B����ꮾ��v�ض4���&��ݧH#�P�l��*���������&�[B��xHh/�^|Q`�|�G�<z#4D��W� ��ʔ��ͅK�6���IZ��5�e�M�E�/�<N������\����Ŋ@����kZ��wپ��(U��e�P��2���"�N� J(X�
�Ւ��Tq�k=����,8�:F�������	A��}�j%Wn/������*2l���� i�ؼڹ�,���W��gB��P;�)���ї[P��ny'!�uM�� ����@�����y��kު��ajd5��,�^�c��w�.z{'���'�t!�$y�Uev����&����G3z��U#���e���Q`n��Ш&�%<A�����`���;dr���E���w�uvod�T��&��v�qM�]�Z�'��~�k{Æj��\������a��XM�p��p+���q�7;l��5±�TGz��e;<���x�&�Y�UX}�R��#V�=<Ef`��N&�<Q�>��5I@�o�p��T�*��ꇙ����-Ԡ��0�K��+i��G���W|>4�PP���?D�x|�V����B��+m/��|Jq��I�'%��O�밣������xݦ�0��A6_3I��.襦��nO\ș=�LA��1!e�wY�;T)݆�� &h���M��(˺�I�|��[~�U!&��ը|7h�����K��d�Z� ��1z��z:}��d �dt�x�h�0�2��ς���%�K
� �H}O����<*hj�g������u�w��	I��][$f��`{ҷ5�a����e"NR�Ǹ:x��~/8!0�l��L��wmNN�ZbS���]4W(�y�0�o$��Mh��c��o�!2p��;�+)--�ѐ\x�/0t�DB����K�ZgD�������`��"����`z�ڍҨ�񓉯QNy����ʋ��L�Ϭ�FIq]#�~��j��7$���?m��h��bf��m����	B�l���ۊ��ztï>���#Ƒ<mAL�}�h�>���2ad�~�� ��i!�gVb2'j��8u�c��P���_�T~¥�6�P�Ѩ��
M�itpv࠲�y�??��}�I�G������%I�%(?c;r�A��}��0v���3-�/&�t��5N9���"�֡�盋�r��+k�xfUп��A[��j�������2�74���-Q)7e�Β7p�2��ժ#v�n�O�L�����Okv��5d����5�$�sN��.�����P��1[
�([�O��U�@Q��j
�g�%��*�2�c��x�w퍱������f�j�L�ځL/?��F��M7�7�X=ђ8��$�C��S��]��g��6����Xh�3-6`,��-L��<%���M��P@K<�VhI�mc[�1n��DK��ȭT�V���A�>�L�Q��%��x��x�kr�{B�s^Y�j��(�tV�?S4Xӽ�5���B`�8z1b-��iYg��AG$�x�D��i���4�9{�hи��J��3��d8�[��{�5�QZ/h|y�6Â6{)�־�4�'�%����b�H�i���oV�"�d�Ә��|��d��� SX2�Z2�����\��^h�͑�T����m�T�TX����!gٳ��o�#wP�a,�O�r�����Nց�/��N��V�NJb�v�����Ɉ��c�r�	�Jr~W�Z�~6b���1�[L�MQ�+��b���`v~%���@:����_wJ�T�D����q�_, ��
�%P��m4�_^���&�Cg6�g���ɐ�'ü�$�n���D7�@��	��T�]\~g���rK�B�fn#���MUP߰�m ��Mr�Іӓ�X����ܐ��醆	��D+�ve���NS�.����Z�*����O�2ZtwyEE��e����ٶ_�7��Y������y�ٲ�����k�p���-YȘ9\4"AǢS2A�c�3s~�v�$q}r��g���q�G +�^�9���NG1���(�|&z�Vb?�a�.��0Dr�؋�]��{��W3�Q���[�������ʗ�4F�)�RJ�x��C:�f\�!Є�q�����X�Pvު�hYd%��u���38�Z�(	~�`0F���n14���O�� 3?O�R��30孀����k�Po<@�Ξ��b��vׁu&��-�g�ϵ�m��B�G'-h�GL���(/��8�=�]����Ih��e��g_���{�0��2��X<��:�Ġ�\�Q����!�q��K7]gHk�U���K��Ñu"�N�r!�(��͛[�ff�|6��賷t�zP��NO��R
�N4�������W�֤i���{���a�h��ִό�z�I-�d����q�A1t�m�~�8���l��M�J�y[�*éK<��zT7��Z��+��0�Ŵ�^5��}�	�h�NP*ῧ�����)�+T�>�����