-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1dYAQ8GJw7IWfzxREwdW6d2hCUG4xqIOwSW5N2bMKkONeLPMr5xBQzHJFGRji034
PkKA1jy0UYeE7dALICzcEYQdQB9vlYETw26+He/rk2bANS5OhBL/kQ0s2kN54wyS
WTgw5vG7BplDs5X2pgaYl0lDGWVI+s7dDF5rxqIJzH4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 18320)
`protect data_block
CPs/73NHbz5j/0s8PDgToahynfRycw+kUBc8vV2S+oh6gcDqQKcYuORuO46Wuq6M
LhqxuSPHnAtq+XMeepuXLNd3d+oWMgiFHeLgfh7f/C4LO/7iKB6Cvv0A3IqKjVmd
ep8URTqKMr91MeKGL7xtpQDgmu33YgKJYrQ+EaVYmYtPwdrHyiKEv9bAAPPeRPtY
FTBt+x5xpt0gff0W0jzIu/O/YTwhJAYD3z0baY3irhW381j/iyxLvY3tdLM/VV9/
lcW1fi1u9vXEgQOPYAXxe0fGFRWfGuTv2KSO1Bm3uXZRUX2DquKt3HxiFa2AauHH
iBbt9KCmCoQKkiQrEhLqElkSzb9lIrNxtsAGJpy9C+CP5cIUcptxM/UWIVd47p2W
T0KRTqZuJWD5EjRqQFiHnELNAJ+f2NJqXE4jr8sxI0HaTGVEtUX933DWd5tYuTLv
oKMCnFEl1geNP9s0npC/HPPNGPPZ3edJexTwa5huP5Ek/WMR0fH99SFebZMGRSz8
6myZItJPFCmQ7KXfoZiYIOrRbNWly0QXn47lkAxEiaFFj3ZrktDpkUsA4GFxLtwe
7vSkx6C0BwcK2FNZtoZenkE6feNUu624PAo+AX3pf94T3SpDXNOmvDvuTmeRs8gd
oF4q7riqW+TMwj1Sb83yR2W/9egpqjpwF+fIcL0zk+wM6P/unwARqclpNcdgWwbj
lbxN18mdGt+DV3siJxxamkhWOaCaB2Xe2/G4RK7/2XJYxgkPyZSNzMPQTym0Uve6
tZLgnGxKkePrHH9dfwzuKTjEv6taaQ6wwyEHNxhBVzauNAQVte9QxrW1tJlONoCd
+fi0mqu0WnkdvdPziSX4VDYc/tGMee8A1bbkOgVySHUgLCEkTmEJiuaTIBkDxK/G
l5qQzRYyiLhm17x8QAqt+F4GIzmWTA0BxdkTE4o6958ilJL+RJhnk0u4sOa2mBw5
Uam0OI+obVGHIGNAtjn3sQx7zHzjTtmhYf+YMgJ38JWSAidQW52gcZ3g86aG6nTe
awPqnyN0hDGKsNa94WHdWz2tpLWS1tgbyCyrH7qUDASvQhSS5TaQ7GF2njNeUD9h
DlJIo3adKP4VaLeF2zWWbFWJ61xHAWFlpBi6U7LDP/cBohAY6QHGHFQLYYjDUhkD
b0KTJRX9xdYrHIxgAL3D9CBm56pyhHi27l1xbgrlpb/5Ud5ZtVlvmucZX+U5Cgpe
QlwUh4bP5ZNAgOlexD4B5slZVc+AoVtJn0gmz9dHxIMNWIAxkPpx2UelzNgtZTZW
/gTukrZwEglxF9Nn5a/xdCCpcF0DYCtnX3/DBIYOQ75fUUfJFsK0QqnyMOwwRSCI
tXWQ8JRF7mic37FHSF+Ilia+QZtkw7ECEX5F6zoXEJqxZfL/e4yLsVc8Y1vGT8n2
LexLr8vuVe5RB/3BNOLdHvnowhkV+TRScIxQIJAxDXKrdsXZ8OUGfVYLW2eYeyqe
5UHYWY5g3GdcADEWs7fstW5xESrzwB/ad59xlIZWSA5HyIQcZu5ikk7CQY/wpHJw
vkQGGlDcvAkYiViiNn18oQIhhCCXUfj/h6Z9XYMmFaB5Z3hZ7Tg6ro+IhRMII0WE
fPhZNDH+5T/RKo3Yb/ZImqwQJvLvBmuUQgKJwzo1ldmaTBwXdqzn+1fgq+Qb12oE
d2K2i2YWfiepqHLjg1UHnXA6WrDs9NZtE7hBuB13Nt64VXNh9L+vwm7sD/WbqP8W
gkUc5WXaVZgFXIendqEHSYX9ChTzFfcYrNPMOyOixgnAPY/ahmLAgiFOSjIIngfN
v0BpLjI3gL7LQW+jl4EcBVImx4aVlWVzfxzWIDDZfHmEF5yNlNCLSTzi0zqLVWOp
cvwdT6QQ3mEk7uOOdal0u1E+X1/VvQPRSop+tgQbB48smfbfUGdYP+zNM2r6IuXH
j6m3thesG7b8ite1l6Z5n2bUvZZV0yV5e2KQ7rOxV51AnoTZciNI6fm5iW8zCoMn
lb8ZnbEfNVmGqWZMp0Vk8asSHGqV40oLexTx9lr0/7SpqUuOV9wIHGieZEYDhzmQ
yLuNlaw5QrO3BzNupvEOpqKTW+D3KhNS6durRRpL3JwaBjMPiE+13iSNrwriVFb7
H/ZXHxFM6ntCIbSmJmXE7K8/l4KyIO7BLErTdXdYxWClSxnk+WLGMsLJt7qphA4V
ybINie6g1aBgf307X5KYZFhd7j39mQSHaqJRfTjF3peZcpTPX1IQVEKLu5kH7ye7
O+fD67rv/+wcNQTahnriqnEBoN7AP8R29dfVJef9r97BSsUal1NHpHYtEIldqnI1
m8cxT2vjUYy0ersBV1zQQvrF1MwAWIjmj0q4ThW926itJdYPlNPiC08TCAX+YcRI
fynhkFt+bJo5jmzq67g4r2Bro6F0cbfHShXv6CHsY5O9Lv5MR+ASkRhv44HUwEz2
B+A/WWnz30kxqhBfRLB2whFfwCYUejQ54Pvpd2Xa2eUFijJMc5y+EfowNSYtWwFk
7xPWMwuGhqUXjnlmmKi+Tp/j+h2Fe5whA4/SxnzIE0AhiHq4LATiwlZX/oJL2soc
fJlogQIu27R+K46XQ7H80ONapP5d/kMzkklh7hH3UTocUx+jKIuVRsy83SCtyJpU
/1PKSG0jC4y+i3Xu4FyqGSya+WU/cApofALdIovshyr9zfORWkKEmWAsmbm/HbeS
tLMq34Tge6Hv/oReVH9UW2olfp+DbJnh7TMvlMa/p8o6ueX/ZJjmL8X823v1dE0Q
E0m6z9kkSdhj633LpiiUaeib6ayqVEjnGWBA1OjCKNZDVGLiEDk+4Vtm5QuOKvx9
76pyoTI1pIIlh3LAokYA88fSX8RdTD4nirv+rW390M0ZEx/nx1nsnxCDCn3BATYE
Legx8HwMv37sJnSdJ64jOoIADQmqYlAT4btOPyx8IEvFvl9eSBRvIsfRYxZzou2B
KdSvvGCoBn8vJobjCBG9FjxGfFWxSlCy8JhrMqmKxo7qD/Qp+/+21xyNfK6a+2/0
b6Aq6i7/PxvBhaFmAnSBIR60TKooZ2OY1eJVJoyrkZ/C9c0OL7SgJgT/AC3NS1U+
qVCnY+5+iqprxDv3wlK1IjEM0lVHdOzQiEbYMS7ZAbrSyEMTMxVLIGxW8kin9k8a
qIZyMk6hJUPzMTnGWSru/8KMz3UkoNBN4WQe9TNI+MV2f3uLPiJWCuuHXsoenS78
Q3eGFHZcPKydnQ+C3K+osjYXq2sSGGkpBdM3G5MQtPbEAjqKbSfzhDV4Oph4/4XT
3/3kCHdXbLyxldVRUWQxvaApM4yDdQop5svHzU1j9tnQHJIH87UKDrN+QlXXnTHk
eLaeS3Oe9C+lSJmXHIOo3QZPMZ8fuKOVB6OXC8XLvlIUv89+nPQDbiCfVBgEKM8r
Z7cRx0VIoz3DtqVA+qs0BEEx+9qdo0xnQk1SRYdjpHimWTLJqQoSTn147ugcTV1E
yneQUuPGKTAXAC6yO4rDhXNfk6VwjvqI3AudT6T/JUbgp+gpJDWhbM2lZTJsZfKa
Z8ByWB1wBcAvYrcu7STdZmt1kshMokQUrTc3B+Z3VK1IMd5dBwLzOXb4wR6kZ/kE
nLkdVbbSZAJnEMz3ELC2OV7C4CRlaMIqA31Y+KrZZs0pfYfpVkmKc6SAeq+ePKJy
5WcZnftfZKpjslI65FsUc7eauahmyVqBKg3E6mXdOxDEAuFC5u2hL2fm/9x8YFuz
tTkh95I4gBzVY5qbSQj4+q3mUBG6Jh5wBOohQW6BjALutXwNZjXR5l5b9opZ7LDh
FKtoCNQLEW3yBtCiUHT4T1C0ZcoLlZsTZ4ELm95wGxyGiYfoehA3p7Ag0VpfSsHs
v0+ZsKB2NmyztFQdv+ToDf59g1EKVNWWWf4XtHV0EhuK6N0CS07b9c6SWPLUsJkj
DS2zXBvS6WTAQVezpBrWOkdVRDYgPvJR/x9fx61Q5lcbznOr7zlkJF+tDKydW/FQ
vsr5ycLDMEfU3Jk+h8O+rdV52WWAVz65g2s02F6Q0WfkjZG8zd1AWjp/suTYD8b+
nvEx5eSe2LjVcnSxle7HigwKXJBqIL1YhNSDuAFAlUzDz66ZdRocNYc+arY2z83t
l/V/yRFLrozN1UR9NXtDkDVmSSm0LTSrP/r/mtxEkRGbmQkeczKXajlVHpv+ssa2
tRXtfCEv+Z7LpyGYZgPTCs6UWJhOm6Gn/Y1/4cVsBlwiohj++Dz+4mOspfGi4UAd
2X9DHAZ0LBFwXB0p6enhvkcM2Dl9wbo5QZErb2Z3IQiGZfwjAG4WoBVM26tLcBv2
yUSjQduh/8aoc9wK5EaJRqmf+vTGBe82/aZko3dFPLgtFKx7RW9vNeWptZpnM92T
mZFkvNrvcmoPs5MvArz8/hlqH5WErdAIX/pZVH+gK2MeMlhVSiT848f9YLnB70Mu
hcZ2yUxSdZeF1456IqDouBmbdKs+u9BAU3r9BqIDdFD0ZMKqm6YbQ61Tu5QdFV5y
mwD7Ec80cnwNaV/VFBQAptzglKaTwcvhO0qJHApBYGzVnCaoGsqTCqwyaz42Eocs
x810h+qIZWGEcZZzkPisTjhLEw8G+Pw4qChOSJnRME7V3QXJMf+pEfxVfn9gkpYE
f1Og0SZ+HBC6QYyux9g4SJOzBjEfjakJOZk1erE+uvNML5OVM/NIyA2s2j6tvWBj
SBtoR6mw52qTbrqRSwTpwfYiLqHO0loPz44q47InElTkQrKYLwYAF2pZ8AqcuLoY
Nf6rt5Jxq2umEsDMhV8yFo+GIGCAADClppZoDYKOQcXxFWtMY02jBAG5PFuacP2C
zc2pF8pQ5c5QVodADtPKQ8BLnNye0D09JntiCJfaKe6JyieASPKvnwocFoZx59I+
H/uDqeYLl77vc6qao3lKIV3bUS/HRXeetInuz6pNacHmTP0MGdfmUkjxI7636mhA
1oqR/TmHhwDm6KtiOLeYabdxvcNrapIDjpWH0fNaImUWrSDUEwodGFs+ggXSYcYn
ncFaS4lsqRvGJb5FfMdc5kp3XqtVW5/EF9ZekM268uR+b09dt7ka0pECL7K7zMRd
/NXtMULTxd2VCts+3MKEpgOGGR+InZL+F3kDlL7CPVG9tTsDYrsNdyHEsMr4wFXb
nTlbIo33bYG7XoaxbWnKJb3qQnf9HQcaZd8RFNeCHNSDmJTUUuI6cK9B7s0H+gKh
5u4NHJYpOLzKeO1OvR8ZR/9mc/nzLKSGYGsazaWZvcOzmJDHk8745cbIEJqohSAg
6/QCFyU7dO5Ik7FWSUxAZmEJHfo/gyasDTCqJmSHyhwiarF9P7Lt95pUMlsNdzmk
gAxNi0jXShtYD++NWkKKwATFF7NwNM0RT6uktLuUfJFlBXxGkj7AfRJbgqt8x9Vg
3zzuVXlbLo4/O+eoBkamO1JF691w8KdeVCh0jOr3DWDymPR1PMbhR+V/VFp4H04N
aiitQKLMZMqAvNBJVIgZ3Tj8mzOuMWOj1MDBYNe6OJdEXgaoaX57vuA5CXO6bglJ
JA9zO9qxGXW3Nb63z3jYO11rBxAb2yqyXXiSinKzQCt3yV6+hXoGAkKKdhzOWDoy
MW51QDkG1lSVdVCNZK4e//EoMlZdmlO7XNLI2QIwNAK8MrLkgXrYsqiwibxWWmMS
YdbJyL7zNkNnSQ/0YOXVCXIwkONrWAp0gDb3ePHyaLv9NfOwS74RhdU2ZDHgW9Yn
sY0HUIqC598zwOLntjKddPIGGVnhARg3i85FnQ5gY6laFuL9GomawPdIB65AZey5
WPwlf8sWxEPXY9Ao+0pHyJ0IRReTXNUT6oYBbRCu9OHx6BZbgCjQI+dj4QkDLDW0
3y/e6v7I8KaPu6yk9T55VAtkI1OSbf0Vq+8r8YjW3DRRqObbueGNb6j5Ebec13Ax
HnUjwtP/dcjazUno6RT31HoiavuBwNkTBDlbhDd6Md49ChVjZ/o8EIcVcAIZ6I2B
2TYWPlnAwHq3l0XJ6NKTrR72rgVCtBibTyubTZPVym4AQ728pz+IZ5PT5kgc3mQR
8jJLLh3njTC+YWwxcmHGMaX5Zs9O3+2wI7081lNcZIXJXC7ubrjR7SkyTy7vBunb
vTtF8D0jPtP4pIacyxxunjRgGk/3HJjNu4C5NXhj6mlOj8nuUidpb8OfazZZrC+W
UZb1SJZGI/8vE3Y/VZ10icat4/ulpUkLFaarD+6EdtgSorAMBayvygE0YuMHEOdL
p3oZYcExc2HYUIwailZz6DQKO/yje4WqIILZ59R5rRTWlA1yk0cvyLiLlf+wkQYb
e7N3/0yrdv/cQsKT2P8J5ck/Mfb+3ROGMaTXAe6An+j16hZJzrgT6BVB+nkIAKrb
O/y8GgGtKXVHzh66juS+qqOxlSvsOVrNTgexauBhYC1Re9PdncLL3kjbWeYNxe3p
IiBaloxDeUVKKwqZ/MJNZj9WUjXXw7j2k96+wZg7vuBp83xis++KChPwatC6x2Ks
NiQ+19+HX1xiFbQvtbcVrXL8CeRNXVgPPP2IYmsmsGASH8UuYhbiRAiYVkRSXrww
BPsR2Z/VUzkX76EjFSPOuJ/g7etNhixHiPgCDOMauPG0EbKEns+w/REaY5DbsCfd
qUFIpdkdq9wnzvaITxbPOEAz414qqUeMa8n4+Ey4oI+wfq8Arl1VS9h/VC1P3vM9
aJm/abPNsedUsVgOyWxAC7P4GlRPZ9gYzn0bAYmlGiPOHQ2ZVCYsm1mB7ltbxuOs
GfR8aMfDBEk31es4WUyoXDh3rLAvnNEwRHcXTBKk8vs1ye+SAKUR3YdotS9S0VP8
DYhdwY5zNTPsdilK/JxpakEZVbtKDB/nRGQ5GMHRR6jpj3+kqf1kAiuflVza6RNk
BGQZJAdcFihc8FnO8rsh4nQVHkich5/fdxEdkBKLGrRvNLTAHRfTVnKDtwseqAND
ANMURxUeiUvmL/j8g9FOHwTNqlWt7Dm+iAWQpjzJ7gQSvmB3Miowm7gKk4o0cd16
czEOSX+05+hxbH59WgiE5bmBgrSIlwdxCcT4kHG03pnvEGEpyoCKyL0Qj2QdwWCt
1PZC3K2yLORoshf6MAyRKjkFN8LQdHOA7XxTJqw+EpiuJkPCo4DEIPVsM9+kx+tA
avnfzxbLLOr9BE65RZtBnmSdqzAxuwtlXEopBAWMktL0nPb8EaYclQb+xSWCb/ue
EaWTCdDFR61f1ozi3jWHhfauQJ5E8pHCzuXpi7/H0D54gJMCAqHCHXEMXTE/Z6K5
TIYdG1RmNVc5255d1nLFHbR8iibemvFlhmNXJCJqiTxbWeq/9m0lq2ULimkDadJV
WF93D8F+ehkrzQhe7EWRYSD5IUFFSZV/RbyPymgWMkG3DWT/qWi6gJnVLVabzW02
5vTFi2Rm4u/EbNXbwjOFOkYkO5UwSr6qR/0H0z2VtV0fHTb0HENT01AuOaqOIS0p
vHQg/+tASCim3MftRaMBV5SH0Nu9zgnxg10JIE95KwICGU/SeP71RmsaHAcIqYfo
l4KxiUHi5zApknav+wANo3PaQfmkA6tC2BM3+LYnqMsrrqartg7HP8Y7tB3rTRAs
YOfZsI2lgBFt0Yl7sMwR8T2nTrFtrWf1sd3YSh6kOSq5bJxdwxOHSqWK3MjXUS60
qpc7+lYBkpXxkrfP6OP8QG+d2IazQWjkgVf8Cxv7oyWPncg3VkfMe8AEN8TUD8rw
P3uVJINDnofVk71UKaXzDo03hQPv6ZS+hx5NQkdgg5UbbP2QIbMm+X/ca1uXfH0h
5U4uHlg2smvzv6HAeVUKRtEPAKkF9mP3EZM4IMCyVwmJsGNW5sMVf/yUAjWrzho2
mDjRFnOcAtV7jSQbTTe9/vY1xWZ91SOivz37iTZpSWhrYxDgBJW8lkjSRs3YSUxC
DlDGLUm68i8KU6UUZn4nFtniE5GRN6xEbpZ44r5wjFR15vxMV83hgDH/W442wpbq
4QZE9tLaM7Jaltj+WC5kIb6LrtLnCJ6hrrhV2ge6nEJ5/ya1Z2wlEZKRjy4lj67I
ZjsC6pECZEDGUuxSppw2jPkaviSRzJfZY0/JrcYu6cAcvOSKjcJx+RWENofMiBXV
NsI7wXs1E0Us064kRzoDLqaBExTqFERFDREip7bIH7cKbl4x+s5my23md70uWwg7
OalKrW1BFeJM25kAcAb467QwVGLoFBASais09Y7DPqrZnfJCmWGMIXo/xGxSoB5H
j8v4N/ZW4X0mOCgtQRH47wjMq5PzO7/QYr0Afj0mYwnqBQCyNxkWc22fc0IALZaY
HLyKzycAg80u0M7EUiNM3DBzgF76rVoam9mwLMCQGMwLKoR463ga7vuu/jjA5Nr/
FCfdhmjjUzA3+LBEfxtUddVPCXRRvwk+tde0wMRap9gqeqEZwZIkka7XA8RhAJ0G
PE8zuTOjgi7umQfHWY8bBggE+rr6n0JlrIWBDSzT0GkpChm6PP8iDToBr4nel4Oi
kXQPMpxziZ6mzjIYYsNSw7UMxb6PX8b90zd6u+p+y1bwQ+GKX9i79ynJsYJfTRba
EH91GLH70oM4QvIJYLfWFaD/0kr/2LwgVVn+DyDZMXPCF218t8XbYs6eGX+VHknl
onimqRug+kYEsPNOW7ujy2C+R2D8C55PdVuVW24fLJcIM8m3T+vO2F6EzDIJ3LKf
/8XKFgsFmtYpWl9OU11deIP4P3GCSFuUX1QRxrjWcQfd4RKHUpknfDTD1t8yjuX+
8s2NNYo3+JPXpr78VXr3QeF6/wU9tiL05BoRmCg1A1gdl2DVmLfU7eQd6JCOkNVD
Dr3xgIqIjHfzHezF9q9JqPyNvk5klGzJI6o7zPBABgvgzR2s+OdyTx066LEJ48CE
1wRqj20x2ldhsD7aQ06TfFM+6FQwTFeOAJjUFXAy1S8AZeOtvuoERQ9xhCPtC4/W
zHmpS4Eb3dIe07+B0lN9FQvHM1D7tYDUVyKLM58o0b5kZltAg2AQo8tJgBWnBtGs
SU0fH9ycACeTkIpEZjh1Ud3PJiqhevImPdLZ+QFDjOvfQF6DAWXxHZnJi1yGKz8d
hM95CC7riaQrDNFZ/VxXM6BflP5Xseu2dE26vYnU9wG/h7YIGGYtTzwE9wSPF/KP
SpO9PKvzprY6z6aswXNjQLZDqGFfCyzilr5D+hGgNYNRVniz1li5zTIFc9DOpwoU
+ws2Ox1OXfi10ZuHOgwpwnNEIKsY/go/Yuh5CY+IEydYty7o1OSHGvSZBTw/+1Xj
XMNNwI4nI32CQAJXZU2jJGt4arISzm//UdtbUmVwh9Ej9WGjlxQi7t3AfNuFgBw0
TRkLA0v9F0EmYfZOfnik11yxRWpNtr1BXwCullAeB+yDTCMrYdybR5XXXxPPFyvO
bHrbrR5Fh3to7N3uHW6I1LjtkJcNa6lic6f+RXmjGmIUJWJdddrYKzHmizXfuvbu
Rupi1cZK7zQIzYMVy96RuA1tVeqO21RyL9B9M6RYT/0BgO2eu5PfFuNB/FqfNzyH
FBnU5ZHVTmITB+CGPr02w5kkhYUzvIvcLh6pPjcBHfZiYpWuZVkBjcoMu339wrh6
27K5CA6jynSW7CyCDZMlsqa3mAZ+D9xS5Qr/AflhvwPd7vIqdLQYK4i/cTFbCQiu
yh8lYVBrfS15J25H9WWv2DaiokGh3dETFl1szZVTBalL7zNHXgU3k6lWY+u3H8Rz
1TCmjy0biYglG0/6yDTXlSe2enIHzSHrSQ1vnbki2weYWVGnTZPc9diTm+eHErqt
CZNVcJsakLtdgTUMwmQOpzRI/3L/ms1EOuap19mYBcaTycRgW7NjaXtCs8EbZGfU
+RftfyRQAflUimjYkayq9lbwun7e8TI/pUlbK3jPV6aPmIVrwGMLhBBIJ9YQ1XE7
5zpjrYzuQCqa3Uh9QwuxzumzQuk1h6tDFB0uqNPI437jDTMqqPW3q/dPXKLonIIX
VHqzykpf0FyIGCi/2+vMMKL+Lql2akT+Ik86bZuP1wCalyhq8nmI2eUXVEgTZR27
unKBxZE3x7MR+lyozvSNVMMKf3W73JSSXu1UA15D6HuvLx1K/7N5XG9xNXsdqQ70
8drlRyTsMjJeag1obdpxj5VtQyQc23GCcYTWxrUHc7I1BU5y+q5Sgh1HnzsuEBhH
4Yjg7p68XAok2Lq4a5+9sTVQfKRw2C1jHH7Z6qQG0tFawDLVRWHWX3d8TMQt0n9P
v3HOpMa9rAEak8ZAB4Fk8cWCxk/+VXnD5pJVaRMKefuVsClQF/O0Y72nuQeOEcv3
vN8X6kHb7LV3JPUv/4nva25rLHwmHQClRswFEAQ0h5yjE8mJz66tWOs0iLSOuwKc
Kzceqp65Y1P5GOjhE+nRfFdY4Y0yOqT7sv45EDK3a2SzQmOFnR3RNbJWyW/suz0J
DsFDlsEF4rLnyRNz8kMmOCnuKG57EkG+NwbXmyJeOmIhxzItO5dYnnM4jlK7mCQC
NQqspPPtFAq0b2JcitEAXqTdXoZ2WZrgqLyQYkj2weJMTRKvq8fqPrdX1JvQ+qJI
c+mwJVqx3uJEC+YQcYFIDiwJVzHPIYaRB3qwOolKT1wUVA6DfVZfpEVJJLEFGG6H
2YThCziZYLZhjAX0pgJs+QDKWiWWy436urrLQOuf/dclT52pHTi031pjcl28SigB
t/iriUtASyZxSFb6VpmtiCosZxMRJFW+Cb1GcsI2aaFaPgwkF48IjZ+GSr+MDtuJ
bP1TFYMAgLb35j8V+Z1mlavqHA6icsx9+w/iOZ1qLWohfSWQEdmpZsJhkO6V/ccC
PzMkwpyRkxeUrlPhhQvV2QA5AHMjE8alTH401+ZJFgIhcGgiNg8lBFYpjfk55iij
EtGIDuaJDjEKnL+CTwMyRsgvfnT7NA2qwBrrQJYictGVJ/u1X4BIZGMgJJfOnxWY
36HjsoavkPngm4kkETFJWZD0dwSJo/sRGk0StfBWfPpYIy4NEPRq9hKgIrQUE5cw
jPARSaZIdtW8+Ym9be4PQFcHm+x+VTiDOwla1glOqPOcL+saf1vhxLXye4ZSd3AH
oTGP+3BC3faIWrxtKKXVch6l/6HG/g30WFHx0BD6ecrPDrU9seI7smQ2jUSCpgTt
/Y/enXpNFAQnYKFOYA9IGyln7QjO85+l3yfZ2+agESX/jceqo0KzykRa0F5aqfen
+6AFoBmxAvPoo8Gi8CpBsxjfz7pEiQu3b66YK8FHDjMmCEXV+Y78Rz/39+F7nAmX
omn2GZQRi1qx1MxMvU1bbMmKv5jeNAblmL2DOE3v4xGLxhHDQoQby0zjccT9FfjH
kKRkYgy4zonafop5osX5ZuUxvStd9Oj+GU9g8/zrk2GGC61NlKHIBkj0kP8zEJdh
L3QsYfi3dIsZpxvA30BgCqUOJDfC12xaVE58Yz2K0GHHwTT5fauDwExeHW1RE4D3
ho4tKCuYMR8lQEKYCYtrFcNp7E0524bl1/Th4yfYPcCcaxCtKD6NU+EP5A59RtC4
KOcR3qHrF2Rnjj2XuAvUsv51sTjHpz+huoXQXZAKvcFCUio2Y4x8WAS6Q+SKLZkz
9xq50wRzTiB/b/wEshRTKwA4MpeAievMS2O5wwy+6KcQA2BsOw6DPCjLK1U0kZ9l
yIj+9OVUftpwG/oVkbsUnoQHbPl2p7tWdGDNFzpozvN26EmT0Hrcu2UZqG3aOsg/
cjdCjBtGWuJiPKBQGcQ9/iPidjiRALH4tysoixTzDmXMA8j+c7KwKg8R5YVH2FCG
nOsP/32DvTJXAWzYWfTqYgHggupApoZAlFEzEu2ExZyzxzdZsTmVe64mnpsuWkEV
Bbq5lV0Ycm09OKfuqvnHbiFROo/gD/tQinxdvCZoYEatMSM/ZviLQLOZa+VXeqHT
tNIgeVaz+k6ERiWq8tEitw8kUNtnXe9cIqEYnsuJCQKQZzND0/QR6QS3R8ES7l7N
zuA/whzDgaPjvC8eVyIVsJmYZUXEt+XAtdYA19WvNDp5BQ+HJ6h8NP21UM7UAnQk
WgsSGiKMJfylYQ7u217f560CfEobc+I/btBc+OL3H5z23r0bcy1bgMObLNmXOU+c
nDDyIgDSA55+gUGscFVqswrEgKBntbqHRWYf1n+awbBceztOYRQP9daJ+KhyrhNL
snL3pughsB6jnRZ8Ezmndzva/Xk4pz355wsHKpYleGMjuG6X7f3GE1Nl16gxofAu
ARNL+ixxY8t+AHXEvU1rCIurD4H5g9m/EXcS3K9FOTrBbIKMsPRyKov4A2yBzsuU
dwEsxaVMKxlkc+ZcFBwk+qzcSZO76UM0pQJzsl5h3eCBrz/Fe/P46cPQ4nzP6ur/
t7PriJYBVpMdBaK0wu+/sg2p8jIhpDoiPoz6LtE7A1OLYlnaAESIu1/dBaWDY6Kz
9AxSztOATHhTksJLe3za0l0x7+b8tcBiu/2JA4D4yt3UDKtPWnOn9cuv0p92mPWr
FizDrpt0+MpGtRLbWXXERf9ujxXRK9JAd1/DLd/sEdaVQ7z5VuZrcv9Orcz106e5
l0v1y9B+XM8ErGYiDAToqe+a3lg67Gr+VRUPxtySAzsDwCmf/3HptR2+XCnyNNEj
hFv5ZamPKTdafqFLpPDLSgDMoK1HYlzmFpZGP4PtSyTHQSdc+EY28XrCWygi4NFc
kENkn/x71lIBfJxunkqXtpquqFLGu/u3S4u42wRpcWtYHeoAr27NKCwkV/YXdSLn
NrAx0IpixnxU3wNRA5Km8yKj1Ly7SsXUlqz6rbPm7zBUyylHK2lm8YfkV6ZQBHIl
6e7r1mjtV3sZ0b/037Ti1xJAtwWD1nu6V0yPdqzHUxVmhULoFUdjQiP/4xk43jHW
9G2MmOwsTVabOT0do0k5IlQD1XZux4HM5G/9lOCGi5LwIedW0zKrMVRVNm1VMvC/
JyKsiaS2pWceLB3rCubH2eKwkE3JFY/rWqO9X3x4ErN2PflPF6sj71JMGux4h5Og
6JV9To/H70W6ktEsFEsOwtfKUDeL+/ihhUS3fAtbk68D2ZVGDwbbCDFJveKwyhSE
KlvqV6vQCvthFUh63kOEGPm6ponCSb0p5+BVhHhsXS5YQbANo+4HC4Lf9ZIvbR1P
PO0ERoAnl19FeBKZ08kh9U/8VNCgiUVgFmaLMFupGn/8AgT5KBLJJ8I4DajI03lH
IG0bz3q7aG7Y4NHbnGUHB5UFadpEGbnwQKchiznUA90pSsez63TGmkls0gwZt+gh
6RRpNpeMaePmhk2c4vF2FerRXd8VGO3918yRf3HFRB4igHLuUCBO7PzN/f+hVAea
aSkKcggB2htAyF8tYduxvVKLU/zwEh8FMZOpAcKWponoiN924hiBDk7QY/103BM+
P1gqdLhR/a1HegLQLRHARyMwDhMX7kn69CHGKcTYtRSc9MMFO0fwiwlseVCURMWt
YKHQ9/xc3M73U+/3TtvfwF7UIdz93rVMOgLmyq2il4TyNGDICIbZYIuqB+rVaKmf
qhKwySTRVd+Gxw1TFKA475UT8qxmyrhSqS7V1b9zTqkVECsoXPUEYZ3PjPtycrIt
Qhsq794Z5pXJNJPfxNUNqeXJn18bl4IDsjL5oxJvjvr2pMbmJ2T1IHVL79HcF57b
daRj+3mWiZTg0BEXsNbTPYbzitDc66fKEdTyMJ5w/GqW6darn4FxUgh7Nm+X3L8L
DT0ZRUEJw1BCkePAf4jsP7xJX+3viL5aemecQfH7AKMG5ZitMZXWp7i/AWYLApXn
u5dCvdVrKBLPtcJqPcDhfu1KVeuav6RiAt7zCG4x/VYdnrEDurs5texbbCjK+ZSr
MMKw0DcKdRMA4CmT5IjIIyfSopDbHA5Tw0WbCUrrCUGPuKQNE1QVqqCHmDABbQ9t
MSPBQGjMbN0uH65fvUtOr2GOB0GlmecYrFxq+Pj7OmBX6gbzwaP0haK2IgPXT/Mg
GBPdxRD1PvwB82G/19B2MiiIxfimhUF7ahsGW5QLzRjij0snsuG3PWyjje1id2s0
s/AN1h791qwzgFfVQRxe7Kerpx1ooofZx2TnNqdacIVKo1fdhaSPUGoMZAcpEQN2
LChtfEKZI+npjB2/Ad1LlXiZpmsRRlvQ5iO1fk4oMaXFHR3y+2g8CPAYp62wmK0I
RxgtoQx8mgceEhO8gImydu61KIVonDMlZLBWJ7RIeujjiIqo8IqqHTQaW2stB7/W
Y188E/ZXocs4HJxUo4U1jG13r3CQ5sU/actpJppcd0nHkw1l5u9iPz+njygolZYu
rEqu382BN5HfYj8FONnz+YIRHSAYf4E27NFTuvu2l6IZkZNItGaevsHlOJ1yycs+
a4PsM7EhdHJr6Nox5OSpAGuwbyz4fNPcvP55dx2DvuTxTdLUeJUqXo9xWjIpx5Bi
ALJvnt9hwIL/xgNrZm1pJxubTEWoi1ofLkn8GzB5oCWw610V/6gPY1x7gzJH6/1D
iuGfdEWrf8JRADoKKZvMz2q5n2AHo2qESF4Df+zPeJYW37Rn2hbvDmXOj1XN6BeA
1OA2I5GALIcwvNv6dUejNdmshMxOjK/2nkGxAo8mEQ8yJ1e+HVOEsjn8UlY8W/FV
wvwOXyI/57kKB2rKX5+KetDE2WR6wetPLo9lSySv/IcOCwMSiZnief8/GDuRxt/U
mtMWuu+meTuOM3ip7GQhf4e4D/QHxVd3i1uHFry7Vdx0p+fx+5S9NPOSvdsoLy7Q
gQL6OdChJdndb16z94V0pGScW6pIgUm6I+yXTGwiTXHS7oF4u3tC0N7KRDMoDJX4
tk8czuz52WWF6GwGJJfs12qVwAwAs8xYdJH4y8YJN/iiHFKneW1qJbmOhwv5ADWJ
5B7hCAC+DWaorRjBc192UiltwGKfsB+rylfXIWzG8W0asIf2cIqSCZr3NZY1FYPy
8lnldA8bzC/kPu2h2PnZqYDdu3qu33obRPUbR/OMXDgXI3XZEgT/DNqHk93GLXiE
3vPjiIqM61ZE8x4OYVJuj8TPUI+MIvunhuDEFnTVSLqIF5DHSCkaHxsQL8WBq9H8
CE/PPwVjAhvNQ6MjOcxl6biti2WDsVW1jIcikAZZpz5Xu8P02Ek16CmPiBdU7FU9
DDUR8MLUnPrrYR+co8scPxgIFQwx/Ww2h8wcKQP2PGu358R7qe8rwcpX7kfnrrKn
MC1OTX2cGnJ8UwYv4Y3zd7e4e9oit5Hjz7MsIxOPSBddukG7swtPvjj0XJXc+hMj
vb6TDipRUudaVulQ5Y/UVKUnaGwPaXQtHZ0xduI/jbBRAVHXe9Ut1NpKbI6ZLm3d
9GyWKBvAt0EKDtj3xQHFQj1fl8jLRznzDlSbvtwXGO+M6DLqFFdtcuYyxtnkDQkO
B15InHySo45V3XQie1tL+f1UsMMh0jjrj5h2rjGcIWOEERsuRaITGDER3R+0v93w
xTACeT5nrAy/ATS5+UP8NqTVlKjLZNgap2rrmrxP1pQyVIXZ1V0isr3Ipir+jh1W
uFiAZZZpHomMCHOjxM9hPZv8orSv7SQpR+hWt6lkbsabaRSo+/C+QQ6gTiAjaihk
VyN2kYs4HbS3htNMcXrHBhnUYUtsz0IpR2QgWfDltIp01ICxca1D039CmJuWXw8S
S7ItWaasafjLftE8f2BU8kyPG/y1yaTkQmMFPwBQe4GUdceWVwwbJzBBCML2BgKB
Ok+NNmjslllSBhGl033ZFnc77TQVaYl2Fxw1nLViGd34Aj/ICQVNyD4F4wa0bVPr
ayCAUFMmpyUyKy7jj4FhwxjpS8R8NVrIKHJzDza6NFMpMvdWzU5DQtNPWUjSfpc6
hLg4hbjZYe2AU2ugnDXCXOo0UOw3DAe/hUT3cmbgZOqhZeLk43NUYHdvw8qtV/Uw
NqUxfMyEJxZ3eI12pK3AttVxPukS7f7g9JSuSOpjJWrzkv4Bs6MrLwJStiHmnval
VF/sjYWkH9p8BkaU5Mzq8qUofFLBLgQtMSIwHf0QEMrNhbFrBwX6pAoP+rgec8yU
+7nikOK6GPh71W5tOSwjhFtF1w6IbjqU/Muh+PH//cfwCRRbfktxRugdQ2SSMCxd
P57BXwFi7LBD2SjZRBu82qz2SDWpFa55/p0w0+AyprQ9xOQES1XnvDtoG4EReG9A
oPy9NTpQ/4kj0wxOXvC2mkXbA5sicnnKgtonNDmLg6skBEU2txPgF3IfwCGqJ8fc
LmnI7RPvXrm4t1vTZmkpggIn8y2Rp2iMBugRB3apv6FWw7XmYKMwgemwHeO+jKhk
aOXJFNhfjfcE6fPD9S/MhQS5TShKkHg1ysjLSsQnQy79NqNz+c1mYh9Edgy3MwSh
6tZ1sJZMUiLnzPI4zYKVtq5UO4FESUeesELsQirpIQ0SivA268Nz1GlGxipvCA8Q
LCU7hE8CJV9+aSjTUVsxxv/vIqnnkjhIryhHZkwthywlU6GFNUjzwVMdLkAhG0nm
TGHwWNa4vpy6IWb9680glFcKtg6F+QcJPjuCJL7YJFhi8RRGYSYyi7ytsnSs+iji
CiYBEvDQiXGutTDLHfEnPtIX2MO6SrsuEnUjWJeI4g5TYFHfk4Trf+R+SyK1QkAj
vNfRGU4ShGSAmkbXls/f80lqDFx9YVrmGy6HnEEBecUovBk41XxJCEliravnejsy
tZ+zsEVyI0YoRpcmXu/UvarTrog6G1G2SELM+/qt1OCnIi0C8kjgSWnoLyn9o6pS
Ob393mOJqzcCFH2u1fgAV3xDnPQlXZHt1/t02X7qCTWTv0tytWQs6SLzp1XEPd2R
G+TrutKMBqYGSb8YcXVkFSbdgAeCvVHkkpq5I3nY6d3qr04yvxuP+4HSZZM/0pH7
XTkLDI3HFbzctPfrd0+glqJCl6UOXyVzPDna9cA70qo9gdPgPumYcc5wC0xTpVLs
U6SE7g6hf6nsxMijEK6K2Ru2E8cOXR3o5lPzg7JTCrUSY8hsspEx97+gnifqjlTH
ZoaqibHQjtEqix5KUHybb98YdlOZSSuz1SxYpTPF01YjxsHVw2O3hPx6PzR9iJbf
S1QeDzbVz7cDg9aXcbNPUh3+W2id6LpmlAiVOCqCtOI7oI/Dq4Vumv22xMtYwxPy
7H37poiigeYlFYUu5uwN3cCRrqD/acz1RnQnEnGAAZR5Ls+czgNz6xwx/eL4dWKL
SpsN8refXDVnCskoFkYhM+YECVwTytrrhajZfVIx46uXWk4P+qjH/Dr0Cac7TUiq
abEDMtDOkrX2w+3mnW/uMlcbLqSEVb8R8MMM2VUsakD9/1ZK0j6iFnUr/jPUht4e
BggSRJ7uKF0N27PCjYgRhcdirwWijpBS8CMWHXqBWOGczriEn4wfGU2zrhS2w371
F+IqkGjOSuUXdHlY7LvUd3ajsWtNPN8CVYP1eMZORWlheIUY/5cYTqY6tqGu67su
aTHR9CMZ63UilwqIRx/0KG1pxi0XPNyrwoQkiU6LLl1Dh+tYkvt9psnS+7tic6Z2
gdafWTbMA79hKYYM8gobNJ0+XA/tiz/R20cUy0BDDttrqAE6FsF3qiAgzVj9R6Nq
90RHW4mVIAzrRe0yTIrqzAeYprGhIk7JZw2VM/zFT0pFtbunmySStVGv5pY3eW2e
JQvWKWY6O3QVavPC8ZeTbTFM52n4+LOTRTpYDuZfvZNleL9qW6dig2pMxwfdrogA
XzdKBEoEH4+3PgUT0cq1owo5ajhZZ/z7LYIfEXGAI86Bm2/j0SPnIG92NkV2dLBu
yrbJQDXdLDwONzIB6POoixmwdJREk5FrzeZEljmy5zAcToExw36ZSAmzzXW7Heqo
yDPFpxr009RlgfDWdD22OPyEuidy54UKdHX8CGCv5YW6ay1n4+RGTV5Ah6Zme1jR
k1gFSITLPOQhLU5AgR6767ZqKISuKMfKALj5caKG6aTAwNlIhyoeDDrEOfdWB6xf
LbZzpDWitqlXncvj4doAuvajmKhYbB4Pcyl76GqO/lb9SR7AYMUYqM2o/xdLUraj
SQlRTbZk8H9kE+O1IOOdbudyHFPJUJcrdeHUKhOiQC99stnWnHCluQFrrFbJiteC
fLpa6wVBfOxp11+RbpjDnFMJtkUP3L8Jcr4PZ2F6TrdhC4/+VPOhUMoBONI9AWht
ED7J/BBKkPhIQ5rcvdryUrzG8YzY5S3CaQ2xz+q0PvjbEDgMVLvhcPOsBPTTfa/5
nwTADglUKqdnnFrj5uZ9h9J7tzrFDivP/ZQmk9KRuA8pPeyIfkYOgz6F7aHhCsxx
wu49Udt/flFoIq48YRygGs/PN0kde8qGkNCSPX8nTtsAF5EOBDzD7QrmS4YzPE9p
7zYroreqiyM+LyCiAA1gaZuVyfRkbdBp0d9CukDpVb1F8DSYH+zoOfUmXXEoTc+A
bJS9+RMCVQaKq15+9Kukhzab83Y0fkyZXRXjLGKsb7RS9FavHvgNZcZ46bJ3q0UG
BHeG/uv0mwrgYzNKCN0mLi28Qan306u7wNTsGGmuOF+m7dxm5Glm2CxafPrpTjba
hhqV+rOkgbUqj6S4a6cfFzUmWw7UmXNtQqX3xNWKFG1dsyFOS1WnN/tqVAa5b85u
1FzPQMnHgd12pRlM+NmXqPNj192owIOP9ZHOWSfm5E3+RP5z+DxMj9UApiyDuGhb
Wxqn7eM7/x3hP5seqSZc9sJza7B17UuMXeZPHEx4n8YLnYc+yg0QNF0mdAjcHGek
rkM28yI1HqSIV0x8TmVoMiJA8x7lDuqNGbRdOwha9Up2P5+eObvCloSY+3NnNCDc
yYt0/sjyIGlbkR3M1jdFZeONeOaj2T1xeS/ordWxobjEGU8g5Mvr60LrN+UH4Yo9
ozaJOVqDHUnqXKZBsQJgQklEmjX5qb5Zk/WY6CwNMOGQD6lgjmdFHa/wk7Prwnzi
7XyMddiL5iLZCfc/6He30SRW868q4nY/jAmKffRKvwM1UH51t3Gnanhua6ZyFMVw
ZRCWg+iMvxli4IgFKU3pS9JH9YjPtii9kDMrRK8c7Hr3fQXQdmC6hKkjS0GfCPqp
JTtBX3DfMGchBjJbdEf5qXy1GPQkbxYmqPCRSV2kpQOjHSYa0Mw/U4SG1nQNToJm
ljg8HNbejQqSk2BoVUH3vEQxEr/StUphiDzLLQB/xgXhq39DhEsWVqS7wGEVDAV4
EGYiW0FZOfLkux5FUlJStb3wKST3wmNSMEtB8La+09qfvnFd6EzfQBJzShvkT1wN
hJQyIrgXrlUjtxlgYPwWTxr2q8aS09dQYY+7lQvBeAcejSNUXuJpHsQHM/uiSam8
ydM7uFbEoF3OLzoTUvT6msotkTTL26sSy9+LS+UkaYyIcDZeypFZHwVZnwe23Z8q
xOJ8TiC6ThlVSOgycNu2hjQfgxfe1Ok7igYaIUbVrHt+J80JQkLfoHtGxBg9rESJ
GYMonLAmMUdt2xlaA4fM1jLe7MjA1HzUe88K0OY0cLe07bG3kKpQYINQZtzz41cM
i2OwKJnbhuX4c7AWOW8P5RXLsydkak/RVA1ctJiUJmUcIl2Y6lBidoHl2QjTe1t8
rCsJGs7cvzbtJmgPvukmq9dvTaJy9lHcv2EZpMvkisdMy5pudcfvRrjy8bhs1CFa
0I/8fwbA2NzMB8nEQMnq/wFc+Jpum25GbwYAfMIQ0z+lceKPEM7ZWVzjv52C9NmE
hVwABaV+WGQXyx2KLlPKGcB/P2tGXlWFpaGWPP9J3g5cLNJd/pygaa5zFPY70VCe
xCpREDfZTOI7z957leaYfyejHMjOk+X9S2Ge9Iqza+PRttTmF+Vy3y3syF6ZNLso
LqAmYvpO8KjpF113ZAZh2TlJ6AV0VVGFWw1KihWTm14GaLM395AABWQWfAM186ho
rv5LUGKf9/50+xSMugXRbo/H7EwrGxRCUTjxL2tbAEUb2u38y7kjPOkprVHIXFwJ
p/pJ0uN38p0FOmjmacrkhUqPiZAoLZZQio20jcmg4x2DJZmubnHZZRdOBnCr2f0T
3HaXglAnsbwGIZPMY+ApPLscp2Ov8fwqJVMDYnh+ftWKlw9dFfdyr9MNJ6hdtyD7
sZvBBhJBO3xw5I5Rmu4oufC5CanFIw1ACU1c1WcIQOvAK+/T1BxdxCc7twGLT4uN
tk4PjDNSU8zsYKp17M85tdLx91V3VN9JYEGrUEfBcovLPPzujW42CkLmQ2G4jLNc
OIUk0qipPonLlT46rpqgcPum2gvUZnrLqnTvD+lIZKH8zfk9NZACqlBLOGfahWrT
iN8Yk5gYhl0vzTeCxBlRG9f9LyCsqZLhgZ+4MkW3BwMbd/jfTY8xriik7MKcz4a4
EvXOFOj0fVhOdpb9IB69WTyxiFGkF3GOkyWQo0r+IazVyS7qcuXK7HHyxjufEQzk
gH2HUSNnufMLGxaJkaH2fDyBmlC5tnI/Jot6XD/RoUnpwPWZjwLEpJ9cwylduFyw
pZfWyFw5N+U9epC57TLQirXjbhRSXWL3Do16dZI2hDQgM3b2iHn6so7mxStUDZfz
yMkiaxlBAfsqO9iPqfx+zjDc1uEKfRTFd51iroW16bq7kpuhMHzy/4WGsG6JlJK5
lkg07byu6DsvPtZNqB5R/9NLl+6N+pr+/y0heU2Z5DPmap0OBegeWH0st6q4tdaQ
haqz53cR36LX6Mholw1/979vdDYoAeYOjAyaBgwwKIkGqO9A7wGmxSJhd+2Al1uI
13xHy3rogwXrtdsmOs82FZIvoVd7i4zUSrvrHUD/4BJj0R5nHwCkb17UqFpT9K0e
jM84dRrFPBC1lQVmH8Ai1PAaAq8bUCfBnG2oQ6HDmkWwZRvSMVgO4Lp9xIVSsmKh
XjZMhMkEYEWIGUwte0fioJGv8/QJCVqnw1cY6iJtArmF8iLMB/J08Fror+MV3dxS
thHRldpDrj6fg74D4NlBW8oxUvvEZ5mTYBR8bwoY0Nc+LtJzZHps1nlkp19Mgwzg
OUGyyKlD0+3HRK7ypiNq2lQ3lmu+QIXxi615AUjN9GAeWHcNJtyuxtWmtqlpIGmz
CILnVpOGNTgUszMKQe4pUQeaWWEEtxOATjQau0LVFcFDOBU2fbdtcy4uy4UJzGYa
zBvIKUDL9iCqmMsPsKmLR9/YHz+W/iVDXrm6uKbL8ZLP2GDIhCz0soB7Ab8qK+9S
P2RIW9ZnD5m2lTugP9musDFxeSxplEuRvni91kqzZwbwoOEhsivrV+DrKak83nld
Dd+yAu4ftUNX0IxZripwGmsrAYy/sPzb9fEIaDYlPO7Azr13T7XvAGWxeXA8S4ri
392O6Y77FORzjjNo2zv1QczcuPXSIl4bAywIRgf5wq4Rh11DTsebrf+PFSN6VgKu
9kS0uRDI/aQDPxcvhpafAfktsf0c8h3pub/CLoCPLaHfIQnAxE0brnh/BptZXb/U
+jDCg/nQ2G/JfDMJ7RXsNqleEejVreYT4Tl/QsSuRPEk6L7+zUa9Tm2RtKKtlhK9
nXvwQN1fX6jCzufFX3F3aowsw6jhmso6MI0v2BodisCmOFyxdqB94hlHebxQo3sZ
FNwgsBnSN2ABhC/e7SBOKWubq7EKEyNCIAUKI5VmMGHyZqLP2d65K2jH7xikc3IG
Ed7uwsG5khKV1Jt6zq8XWN2WWuThfOYu9sY2PwjK8O4c32xL8iRCyFKcvYoCktv0
K8nimHrtBHLaYnyNufleQJaQEN0vhinqU27B1nxk6IB8BLTE/Oiq42Rvfi/AR9mO
daMIcHg6O+4nS1MB6wjuItpK5a+ylEzez0zegKG+CDyxouTBdWFv/Xe1utAGiq/n
ZVYKPGAfPh5ZbzimBDTkE7rdvgy/Cc8gMSUCTcxLlheViXq3A3jZJzT2n7G3oYtg
I9xh0m2BL0YnEFitjtW9OPETpBFKv/Ezr3nPpZcl702uaD2B+zp9+uZJsrhB+5kG
oOYSl8pqJoLXyuOeZodnae0Yr/nQ97AypWAtqSD72AAVfS3/go/awAMtk+p5Vujs
HEpDBjhupodtbc3k5hDnC/vDVghJEq4IG5z0qtxTp6uqHkgcpjQoco3XdniX535i
Alucv7up2mLq17Lo5AnPWNA/9xvjBfymNrdnl1/HWixXJlcuFNs4cjquWB26lMz4
7pKvQXMvdQALH4Mn28H1yI3VdOfXpSl2Jl5RUpmPXm85/jX2ewJ+BdsD8IlzXAQL
55BgNRHlMm7Y0y6aET3Rz/lsrR8bB2xxdoTIWO0BuHkoI+zxQi+CguRMqvpGJRMj
qOEDf+jSMEzvfZAeXeeYoWQHFxNUKK7Ib2RIOjwFUsLA2OZZgcVDY9iDvYOL4sib
Qtcyl0/NshiID2F1SVHJt/bOx/6Mn+rOfr75Jsq32SjEcU28Bt+xPwYsUWM1XOkf
SOblLo2qEk73pBDDL4W8Rqcmx+QHFRaJOnfsuSWImwfEGrVaUNd75UTchji0OGDK
oSY391xNSQibmUoEOTMyiKw/b5CybiEaCEZHR2l1PxC3jGjZPWmvQdvNSccuW4UP
5KfynaQJHfFsXvh5xD1uxG9s8Zy0U9+cG36YzAVOGnNqA7VGvdglUG0VfDYLzAl6
nlwkqghG2dSuYgvRtO1cUKUtONLGIy5y2F65WKquqJ21ZuN8vJbnohne+gg+aLoO
+SIIQB7MZr/ie0G2pd+mRHc8w/RpS5QKjw0cKrUEhjhljfe+gCeN8CBhtZYSMknp
Exlx2DMJHvcwx3G4/CyfgSJ7Z7iOFtU1wJWBjgWEHdHoi2aw4t3nPG5NFTncEzk8
aM2kciHzQfXy9CfzoIOL6PpTHUPiBzI+p1u4z8y/PnlYbkmZ/kwCfPVBAs1C4hS5
ki5kgQfiz3UAw1zGSvdaYU2rQimJtQh8CeXzmgpROqqg2E0UptAVRncz42sguI+r
pFJMRiqYiFiYdodpj+EGUFqcx/BTMt9RAiLLSIfECPaa1Nb0RwhVcMugTgnmqzt8
XEWyRIoM8MZkT+KZ0sEbwlBZRwgm2sfY1LJzN542apqy2h2tPKsFhBIJL2+5V9nY
ReNy61z8F+VXBv4Gm/JChuNzXn8YDVgLgLBgjW6p+Yk1+4iZfRtjnR/MgxWFjyre
F2gW2JA7W3oGtlrZzbCQY9CZ75nykGKhrHfJSu8Me1VlL5tq5tr+wKFfMmGtmK9A
eLzYEbhTW/lgdIU+95NHbKjiZ1Sg/SUr4z2IyqYINA7GiVuejJG0fqCCnrP2fzlc
nkh4OJlaDWUn+GQZG716YLCcqIiQmCYIMZAWV7G1h/fIHnpJ2pBpXsYpLhaOIa5R
BABh1aharc94/Uoa1xlY4yd/In7LKcWhwvhnli0hY38gSqQ8bqecstgQ71QvT3AV
EAd+uMkC+SJq/XsLlwOU4uHEM9CwCGPdqzREnYtUB4UKhuyx2vEAqC1Jj0l2q+3T
sft+6ac6IEYkgGP+xAlxwpadvX04jN2iTQJfy88t89tbIN7s++fEUYNAHBPnonj3
awqEAZAqKHo/Adz6jOH/mAp2aHecUxV9wVpUO8FlAhFc7NJ118RhcbHXs+cJ7xfl
ikLiT7If+Ix1/9pJaVBGUUDOO+eTArnH5EJmOoM3baGaEgxZjtpsYcCEOXrRu/Je
JrmWpUn0s8ED3b8B/tnCG98oKZQ404xot/uksR1MkrrphxYjACJ6lTHli88GieyB
Amqw40hypK7MVDFHxslwErjJ9Ohx1YTaZ8Pp+U4bRnZF2ZJ3bBQZbZt66RzAzG59
h+uC7sG5hWm95Pke7E/GjLQE7GZBBO2DDCaWAg0nbe/J1NkXXUPLjOxcbF1CrPsm
917lvqzgbUZuU2mOgVo9uPOXrr49yQ4ZEx/aq5JLWVWUdIXCVgCL6x/fwYmTetJV
+4Eyfv9aQ9ige6LCJ08SIc1BWGeA1HLIl+04QHqIGt+mwwuaJp4nv7njDha+d9vo
iRDYRgvPiPlzPAUjpnRvfxN0rIFEwuxWztCNZAGnh1Fv5GWAcuAE+a2YRZwobpmE
nSwyzA6prNT9n/CIkqpypGEoU8a8l9c/6AJ2GDK4qUGASAKYKW26BGZosC8XQn5z
Mas5jubpd9NvV5/EMv4yklkpT0mdhgHsP7gsG+SWxegtErSpPu2vhVCTuP0f0S0d
YEh+MUoza2rKYzlTbooXIFC3jimakotCKvTVXKHyBuhcNu0YiunctULGnfMTB+/x
t4WiWCCfEBPI4gP/sY+ipFATr2EdcHxeuJsxfEQStDVgakInSh8HTCi4cTPy6A4z
jpx5K2EuTXgRuANrm+GGE4UyRdiZe/X9tH/pvZt7hrHdywcvTPweUxh2qJiKg6+h
GJK8MsBKtgdXfGWDxG9b0S/934OeLpUv+5R1cGdFS4Vi2+hbWF2TekyvbuSo+DKY
KlzdK70RS9u1u82ESIJP2D0cax/QT+vQnZ5YQX5TIbbIghGvl8mdU3NnPnjQdBtX
QH/cIIqG3OF5fyR2EBg/sZ+ibDi0lQDV4V8FUnM8Jy93KhamCWaU44JeWhX+jRJU
B8KJfezW4VUQNnA7KlaKCF+lahgWfTzWMU+p0Y9MuHU=
`protect end_protected
