-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
KCavnpqmLVmqZaLM7jLz+regR0mmJKnh/3DwJA71CYw83uJZBYFigG2b++GmU7/Q
HigPGlk1+25mqWBW8TjXfb9xpqKFN1kemcODY+reCbUdHRzrom+aYcdQ1JnuKUYe
lhIUhcXm2IwdQTb9x43mSxjTPd7ki+5FLLMYDGcDT1I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 18290)

`protect DATA_BLOCK
U+EXf8A6MXq0cguhxnv/ZfGUk4dwnxnOiOsR2LCWyf3u3/PRwW7YqHX+7zb2UToB
NZ07iSULY70qrAkOZ6SzIAlEmTmnLMal/d535Bm9jK8wriU+cuh5Lj967MmZNywy
o7QApgndfoyi1CQFOODmC6rbJDaO0wgSdJxLpJhLcplN3sB+MJWyZ/Fp4WB4oC53
d/WMjfjU9Cf91MPeP5EX31QX9XgDoXd98Jyo2ehf6HngdGrYhffXhGXCvgTJEu//
3kuvVaIppTU9x3NxHqvsuSyiqE9W7sZm5ZlR84ZT+IIEDg2wnH0EX5uuSSRom7cP
Wxkx58bGAv/aQ3Ol/HlIgZmZMIXGH3tCUVLJMCOFZKx2rzHRaZTlr0VI4x7jmfNK
ScMzs2RcJHsT+l50jMCTpOx5pWkgiGGddHh7n9c+V4c1VOF6Qs3L8CyFCmKzy0ZZ
CfTwep1dl094h+4QSpQFyX4y7I/6q2U9OtNZkdut4+Ez1z2uZqu2baDIBU4Mj3Td
OOxLDgwY5BipyqOL8BFxpXjtCvpIvV3jBQpzmP1wvMm3U23xWjkUanpY6XVUZnu/
sdj8qb7NcZ/ebgD3IjDisP6rLDfIamDSaWX8NYQGcIyWtly0LzpanBqSX4V7f/Zk
iwmOg77oJECQ3H+OxIdxPhtb0o8RzoXCSPzv2l4ouWQpRxhB01HWtjQa03nsBqC6
TvpYVnOmRfL8AvK7v7VsenOFh4oN+lYJMzpYS3DiIUHP5TVMmpdbJQMV6bisbNDz
lt+QmjQ57KGDZ9YWJXDdiv4Qhhql0e4atdEciu/tI8oh79FdF7PQRrZRIqe2SfFu
rJnInMpnnxnRLsfPes8ECaz7m986eaOV2BoFvi7HmSvj2URBdw9WOYdDuUm2sMBN
V35XqVbnjI2awWTFCdG5JdmA8O7q8Qt8/TxBoHqpeQtvI55fAqdl89C/damGeQxo
yuATEPIgzEeoyw4rdEtD01jko2xsA8E93Ka9xAPbaRUIN7xUE2HrN/kiiCYLBwMf
PX8BQXqB4eJb/yO9AyucU/FMcBlJzJNNPXv3xP7gNMIHt/4MFKAS+UWQ3wFFp/FY
ITkYCFsajvCJAo0uqzmJ2Z2orpn1SpnWBSVbgIv1YWJ4aFevdPDVf+McDqr4IHr9
YWVNdCx8ERAy33+O8ShC9HEerrYRehvukacNZQZSCcFXGY0SAKmdkVi7QT3OApCx
CvTw7XXLMafQgcy6vHo9iQ2cpvzhkPMw4L8hDLl7h3hsQH1u225KQRVuIjChDI/D
Kx5J2GuM1VfEYYU3Qm4IQg/gOe67n05WQyY0kaLc0HBtigvGuTokfx7u0incq+0L
USAVYn8rfc8cTsbi5e6ncV+PvIeWyAtAtPoOzM9ZVd6xw1k6EOvVNq7HrDGBHmex
MT1AOqzX0DaGpRwcZOkxYsJ4Ia24a9rClzkkfQRBeLEgU0w5nq+pQX/JnRBhbMn7
6Oot+KRJcSNQ1pE5wN1OitSFwGjoVfCOynjvrAaXAhKJ48bxakhkg2dxoVtueSKy
8zqdL/LeL0MOzBNQcWCFj3MojGrB8vmPjzPWGg7XZ7ChBwZ2RzEL+FW4hbS7kitG
qxkQTuIPf34TDecv8SptWonfjudA6vU6Dq5g3VS4FKpQeaX0wBxNyoRqd+O3ahYF
0ejtNoIYTonqdcXx6yBEQG4hzjB+d32LegLOOrSLiJJ5qJV7Q4rAt7c6Y9AHSG1G
uSCIsTfCwuWCTR/OVn73jVtmN0SIbe4eVJGMmRXzppSWgl1Sj7BaGPW34uZYOirj
fseilNwGlJGXn1gbFExWiyRub4Gva8J/+kqct9fm5ziUU5NRhAAKatMqXpYqnpp8
any8Mt+27e08+qxHfmpImbLAUm9GB9IqYH+xXOWxGP63xbIR/8hRKC48t71fSDxx
AbXrRCBzlx6Il7Mh+AZyKGUwn5e7mP35XejuVYiwaBwTg7TzVTnnxbWt0D6neAM2
ayBzgZVd3+JDEMly4T8DNBVwsENTtP20X+Q47FDfmGlHwQOq6uIC6x9KLsv/RbOg
eD9lfUcPQtv3lkE/ezZTaj3lP7SzB4Bd0Z8wjESUnjpdXLNeBYW5rndJ4BrW/eiR
Z+Aj/tE7WZzvtPdxO30sN0wIhZjVUL/Yj18+oSbo4t6YyPIt1EfYpqZn+gMdbUWb
12Wo6etX8CqhzG8cndBlG5WNrBpaXODtWhovU4e8crPd0udK7Bn2cFRPv88R6F/C
5nIefJnYMDMdOlt2ewV5rMgtjOdLy1KlIUToWywbdb1ibLBirySsUF2skiD57AH4
uLHFnOmSqBQldnDeEUl9tAyA+hD0HOFpqHVEflYIUToa85XwfrcfSh+dVh19AbqC
rSF3U0gQrQgnSYS/plmsIi1QrGk3gJOuOQ554iXBonPDmVnvkgTBV+lMJqox/mir
eSUjMv6u2G703mQ6jSP2CE+YtEuvbaKoXq+mHmjPlFR+HAkCUFpS3mINZzcGZRys
UAIXAx/xjlo+egzO7FuDj+HNmHFVmKGGUCXSaWPCSkDSj/OsjADCZ1r7KD4tqnqL
T34WZ0hN7H36nE1lGcqKivsZ4kqVNhG4XqYNIXnRQbN5zhIfuwom7tXm2AqR1hH3
AFhq8a0ulKrsCgjgU75uI4Ex45yxpfUE5Axl96HdOHmZW90+MHuNgW89MwToHDiY
FdOfTL7WVObb+dDHbFfoQbt6oc3YcSsVv6/dwSgtIZIlGtmGlh7nZUhZmxuppdnU
M1JHnYAx2v7bGVSJfDl1R5edMMkMh674oiSXSUhT8fdv8dprapJJ4Q2cXjADPmzh
0OCYTe4rndubNrUm77OSpOieC04YSVTTrFDK3zyo7F3HRytxBuSuABr/LBKnqqy4
UO8vWzQkZxTqQm6tGm3zA0hCPl1kxIueR8rgLG11A6AoFdd7NOPTnxDU9+nZDOf/
d5qj6MLzItFZq8JtLXyRzzZnCCVwt75XIS3jjxhHbwTJKTSEvt+IaTiUIWiXqAFB
iOSNH93x5penhbD45o9EzQuFTeepf6Vcex5R/a+8G9F9LVCbTSZmMps7ZyTHnadG
R+DWjkc0N90zn+853zbsuHK3HBb1I5gPs3mqOpuM2qfY2TwkpdEGkZ/SNaYZ0R3W
ANr0CY6tMTT2ICJ6jWDQoXwbrL1QMdrw2UlGqZkHYqHzdZBabbgjEmd9GiVqpjai
ZKFWqfWQoQ309bGdwdkARKaK+evKjn4bLYIGmw77T+GQy1Omqei1ZQ6lPpytLGL4
E26CGKhPqk9tfvoLexcKa4KeVz0SZx51JZmT94a/aacBVly4PqetA2qZM4yMIjB7
AY4dPgk7C2h6FpPCeaH5MorZtwq1LM5CBAcBumsa+Qr0qmJS9f64+AZHxnMRJHxm
oVEJooUWdgy7shidlkgQ8ChATxZqhf6m0nYrrUgr2F4Us0FWMCwwqj3m6Ads8V3T
eyRp3lnoSenxH2QzLml3fv6Ua5Fyr9H3O2Ve1HqNhgofW59CRAuFtbLokvIggHpg
Vh68/UD+Kf2zpBYPmciPP5QeXF1IfNLnmd+vo6UaBSRzAxz0udrsgzhV8CKpE4OW
964zZXJHfs5nMlvWGPtdWDq2Mkz2M3UPzLlDdXSKc22p74a/UlAk6HGDdToNjyyj
73SOr8YDHkmpF1c6yWrFwCc0ojWDaEHEM/3PMXVAmAbAKRYh6NKqjR/FcpTlubDU
vHiPY55Cc1/BzXL/xbosxPCBbuhhVLYeC61SHaVYN+rRI+uNqdX1Y9v97/MorYcB
zkEs1m4SXpfZP8MxmNvSj/YwDKbSuKwchQZ9BJ2ol5QFZxE0kIcw5AbJF9qqr/4p
iWlsMegLp0vhgd4Hb20VHJODpeUy/GfM6b1XkQmdKP5XvCOiVuKlnKYXGGUgfQWX
32XjyljSNJBHHNAUOCzR/l+VWZNz/ucoAE7y7nklfmHVIKyJZrucMkarU+F8/uVD
1PtM8uxwD1k1nagmdLmivM9dqmLafjmtUMSoy8yiwPIaODqoHsT4P4YcU1g12aOA
M1A8A0/LqECsjCLmWchCuD2hpvn36GqjckO8JMKle6chxB2B3mNfWIXrMit/h9tM
kIlHtroEoEwRMAnUkztw82MP96JM/RaXQyOM4ni224Z7kFFL892oXLpN8PSJcnAK
1USxUGmNGXDy+qVslga6WTexrPX8NfW0l0miBrB5fnTjRX4JFe9v9b9VFp1WGaRp
2Jrgc4Uyd7HIfR/RKf7FRML2eAEj6ky+UW810zndphUfsQAolnCZmYlz5SXug57v
G4wDaCRN/C2KjIqmxXZsDMU01VnYfwokxJ2nbnigbDi11jAgU7uEvKfpa3sTG/oI
yx6oYZ14PqmNM7uUeQImCPka5vGO0NsG3PkdMkm2BP0WrX15Z2s5QwrwAPdgWRl/
TrIhPJEmdp0TlS01cjvyUcSVnP9C9kWZi/Grb8nCctNLN6jFokLOQNciKfB8aipF
7cnQgz3xS+3IdG3ts+AoGplVGW9cK0MnJ6cbtC8T4jBlOwKB4v5KOWymZuKXREEN
VH8Y3pfjUu6UZvGCt2O/ITsmyzC13X0A3rPGKWTHMLzqO3otuqNOacDryrbDBZNH
nSrk6GAe1QLgFoFRjbXXVUIvCvDk8lcKC7EpncPC3nDU6qbz3zjtNeF394gCGSQS
JxYidNwVwzFaQOXNWayrUdT3eByYrAIOSVNh+z6MZk5CLI8RFNiFpkKt5vZNWlmM
ScueBxxJEwCMwbgZWie0YgzGW7C2/sYDfJozgGEraM6yxlLU4jMmeIU5XiAcXE2r
sYey0BasloXzOn1NaazTYcwmT0YmBPxhp1Co0YSqlpz9F2MXXUwdInudo8gucGvQ
ftN5yM0WqTIBEbPbJb6JXBHHoJkOMStqrNtWdYphcvllcYdE1by31qpPl5flWwqD
8rx38/g4lXIFT90o5LfbLJH4Or1WD/pXAdgcCOd6SaElmSmo46UssoKgV+NzyOji
D25SOjIBwuZahfM5/eici9m7XFa19XLvF128lHYuvWjfCHHm2r7CzkRAvYdusVL2
vq4HkciipkYoSlUj1MLay2JbZGp+rufG/wutKQBtu79acgMYTCM67K0pYY8LEr6T
hBYM8OJQkSa/7igjVwo6jN/vrbPxlM2la/NIcZjBdC6pgxEnvDdn8NMCbq8QS00+
cqiMLWGSTC4B7Psy49vIOLlycClwXNc0Caa0Yc3bYpqjQSfuVffCTlCPy4I1y7Ei
WB1voNUgOj08F51NQA+xDGis7iOeHKMNJQEWiX7bW5ZsFFEbYfQMq8t4gr8sol+3
9zrElXSNQCy5XICn0f6ZeH8Fji8XezWuWSP3gdZY42ecAAkgzharRrwTDPkYnOl3
HVmWyO4JTBJWUConCiWvqpBQDyRpJBwLkPdVyMGerrF101Nrhg6bGkmRml9M11d+
4E8YzDL6nA6IgvWh11+fT1esjBukoMDu9wwonozijF+IC7Gq6giOJFk+YHJn+X39
vaTfEpcKVlU4QELerP0WBrdVvcA4Umqa32Kvh1uYucy2NwN6mswy/2V7WC3tbCXJ
Oy9Rl3lVoIBpUlsgCQi+UAM2b6Gd37BFNuX6zFj3YFwM7BWH+wgZM77CF3Ve1Wgr
I8MJKHksKtTtLVs+0PBeObIBo0ijPdlKp2IsPEz18DaHucugC+jxkI/X5aJ2czY0
10c1zOHn2wklc+AfKxN62JGRWye0rv6HqfehZT10HH7yjjjxuz9Ica5EH+WGEf82
AkePmcu2PllgUtKdbxFgBs0F+Ws/p7Gh0dy+jT7Flb350O9nTXXm+ZvLft/YfCRb
bDZ5t9f0RC+N8DJP6SLYGLY0rZCqkSbd+aXrsX8lWBhVIJ+fFejEHG5ly0kKgoWX
E2jp56aMznOmN+QtdpwkiW7cgv+hiI7ccpXCZxCQpLaSIakVehTf/VeJZ23jBg4f
otL0WKrOzxW3m5aYKLUFOH1bFkN6ysM3OaCRGG01sE16Ngypg0q25ZI/oG8C+cwd
gmSrcjpOuddZizHqMXKTFAlg4AyTCr5dlNeVq0t4QjsOhBe5qUZg5pg0UAGdbU2g
tpYnNlWqSlmSwoDFM01dzErMGTFhIPvun8AYOGAeEPlSauvLuwG5NSgqM7ztWiSi
ZKP5LIbm5o/PAMeu9sTWMvJyS3le0QEfGNeMDja1IvzV49uZv0StXQzXJsQe5pKT
X8oZ9uiEjKwaHLL/kbW3lS057e75gNc9uFBTYIQDrzQAKgs+fL/eYBFbj6ZsD6Zi
IGmGLcA/YiN3nlhJau5VXZHOQQD5ssREl2hWRJN/YV75DJ7ByYuCs+OuCrQitUEW
Ro9lIWbPYMrp9E4KTvK+24WV2esh1ZlKc+x2KxomwuI1IguOSOF/i1G4h3aW7oCt
3I9qUq63EUmHSNVZRYGbNDzsFPS8MmsemhKh6TGv2so5q+LuXy/jQ/GZ4MYHU4Er
S6ybTQYcAXEz1WaO6VTHBWUUpRCmyYe/X42wWnkdQ/icg6nhQMnYZLIpiJ/Q0Pe5
R0OlWlM+9gzCzWcUiNnJcDH23ETBv5YprRYh3PwEru7JnI/RBppY760CUWPwW2Yn
KsgRKZBbyHkNZ7Jwv3cHCQv7eN9cUe9ENhbRsq3MkDjTeuetUNp7Mv01clgh5Ul4
xHtr32vemLX2sK5ouClMGmm94Xog7wBqVHMdKirLdYTlhTWO9dUjOBf9cxgdBNQq
NQmFRY086Y77LqHHrOibf5zuPBb8pR/qRkVndYWza1XA7oOP4uWI4+83ucv6m6/v
bgHgDK7/GZ8OARhu2DvRke4xzYEKXmXIKKp2zcSTKAAhnj9sep0ky87TfpoUut/Y
pl+nMKygFhxvexi01pA8Mho5RtOvRBCaN5QA1M2UtD4Js3XYAamgXGkEJ00JTRF0
GWLFEvDUTu3hvTnDru4dYNWOfS/WsZwmIXPerWKcBSXm2riwXXLHhWTjcHdJZRkU
zIbN/kTeL3jVa1Vv7BqDYduor+gFpDy1Q2YvePejKWA9xa0fNLLgmQAL47KmNlfX
yyH3uIqZFAmiqpKroIfaY8wJT2OMPezd7/6Nk0o9QG2/XTGs3Hk294CZIyclnPNt
WqGlG3qk31d4/Koj1EPMXeZofELH/Afy+dQMqAgRIv55JlhT1bkQzhMWNRloTcuf
0CliQlcXw/sknG4nIWiv6Ersz248Pk6bINmlbjNk5TH+w5T8oD1Zqx9fIqFJqsPR
mIF8zfyeHXcy1woHS2CGiyAVcJWpy0pkx4/m5FAmUOyEQteIq9HYXRyaM1tPFWQf
2jgmUTI6G45WWsYA0bbbwmz/3ObkeMZXeDopvXkE3aK0YYAe6Q+y58m+1pN3/mHx
Q5qwdfWa0ssXv98Q3UPjKnUPT4+XICQjGluOY7DzhwjMRNo6CwmSQNQsC2D1ObWl
YGSDUCKwjXMgST0XFLGP/4m3JtOrgZDoLNmp4Izt5dnGDKWuSySBrxaOIQ7wXUtj
iqhXHfvdoHmawsQwu+HHy/QN2eNGf8IZSslCqVajGWNa5eJzVi09IbZ2lWijKi5e
VJ2aaiJo2TxjlXIFG4oTNya9KO5e8fpic6iz2g0rnQJfdlh6fkXUwEI0nWHE4Foj
CEjVB5UKEjNyfFH8uksnd6VRx17Q/bci+rZJXYEjm8k3/IMhuSMASCJvZiRcZjuN
wvTNodfC1TjAG6ik3RfKC1hvKGY3LTgvm+AlWLPd3JZKfurULEkSHrvVcI0B/dHp
7c9oSP+4hoYNzS6WHxJOJhuOgIROc0pnVKY/t6sPEwnOZLmFFbQvVOexwCUS+P2K
P/F/d0IHEbYYd4D2T3vcyM6kuVkeg0KG5xkIv0tBDwxcsnVFzjUlrHMuuTqQg+ah
ndlEskvLE2uRtAWxtZJZ2cr4Ci3pzSnsgF/YqXOCjL3yqaQgZuV/cp3tGmdEfTb4
Hv1Jgmd/pyt+4qBOq6FcL8aZCD5aIscbvCVlGjStMZJljC54p1PBEfT812ej516D
3kCIg83j66q+axRoZoPN2Uz1Si15dMesOQ6cuI2N3fzXXQ5V/9fP6ggUOUKIZt5K
3zL1ZC5Pf+3gjFWB3N4VS34y7nnw+1eLRKOO0+4dHytURPP6PSzFF0oN/ZrEqEtX
kaC1T5vSZW6G4ZNFzeyOfL4jAtKtG4rPoKrZtJX849Zbg0fOga7kduF+2oPPny/t
9WgWMoet7F8yC/jyHaHMVHQks95GgbmIVLqmaPLete0EcmtRqNWs9tMVAg7d5Ysp
rc/2gWOinpBxMlkyCP8TtoO4Bv01rn5yejoL7IC28TGcy3NpsGCsDH6yh0/qJzVo
alLAUSn8/zovNgwv3zZyUfds9k98QUzFGjM+uZyWdpNUo14G9Smj8Qwkeh0DtxD3
jlgZGWaKV6RUaVkQPxBHD1QOHQcZ3LVMo+t/H9ImiLwHhMdoKmrqPcwekDm8jUld
ITDlK0dvfrpqO2+4oihmwHdTn5TQ4gX2i70u9jl15ffNLkY6WOiEkxJwZCwQ/n+4
9tmpSM5P+/uQyOBIFU29RikJTUUkBLKUtXHRmzmGAxcUrx+sVML2QGLpYkCoB/B9
pQc41+WuTCRB3UoSBaYFsMxnonkOZrQINHQ++tOl3taFGByPdFWV5OMKxdAXfaRR
5AFVMWSrmnLLJVTBWr1ppA8xn+8ixMJQ/6gap0+ZxDUidmf8KiwBFn+V6fbr8iHB
grZHo70fEBHpaoGlOI3twuE9gJ90EX7kR7cvLz7sbBuQ3Rrres+IPre2fnNfe0dj
zBzmsbzkmP5OXLgT6flgEx4RfwsThF4AKvdsER6BF2u6rQF088ZYdADpLanKJNPW
xsWwuMUXHxJ0Me81V+n/hYS6pHUFHcbimiF1/+Si4VHtBu+hPNYIbyo5OC/51K/4
QJD2Az63XiGr4IEL4rCfOw0C4mYriEnBqF3xtRKhvsU1wDKQkj9sj0M35hYFIS2E
bG1LBLjMQ293ZnS3LShvwpVgt0k/Q1xEAWmRULh88UX1lfeTH5xErMGVQY4t9ZvJ
7ulEu8ZsEegou0KviSzoEVkXwCiQ03c5JGqUKoc+D9FZW4hGU0sBORJ4/0+85S9P
uEg86PZMe3q7OzKmFleyUrTW3cOmv9NmOKcuo53EdxSWrpZZYK/MsZ5mdt7svq1D
YL6k0H8IXOC6+7cMa0o9R/LnHX9A4vCCny72fOk0o2RR22kTSr7oLwb/PWragNaW
bVBScGEG0mA52gAOCoL7DUKHDHycHeE1IkJgUuHHAZ43Fvw1pJCujuOYmLzA5+Xh
mdNvGFP5aBdKQFJM3M20mYzJr7IkuEzcv2blUZgpPCUOgyKzj4nC+nWiPPeViLZ8
FRJ6k7JrzvsS35QyTE8ggIpIP5cLwSZOCm/D2cyQ7VdXtX8f8lzlxanJvZcPdQY3
w4J3seX6STnGlAIYjb0Rr/LwG3E/KwXsrmGQGn1HO8AEZHPOZysnSYUG6YIJ2Z4o
N1nFAypyJ/o08ovmxvFCojttk3QKZtUZyoghxj2tdoWYr9v641ktsEWosqNfVrD8
X06IbehGpmh28kCnuAlS35ly8eJsNTp9Lob/gjwh3WUWO+cFsp5xIcrG7l9P9JxM
+8GvMd5dEU0jqXH/esQ33ckApbCoGrB7OnOHnf36rUPzQ8dSa/dYH/vtKBnBhgEg
G9HMrzvy46SSzNMx8oqL3DzwRX+3CYf//m2BgGky6yKGk9NiVXwFKE/R7W+3R0J9
8jxaWspoP57nQX8YzL+2H+/z0gFXn9FWs8skTEbyvzCAKXyZe+KakvWodm0qcas8
13GA65lWFDJbsRMhMvJr86aB56lu9i7AGWDiwU7tdAr+mcQSpSSeoCV8WOrn2+UV
iAn+WDgO55Z3ALwcVguJD9FQYDonEA1OvERYUAE99Ji/OzAAkUExOtLqC7ibzPb9
tfsq/Vv04Swv2SkoWl3AfFglYs7Ha8hhMN6UofLKgm3dOP7v4xQhpX3CaajfKZzK
5kKJiCAzdGg2wJA6Y73XQ/TCZp6t8RkXBT8ssQSOB36IC2aANg+7iZBxddzqcya2
Q+V/QcbXC+uORuUh+1BupnKUWV+4/MP0C3aDJ3ytMsNPMEg7yTRGB/QBflh3qP3L
mhnZDkb8d96vDqPNZ2Lv9a59WZd7AvPVixzA8mvku/d6QjZNUlV7ATMjR79UOO/P
USPANXDGFzIX+73hXBA7ko3jNDdUoLRsX/luHJm0eCIssuaLtRDA4pVac3D7pB+Z
GMaAgQM/F8pCJGlRQz7TXlcqrt0f2O5wQFJc9bU3U5izzXoL0Y2RjPhMFTZUwceI
SnUu4JfS0w1fosZA0HClY61nC9bCCFMh5HCWZShvlFzcfMpSB65XsKMbRbVGospk
qErrqEGbuT30X2Kwi5zXDqCWujB1lLrCF00XLH923cTqnpf302r5xnEnvImRRRpl
lxHJRDoz1qFs+7sDsZByYKN6l4PMLiaxPnJsPXsAe/ZUB2sSsZSQA/SP+kzFrgAx
AVYNdY7h7dNYwgMOkjNGWFEXwRiHyBOr2cpstycf2QWcl1vR2YZRUFKE5yf5yiMd
BGTrsmjeb1+Z3ul2Yvn+fevnE3zKRkJ6gZrf5c98OalsuOO0DcvLcUpvxRfOq3z8
zfw2DaltDXyMA6Qf6xVZFSi9lZ8vwFyLyH2d8btUlQule+fZDRG0vaf0Soe/f22F
NQZHDar28VGqaazVmA1CD1P5I1HYaHcZ0VDO1YjgBy02o4leNjUNXqbbY6kT1YgN
BOWdGucpjJlkkwRGCR9j1LmXJzIuI0UANVYuTAb19VqC1982VUN3JaSSve/pnGPd
wcCoLW2NCgARmktQNE5s4H5otajgiaRUObRawzzQ9aKf5nU4pHdkOvHEX1t8jM9N
6xkfwEBACFa02T+ZFewpSzQeKL6tXqH/VzWEZdJZdB3EoTZJeGXL+79mvYTlJpyA
VSxMZBZvGfOsMGyCdBjvwgyDAaJsLY622JeWRc9dAmEhdQokcqaVkY1kcW9KnaUc
47mfs06+mOQL8J4C5hmEJTHRrI7jaavwgREQ1a5esJyCOBJioGW26NNKpgBPYM55
bwVhByWH2wgcZHUWMB4cnnpTEnn2wPbubSqwwq95TYHWQus2RdAFZyGI4eP1mu9T
DbxDegE+xg3xo4XtRqoxv+zak7T7HbE5Xd69jWhzpLHF7fobtP3DvJn3hHKZ9tv+
67lgK8+4X922WexdRFBaIluFOI0+H2RvYGbwREGfa2/SzGAkC0JcGa81U4KmJ97l
PipITZALR74l7XxDR8Gqmnlq+96zs14wriRhWBSw9t+dBLRKGgdrWZzv9yKe2AYd
wHpF6GVhOTVZ5tp5B4uzznL2X777J/AflaGIYVKTnnEsXA23B4ZKBaHF0+0l7Pju
UjPNzvPCkIIQ7rSrDBff1EYSi7cUDXU9iB34Ykt8+mFMuY4BBo/z4JYSkahdv2Sz
QWG80qREuIpaXCx3k7u18Hg8ALkAfRT1zidcnZUBsPh5Q/UyzGJWjGHIanLGHBYw
MhFBzJbw0hADtoyGisUT4ubYOqKvTMH3ASvz1lmc3uyTcVkJNPtHXfVw21nSTIhq
7e3oPDYLd9Ay5ZiGxEIDp2ASxTGjx/XsUsTDLM6KbNYUNixYYnk28w0XG3ZF/qQ5
nIcdjqcHby3bF2j8WX7PUz1KnrzACqyjvuw5H7w5bAG3VghTPRMEETAb+SzyHC9g
/U+Wl9TLsbf0F6y3FMG8ge4DNq3fGwNwP7eHMoX9UvRPY+nHkSllc813Bf7XKNie
GgdwePLmgC7lTyTGJRrvfcU2QRnT4U/nPuL4bhKJG0GgFAyr1Fm4hIx5FwzaJ2wh
hklcJQUK9jVPgCFGBvdQFbgPPElkZgzFd9bJgXQKTd1oK/Nx/yKu6c+4jy0gRXBX
JIayTq1cmbCtRSpVHMz6NFGo6dXvLa+/ncyoIvy/iKFtrKHNGc45wjFZkQsiquu0
LXDhLLLvG2jdJbz8jCUWp081cPvqt/MyaYztviYR6UVWj48njm0HC0jDXqpUmsAR
RpTm0fcaFWPPnVPIVC8hj6E4NtmWA3pTrzjbJNQAifahQOUbha48/2G+XVWhfens
h+hXWMPEabae1Ft6iJm3wNA5lJyZESJgmy6QwbLEHdkrtSG7hLB+Ft+Cs6KGyh5W
XiHV0O1ngG+spfhucIa/858JiAmNAWErlLNWhiutWRevDGH6YQbFtK/zbSTES0vy
bRvJacGnyns3f78wlPerXDpFFYr3wLRm76dIM8f6oOWEyIK/opFJ1zfwW6WaWXAA
HxvV/b1ywcmoWHF/8C3L2n4fpX5FeSwpkZV+qEJ/zqdabblD8OJlM0pnrPeA2+0F
Bq/cbhiCekQLgXdzU3AkzItQx71QHidsfhTm5aTbo/7SLhlNIiKr9w5n8wkXD+wn
mGd82v/0lPGuL4XEMgBquZohhCoKXkmz35tg9koTTcXXVYgBP/dD3tOvX0kIAhkr
0NRjR+luCMXefwG7f8RpMWQG8pkRiZQMw1qJM3YO6AAfZLSR2V0E0QWBPZAQp5WI
RdDNfFcJSni3ximP2/77bSgGI2gPzWLjgwgH05deRFD8XlXjscaKFpDybEiY74Tp
Ba821kZ2bZd7g8DcUleOOi6U3L1tm7CVsAakSstTjuDiceWzfD+mUhuI1BN1toki
RvFc9tffbPbXuKiVPPBa6IOmiqE3LcY4Uit2xrGniI/3C8BEchJyo+QB7nbOs3vu
yx1RPwHxhx5mc4+LaS9xvhUpsSo3EL3yfY+GJm9zB9AlOkVfWGtU2uOKpejc7TXx
j0cn5hErIB4aWNSSvff8zYzNpnoJ6pA/srMpkn2QmZ6czDgpYx9gwkNAj7Y/mssT
7vjGR6nvKKy2m4xsrEbbDs3DVwasRtL++9dgen3EdCzloEMSnx03RxEi7ibf5b9j
ULYhVCkFZLrv/vlQLiG7Kq00u1zJoj4/0UVl6976ZPTWot7si9bJH6qAQJajn7f+
9OOtpVmkF3aZTP8layC3kOztRVEnUFM0nEcm+Uh3ba/U8+dfsC+YYCV6AOqOljWh
54+QsGbOba/kTmZ/Pu+r5kCijRYysky9Dy1Eyh93G7iJSavsuNUs4sHiWRpCwHJ+
nhsiFH31qjLjodS+X0WgBZtJz6oYZphRGOPTsXG8rd6+bRjWh3oqq9Q1fard/6nO
kDevV/TmJEWb0hXR+VRtxMYJ14PrM/iLej+xqhOBcFFOkQjZLnC2P0dAmZsb3yNL
1S/l1eorRIbjgf253hXlJRLX0B1Sz+PjjxM4O/lixf9EYEoVJl9CBJK4ZT7NBY3Y
xTtOo29pSlvWnEfkZXSHcAuo3/ZNisQVlX0DUYsmQ569RW2lLFXbbeLVcavQl1yO
sIeHTqgb2h1Cd5PZ3lm2rumWYi1RBhWLVQMPHC3z3huRTAlYANmNttStoQtZNpSG
z1GoXtIIzUlwkwG9LBV1W6bUhEutz4xaEg1jryWNzTxVEj6y1pR31I9ui7nwGtED
BvdeRsstHhY/RzvCSjsK6yoNw0QIIoSzi3Sw890fMaSaMgLPqEQ6444HZ0kNUg6W
jz7pXdd67lZ5GKiJJpQ/JRG+sOPJig7vCOND9qVk6NqZfVu6uSLT9UMKfpXgTVtd
jDtvHjauKT1skcPaQFTPYFH9j5pS5ScCeNZCjwjxL3L0+gQIS1oa6CA1j8zj1yWU
Q9eAlnYf6jrKEy11wo7rse4mOEwAK4kcl689olZ/XnhcuCc1g6z+wegbpT520C+m
xbcDICAxb7MSBsXZXh2YEo/+2aIlXvJ/FY1O3dX0t3ctj+zbQZXhwR8vPYTDcQ8p
lJzaBUuoyO3oQ5DsPXFzXckvnHNbkjr8oJuROZ9PYiDkZwxZd9GQsNA1F1iSoy/W
nbFoi/dMIJ0tHo/1F8KssMTKYPB31aAv9YfYhd0qLUQlbsj0WskOw5F1rtV+b9Aj
pykpGTkkf9IMG7Tb3HzBlV9e7b/ulLH9mWwCynpamVmaA0ffQhpS5xKMXQDBpX7O
z97P9djmZO34h6/hSAvc4Wr9oXknG3xcJ2UMXp7UP5fj5kUT2SdjGYPUWkSVOl6k
eCZ7sIgHXpa/svKs9m0r5J+fNdsDzQNxYtvYTQQey/oMY28EM2bE3+AT4I7IfG3p
NnO1HcCEArDUdr6uoXJ2VvqSKabs83JA8MDp3WqX3ESuhZ2qp5AkZPzqBn2oF0Tz
NmfAM921nUyG+2iaLvTI7PInjpewRmj/xtw3k1TC4XVul5SBRmWHb90KRI5R5CxF
koef1uxSGXw7royu8uPha7feuogplGmDNhFQT0m9ucY8Qb1eNAEjnuwVbBZuvLWY
57oiRWpm7wUFugF4P8GUS5fZxhe+dO2AMtrKwXYUaWM7jmh9oGsXca9yO/V0Lkao
c/5+gXj5ISf7bX2wvZ+al6a9TXOzgoe93fI/8CEZhb0w3jevUas2Z3+cpbV/eim+
KdOGrxjKquECdHdkDXxl5bbV46NiWx71G7YXZgW/ujzjHvm03vEwmV6xixLSVoRa
yhSTyFxZDlNqQhGi8dh2KWjyYh9UGelfOjgaPaC4Bb0rAHAH4oKuAVidk51RA8j0
yuUnuKAr2MCCy/3nZAji8DNImcZRzbVCvmzLJR3EhtsFu6BrV95pzvd9JXHlOy86
A2FtD/ZIJGDc7KfnuoPN5EFXEFNgQY/5kV2CuJ3sWwkgPf+M6+RZFia/mFVZSX/J
1SOLOyAkI93YjC5kYfBFxG9ZZFKdwKbs6LCBiVtOudBfLbD2tPaGYERTr0CJX8eH
kVnH4C/SEMi2VXvGYmU5orXABYGWFlodNJNzijqZ3XG/YxG3pgsjtVb3X8CjfykK
98+c0EFL+H5AtD1MpAs3NXHn0glgKwt6xRc6Yv7/72QcPjcJkdWyRFOWt3oTa6/X
m7Bb9Q5bVwUbo26+y1dXUAwZnh206/rtJXni83rcwjk52vzUB7AM6uBUIhqXnIpx
eR1PuZ/zaQBFkFNz/P8zQ05MI3yVRqHi6KAyCaC6wvSv+cjhjxdvfBLfdLNQXieu
gTqjvEzm7TENEHVCE/5aYLREHGddsUWcMHRCszMNjj5tHMGHBVJV2UhNfSaKmNBP
VrpFiPH2Bi1Z45WXyVLUZM4XahI3HvcWXcHVo7W2ew7CxU8kcypPyaBzyAMhv5Q3
aw67PCbRO7+xIXwHnQkurlAF5ICd4p0TSPZX1zmK8t1x1CY4qR7Cc7n9vimqo8L9
HxHs1eOGF9/f9j+HLWhHgja/yUPXhXYqCcowvbk/UNT+qlDEAyibp8TCCmt97Rl9
qZWghgL45t8BulipozaaEKecWKDVgsC0PUDtfI6NnA9fX77Cx9w4v6SlcowC2dlJ
yVZXEJw6OI9eB9uN31zSm0bu0hGJBSsr+xF0Maaiky756OOE2hf2cDpXzPCpz9BS
dBYrA8HF1k2dqVvJ2Gy4Zh2hft2kms0QQY1b/BM8QVp6dwEfoofh+rtscZ7SGdCw
SM4dRs5LiZHyxNLfMBw4kbL9OFT8+GfFOSKB5FTg5igakK/LwLWW7bxBkhxO9mAJ
T0ktiMt0N5NhgIJymFmCyvSM8f4d9/FrEVVWW99Pi5//3kod/gNrXqlF/fmh0jXt
ilW9uTuvCfbmr+O6lpjIrj6DVKkru+/ObKoqSJ9ezyVDwfceo59uXanQ7L9YQpWy
oSoVU5GBdXvqZy8FnFGH+fhtgrGInpGwm1gPvYXetGtZ+UIJ4erLxmMs6mGgC78a
r7GY90UBYLSyAV/zdS61GEsVTl4uH8n/uTJ+77eNc6IehI7ezs3mgkd3A6E7S1qA
eEtShVfo0KJIZlVjFhF5keIqQJmhwoY4HxTK+gB/J+SNz0me2F0P9ytSMdOyAaDm
L52T0/PCXOEWkjGOY1D6uZW4qxjJ4P4s3PKSmsdDD/Y6oHdHNS882a9zYLQeAgkN
wvEWJVCfuyzqLqoS7HN24P8pC3rIM1NmtyJ3EtHDTBM2wVThfVdpPEPC2Z0Ub/YF
SagiRAjcKT9wSC9fq+9W6tf6qZhaYT73+JCjT0sRBAzfsz2uwGLpIUzE1BCCm5ww
fMr1igaJ96B4UGxxn5aTBxMFnmHyLQiNYBmda6xLoWlqh3SVwTiDn0zQnV2i3EmA
MavkgJ3Gsiyp/xdCa2grbnyyTr0ZxGwjoyi1bQ4A9M666FhBbQHZzKdW3U/6FVAW
mNJyv8RkhXkqkFB5xFUQCfOpoRHNVEzztoiyMlPmjHNfcw4V7VgnJ48ubjGkA6ux
Q+epp8rXRuSxie9jTxhN8vrjqm373AviKp3zrGP+eJGvqzFuaiPkweRX/XTRVXHl
TRj/XRh4keq4sX0DW1sICd8Mfvkvk4+O4LdVKi4hWRmIAVhMtn97tg28lXPVUxw4
t8IDYyUk3AlugA7UPgdmwcUwnjxUnV3HvB8P+ZoWddLNEjB5gOmoARakOjox4QH+
L0RuXdmfs1PKg2AgKoR4dp3QVxetDULbfvJ5zkqksT1VHzEuDGr1WAYsSTFxYkqD
Bq4xYHhFfVnOCSfYukYEfMrWCwn+UqL9pDCbZNt668LvAtTHxELrx4eRv6zYMu1R
2nfFS0HLh+2bmVKLWmv0Mn5ckme1fhUxsDnm7K8x7ABaOQbN+UTYPJpVUtqe74Vg
EikY7TVLZynPaUR9JdKSRelAtmbSIkU0/N8l4DsSNT22fkB6DUHntKYZs9maNP3O
eNLJyzzF6VA6l1fwRmhMCmz8LLKRFdgIWPZ7T2Lt3Yv+Vj6x5svp4LQ+HvmoV3Im
PMMarwGbHJADwfIrSAFZnN+7nSTbho5rsxeh1LYnvh0EzyPYAzb9lTfyvW2ykFRy
T4i+9L6P72nYu5KDFrnd6ZBWDFOcBAPHNA7ZDkCVpWcgKdHnVANVw8tcinNiLYiC
r+5twM9tuVCFA+1Qn0WBmzie63IjJEDlMKvNrs0FuaXJy3zy2qkxHPF56Sa0/NSK
M2Z+odiN5CHFzfeteN+5+kGFBSzKYcvzTOWz0OyaYAcThjDo0a0A/pPVEiPk94OW
vaJklh+L/pPFsL8QMVDZDs6SkI43WBPrCLtf1tle5b/MJgKGL5rnlFA4QwYu4zXv
NJD0gEyp+eJEu9t8wn8b50uWGgB/nHdOteV8cYpQlx+Fv1pSBiv8TIJ1dxso2IXe
uhDuYpXKmnTSujqUJHbhT9vlnhg/2GxKyO74/0a1QXjCoRSj5xT+VWIhuSoRY/TB
lt6Ail3tmZn/btNjsDjXcCguQ0CHttKsj2zZBto0cI1oyuHH3oom3KP1qHxDwEJx
Jfl0Q5ycQkzLUSRd2VY8NseQ0w15d1O9kK8V5LeU9jZa0guS14yyCYr9W88VxekA
hOun5tYjI2QWPTkkMWvnkh4oQw62FfB+ZzOxTJy7BT0nXKwLf6eUOZTLW3Hf6CUm
qWkEfgxHWEOiOJ0iCpMWQ5byHkFeFAduxmOO6Cd40g/tg14AX7KhJ1OPT93TKueL
jUfrWdvGCX31Ug5SSDR0t7ZMx6GMplvErX6YrNvkr2AGF+6CqfLnDyGpBg7ibfOC
L2HwuyBmdblxqoBk9A4ViruE9zruZq5x5xv+luyPK8evP6KFLNPob9nuhzpqACcJ
I5eXqH18/m6FJSa6jlZ1PtJvTybAzDuVbtXeO2ddMgS+4EWl/x4osq0BLmnDszMT
80at3tlzRj7VnN4bQT9gcujhab0MAYa29lNT2ECjbogKGY2z/dpXWlcH2doijyQE
QXfC/ypmAoHwwqjNktUuz9I/zIKCpCfONhLit4Hiy1QZ+k/Pcpp2FAJKSdCo24Fd
9ou+Kw8J3zFhYokPsMWznOmbZlpaU2L9E1tf1hg1DmqYLV5qmAtQSnLIVmjTa5gT
2V7fNhopprRmrHrf1pGZxnhQChVdlR+O680fTQ/UYvJOJxRh2sZDmyflJzf7o2mq
siP8bTj0zoh4gWYmqk0CKtkVAqbfjEDJ4Ixsrx11XS4NBkaxwVprVP9PTghLOEym
nvO4p8yAooJ4ukSSjWPJDzC46cvEJUrgIMaSRY3Im7cP9bN2zVOEf243T61apawf
jJTWquzxAWY/1dOxptL5Qu8pBObRkdEJh8q6J8dmZ+I8m0VO6JEowXNFSh2WR5wj
m1o53bjLaX328GcpsoPZgTssowbgo7JRdO+36AS9OOn9awCRPGZz89IL4cLGDlnA
7c0q+7jZ6W32jOvN3Qpe1gCLaH7stLPGz7Pj+t8mThyO4E8MZUUDBljQCMn+v7Vq
wpP31FoB7+hHYOO+MuJeEOmpHonJ8I4nmn7dnTJwyJVef7qX0NaIaZhgGoRNirzA
+5UAYMjGJmvK+q58TKz3PoEq3eTuUpQ/la99SdEyuFr3/8TGUi1TmvgO5TQBfodz
laGUrAGCqMDCtyrQiA87vilCtjQaWQ6ZSueZabHAMfw4eDpkcNfXDkdFcC2IMHWh
Ub7XJtXg1GGztgO6/00o1/jbOkpILih+Ay+SQcmpQh2RC2NtafHAVR7uyFRGEDyA
jIDeLSfVrWzXUfz7y8qtzj/8RXtb++DAfmqmwXmNUbluZ3JqdU+rjbYl2VbYbTxW
1y3rr3syBic9FMUqsNFHIzhfqh+eDg8pmTTIJyqpBSv4aENFmM91bvTRU0ebmzq9
GLOeHMeMkvge8iYzIR3brmy+i1oGJi8cijCcKS/ID4NXn45e66k+P3WRw/YgiRHC
9aCQmxvn9AOREFBtsG2N7hQqYUDKeC6ZMOUE+LsjNoPEOaPcNonZMPR04/jnMD8j
kc5w7fkyYkOAn96NY84eNYR4lF4oKVWYgRhkHWZz/IyKOWM8abbRT3iwRAvbSs2+
5PQPy+OvzgZl8qxmSY8Dyz4bF8Hw9LegfbtUQRy3jgAN7smrSvtfyXu4ZzffcH5T
oNJSIDwtCU8Yb9jSnqIVBirqoRvsRCvzur04ooTasY0f8CVjUuB21IvwDA2zpJnG
X4wv2K72GQfWuLdX9BooVsx8x50Zelpn919RWScQ/qqzhwOJaSyIjQSzCr1ShJqQ
zupNKp5lP256F//CxDVn+v4e8poGaSM410RtObnv2Bkv8cczILpeUUFZSybw4Z7i
Z37j5FykiRGJUSOQJ7s+Bkrqir4ieLB2GFIoaM/s+WaHSJTVWaUmddfKPMcK0fmA
H3+pxj91a9LhXmP6/MrwNfRJEnYcGSZonB8dLpFIsKnwwMfPHPQP/unB7WHerX0p
QpnaKeEnOUpGAwBkoT68pPBzKJ2mds6bNNMEuI++VCp0CCgNIB21iRlsMAOaZkmW
N26s8DXafnn9z27Z7ziqyNtZma1WQup1gf2PsRjT1+cqkwbvfFMmgz8TiJ6pZSdt
KfwtLS/Z2IBs+tUvz+cHYVVfjPy4VbXY1DlDN5+0lInZ6xiCyHv0QaEsveeQ8yC1
s1ZpDGImq9w+E5jDfY2cG11Yx8yOtB2YCzOLoVlGPNvljakwuWf8ZyJPC3FtRlv1
bmB+uv3+1hmf1v6BzclgsaalOkJ/YBS+NjhHroh5c86rbjhvSUotolTybh2la2J0
eXHN9Mn91z+lDLRc0aurKzWcHXyaCJF1JQ33ovWcwr9C3ke4csAz+WvNeY1FoME3
8xkayt8Wh2SndthRXke3/4FxKEB5HfhvTs0+XOzfAAAvoaazFcn+EG61gPXyj0Cq
QGl0bCAQ5lqA/wakAtUzqIpe8U1ENR6521UBrWCfhX6nJt68tmcOzrFlV+nDZlpN
dy1BAdoEzxWYFviCE578dufG96KcicrjOfLcUwSS9xrk72ozqJhQaZ6TQ0tW47ej
BdQCS915aq/IHamPxr87elLcGEZbLe/nyoTBhhHtIZ6QSM2EZJjBBWQbI8neEG23
n+Amb4N5WWCAhth1hUbI2IHQrFCp3axBeG5o1ewNfBhuydz5sBXtFzQONtSQ6QCx
YKwtX00q4YiA3LYw/xL8wS+SuAr5moaXKwsxmj2mn+EcNh6UnJQLlZTyfnvcV0wr
OGS2D88do/YCSPEdsvRIEoMc9LBZl9ip2L3n14AnHHrZ4u9OzPnJaBSx1BPidrWS
epNeyTYfbVMjaDopjRwbMdvDjvYF4EEZJDX7t5AJgPJ9nJ3Crl/oQ4JK+KIlb2D7
ySrC7SbKgTuqJIkI5MVf1Uhon0CDy4IrYt8keD3xG6llTNDBOdWMbqPvLLDa1IDE
9Si8s87l/WCd8OBrEsfzgcjNgwmmRaoWoQabUrWXK2g/y1y8cFodQnby8nBNrmJV
0VzCeqF1H13vcsvVOzrKR+JcYfGk3n91qjBLbgdhEV6VNTSCNM+97vIebmHcGJFq
7AAYUcwyd7FzkuRtvxXpYj0QI1fkSmtUlNwef4AJRxcP6UW/tTz1AfAmfTBrm0go
qqlxCnqXgXH7+pQwtQfLOOODVGs2FndthJvCogQumywFU3emh5NH1bCe+OwUz4g1
m9tm0WCaQTz2kRwgUbjeHqU/XqKctceFVZW41rxLNo+WIPJRu+Cxjr9NemAM3gYk
yL/DqW3TDickYazYd+Nofim+qLV2TtLzjP0Kzx+qCX9X278rC2VQxJqjLVuPpEw/
x9CHlbJFHvPPimKc5CTIBCaF7bDJD14+fma9sDMa8L/WeILuaCZkdPHk1bl81PnD
Tw4AC/UgwTN+3sxTR1XlLaXpgMZRoTSYygWuVDj/hpp8Q5zJGl1ebDGaemWYqaBH
r6JWFYl9M7NVJvMAc3zA4vUZ/v6yDmRRBjw6zQ/GIM3Lpols/8tSwjIAQT+Nid4r
0PLnpeEBldhrt7Ig+Z9eYXAiF1fZkwQwHrePrMxs7R+Nk4mhI/QdIFEqApbheoRB
sarp5M85fu1GtWtF/SFW+tZrWcAGFMXftgZwtAzqjU2O28DgJtf389IdIMlx/vUt
MCGTI4Jr681RPUptR6La8mPonl2cfvlqrT3sz3mhd/vS9K8LvgtBO4iwKynM529x
6d6EXKHgSi5FBEeEwFFlRIIwKtXHE6RuBy3URZ74bYjuqtbFs1KBBqy1IgD4/9UR
WctcXqR2OLHomLG5ZLNmG53DqgB/+3gftWUPF773HzbPR12uZ8EsVJ+/uo46XhpK
6LWHSk8eyarOd7ct8+YzT2YwAJPHLFmETYdXyJ6rV7miOHulWIBdl69KR1GYv/j6
sPBs+dHktAcgxaU36pYF2w4byXmYx9BJqbWUMhVK37luHZ2i1GSUqH35Gn3C/5Pj
OAdsAxYtiA8bXctvGw8CHNOfVJgkxgRUbQMUwfY0lx/GWshk3xGExQFVzDeLYUYS
pTEoNNwJ/4qikYFoHvNBsepQFdV+EVXhn/mxbWnsq6XcMzsfjPffmqsgbfrQ560a
EPJk5/NN2nzV3UkgCSkpT1xehhwkJOKoP3m71EYv2Cw5GAkS4Jb8SUGnRhOUIvZh
itjV2tnYleVnzCDhKUWQq3Qve/2WUc+aud5HJx3vPMUHVLaFu9D5iySzk82RGpra
2S/adHeQVz9D3CAvy2JZ2XVCOmyM3apROoMYkzEOLHDd1CvSrCFOhISBVoFZl5q2
B3EPIrNIrpCn/1IjCXt1oEQiv5A7t6bCmV8cOAjzTsDP+JGcJiiI3mIthudZEWWU
bPkJ59Ifr+FV98KvCiNBSeEONDzSQ+k+7zJbODlmeyr1Mr6XDF6IBy6QOSV2nyoI
4ysV3xtKI6Lh1uFIxAUPXLg879GXwNBpI0nhqGU1hfCDbR2zNGCI9x6/d1oz0VtL
udXHTrXtyAsDB/7zJ7irt9+iLzavNxM6mCSYGiFtp+O/NMRKfSghqHv8yVniIWrI
LwQ0KfSWuPSkMvIETnYyZZYamfOWj6O24jck+ibPvuL6uS6kIw/2bwzYqh5qv0Ge
jLxRwQ0K3OImt9L4Z8XVPMt/iyh+NPHrbOOCmBB4Q3LS5opYWuFKxFk0z/u+/ZdC
YYXYoyK2yAoDateEq1/7LGPYYoad0JZ7avqLT3RpEG6qeNWlfFOCUf8KO3ZbUtZ7
PHuHe1wfZki4kQEgd/kSGG0T2RlmsMJ830qpK53OrjjEqGhKAreB+0YrzOMRqV3c
2Pc2y+8YPNiiGxZ9Eo4W510u7m4+h1NcfxBLfixMDmxD/e2e9/xZwj78DCFlN3tS
dsd5c9Ne6bQrTyc/c1HEnAY9pnUNIMtQAXHMbqLJ33qg+f/3Cu54n2fh6xTwoiG8
i48TF9JphTnazWD8jgV8D6+Gbrw/Y3Fj3ZPw8aH8MHVG4I6ziwgfdPR1PZuVhwQm
+lzxNACZJYmDaVf5GHIg/KvDe880YbhJ0uCVIqWR1BbbP8oZqOSbnME+AwY2l3Tl
pKGx0oGh6msgl87do6HEBSRcCMQjhC5EdyTf4FZB6IzzyBVdPLMwXYcfaQAkN+Lx
dKvN+lHd0Rd2MplOygpMvMRCchcDJqoYlnt2g/CyPA+DBRcrvVEOeLNFHXZ357ho
QdCnmjIFXRfCo8H7m6QqOuPGF11xgh6qF2z82KCniBUy61776+7F87Bf39E5vMQi
aXon0NzeKnZBRoLnpcIoM/etzrtHnjJOiKrZjX5OFEZ+j8Ou9XBdzipMTwANogtV
LbZw7LKsB0EKysM5g35Q24TtyMeZ9Fw5DcYPCLmXNJLIm8Qt9xtWHFi8VwRK6cEq
ns8N2lByHkCY5NocIQ31idNBKTMne3PPYE9RNK3AjKHRvh7thYo3wzuI/5MVqKkj
uVkV44NJzq6Y8f6uZcdl3OkrCn77wCu2Si98J6CykEHIyxZT+XQDHUjn7dTk86FO
Pm2qtcG+jVqeo/xGo27GKrrteINgiUdDo0qIhvZ9t7JErjDq63BVPKUsqqgSicwS
+BCVxs6f/7CgeCpn2goZhH0jQgPgU7bKWC3MNjUnbY62EEERKzCXNqd1WG90Lm/H
TbMdF+pjpRIql7R3zkGCmOp23Ybf8Bo6+nt5wNQszpIMkNP+RrHyqzreHNH1dfKQ
dvraNuuedsZZoL0gHO3tW8vHWsD6Yg5PWzh+eaNkD7t7uTJJO7Nwj4evWCvPSqS3
cU3mjjV09WKZ5XqK8YjKKQRfptZ7g+9m7kSvhP3TcgTndu7xr2/Iu0zs5UaINh3W
2nw+PaRX0+ZvmYksGgmioafWhZ44WBF4VZd6PD2CDA5d0pqbNN/3t2j6ku8YdQkt
JOzU+yCy1XqhOAyddQh1/Q9EGvbq0DZBMzZ3zA1QY1ZYLM43OmQlAXEilM7+Fwwz
YkgY6wxrRxOxBP39sSYLGygojx16/lSkMbHAZDHV0cS68tM3gv+YPzpAjszswIRI
LdrfLDjf74BdNC0A8lUEG2OcxLUKBWCHCB0K6wLlWPbY4DxIvwVLSNoU+yAjmtXr
lamagU/nmTZzjZlOwem+ccH2475HXPc1eOWHz5dl2CjqbeOdO0K3R9tyimG4cTXa
ael7dg2REmmZTaZVxo+c3d4dW1/Er2eSH5ah6OWZ0NXtTusmrCnqZ8qBLzLj4Qcc
KThcVJAna1uD68FOWNm06lhJbJvWZNgyzoiGtgH1lEWFShTsAyHhLNF7mAZNBl7a
oOXlVAa7CL+VP2KRzQGSzH4ec9noyYbFIYG5O0olwv8HXr0YvS4+CC/8/hOT2qkc
Q1IyP9kFJXif8S55bLsqN6cK+IXaDvTmSSqscdtzRSEvakvq5ErCWUiqog/6ufex
IGkRcfvKcpHKbFrIco6FNbqO8e4e7qB079LeRqIIQzakz65sJmMYQCrqk4uXR3sQ
F/i1LAXTgSo10KemgqYdmuQDA07ONilta2flhrKYZKS0bvVprA7rIO2UY7opOiQg
/KT+zdNg8Nwn+P8HFWOut9JLOyOOOarSQrlbMNX/prcpmJpv2beSOKWaxc7QihL3
Aw+Uc8rbOL1Z6NGG+IKgmrtHUvufChIuOvWjP6tnTMC4veYb+0PIjnUOte0XjdEj
dYAyfg4WcjPqLUH1UaYWB8ch2D92zlqMoASiGwRW7+A8MEu9IDyXBOiFdBj3Nqqv
xaLqE0YKyFYPrKGL8JByEeIyZjwdTIr1SzvmwBpQQ6i9BUvZjikU+zYmHVYmcjEk
UQCzOgbvanRWyOupwJ5Oq1QwImtj7dMol4xEkw+2m0OnY4LuKGpSMvqu97VTVDCv
baTFWQTszgJ2FOp+hMUlws1qaCKS59Qh0B1ZYDpPb4atVHyD50U4ErEJNAPVK0p2
y3Y1ShGm9TdtJ5jyJ5aY60DHGRnPSbvDudpDU8xa6ZvPNk5jWN5WNuSCV4PTZ2xK
RK2+UvOTFoY0BX4nr4M3FBpQAgfV6F1XBmt8+R/0VBazXZQNX5J+aglf87rIQgRo
+DFlyn4+qPxxyUjVmu+i4Fe+5kSyhy1AXz0Fi/9DuLTcnp5jIVMIYcuNdKAsCNO3
L4obQ9TnOclSBo3hiHQQDV677Bwruyf/CygYz4Hm46DsBRon1bt8t5dW2/oi1daK
4GPHtoovCKru4ddNe5gi6HYzlCc1KggohubSaWprJJ4=
`protect END_PROTECTED