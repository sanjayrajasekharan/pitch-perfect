-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
aELPdEgtXQ6KxsDn4Ze9Mo1RxnqNZhRmtYdU4MhsKOVy8XhWlifM8/ZMKfV8kt1a
H6OEkV3wnAa62yjxBGvcRpGZsd35cFJOhFXhzTijIOHftfHZKaXaLGmK2yW2umaD
ONUyo9/0eRlkq5BRAGdEohc1gHQHU6JAjUeeU7qFjpiL9tTn7bpb8A==
--pragma protect end_key_block
--pragma protect digest_block
T04izCIT2/q/UyedEL25+OD21uU=
--pragma protect end_digest_block
--pragma protect data_block
KTwVTX77jZRWUIZsiCX2QU8YVkr6I9fcSV9sPA7y/1pT+NSUkHX/UAYmfvqyrlC1
Bf3zzSZ+5Q3lLcjfgajBaIq0hahvBMNA66dqhulUKKst5ekiUtNyj2AqLykGr1Pi
qZztk4TZ8WhK+WYvlXmT6UJuepxT6B12fptADEZD2S/HRVsRfzD5VgOvqsLlUSam
ux3mwmtKHfleD1smMxTVihHztx+jeiQVF6BWbuzJbqcT/aVsRk1VfEOvHReeA1Yp
u9uWy02tUTkcoyHwiSrrXvBGtdFg3pbFFikdPbrkHKzFpFTMO+/hwa/NUxZ0RLpN
LwzqWNImbkbQwhqSamvsaZB54OyFtwmihp0LHuYcr2K92GVcEyqlNyKfktjgybNM
YDgmw50kPYcIPorq3aMko40LHBQMG79kMgmc/CwcHAuoTdJimmM6FToAx4MitOQN
XAo6MyU1nDpsyOsud9KR0utS5jl0L9WCqlUOWgmMdjiieasZIO/YhJlzKlop3oVE
lIVVCu/EOUbUktG4ZZLhidJZrc1lEMlj57719GKheZQysRQy63/M07wwyk4fLamU
IyPaoOSF/vZA5BnxP3wf+h8640F5de3qz7oZc2Ow1vEVLTzkFEHwnfR1dYX+2RBB
oljoRw+LO24z7eewiV0t4sy76SLVeiehw5OOLUsgdG/s1xKhPocLsKhWfwX17sx1
zF9WOVRCASjvUl3zfvRGLxdkdWrjZ8+SGjjV1tOdLCTkWEoeOZWwthlUNlYgSWYk
vlBCHd5BNoq+pty5UpkC97BEO5iMdjEr7x32Uwfrp4XpHWa7T+WGoBsCyCLtTtGC
xfNq9KxI02P/oomafxKPxQbvdg22TFb2V8bnzynq4Rnv/TiXhc/m1lEy/hg7y6pm
5JOThQ1bToYyYEuttonZOmk/EsaBsrxs+YcKqfXNwdwYZc6zmHrIBGczcEtoXO6H
nl7h7snMy1s4Nb9XfgmzZTd+EQG6df7EAq3bUPFDxim/lnmApBjqNO+/5LzQ3VGh
IOWIKIp8iQntb7h8jssqMG22qM7BuNXGezSrTFM/DRqy6cOjt5HKz8ksh7br5oJi
zEEyZcdpJgCA0qdgERkIZmJ+kt4DqcWBH1UJ/Gzh2VaMdwJSXfNqt0f5sR/4mhPU
ITcfiscFFadECtFHJddGMdF/lJVzZ/9cXr9escHJZ+7wfwhypNPrRGLLDPjELkeb
qVj6S1fMKFRT/tp4m/QE/W2uK60Lhr8asSWttEv8rF2V9IRM5Mqm60Glxc6GRlSx
ZdJVfkLmTaa8COLGInruYl+4fGPpdZxVNk809ygifFvvlpp+AaLYBlYKFBIvWD4C
KiiaY8/dlkXisJVC0xl6uRX3arGkYB2+/o6axIRR1LY6ltbEn9GOvB+6mpvadUhE
XALUtMn7G3Gm2xQAo2IAL3V2sA1gN9s6F+PTBUQ5dZHFD18tyD25ztmLCDis+28N
1VpyYwu0nPljNhZmE9oFMrKEPkxQEgA1MQhclB5YBvC9nX0/607WaZFO5CxMXX8t
66HfnpVBcRTDgIwrVMZc50XBP9eGI07jceU9wT1Q2Y9wU7Iw70rM1Z2lnqMhxlEP
0p0Kloy66+Lo+MsIa0+qz7lU/P/ydJo0tulMMmwlTcbUoqqXvNdjMrP8oDTbj8P6
HQlBghleOOnAvxgnETsvCcMnZuFGGB31Vr4/AGdONKa0jsKPUlPp/PjJvH3FcTnk
1K/iDyhdwIzN9OKH8T3YLxqfMxLWDZcUW2tQuWvWHsauGiex5Ju3Kz9Q5hRTjZgt
JFMrJJytr02YhxVqVx1uFFlY+TPBUeK8OmuQhDVUwwPlOzk1HQ9ZPR5uYBKfhvGO
wX+usCpSc+58E/GVXzlhy9zg+6b4oBuXkLeDR+40lEMClraZrCzGQow1rJqHlXgr
+YvVgSqdurWPCKEHe6THKBijpHquqyUyGd9ecjs1wg9P6srpVFIkEoBCSjDQ2uOI
ox3J115CTrJaWHw11dT8+RqtFOq1r8a6CAGFy7zaN8TQj36+V2OMa6ycw0+gnj44
FfXQvpqMlLq3d9A47QR3cvR40NRnfuJbLQ6Cx30rc8JDYdGiH/31WqVJepwNBWjz
AXBF/UTYHlTPHHUK6Q/TgsCbDCOOsA1YG7eDrUSPf6gMr08dqzw7sFfZ2wp+CfZP
vGvdzDRl/FwYBfFsMZyd9zFoQ2OF2vlJmubtg9mq5+MglGbBYYZ164JJxW5pEjtg
u4m8JWm3TK8hxeSdkbo4vMKNayLEuZucn09bmCwH690L8WvxW1I9EeExD9XKwu8y
sdu1yC96IMNhRMSHcjlPbQ60ZItbYgA13KvZjxMq8eWOz0VESv5Nja+7VYypuczv
zwxSm2NMwFqZnKJ6CIGA/lgtLssnEeTLyFLxB332ObhUgwSpih/C1CGkBC/WuDBN
8236VZZ6W1yPVYOjpKkcNJTOCy/f0cg48JiqiRA7s+PNtTCwfK6xJv8XWiqLkvQ7
7LT8E8nAlarGgWMADg+wvQnSeDrDtKqk2jJ0SoFjXQzgVBQAPgYJzKNrSNkA7dJN
GJ3RhYHoe15UYKD8cDgjudpLTJ2b59Zfl9a8X/Gl4v99Epdd3Ij5XrOJRk+Iq/0A
7wBTjmLkDPXjtKwPIVUkLNYL1Wtc9qWmN2YOG//nawIF+SHL0NVud1BGFlSq4Ksm
LtVjLlYktiBZt5JC8yo5TY5y1NdB4FofzndZPVRj/JUilBsVZaoAqQqpz6F0SWtX
JOTQrIuQKc6XQf4N7LM2Y2CG/pGoGPlSlhzH1ZKeORilSHG7JHp2cY6XsXUfGw9E
neJ3LcAV0JPYkF9fI7QPt3BLGc8TwgPOYCA1eiucYEciVcdD4mDTybGiospmG1AN
w4fZCKy1YeOrqRzgGurpwOnGa5CFQ9MZT8JtJnp9+IROkdFLLLMxERu1PR0xoDfF
SR1RGw+EziqTve/wORJiB+YJ68xjTJni/bX9+6S6LxB1qzhame4ldyLB1KGgJ6Zj
yyOA1QwcqM7PblCWYfYHkfX9kB5D6pUp5tv4q4thxsTRojkjHMPwf9D+barlXOYG
d35Abr3bwNwJ/5U5cSqaGAvyLhfpJobVxV7DEntm5uL0Ai4VEgzUOjgGqkMGtQgC
VVlk35bJh/N+a9fjlClqpa4eRUnMPT/6iq66/9K5i15igFpfTLhZ/kDhfI7BYc81
comVR8AWfzlhLJMcBSIqrRp1VuKWh2QuCZ77WcdIy2ND/slQs06wPYiN8hJ+NVhh
V0Nte8eufqe8t46nYwwPH+aCpUN4flXEY4U20MM7GyAPDx2ZmdnJK/t8Xxkp/JjH
KD6CA72x1/YRrBk61wPmdpFT4GJvOuvjE8I0CldKWBSrQGIWQ3wxzbh+I7pQ/xUu
PWrkRfP3rY/0K4M2U4SK6tLRHo/snOJEeRV9T+JkHKvbOxHC6qvutydtXdl672Lx
OLPoTxypTLb4FZVT0NEFl/cOqgtofb/xeMoMV4CtPj6euprUIqsXGU/wjS0HL8D5
9KlclD02EWF9F7A3B2irncyndYJlNtYty5d8P2KaRr4X4/260VrNbXMYBQvTbh/R
U7qMSb+/HMtrLPAjVRwzaJxA2jzRhTAyMwFrqyTI7SM8NTLtZqdvD3LpeGIOl/8G
sHAJyuAJnGoqHmGdH2Ah+gYsd78uUvPGIGLekgkcXZde3QL6sj1aaropOdZv9b2E
hc3JZmTicQFacH4R4eLS93dJDx8S33eHliEqhY4DXagwOOeLCPB9Je/2v84Hfl4a
2Vz204XWau/yyvddjhjxtkeZKs3ggbNKojS3ULjs6cswfyrSFT23UdOjU8ggtPr/
urZ4HgNPsGbxYx+VnTLXO3aRM0rQ1g4e81Y3iDvO+DAt107KmJQ+xstI9SJbJUcQ
mENwqXxwsDQ0oO4mYordgXHmewEX09XKYQVpPerORHiu5DotXcyZTIh6PLTOjYiA
72Ip566Kw13nsmm10ENw/jaJPDBV5OfeEPhB5vGYH4rCT0YhO5mwfMbaPkkdYRc+
ishkxcycMnmFb6eq4bfg1eeuqePa4z8ce3teVCfNpYZG2cX1GxEeNRlPXV7CBA5P
Mb22G4vKE2w2XpV3GLi8qjFTeFtUtXwVFl0kbmXlhjkXqb1ZqhpU/xBwyUvJ3BVb
xKXtUJno7XhXtsE9DRUrY2UP+xQp2ml1LEXcoyaXkxGuM6WcxHZ9ItNcydIarmOa
iutiqapsVGbRSl3xd6pyWiYbkVYjUl3+rLsM9Z2WjW3CG/D276tJppQrF7Ic7kZ5
5FNtEyt7tDrxtaFHCklVOEwwUbpv0Xk4/Yuw+MVvCegg/O3OGgmC+B77LQUc5Rlu
Qv4/8xV/IXmqLof1p9sMf6joWsfFCL3/SrcAHIxGzQiH8IoN+R4d7cB/o22wVVL/
aGGQwxKSkP+7nafPyIfIqgff6pIyC8PjrAVYkcGsPc1TmecxZAasI1PFK+RFI5XA
Xg7ENMTZBsnOjCdT7dCM8CcgxIvT0X8V1j28XSPUdiIjPm7Z8s5WxibLFZaPkcMY
wK+YGfl04sgzye5wN7ZwHOS6w4rIJFUK1NJiGOXw7E+gUhrKcS+uPyUyXjnzV7ZF
/j/u6DjaewG/gUfE0e6du2lPY5WrrB2h35/BI9BwvfobPQPOwyuHAzn3WMLytM7L
QVUQVXCAu5tt+E46gLeVhRsnhGCA1MKSHMHEQP9+3XZ++6Qp/LfW6RmlWhu8vx46
38W/PK/lXYR+7dpCrp0y1UIoj6XQzeJQCzvvHkSJDcKIzrr4HPxckvA4Lh+tCqGR
odgFI3stCHnGC8lnkPB/3JI77GKfiHZlW8TgZohR+YBj6OWUPNBE7Ae6xOztv9iY
8PGEE6cbR2E0Bl/T00iT+dSbIOjGG8ZE5X7TQO6StyDEo8DIgmMFXdYvstJbeZQo
BrPMmSb1o596lfBSnP6/gkndkb3AguSFM1Go0ohEoN88fzc/1ktn4SIoZb1XNCUr
ezFnkQwOatiYa2fIdRFHfpeA1HlKx32uXz0RSYTgwmFOreE83bzaa8hzUYY/Gazr
dFkz5bp8I4w/YdFlaRIL0Te37s0W/mCPgp9vvNKRWiKYayY5Lh2cd7sd+mLmojRc
hvuXsTACDzdfEdFBuJQZfiCHaEWazsnfmsjWn71yNBNWvokoo90c9lhydSMs7shD
hYERbgVeJgqMKk3hsEtgKk6HqjwoJpOblj7w6siYu2xKOi/A8GlhB/5mG7xSP2Kr
lNkdDqEhKvBHgjpG3gcCbHC9vfIBmgeoj5YkEaVomti3VkbM5IEfhOk2Ko0gB8IW
ocFL7DKGtVQxBM9tSeHnE4LxePwcuHWPQ0bITmosC10OAHNGIIpaQEhDkvkWYdoB
Sgbm5eEpA2d5R0H1MkWoJhw3lG8YS/DU8uyN1Hq8DmtEg2yuWMMXfbGTxHo/3Khv
X407sWPVbj+OdIfpMClye1n6Km/KWyKc/fMQM51AuUorGeyJKY7qI8xijgs2tLhs
L5dsWZwPDXFd9GzfZJRqQEcVLRoQmJWvq60hH/JWx1w/sjoAIrdP5EATLccpCdZV
cQNyrBtjLQdoIZeMb8OOSyMxPVI3jBJaU+yLBjp888OunpAfl54+ar6HFnk3IVhP
PAlQuZn0wf5NAONpQq38jE4281EhzZq24plAqQzi2u5BhXZJtX3hGjRj8V2Hsek7
waSTuM9qFLL1o2FoSNbTnVEC5UIIhy9kphRRqoJShe45bh5CKJkprEWXj5WbTIpB
ZgKxtdi2hOvG0yi7lWQMGNHzwg6Uc/RsgFkZAZOlnU3vBXacMcjfUwlgJHmZZJ9p
eE6iNRQrLqZenY5l/t5+3LBM7eB6AZT363lpoI4UTW0cbaYROLQjqj6hNX6FWJ1p
PxwF0rY26L5qLmEUAWGCu4joktoF3Zzbes+WZld58SKQX3rDZdD5IfeUkqeNb1oC
h+58AvxlW5NaoB5xLv0dhra19sdfOly7JxP3fNl62Cw5+uZfYYHkXw36eQ34fUl7
PgZqvn0P18UgXWKqftIsbp2HXnXH8iWo/SMrUZO8gzoVHVzJGPh28shlYyKZ6GPM
CVV1oV1SKRoOPnntwrsrqLL/8cZZhs59I/Cfx8Z861B8Sbpdgfb3EpfkJksMrQF7
gRYr824ceiHK5X0Yd9rZzBc8iCQZky38y2xmfqoofMmIFp4BHAHnSKEc9ZYdzAf9
5BpMOZiKhU0iKHu3VDzcRqKg+jaDxQBRgvDrU7MMx0swe/PSNYHvkn3FJwNPjg3i
8+BMiXQogL1abGkHqB8LXAmLnFN98ynfN7AsUwwnbOem4iZ7TNfmBOrmt6znfCtj
yFsjAGlQKWEDnvdK6C/gywqoUrYErvr3SdelpINjuCt/o+2XrPsumvVS58s+YLLs
ue6vanZh7ZlH1D/49WyP3poKRG4ucRLt/nXSwQ59It7hLi2eHuevEGG24NA0roXb
iTKUxW+E+ZBVpNOsjZ9dTXVJAT9M7qMlFrLUuEMgv3oiyFt2R75r3EGXQyRYJ1HV
U8WY/pXSD26qOIRcm6ht4+iWd29NA+fCeL7sx6sOpMklmhNxZwAVPD1Qkn6/9qRg
scAJCjQZgV3zZuRdZ9WcZSTOnQKGRXV/rrZ8BrsOJCLTKA37j+G2oa12G5FHjr9+
KBPFxtmG1TElP6mCI1Bi/jzPuComeIIVNeKQMcyvyQwZ0/OfXsMm6TFrbvRzknin
My8Dvd7/mUNo0Q17hEToQ6B2EzpoEy/EILyY+79V9SIlBc4D3GighsoPtNUrZIsv
csiFh1TQkuBeWcb9A8fFz1i1OPXTKvA8hG9sHA7PBy13gYdEEdWOcIyK6YA2W+32
iEruCY5pOsletxlgGcRvGSlyi+mMaitBSJFB3JQQHf2yxQwj9EtBWg7JTIigXPbm
JS/05HLsDiBboS33WAQIQnxfXrHJ8Hro1tS37FdqHlKW6XKsM1AUJwp3d/tfo7tt
YUJF38FguhjvfjDCuCdKh0gZ/Yerr6ovJFrwnDF8o0qGe/DzsAQ0j3tdLemLepbr
FSFgRKB86WAAXMcGwADfS5mphCWZMM+LVpj9IQXQT+iFYCWfhj7rh3Eg5rqzizIi
nV1Cevu7e2b1NPTJe9z/YGrjBV7Wsw0tCLtry6mt3Xmi61Hsf/1uT405ENriajKz
+iSOW1kWjiWwHBNL/3hXWg+0rqh1uh9arLFUbPf5q91lCbJH+3uPtzxi0iHkMF5Z
bz/czU91rybEe3CFuFG4/xQEyjKzrlCV/zlVLlJyFFwaNiDNulKt8fPZNp9zyE3H
hnBsoDLbbRQcGus7yBxgkrbHfZDCdmWwfcnxSPGvVCXOzxGhA7WfimUL6rtP6ZMG
YQpmCqZ414Y9WBulxJFIRfgAGV/fIyIoxQQl3xGAhaKj8Yt/8wA5aLxakx2Z+H/7
thH/iqVt3UvY7KRXj4r5e1CWnns7033GyYmO/0rlgLLCkmYwPv8E8Rde/Td7DHdb
Y+iXVJXhDK8TYchLMEDpSbWXQcwIpmD6UZlTSqMqCIWiWDlHoIQ5tViKLzIo+hBZ
lR9lAGqUaYHXSl1eBWd6WdDNx7zJ32igfYSIu0uLTfkaAyycOSyeE4EepQODHIhI
lfnMWroaUG3sfx71+u3T8F38LU6P7jY89DDSekI8DMJqiXxMwfZ2TlP/JApUMd6Q
G9yGHHk6mzh0UTg3MyzeWu1Bz5LiHczr7kZwW0Wdkawd6sv6Bbwbbh9zS/e5pwMT
yH5BGiTDVGOCO77fPPBhNNg0ST3x30/tGB0jiYK/wx5OzhAoGMMSnej86tb0AG5f
DcSpZTZJp8oO7MbGbUdUxsEnD5Wzm+kS2NLMCr91/jHxSrnr4A8tJgTPlsWLKaLb
X/EbAn+CFl7j+5MqQL4KAZT5Y5fE/cD0l2Fw7+se+whpubaFt6gC6JLhUZiNpToo
Vi05MXs7w8b0J/oRhH/mzpnQy7V0js6UziZI5D7WNWYhhEJv/YP3TY1Zm2tH6SRx
TYIiv2SzVUVxbwm8eN7C6nPd36XvO/CFTPYPrPOgZ3fRppyt09+pPKFLPHmbOdOq
pdkuVEKJ7iErp0oe5yiA4CPPrd0HRNyUm2HTASalhUb55qGhC9bIl4fLNOTufbYp
rNFsOLG9GO/R7w9E9JY+weLv1QHyp77Sv19OrGJQLPi1Utc+R1I5tOrivkuii5uh
iEWB3DzDN0jZvNVQ++G72EekaXsqO0G/5uIPX17/Oz/tp+G3Z6qnJFNNfFqnUHnf
+uHTk5qH3eBGIbgsJJtjsABq2vBvcqIG5+JsZHEHaQxv+EVwzE/W/mE8ut235mzo
dV5GEZArYZZxCpqiBpf/ZBeccYMMr4QXApOR8hr2yt+sdXrzNjm+9oAByCx/arkc
XsWDwIAmQmQsMQwi1iMZYy1LuQGuWglI3kFc+u7brzKHeXMcQITxOZ0lWSNXLfXq
aKUY0OusU4R+F/spruBLNCtfqQ6qyOxttM16RBqASrEA3g/k1yecJxtr1HmDdmOH
LVe8P78YI7219D6Uc/6S/Lp5KaPfF3OS2bGZEDAFHSji9BFzhdYQwTm1CWQzQz8P
UIW1a36aXFESNpTdJvTAeY32m9hwZYb3xry2u0/HG57QTDCPaxV6R2TwMifLTpkv
HuZ8/g+22LwbUM0zIvqT6HTkAgCpN+5+CCqPYVzVaPi/gJ5KeLmMHXuCEmC1W1FT
6Xv2a93WkEg88MbapFtH9l5KKlbC0mwExGwDZ0kvkd5uBc4NvvyNmDiIwu67CToY
gAXAvu2niQIDuB2+iSBoDRyh/CxNEHsi/kKrnqRaW4/Glemxt4T0T7+Bel5AHX8L
d367c30gYQAoIOLRBjCNcd2RWkwLkqdGqPruP9fsC5w7PTOI+79CxFb2BgCRiPFv
/CiOu5pOBWogZiEQm6JTUcmd6sfqEfOPp5T54cAioml24qFSm9QkHcALI8KrjAvY
3fipMCCqcW485FtVF3RNdAI54Bjr35Oq97I4Tjemx0HP+3v+mXtqTTl05ve69b1+
nLIpypk5mnB0VG4cHKyA4FPNdJu7yNppsk84wdnbEdbEqoCeENlNGbsB7Vki7c0X
/zMnwxtEBgtmypdmVl1K2S1V+QCS9xLM3kMIQGumOvuhPgvkmgcxjhb9z8whS+W0
0ULW6Y85XM9zVFWPWiDcifoeBj5MBAGMZNPTCDyqJwWivnoyaY1aJf3tYk4Pk6Fn
gyKeB/IN7H3r+f0UD2vlF4J4KwMxBjxUpVGkR+1fNtTbeUZ4j8cAZiWaMnMFFPG2
GbHS42Pvx05DS6m8A3b5UyHC8RELqIeWHNO67P8VYHWbJO4ZzisnvLTnYJD1nOVS
+OHgVkR1Y81lM8RtkPpp/xZvHyZP6UgpKhpSHP2snpIUPvTQiRA7xWhK4QPjZEZd
1Twclcp1ZBtO855091EZQ3Wf1iixg4GA9PvVQqslfwAnbOCYRFdQLeEzpdjY6plg
VFS1fJZnteC+3cai6BDu7svUK5j2djX+g4HdMtc4JR3CUq9hwNWBQ/VujjOrJhta
QZyV1L+jkNEQOhAd24aSJnxcMg6Ux4BCl52bndwVp/M0p7I498QjR67zXBB4pj3H
cnXI1vZKVJ7/IcJLQaHxChkty5nPzDCZMCC+Q4FDSf4IJhYHcV/QrybQi0JZdNw9
jjbuVbgvFGIr41Udprbp+DCKGMdF4T6hbKvcpfHTKJpvPlEUcuFODMx/W0B8uBcP
JjnU9L84UDPhzfijsz0obF2j9Nvp4lBkB5et/AcgpTYF6sayrZ6+jqWpNgtYq2kz
lUzUgm0wSVEJKhaGIKTGdmQzKgT3o+m8kZ8WNd9EeY8w8YVmuivOUjRXOWQlGce5
/+8I4PKAmEFnaSlqWKWyFpdw6QrTbsYXKSTIe8ORQW3j+0foneLYfobtA/GHgglf
+SIO5kAzASAqJ7jZ8LpLTY3aizlPLhukzMdWdDniG/P3FsFvCwDYbZc60VBOAmrj
R8SI/+0uiIoOfR2zyRbQ7jU5bvQ7WuggYqZJBRuZKNxyMCcOA81/hIMdPSHz/9sj
/DxUEXjOoHdCRv4cKHiT1uaBM4HMNTeaAHAIbMZeCIBRDGY4dshD3qpoo4ixIo/x
ohER16KyLutVkuGiqgQn5etcvInSm7Pt+C2BBh9uGsb4uI3Nj3UcOWFVi7ALbu0V
vFNkWaENULp/RuiCkAIyGXnAbeDrELaN+vsC9ku3WQGliDh+eIOuIZT9PmUaNnm7
gW+PXabh/aRwNYN502jc7g8gYwG2UMsrVh9CeddQ+l6mcF16sMnSLwYSUcOl22ur
2nhznr/pQc0k1BqgZvzCMz6xtsJkchYG+TXG8F001Kmacx0jEJKN7fy0pJE3H28W
p6PwWbgOSzzznyc0+Vpr03jRYhKgLqAPhTBncPcPWfoWOADANAsKqFL8S2G5lqD4
oSABOb9mVRuxSiw1qfX/xzhhY1M75vafW8LzpcFulqTqF/Qgl7ut3HXMJN3PPknh
rbdFLT2YRFMg0BYZznJfJ28L8EO/TsfJH4T/674fC2TR1PcouFYDgW7VsTkakSfK
hCUtrKi3+ZopbGnuH/KuCKUxV/JstTp/YGGCUEFuqbS5IVBFyaLnzwlCdEIzpONN
2KS3NEFRglMiFJeqS4W399ZaQHleSsgMTwWaAfptFndZTc7d+eQXh0gSmomPso7B
YlT6u3Aj+el2uCcurYjzj33KoldAf9uQv/1gq0/mC4gIg5H0wAyrN+4sfXAZee/I
4d+3AJ4kPcA7lKCWCbzCbxXWqOJ8CShQvTROHYqAUSfLn25v5CWcseRvxK4yDQNC
kcXRKuCFMsRaO51yv+c+WgqO76w7fxPSuFATcN8o8E1WrUTlQQGTuoAn1gEt6nRM
SR6xMW+z0K7MSnQ7UdRrsiT7u/A9afY2EkSeGm0g6vhHsBmY9rxMzv13yfrAJhcZ
hZCBBVVrZS+MaWVucAau3pj+4pY7sACWV/HksKCgnwzT8dIwCNjA5uaqVSJS1Agl

--pragma protect end_data_block
--pragma protect digest_block
FTc+D+M99Z5yuP6OO2602tkk22E=
--pragma protect end_digest_block
--pragma protect end_protected
