-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YaRW9o3lpTOFCeq+bhHElpmhGAsKq5SVbGE/eNcpKr4KvnNHM8Q+8L8jLmHI7PFd4pUpLcHpkD7G
N8M6NWDH5KAFwIjAnRzQwurO42xapjdpdTgEjA7k5rbmdbLet5VWVcJH54BtEHmGWpMV2e6k1QOP
XmOL+cAD1IJfYKJlMXqncH0/zOBk3IbLCbkTgbEf6WQzM2du2n+scsxLA3B6HLUCcmROMhIHI3qA
3c+10Lo7e3JevwLzFlP25vwCqEhFhER0o7lAw2//dRZXJjnY2lEQTnGF+Yq1LhJJ1KonSk3fFh5e
yThdWAAp+CmFXKUT4wE1YIEPDeA5pX5YOZxmUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24080)
`protect data_block
dr0FcWAsxBsIm15JQ12dXD/4T2WCZZqltDHqt7e9R4VWqH75VmU6sKoQS5L06eB8tJA44VvLaaue
CNBMgo0K/TEIG7oisros0NPU79CuuYvcWv1Q8CoEeiDccdynOmmVMa9FjHNkNfD6jDFAyuE73yIf
npNeZ1VNXoqXf1gpGWDOnHU85kVJDbYqvPOB9/94FkVymOL28Om13JijuPKa4+KzMuXtFOqwtMZK
PQp3NhyncfbcUHKVWwoMuQJx9zJndb9ZPKFV0WWaec5IAo5uzEWxLHB5BITKa8FA12iBdYtcUnAp
P3ht5kQZbA1gcddgZLqYgQI2nHTXYtOoehaleXGeiBlYRO6KoG1lBk604NjfYMyRYPAr6w7IIYz9
xbVOHJskRyRDSQfWRrTB8aI604ydoEJA47/iY6AUnkigaj/Tyl9ZKmt3L8dIWNb8HgrNSKgMbOBR
KaoxESbxace/ZLx9eUXQAeRlOIU9BbyQaaDK9MVNVKb1kIyJ8l8HKfxvKIFR/MsaPHBKtLeZmah4
TS91muEyT2nc9wqro2eK0B2hQXD2jhftzEqKRRpW7da51yJXUdHY70eZ0rtBV9uumusOEA9MYh1W
FMkntKnh+KgHwuydcGCLPydWws1HQHSDOVUa1DAVbmehkVHBsAi+tKbzlxYQhFumTFI75j0C1vYS
mqZdQ4G5ilJMMl8sdVNGriQTJbu9Om9MjIZOFrEm2RqZD9bJt2mHfgzDUkaVBt8L6kiJBv3QTCJ9
2HKfcl+X3+xxuipf2O6PIVu16O5S2+mZ/fDWLVzf6HR2398PrlMoh1etgs3XlmqAKPPVCM4OaXpM
dtPy2Idp1tnK2VQlMwFXpk81MgJVKIsuAgBbyd0ETgDrmcWh2z8AOKX9GTTQrRguagF+z1CreXVx
RTifkAaxYEoNCRaOSP3HPNlrsbWToroTqtY5e6YzIoSTLYkyTgieo5anLLGn7zJ4SHr/PErzRKQx
EKetYh0AGSXGyJmKRrsujJB/U80s2ooF4BrKnOwCsk/895aqTC9zxN74XSgY5LimNdFbG7QJV4+f
pvtiK41FDRSZSN/GRPOKHEc2imyY1/59/hO/C+7ACab31tNb1Cts2+IdlFaSxH0PDatS+z9+jziM
hJEsCc6tp5ygs40+DzBvHuitlNUJs/Y8p0GCFxmVp5P1PqHlAaRvSn2nvL0WG+RSJ8tdZVTB8Vlx
DGnD4k3INj7NI8m6kwH8d5vublndms0JieMwE+yuzhiU1bwEnWaxoKAv6KRIpeJtjzeytyfMiv98
Oug3dbob1Xd9xvOhBUZ3jBzvJsPfg3ddObTn0uCxOchN9F74Ofpi3rkdJuzN2Givw4Ni/OkpxBpS
rNXKeZpxhVpTUFXpx5MHzNClcOgSMx+XvkRrgHMdmlWQ1CaeUVk3ZyRkG06mXloqJqncETZwWkkE
g1n2kxa6IWMHZY41ZoShOe+Emgv5s0ApfF/Dv2C409KwmW8+mMy5SDhzeGaseZygankdKn7LMHNI
8YXQptfU1VwpuvXO1FVUNw3AbEc90SCP4ANa6Vdy/C1BWv4KS1WkwqMhrRxX72z6v0SX8kiUgEA/
3loXqWyAAQTb3X442d7BHe90qlyDAhTesbmYS4ciN/IS9NWgKYxF1BOqjCMmltpiV3k3j4GBVtwV
f8bPeM6R3z4GepLdgLZLzPLzK2nQ3LbDGTeSfINvrUnIFW+C+gNQ+us9xt/wlRAJ/vPIOWQU1sSn
z/P2MMcGtHAwJn6Uwks48wt+SG4QXzP5o+lpkU3E7wk2Jf1FgNytCc9iCg/55SIm62sDxA0FeM3t
/vCXa1+/QKVyS0TsdYWTz2AhMOrKq4roqljTcC0jv3nZbkHSGpIL99iyoaj46D+6bD1bhUG69Wzm
ZxgW6EYywqWc3AkfNh0s/H4mKFX2w+nGkP0WvyKbMMYL7XoOOP1kf80vdD+GUn96aaJF0Z7bY4JH
o7Ca7T4Ukuz/ZqIkM8cW1H5rdfxb7hWnUXu5RzrS8cR0DbIT2NnfxiZtrCTWN3WMEDM0tiZ3WQHR
lW0iFakBhOFL0llx5pSSJl2eZ8ckX2EplXcmINqkVqZ3uDaws3Nue30LpvGzmxGOEuyTDnyqslUY
8ZcqbjUzMPi/Jr5Qj9agDXV49swdNwMwsnEUyr5KN9k0ZTVbAEmBOk2YnfQOmWfxltk7h9SsHx2A
gBPNr66zuD4cbaDruruH4mKvGDx/9ej1GHFVnXi96KgP7voUXbUtwGkMFxTr0d5Vs1Bt6Y2jm+G0
Djo/PR5bZ5XScEtUoZCXeHgKj2uJI33axMfPTKRdxMHsGpfyFjTLOAbHKx9hHa+Y7kj6pUiMTL64
fS9+eRNa+FwpvI/N1awmG1HNRmgq/WPBoTvL3ibC4p7NIF69lkjPRehm8OtcxaRkDDFZo6WrGZfw
xEogLcIks7rdOobt5G+w7PhnfVYZHIeS+N7WDIqgjmLMa13pbjacCMCJk0Uni10FTiay81azfwpV
aqQQsFYc+CqrRql16frSzOyxbJ/DGdEpnyOuqHzvzkWE792dRzwaC9zdBsjZg5u4rtJ7VpeaIAco
f/sw/4p3idv2cI8xrAQyqvkQ0fzUaFTX+RfFjYB9GV06ABnfKIsHEGAVWYIxq/t7abymdkDKlm6A
Dz6568X81LMH7M4QuDYft/6fQvNG13tcDe9u0pLbpgchG1MkhAbHDRhPTdCQapqjLD6u43fvhSYP
v/I1EdJrXeTi6uPPh6gwHod5tlDkCnTm0s7vS6zlC16uflfNd6Abol+NcNduw8J5sUPAKn2cP7YL
ZlPVfNGnm+LaeAiJ/JqOGt8jwYg9/O5dDx5AXyqaVQyOF5qzq6sEepjZxH/Jc9eR3xwQ1xYD3uVn
nOjDKZXmKlC0WWpFcInMAADx8jIZyF2npYoaYdboQH4c5UxXiJS/rXUQhfx+yLnM93wQhEgz689p
id8riZaafLoMJmQisaL7glBBPHam5/ePKONc3hm72iazsFQ2UqLBwBIazrIS5FEqsPpWeM+4VRGa
5jXiCv8nuABJCCjmetz6jZFXjJLOSUrEXlhGJ3uw9HtYyDR/8XT80ZEpLJUawZcEaZ7lUgK4GE7C
NEnS3IQC7tn2WTrmbV5o3WNfgE2+tt7zOvELeo5NoYD0qxDjDKNiSMLDPd5tQCaos911q3T04xOn
quC32lc9R2bhl6s7RngQtrtf6/U494MzyAdMR9jC+MrBoDXZCnrx8rnJyOlnR4AsKZS8dsQGcqlb
Hlp6FrKshgJWLxLIjhgg5Xm4KUMhksqZOlo51NH/M7MWLwLXmJ2KhEn57bv/n6cnUirZB+/N9yhB
CdyBLwv4k14BSTVFRpfJTSQxvL+JnSIE8aDZ/Ssz+BhPZxwYH47uo/QX0Ahw9jl6HgzwTO917jqx
o0q9LFAY9kTOzgKTZurVmm7rjHOwbhkXm6SLA7cPWZZomZKnlJzB4Oh3EE9MOZKHcSWeLLJaquRK
Zz40et4lenQtjMVYjZSo8iBDcOp+/CVBJ2iLdPMtrA9U21gTyH8nUQ94vLX2YXNZXqgE56oPtcxZ
NXzWvE0//5hctJzvGGnt2jy58NOu0UZS5R3k42YDuMFuhjLuNdYQ/PWENNoqsnhZOWOn6dq++lAe
qg8cFJKj2XT6usV4RYLxcfAol0ew2eqDjHLBCMQ8vDPIcoewZ9wwI4Vr54fjxm3rGexkaI2OK0TM
O0i9IQ0HwK36ip83g7DtpYaubEmQBZHXkKMD48pwQP4c+B3m357kg2D2XZFJLbVgIgqivAGB7k9u
bU/QQLnDDaV9y5FgCnKVTPkt6L2w2Hty2ZsLVFdwPRyimabQl10aq/FlVbDgK/h8EjbckhCPHiKu
b7dJGVIYtG/FpzOed9m+sxicSG1x09g039bAicTar763utg0RIlOVnKRCeiyspOiphRbJxbube9v
v+iHHoi2GurLA2ajDZgLqzcBeb+657r55Jp7Mg5oWsL+IoTH5+kFqpBvOBBYntrcJlDElq9QFsYP
2chin68yVK7q176q5uIZmIVyBXMynmOl3ZmK3/uWdnJxerbskDwUbLnyHmRq7OxIrd9HUZoyV3ck
iOsp9d3jG2Dv4OlNnFAaEukZApuKh4O2FhEDR1yZ11hu6MkdSlIqzpVI+H7+TferfKR6l+5ewXrE
iv1ACDAQx8WsE2P5x21eIxcKRhQJsADGsN2wrmV7FXNYcB7al6M+4GsM+urGTpR8xk1fzsdwzl73
jnn45weiHhoN85Rx/RedBLBmmgwfJv6w6SKRuTP+wABPTP0iMuEwYZYFaXczV7GFBs3Z1G7X6yZe
0DgPEWDWJR/SNG6BVn8NjiM10JbsC6KyRb8IgmZXps/LW/+O9JIHntHcqi0MrUtvW8BBafd7Gzk/
n+v836YQoWBUSS70UolES1hwD/EPOMcTikNQ/DhAHYnH5DzT+zuynQQimOoQ5lgzvYVQ4YnwGdR7
F80WMh9OIQYw8NcsEzM5SR68ddkdjhSPErpYZtErw2tXomVcnThr/bcI+xIRwUW8bQyz8MRcSQOp
i3U/8aVhtJJc8rhu0n6HeDE8XKKAVdHqD6jzNK4bm7RXGMkcJJ9bs0dEIp2UTrJ3CN6TZVSH4Duc
TLzVmsv5zwNhFL/pI8Dx3MZzNEcq+dHtOzlNGqNJ255koRCx+AFfnUHMDO04gtIKQkO6sHO1j8v+
/cBJAWUWBilbZH8tqjzStHG8zwic0XuiM+vIEqnYEubhYFr26oEFR2nO/qLSsCSpqX7G7+hGpIGr
pA1eE7pvZBT8NVVXBtjsbdmuld/hUfbp3GZFjzjWmhhD5Ipw4iSL/ZBodUdTIrI14Hgh7D00D5wx
LZzDvgPipPZ12ojeOzY6otq/L5mJZb06jS+am7FwZFbKt6evWeijwkRhm1mtyq18jBD2X4bcedDi
RRgHYj6rsSkrbnBStCcYZzFPChtqBhBSGz8xav8qX9MVe5ffXg05xapTfzNtmjSC5aorQ/2EXTEX
FMQEk+UbRidQA0S7hoDiNBe3MIjhEjjnal2T5y6QJMYARi0KFVorCE0G61/ljcZw85nYFy2rqKVX
xALE268jlicTmAKOCsfFZStoJK//OnBijffcjcNi9cmI6GB2UOcf+u8+17jRcrx/kEVj6po6UrJW
DbCaTM3xPWTxe+452ARr3CxrSX32ZP41UA12KFtVEJK5a9oZIM5Lubfjvsww+zicv8Gh9octNQ/g
HpR/64YQwhOO7kK88Ld5hDW6yd7oXvIDL0ax/k4srfQyt6R7JhH5/PH8iTsS4OeDToHjpH/YUGTj
C5z5qUwZylWueYW11vi7bIyOpyY/NvyDJ1eDcV02gQK9xVosgwUGO2tgqa5PpPEC7s25zdPvlVLa
7hSGNAwvvUko8OZ6f+uLLGDH2PYnjSqG4GEN7rjS/ht3yNYZHopGTVpPwM6nTZdrFtEjRSIpsI1o
Y67NHvhWrPdpA7cl7xxuxXsoSBiskJGx56S3rs9ziyKPqh90U5a4eP2eOs8ELcYwslhaAGT7CsvL
xiqDOxrGRkoNFCp5GSI/QdzGZOW9gAHTY15cQ3IvOAhDF9QeUzqCWrDCUJx4/1ETSo5G3P/4IkJV
mTt75bPhPflRxwj8wfZ7O0U5jTwjeYodRTCEGPxk5J48KsgwS5xLQ5BQCYL7aSk7SHXdiQbfEEkP
X7gp/BtYdejBVrOg+w7PIHO5PwEb8/iY8qo0WIAP5xCjhkNWqGBf8mam9afggPOJMDUZzaYaRzJt
GIvTva9VhQODgLptwho0EPvi2yhRrXA488uej6aFS3mxjAk9Ya8vOy9S0MHJ3rxFvSoooGz6KGVH
h/H5vBQDb8myiN7nfIYVMtdZODgAIkkfbFWm3xGCDA8JfI7V4I5QBucypRNx0FbLuZ9RjAW9HFPC
aRwBqGuLR7BYESOop/Vbkl46f8sA9hrJ0+n/hxXf/ZlyMid+WiiEKCpbgxYwkbY8bYbYb5sGEQJ4
Pe61ExUbsqX+emJo1ZoaJdgtYWqpE2qgmI1iBt4mbqNrOv8ovxF9QcyPJHAAi3K8kXHp0Q2k73iW
/ALGeui6xV2njHbo1HQyxlYImypytGummuT2CQ7AidwYAxr7UMViddPlnA2RVpJBv5IuEanUComZ
zIIoDdRfQw8yytd6t+9Wc0fAgAeNfUvwHP9VwWOeroXn295H+FJXjf5OSEHhWJlR++bGdeHqHWtg
yw7fSCo3ZEikwG5eMRK0NHPsnOEsBCSMjX1m3C8zsaAbqr/FvaeVtOITHtioBbl+fiyvcTkHWnO7
fSTwriVsXr3tXxVagxA+UZvuOOdX2zI+hRSzhnBs+sGh4ZeCLJ7aviFpWwrPE4op+76QSNEiVwdC
/CywntZLUS0ulkofvoTWRB/kDUzKCxPCeXfJRlIBNbOQl83n1IFxy1zODESBElfCtwlfQPt/3SHa
HLdacyLfOwDJXragOoS4jU8pbyWboBdUKZ24m56+EaPAQrdDgpu5lJfIYRUI9ckb6ABwwNdpEubk
AyXPjlhgo2EnI2xsR7UbtfctE9phiY7o+7jLow4Yz79ECTSUlfIuFk8eNN9i+cnqRYtnFscU5iEu
EPrGlcxJvkhnJ5Oyh3+/LV5FxVh7FbVZ7U1YkLrS/AAhAY0kyZlf5K4gPV1CiNp5Ope1P0fJu0Jy
uCPDJ9GKs4+ga/trSYMbj511YRw+8A/rCmEoWqMX9ewzwhU9AOrZ40rB0Mf6xSscIuYVKKgqxFQ3
4q46hevwusGco7D5T+UkPjtVePY1f/m4WQF77vs0CRwU/KEcGGjf/w4I9JQZ4ufIvNb/55a2oX/v
uhzf9QlNzhHlLKoBNEsWaMsn7FVPxkdHXR9n1JBvDN4Elmx8oxDJcADKEld3rXAXDC5gknnMEAAJ
OfA5nVk319LtMW3ZJEgz2oqRLgLapyNvML/XeTKXWU9DkmM1i8GKb3qrCoyH4Zf1254Na0AUJ+QX
FzD+TGDaU3IwvcOjemvcxg6MPwsAAAzpFdu891/K65RLpC/0nFn/LcUinxRdLfEVR9h6qeOfhe2P
630Xe5dVUvayacCSEZzb++LeyRVhxgKetHc9pU1h8iDg9ZHpugnDP++W7OIuscZ5pfBTQI4yNSTB
78lPrJG+byOcHRVNk73v9J9YDiWkz7GQtN4+WM2fxiYcRV4MmDxMDNWhlDPXB9w7BNhW9dtqyT41
xbWQWzu8RAC0KlUlFqziwc8CtLkLURFqk2jZQ97BQfIWu6loFtchNmwJHhr2VKgJzJ+Ip7y2+6Sp
J9/FXcqAICV+2cobRLWm3FVi4tPYe0VfR+tP2hKhc0ekJemau3mTNFhtTxEIa7Zcfp+ymuepdC0F
TNNpY4lWl5GrcH1OLr+rb5Dl6vi+uGCeY5IWmJ48CJaAn/AoOshxNp4jh5YFrSfXM0ALY5tX9UhG
QdRJTRrZD6BvOYSQ7eKwImVdXzEkLkJJ4Hvp4aq+yqiB7pm8gUSXDTRbxHzXGN9OUL/otw5CCR95
ZNRebWD9uCZ4Scrdjg5+VEmG2w9Lc3bqLOcM6hxYCzgHX12NY2jqBqxzy9OGaIC+GwV3PPOcdbIr
4xbGzVn3As6a5EMWZi94GqIjG+vQ8vLS4cBoyNE4CPtR8PUAHnug5Dosd5HiZoShuRxUxdJaXLYr
gEgBa4CSjKQOsBPkVC6v8+ZFL35/ciolhwoPSL0pomjoLBLV8RJ5AsZo5HasB0KZlXPz+K66RN6p
HZqTGdfNZmqjTsp/KNguXHi9nbUalOey9q4azHyzCM2WEoA+ZHIeN7TsdNHxuOp8TXO+5BYIOp17
CZ0UhKFDwi+vGLgylDHbis7X+PN5A9p1MwFy4y0TZMvnU4mr4T4+2U3QTGrWRA2pE96IpjCYn3/a
Ndk2WLbUkjsnl+m9net0gMnA+F6NrArTkkvoRTZKOLvKJmZbs2/yk6nPD3k3GI4uW1YkACLy7beM
ZqdXf2IG4iBapzx1/4k/N3B/mmVLnekbwhSF23GLqyczwdYrE56p1Q2JYEBOxIGqYn6d2pf2g0E3
ck4NE21GuMK5jMjLUFZ3OD0FGbe53Z6WqeMMbtgNqKWVc5AcKUEJjgxtteX/uAYAPvZ8EhbTY11I
oBD8mPE2wT+9hwCif49v74Ip4AX6EICQAOaUCVOCkGwK1Q/ywELatg4WCj34eXz+PqIHd2iOQdqX
eB2ahtxsbPito5yvoBsf674flsgZrl7u63ySIR4TgmlW9zG0ZGYQJsyAu+YzJsHty1a+NyXzCXfh
d2qhaDb24BJe1TRspS2MUYjxyqrYXk7tTM53VfK0Z4p1GNwba3dR732ma2McqwGInuk/CbVUBze4
ynp9UbrXNGnWqG803pvI0eSxXQqI0kRqdURiWm3/gYQpFqqaWeuIcqs9deFmhYjTI8QAVZHkSX6K
GkQT/pZDr9pO5s5WDa7oHgorG/kucVf2D4h1qjVQ0G5RMt2IOLhJiGNWXn94iKZ7TP8oriYKPUAW
6LD309OLyXf65hfsxS286i3n2OotGfxiYSOe2BFDRZina6aY5NGAewkqDyf2uIJr4bOZMxmxAAUo
CINtTRl5MIs0Nq7CUMcYpx2FtU5yRtLB39rOuzKDzM2XpdD0Lc3fDasXANJaFhNG1BYAO8PCb+aZ
CvhAJcwa7waCV+XvzSvYzJP2bQ2jTSb5R8rbrBfrxTlhNMuETSBbbWf78gfq+e/bjALHQzGSQC1g
nGFjb2bn19DiOSkYGRuHvf0xKmTwC4vafWgk+T+qZPC/BSqgv3J3/1Y2E043JiRCo3sViOlnqlBm
RDNndhYXzK2v45Pyur1XYW75LADLhrePfmrvKqHkS3brr3xRyVCSYQUZcQc9gRHCI2Ng3+9ay1KG
GeLH9dzfER1gWgiu9tH6JCb+Lru7458ETQaMkpWobBV+yffQ2npf47e1GEjW51GCjhSEzirdmTmA
kWAqJnzcJkN11k20jAPP2aOPB+e7ldu66IPOpu1T9CV8FSlKzQfPJL02/VryXepi2/xWy1R2e6fY
Tm0guAZP3qqMZSxKOQQyCGNf4DtrczivpzqQkFbj/9PUlNl3luMiloa/5tYUacxglF1Ssz9Cl/wx
CI8zTUO4g+kMYIQPTHZbIA7HnLyT/L2eUm6iiqSxzOw4hzROenRbRsBs3Ov6++V5Df2ZowVkdCQM
1LWRr/Nw73d7D3rlWgh8SysHobFQh7PhV6Y1aoR3mDwaL6DzdtL5A+Y0HxOO6SXuXNjt/0y0j5CC
kjFcX8cfcPNNIel8WBA2J8TWfL/MWQRx2bpCcB/9Ky0/nP+kj5V4G2O19njgu+pPb52GUB6ocwqR
0BS9USTGTZe0CqBDBnd/XdHKLLHxJbGob5mKcY2eFC3VlzGxPrX/jxrujv7H3uGuvqiKbR3rpakO
F38kxmVT7njKiLs4m3T6tf1Lg7ywX+B1TMqq51cMGXefS3f14FtVcfkw3CijnoLOPVXzIaEY7Rai
N6xiTuoaNXU+N9skwlaob1UqRGCZA3/qICOYbNkABIxah0b/LluMwSwI2oK9MXnF4gjvjHOkDkr2
+bTOT8OeGciOAu3+kFSZfBkco+vRnOPO6L+SmUysJh5iVE1Gi1vwcoe41PPgBMeEe8jTMMAEVJO3
tftSBEh9OrHs/W5f6mIrU+SvlNayjO+mjRcXaADExFTS8WrbNXgttQI2QprFHA3hcGHLqBzeAm7q
cvMAO7mAOby8f/2gOoQAbnwXimwxY8hQJSShhhTso/YBhXgx2/rAIEAuH0Fb+ZUE8C+EJ2y1CyRM
cX0BhaKoDSB0WSLSHiJUqINdd9QlEN+gk7H8Y5w2f8CQk9UEF7B/JGfRXSJ4SFxvtXZ9Q6sPnpsQ
bH+CDHIwGvcUhqxUMqGOnG8WP47ehophqwm6Zi43M1QK+s4TQqi4ulTKHT0IXCx16cvXJag+ZHDW
PYEqOm4lReEytYpfzlj9haoZ+ah2GJdTE3E65+nNJ7PyTpAz5PsS4YzY57ghuWwtQV2W/PUwZlhj
QZjx9VObLtCVXNTR3im4gRPH2NX2ltBVPft/Eaqsi83zEsw9xHecAzbDrlK9RksE4zvzdEUShHEA
kBXQsfr3W/aEx8mp4OkRDjeAXgg5nXM5ZiLx/AFgrPbCo6fDx0/cusyf/hutYtLS9NZnH56zNevQ
zx398qXXyoVXbHQECsT0iYiM+7cfmt+2WVaVXblUwmMZqehbUSiGD0SBrWW1lihPtHmi10Cj7zDq
ClPxUxiy/bkuUaD/A1noft4Vm843snUmf1fLIvDePd7vkhhd6DdCQQV1ezoVIT7skA7iu8NgPFF1
7lz6viewGs44tUOZCxWDl+4mILonXGEWD4Nergh1vuPBPkMNzCdJom0FcNV0Lu0BRdimsG98xn/9
5uSYYZZmLjYBvzPr0GS8gVCK19SOySSEImuuoD1lYtO/wskc3QxFOF/rzqWxHrqKEVdX6rOgyJoh
jGrO6eTrrgJhKMehYdk6h0x+R6+4MetX884+naEsMjgaBV4aOz+IUuP84HIDoYNFSsicenlgYgJz
pFdX0RUqCpNgJKOU6EqjX7kNcKGQHH+CzKMVmrM25d6Nw47YyFqScDAlgmDnaGxS/Um5Ly3t0iWK
GB0Q5cmphhy0CzsCqnvSgxoROpzZIY97mn7umDHIGllUbZt9BBu07PhSKaIUzMdcj4MGz3Vk9QtQ
F8hZSy3kcO/4QLE3RzZAxM/s5iZmtrEGcsB5lyQivstHkrHFPJsEtX1nAwwxQKMvr9DjCXIpixzO
CEojBsZwMyOLp1Ta1aXU+VFAzdCfYdQ8VFDacp6kRrgmBvCOSUlqoxNzMCAKE3wqxczVE4WiXKl2
js9MpDuZwO3/lJFcsChANpGwz3bezBGBfVHkG+8dogfWz/ADMOgPxxr9UKBrpAE5KBaQTjJYEv1C
t8XWvmMCN/xz65LFnuY7vrERBzlMzdBwbLBmyhNEStYu+LPecMZZ7FwhVnDL7QF7vI13UzxEiSeU
FfOx/m9nLSHvns0pP1AW5+0/AEhLasrAVsEI9iBWKy/qBO9K72lyQXMhwufQCkQkKKSG3PEzwtew
Mr0QWh5LFx1PbyBFt2lreuupDB62qO7ElgLgIYMo52BZ8l4h2Kmnxh5kpuyyQOrKH6NfTq1Qw7B1
c29v5fghoG2XXB2Ck925cnxrDwbJSLXQOtY40VZUvxsnlAq6nPfE+c+AeVWIeg2sbIxL2q7YriR5
xigL9DP4PwDRxWy5XxCmfUxm2gP2ikOS6Rcu6MKNFlV3hm2Xsbt6PiNOgjB2GL3ESiPNNf9mq69a
/MyvvHlY6br6poN8D97jVuOKN0DjGDsUzupSMx0sYEJMwg3bLrbBPpMiovKcOuJNxSvqgou/BuSv
Y9GcYEush6AQyK+a/X3zhGWCMedg4TW3fLgeus4BC/6NL1XxuzWzEmm8/YKi7iCeDNetlxHlzxNS
T/eufrKZ7dFVdaf3vQbu1mQRV9Rd6aKxnezLZpy9kVBnhmTL9r6bPVaIto/Nxl1A068PU2tbiCmS
fp8yLWepOI61fgDBjIpfR5Y3CbHTKI8aGIYygUtCjI5X77uyxQOVyuhRSdk+gsKadjiKF4vhYYv/
HAOG4epzY6C7r+vkl3ilRXuGTkWy3fbxYeB+B/mVpJr2kg+Xd5lLWZxBYCXdeZqRD3oVYJCIvIHo
liu6d/pFQ5tMwPpzMycvNDCPSdWxCMxtHVEEsggYXSsxsF6g9V0xS4bWO3glK5qRqgkXub/v01ME
OlBV5PBb+Or93/PC5YngRYHU/gDUUo2leTb8t+thgSkDlep6ZFlUdf6DDL1CutmdTFLkyUwf923O
vOv9rn6/vW6FQ9o1epFYryQUlAh5Aj+cWOG8DB54rtxmtOuEn2Zxlr84SrRTx2+GaaxdLL2GVv9i
qE6dhGNiRK3h03vEdQk3oN4/k6G5IACtpf+huD8/R+ojrMHDB484eOPyLIgjg303c4/q5tKMowEh
u/AXmLvSLYjUoqz8W9tAMxKZBPhMDbUScNW56DzPLzRR7ffiw6eCEvhVDYev3xzljnwqlh5tWOxi
k3MwhniXg171AZaA6Elpx6HrHCDmwY6ivs+yjp5uakOjdwNGMxCkrqjZrgovw1rskDwt8gW2UCJk
N4Uk8sSiZxRl/hFiT0p7AToP1qKCg9OZTa/TPTuXaZYGHXwckRZLzJXneV8tPM5Mi+vHTVH0/DSd
H7tdP16bhUNrzY9F3hx8jDjeej9dQIUp1XkM1RsFSlY1aUj64AsX+3kpMK5Oji1g3qGltxr49aAm
9PrWokpe9jp462AsIB7BnZQYOVti9UJy0x6Q8N7pBrhd5RhLqZ4bYhmG88c6ScgVj9Ak11unm40q
I7O7LDEZ58F5PwL8z0Yff/4ScvLHg9xzFHxbF9CzMyc3bsyu7VchhxJZXCS2P4z28Ptlbx1qnZXf
k6uCJiJzgJ6KpcVto6yyHAcZk8UIwOW7Gw6f54QHQVpcr5r3vDwPO1pujzWct64PGERrfr9RcRfS
AnEofa96cFbMYUgRIPLIQAq5W8fDuq4/lfCu4UdxVwc79BCmVp1O/L/YbXjxoOjegz8zGFgTMnRO
yXfDfHHNetLWk6QLanFgj5KSveJf7R1hvuSVv52JHVrHPaJzxlWDVtzpXWQD7FxzcCTCEfQfcggh
hk1iA+W6rG8qLrR92fCpJdrFsLjD+FYacqUuPdIfOTrbYt2YCG1kKkseQ1ty5mUkWQ/HzJzLOMGw
+sNZ9wK8J2KuK/YtPxunN0mfpUMtb6/ym2Yts9gx5vt4+AdKSne6Zlpeu6ameYKM+0YGoU6MD5kt
FvsnSwpIkJoiUBwB1iYC90B1aQ+mPp9eDdDB2CLbHmsz/Qo5b2uiMp4ta8DSEGuXmeJ+g5QZi6WC
FRSJKhQ7W5eiTFf0+eQiCIz+RvblZxBmV9tzl6HJOZBCa+IVRfdd0hQz/tmisX4x2zXoNgL4FmtI
7qaNCT0VMY9TsGfnlFluXOyWL2TQcQGRZIgt0dUlZvPA72wJWQfSfj6b5qAK/eBS4csKdrXWj6Ln
1cs6Wz/PIIh179iZdTCmmj5C7n9ywY7A04Te3GjB6D2bzSMPnMpwuiUbtUWDS522xzjhED7tzhvM
/tMkLCF/MKsPqvymsa4kvak4A/vGxCoYx3nLW/sviZgQgJaHOJ1BH89iqxrtkfrkPwATLq1yeIiW
vPLNN0P67yI5S7O3po4wMtrg6kErlpGpeYIpEbeo2vU7/uP9CGDkDaIuTnreEZ+gA6YeqRZ+X9d8
yAUk3oOQI125nwnDp/vm3DCoxy3S7HOvyBaazi0CPH1j6zWEmBjTzRK8KYZ/LYZKwFbspNRt8ZOH
oWSOvkjtr9joKciZyTubqiyJr6ogKq0asx2gAk5co7ZSAplziJVAji8qSFUYuQB3Lr2auIsy1CrO
gKRLsBSKxxotG23OwPdFTXS+jhxaWzFDFHbzkkcqGWiqPxw3fGLkQMzYJMnaodZ6OD7eGTGzbeTu
OmHa4LBWAUsNZLPrAaoxN723QqnuaYqvoGxje22RzrfG6gpwihYR6OVgmEzZkcfVyqRaCXjLsAC+
1UY3agRC5HdVCTohuUbe7CpTBM57zLq+6GMtX7Tm5orNfD9H7aVo1t4weWV6PBDVieQ0jKrJr2cj
t5q10iTW04CXUPDwSIkflrGS5WINgaOWJntD4mmWffdH79g5Wy7Z1p751q2R9kdIUEA7dUiZd0ZK
E0xNGWbqMZqRvGkW9APlW7WLW2IJIJKR+tsw0PjUXc2PrFdU/apXADUdhUFIiGFPCCgL3Pommq0y
MDRlCLsE8lkVC28tidvzbtuflq0XN3lfrYExUlByUyynDVssrjHUHAacBXqKPHTDlBP2kDRYbxWr
9wgGEmRsAOaKBYWJK+PUOVvFJB/BSBJOv/8KVKIn5eV7GI4xUSkOj5U4rLSR+dR8QsDIKbY+UdOJ
MMdlLjNw11rl7qaoCH5rXY7qtQQN4WCVJ1b/fKDh/y0qaNLCCJtO3QgTD4dp43hadDrHsRVTTBYu
ypjy/ehCkV8Ozxukl61nX4xsSdJ2acZqTx06F3TCtuN9Yf/u3wyitc/sdvZylBm0UFaXtFl8oxzo
mi1pN9f47SN3cKM/a7aBVEaY/Ewi63LdKbJgEA8RL5GxmWkhQgGosw/GKTFw9y+AoyZrt1ZQes4l
ytOqg5z25zNPtbC8eyKhdRGVuyXR2CcoC5QSKd+E0aUTqOjZzQ5+MsAyIZzwMStSIGbdv5rK5ZLe
kk0cVpHY1jGBsu4+ynD3QCgt0R+NCqLZh8tQY+Rwee8u9ZcxE/jEBCkMV4eMm45PpRsCDN5WoarM
J+dVCDzhociSlJW3iYlJjwPHAsEM30upk6t0JQuAGWTlbq1WPu+Xb+LLHVdICRGxOL45V1kfAW3i
iI2c7uA3VVaEmlLOYwZJDf/wr/oPP48RCGlpYkARu22c73eRT1sZ+ZcAM+7MZuadpY45GP9Qk53o
4rev/EtwwnEX5qgAlL5/zbG5bbPooQ4YlQDBz0h1yjt28CeBHudjYBj/Z/a4mBVYXcRpErcEtmaX
SQvcKKuMCh8Xx9cBwo8btGhoy5N4J8I/tgWkTFLnTv99l32c1M3mr9OqklwletGpdSz3R3qenLM7
i6QTpuKSbN9r3feRcQFY+yMO0daliYjdEFb7MNTWel+QwhEdTausnLvzmG0dHZaM+V5MS6BFG4UZ
7MF4GZk0KA0UEqHr7oQSseilET82uzfQFjBOXI1fhfDcg86PTaOAo0Foh8SOEwdMoocXItVt2akk
AFdRKmlHHG9ZvVDagZS1nTeaTLowUqHieHG/KOztFXzScbxkEZlYdylMAcFGbm/aCMKgV3lKyxhP
nrU0w9PPJ+m1mub0UFol1O7K+9MJrt4LQqa0Afi4GDQwktJmZzznClZN91oirHmJ7HYZmMLypk2I
0rqYy1UCCGW7GblkHkykd48qfgNy4yAicJ1UMkQxASbjx+sVu34Ntfiy4SAw85ekZ8WJ6ZWkVCPn
0yBwLpe6DvuOJC/bdhYWL/O1FEYfMP69PSkTgMGVPZ54i4zsl6Uh7xwFXapaCvbLnYoZfSOTEc2X
GXAVTlVxO2bEJVlyt68AptcoMPdJmCNzfyGW5gnUzx38MLOAcVkkIKA5RHPg/R9MnMgWkplXORvK
kjGOb/ix6pFDcv2P3vBMyfin9lsZZWY0kenpXuYB/shgdM1+00HTJkGarvTPyp4AlJvvqV4LtZWw
+NAYDsCggu0ydlZ76GOxaCOVT0O7tX5Y7lrrfx53Yn5e7gVoZkviEJK325Tz87EfoyXNBrgb4BL4
zsnG5C+KkIu/XU/8mi4iw83d12dO7ilrD1Z/7pJ1+O6f1BwVGdTlOZDw3TnzDwV/AumS97Ewj8FV
gowLn5BeZ/Lr1YklZgJHaZMgrN16PfKsCI7Cwx7rPgXS4yyW794p3A46U4dQfBndQ3Xrw7RDnusv
cdRSFFG2x/7LYROLVwm0k3XMoZbmkKCmdmLidsJVJS74+ypyh21nAaENCK084my3hvtTbT9lBN1A
/KxTuMzSpKDAnaoKgWvrz30kgABs1U69mYq59cAeTsOgDRS9XwXw4LPFDBUqvfx8DojREM+/ppW3
Q5fzV5hDRBIhSubPFTEvE/kfiriuMezMAXaHPhdMYD5bEegUcY00+HeghzeFrlVACtbdk1qdWkig
il5LKQlAgC+DsvpycauTyke7QNeQOglX6ByFJ0kbiIG8irvakqZ61Ktf/Brqh+8zenF3Lx3DcWDd
/nLysQjBA3wTachChsG7irH5JZPCD7UGxFUqNc51ZV1fG5dDzAxKEflXIiwxTL+SoNM9vmKsUyl4
Z6hca0228xtwtCLsklMgKmCtHQxrJKOa8uvLnw0N8wdvPmtQerHkK6EXwLcxnwuSrt5kaHlN0zH4
vBL9EaLZ/q+UjU3lTriJE8LvlIUJlTzh0OH7TPskFZGzNAEkQtl5Q90rDOiOctKiGglflaBJYb5U
dYCEJsZbqXMtIBzxrLE8wFNRvAWU9imQors2EWnzmC33/WNYJt5f+I/BHpi6UVqLMMSDFYeULSDn
QH6drDt8gXgOjnrOTXjKbevd7s3tb8u6lBAGTS0rYfPUCumeB+V7uVfxEebcY13iXlF6zVnZYMMu
etZRkMWihd6uZvDvLvktV2ihce2+/9WQroawE2PUrRKdeMavKok5ky7PBi2PXi2TaYpk5yVNn0cQ
j6b38PHdCTkKv+GZyXCCAOOXTKzU1+cN8lQaX/lUUJz+twuOSA2DoG7cMeMfPfPj4xbyPy6LhAFl
hjeroyxtcYM0HGJux1OMCMTEZAOVfb+liHPtS0dToNnAJ/dnXrzE1CbKKm6qTTBUdJTxfFEv2HlV
jXChVezOpL1IStOuAbg/QdjJtoJgB5YYiKDLqCE1QrGEOrK4KSApPBPcd8HnF6B6qIIvABI3PCLc
pbEij5CxMbKcIN4ALKCCr0atoTapFBGV3AwYZBJC220mz1+OIc1r4Hg/UazLrIE9O3fxJZDWiUNa
x7YAaabNTQa0ToiPws0Iw/9TVxYYadTOOAIwBsQUCLPyVVx7lKH/e9tRc1ADdRTnlB0AT6kcnYFz
2dhA+nMTtYZTJN++mKqM+1ESKThgXZXbilP/4MP4QDvran49E70ISWBfGB/EkIYR0CHeuLG/92ll
Pk+TJ/4CX52oB2yGExhtg80MGKC0N8Udlbl8KHoe5EGvNR/sRqkfl4faIetTyR9n3N0f9DGeRAk2
KslnPO8jUWoJmIUyxskZPAf2pC8l6pOGmaz/y6Y2DBbapoNHnTMvaBfLY6hK7w+AlQM8lsZhsiB1
0ULK0znDKyC3JbCAg4awuKwYz0dVXnrxd4VLrNGcXY+ie0czt4VjkktFSwpRE+djEHPQZnV3tYG4
zz68J+yyT1sKHJn0SjeEtfjFOCvATUOF6fppPuCJvtfYhv0gV03Gun5QVyDSiOjSw+JpiuyYILU9
YMDlMcB3zdJZfo6CSf8rF7uctlwk8hLeyi3yY/g9OuuWT76qhQ43GdRBHGbDmc+13H5og9azYsDT
BKMxrQOuUN39t96uo4za4UQ2pE9Zjk9QCJW14Qpnt9SpitURDF5M++xETo06wm/NI6R0QiK7Xbiv
s6rkl7M2iYauMNok88GSKsygQkNv0jAHGMYvI+PCFBNtcb1CutPcSjDL5EeZEWa2lvPm2ActDCSS
FIzn7HDe1PSpDZ7hrt3ai4sj1aoFrcK9CSXbPTinW7UNQT3voF5qVN8iFYXX+DbJljWr9eeFDC7L
84BBTVyeXFSts5i1NOKJ9pldEFfFfoO3lDKMd8cUMfu+YSOW+YsMo02RNeL78Qzu5p8sxrfqFYe6
HLSDtGkgeGAxU/8vOhx8BT0MQlQGhhm53Fc5Od965rhNbU1v4/M3I03ILH1pyeydxoCNPSC9jsk0
JF/2yG3Y/+ePfyt9NU6h9U2joVCmVW1GKFByaka5ZT/e7SXacrbNJ8V3tWMR/84Qxv09XaYBg0sF
HWVnyxMugQbhtQfPU87D4DFG8ma9wdf6mmKoo8Jqnu6QckuxiSnwW+VkCpQC4LqKzJ2pzltaJhO7
X3j5JB7pncmT8cwqEh2wF7k863nPR/rPk+2eJylFhCFYnqXRdpFiRybh+P3xWeT15jqXvUur5PJ4
KFcqCe6dQaI+LoDmjchFnGu6fVECgzlihnSc3zGyT1519i5dkdo8YnsJG0dK24HinGYO8H5xnnU/
tR7Winn+mM0zt4AWeiqj5MfVcsCaNDKHlJSqmPk2YJL6Q0wyqeFirUzDb3VKwkc5DK7bty7lX6sf
/4xJRBKsA+xAa4K6PoY/t5gX3/NFm3hjx47GSRu8V3VfdDjaVWPzJDP0PM0KnBbM6fEAhQgGwmmM
dG1SdZs7NP9sZFr3zHkLimnldQYByqFxm2B8EfBY7XiHThUa6TWyl3GDebTrnade+Ct1flGMj3LR
+HPDjmpHEh7yV8PpmwZIIDKWlwYm/mfzbUfRw3L+aPh0dg1ZKo6JPSsTaFlKVGAULLUa/ed5K/fi
kjnasNPqOZeLUHxZwW6NMRZ9aoE9h+rJTuugTZ37BND5XHJNu3+g7oYDivKp7JBtqq7LZLlyegS1
Qvn3zyCi8uqwJG/20QomMtEHV+SwYrbGNINS63nqiKwdCzTXoC6jCQCwehJ/QmMjQ2ljQjWyHTP+
/ZHqDVxFq1I3USk2K7dtH7dN9FMSHyQ0dtLH1ScsoRc2/w5vlrR7+h/nMe/cdE+RXezLS0KI6OWY
ZBm9pttsIAFjcwLoQzpTSBrzcOzjHCV6nTRr2GR5i0b/s1xPFQaVHMucRUZZ8OdMXI0UUhBn0SU8
Cj4CaUa23VVFvJ4A3zjHQ85wLi2GnBEXpOfacft9Ti0sQN3mdWM8VcdZZSQUofDywa/F+/TKkOZL
4+fOorFV4RkgxmLUmfBfJ7918oYc5QYx3PljVjh2FwJI5IqYtDAret1NGOkjDRiaD6ePgoY4pBkX
c2IcKTiDVLJpi2EfCag5OXtzi1Ojoe8mvOmKHCvQe0D2mpAmOHYw35BXdjniZJudbfHJhLJOn/9I
9Dd5iKaDCvCdhBs+7cfdRromByrF+yJ4JEU4f4MpGDlN4l7mcKvEcqKAAzyS7se/QzWGghNz6mec
79knoeVRq2coxJvNSpISrjqo9wnvE98vjsvfH8EiZzrSrTr06s63Ajmj4/GHYuRYW6EOIBvpIhq7
+7Fp7Kyxo35d+OS8sgvRzq4wHtpQKI++KjrtsJUnvouhk9QqD1ld7qU++aqLFEavL0KlG15ej1UM
AqO+HIwv3dfCPdwsYVuYqrLgq//1gSjd+PWW1a9xsN/sykAQfbm/0dI+AmJYpo9cvf2yW9M8tXFE
no98MiXiHfpOOMf6tW7yFpiB/vrenWuaAh/dXWGYzeIMXVanBE/2DHYiSRA8C8Z4MM61iSeUrTlF
bKJ780RbxRLGMP05yHWVdLLDcyoNSyWOCSEkCXZ+WsJqKrMjwUWg/09vSz6NwJ03GSPNWN/Ywhrs
+lrLr7uVcmnR1RTTMi3/LLfPjxzGhiLekFjlifcW+VtnuKynVYFOKUc71f/Yv1s598PL/nXrFvU4
DEICKEhjJCiroZKe6KynIcG7SdOrPM6wQeaPuGJm+bqFq5152KTYWkwB86gzV9FktSIuX5A6oAlN
6bhVe9jKX6KckU1qKuer/t6tJ2GqzmxygAMYMqTB3GVb30BdXNe/ba7gU1TUAcUfxLNfsEuEhAOX
t2bHWpu4US3TGZfqn8oZAXRzjmVIgZn8HxhlniM20v9UBcIdxRnDCYyzl70+STMfJLrwc2WndvQY
FsbjWqZVwzeK8eciXfV0n859Ux4s176QPaJA9TOWguJXN+OzH2yYZ5dYETNc70eyqI/bFZ9lXL/5
BXyM1lxAf9o2yBi5U6PVRI/fDgZ/nyALRl5r+yL2eTG6m5jxSoHxqIYOjOMNWIxFuFaU09H7fvrI
XwXo72rHEASwPpQfs1+sAoWz1YfT+KZGVYwhiDfvuGpDfK1UiYp5RGt6eDsp++r0Pn3Umj0hOLbM
p1muO6m1BIAaWJer6G/lKTYDsGnPo8XAGZq8nlCCe+OTV7B0OFLMFUD9PWLgkxCSMasZB8AsvGZ6
gfh59zgB99BC6Ynu+erx1YF5GCLoEu8/aIgXMP6iM8ydx+leDTMHninOTJ/KekDNYxdQcsuSmTrR
fzJph9M/ITDZKCQFIs0h9UcISJkJ21ZPws0StHDhXvcDUVQ0eFLhvRslB5twPARo7nEucEFnIWmy
YflCQQjsMLYTVOWohosIwjIx+JlOCkeuZ/wm8J0h8xwRW6E4kiD/cLMZBnVE7kIY11vmvPPdFIjU
DK4HMLaEYj21nKVXYUPantHsMRhWBHAonXO8fyiTKzl9uVHYiopg6brPozPwhnql46XZhPcBwzlo
gChhwopRfqX8sgy9m1sjqDOJDSlM9zPzOg8h0Xny2Pzlb6nD1Af7UYEHZlnABTfiw/JyC29RODWx
AjKSgjRsL5J1Bt/wj2rbHYslomy9nRKQlFLryRosM4KBJrux5qBXNl6qGc1Lt0jmBrNNl/HT0idA
3XemuQiOh2jhcTFPLeM75ZmnAqys8DG3LBKQ53us+Nv8a9lp2e8V8rfaV+vVU5NLeLpfeenCqnVw
vuumtnUHik89V1RnmvPjjCvRgX1EFnqMzslqN8pCnqP7GjjYMyuQ5VDHyo1SOfmR3e8LZcL+uJF+
qYjmqFttV1d0d4aX0eOM3tFPuQBtrEDKw8Drma0Z6MEEpf81hMz7sXFmXS0qnYnGs1eM6GHCxtcJ
jbdgmJpl3y5R64fxOuZ4IS7QsKgihEOlfukm4rqcBFlsB83SwT5xIAhF084VNc16ZUAzodRzJ+GL
Ul1WY3cBy6JIFlbhqAynr4q8H3ofNf5+hkCKprae7YcWLdnQYWD4U/KG7kfB0Z0slqFuyreOX3RT
mVR5m3a5akMqErzGNsf+4qxF+XJkDy7KT0Jx/YqLzrBED32PaU1Q2wbKsDE4l7+2azGxpYjzvt6z
F+B1D7gI9Ga77w6aYHLnPWnWhAtmr/mUzQdpyox9Qqu62LwE29oAq7Y1cY8LkNlub+//X+tA7Nu1
pPm/RLD1AUMxLnycWOOEAwHeLrU3GElpqH48rzo5XpjXy3RNCSYa7/B5xV8CgRNhpNuVHzdbEz1u
NlAuWdcXocu9tA05vtpHw9EjaqkA0EaNypZXFTNzjxd+yssgDUCbrEZZlauHG1u94JSBoOksqbTV
EtctMqQ7xKtmT6ibyjjbXT56HslBmce66w1SW9461ihicj/BVw23mKsmJmguW/S2oSUrY+v03bKd
lErfCWA4LgK05t8C+F6+HmpWIxDqgF9Fhbg63Dh8pyG4La9AKW/tyI5hM92WmIhOKnVsCuhHmTqF
jw+Vs5p7VQd+kVZxEe6s8l8KuNi5bvoweOsvMpR4YIymlr4VqF6ZCWwLdsyJsYH5kN/67fymwe3Z
Lw8G+A3R/4TVm2bUlg7bT2ZUNxRSfIlzPWimv+io4kUHBG9rwB1FBQhLC1x4UnUns/JPw0Wj274G
/T7uRlHkH1cTft+XzmvZ1/qfwO1L7d9U293DNAf5Oqij43uFBIiocWgygxvn7QgM5r0B0gHa8vM7
cGgpEnCuP63s+ht04GuXiAsz4JZFdI0rRzU5DLEcfFRk8vlHYcD3iZD7M8XvFyua3FW6r6yJoJnn
YyMorHGwtefjLDocs2BDqrfZsJrCb8kQp6cEPE1SemKySpTg++XoVnasFHZcERM+yGIav23DGYsK
RdbTeax1lki3ARgVcOlTwyY/QmBkg+9ylC76vcRoc96a3uK3BQAkGyFAlT+Ns8G2zy6c79wvh7nG
H72l1DhclYQ3dKBNd97BPVcR1NnQ4CR8Xxm/fiI6yKCHhV7NBVI0/wC9bs1dD87O9LBFi95nSkkR
L+s/q+Ypeqk3l7f9t+68eMQNyc/h5Tk0RxQg2BPgWXXVvHBtCiKsQGwLekG8XKyDk1qP3g0PNQOp
ApKte7FcmkBwtbb0C3btIk8g4wnmJfcGoMiFi92ctgY3bnNeLcVfkB6NXcGuCbouP0+46i3Pf5LN
YyV8naq7wpJaddCd6j/qxv+7XAdFWDeW5Q+cU8vrUKaEj7TEKxbnETlBPogJOEo+ED/qUY+o7PwW
3Vm2kq1TRAlqZigz1X+p86/Ty120PK/4KTIbCvDoOdgpiwWIWHc1GNmMPDXstZavx1BzrlkF2Wq0
ehsJx0v/kyTkf1fk5dqFpkHeYT+b0xX5er5G6YjLvekE6IByCg3o/O8xMO1wACw3O8t6+Vau+X4o
Ybz4nRQp9W+nNylBIS1zgdDYzg0WpMJ+m+uINjOAYyo1DnBSjlNFpHBqmZyGdpDaXHs/MV5KjUrj
fF/v/wSfKo+6aK+ukNzxl8K5qXRdEHP8dld0ZMy7fPns47VwgC8MVsL42h+0klq2js4B+eegn9Qr
adqrUuMPA/eaSKR93ShAvIqt5tO8yt8IhujDPi1gpFbcYgJDXn4j1leBUKVpIKeJorR53iwpd58O
t6bqVcFlW3gSMwfDT7eXMJkNGxf/WeVYAKu+NowN5B28umiWfMQ2qyRe5M1e30eDjpUfm1LB59f5
6dx+XQF7gU26c2PC7Seyctm4MYOmenP+hVwzW1vq+b/s8lmX3c6MqU3Rnc+iBpZWSX+bv2gzuxET
12OrWd4PV7ll4iW4O+D1pWWBE495g9N+5h2Hl2Y9EitTd0ZoWrlfYXSB4NDl5CSl6hp0jW1KcrOm
0bGUTf0ZK+yMWNd1rrt14ryp2Wi/M6vkstlgawptxbNvF+FvXPKG/HfL1Pth7TVceZom70xV4tBa
a99VySsIo6jwNX5+5p1keJGi+rtM/ZAwe6PALMYgXcYG5e/z9OOMhjn2rSCluaupWmJbJ7YkeetI
ETL3Gpaf1MyUqlJcO16wJubDdCSiPBNC7YTD5Q8VfYrM9spMqfvSzfwChSZNAt9xILh3H7r4fIHx
mcQfUKET0j72N+LQHt88rd3hu2ju6eqg0yvcSTrxIetHYyXTKdF3du0PWPR1LwhGvEp2Edsen6cj
xGtXfft4oYYHthk+XteS6wyJJfG+lmwlUlNrOVF4o8vyKO/eBLXWVLNJfhSYWIfWLq9ogK0k5qNd
Itns2MRdueO3s3sBvRzbBsNE0nIXvK/foj3SerMKe4nZuIVBOCbZVlriwBMorHAVPseyrUOAmtJb
NLT3xFDdAWSYan0nvuyu4UCWBxRo8PQcC+6S5PpOnwb42UiQCBTNMJZkGsRT0MTkFtTP5RkxTUur
1ghcabGJGbceLccHccJl3wG8LXwVhz2K/G1Skb6G9+kAxME1aMNuUuAlClCCERGNkbd0NXVf2Knv
L/EF763lj++OYxkF/pSx12E8XS3UNo9ybCj92EayW6GEERb+OkCkTvTRKd6+eIxztjsucLFtscQr
XWAXWABdq03FoFV0DdETMYiigTXNhmkmKYozGiJFhdYJbTHvhSH62BqctAIfLSLH4Bv+S1+//nEc
QAjFDTRB9dyqdYu2F2PpDuVjYb8yY0jlXi+f4Ul/ZJMfQs1fbB7DCQw9tqy1H63jOmKD4ORJ9Gk6
GuSzi+sfbtfWwPOjR5Jfh/L6Oex4rF/HN/uqJxW+0Pm/S3M92RDimmE+Jc3KDBPav4jaxmeXnBmJ
AmhN1s45abTE9VvOd62ivnNXvJqEdCPkdlPQ0r21Zn43BVmvIeW0noyNxNdIivPjpfaPi97aq7Sw
f94T+bOKC+jrtLyCbg7Pp0OngajMCcwU7RBjTdXiP8kdNA2X9BIUARxbqt41z3xusENjnk05u3xb
v3PS/amZQeiDDhP5Ea6U91I1njRR390frQSmTmZ+nM+dDClJMhUh7oDkBiyGePFqTVwL8JAPnwL3
rxcNX/vOFNEgwPxGWoaA3b7F9+SRhgEM2raL2Oi43JPynY1UUQfiTBWWHHKqPtODx+RjuSKyGg+w
VaDfDFV7XACnFxcfbIGCubt49R/mrsMlwmK/qiG/rejLG2tj8CTJ6uwYnnZjs/Gx5mmpw0UcR7Bc
UNml4ySvW+qKNe2tRmpS9kK81yLGVsfDFK+DkGvlDzpv0YNSYgkx2/1CYH5OUyGdzZoykd1LkQjU
fthzeg3MFscym+IEnL+JCwBxkstPfhuzcOKW2vYUdI6AXgDrn0NJhGOStsXuO3h2jaJy5s/brnsQ
tF5qQ1wEt/sREziVnFrFsNeS52nH/kuayskMqfgLanfRxTAubh2/dGHW+4ixtgceFyFKe8z1FtTH
rJ3q0BR7gGUMTUuM2q++KMBVUbhc6vljkHd+WqhWCg1Z21ttys0v6xuDILBQ5pzkwgA2hyaVJwN2
JVuwScPuI8TdE0snrKNQp8wTqx3voBo+eO7F7cRKAXRlneTwkUNFXWcZ/gLJ5ElTaL/+3oApuorl
+Vp8AKWCw934IKUewKsVBMy3/WR9refM8G/SzI34T0q9GsSXeYcYTyqP4Hohud+xeyadpKdVVckQ
69R+wKELVTAFjIUtRTFVURryQIZrqle5BOlJ24qMsDpH8MBLJ1ZfLFfAwqu2nN4vJBmCtnkrecuk
LtNWoUk8zPhFd2F1SskpZbcEEIQCQTrdc0tvkz5/c6kV+j/THrOoPZKzDgHc61R4y2jgtK84etbJ
BHSE1FOyjQIiZ0BXlDVzw83FEP6XGqy4n9MnwWFMAkTK0l6ozsWfIljeVL1CSNHvj3vkaytdOsS+
AMKWHEefZzSb1XqPhByTrZO4rtYeW6xlStg35ANIMhrlBwUQ2CPj99xEJ/9X1q2bDi9Civ0JX6uE
NIp31WWBvzIbSHBTGSuoDLHHk05nWFZEQc+upCVl4NYlGXU+Udjc31CnkZA8Bc4hC9UoYBOdJ10b
snfJ/QvmygHQPp0OO4WUW/fEo0dDzySVpZBDCmwFXwKHhyR1qfdT6zmcbjv3OCMCo1q4Wnb2XL/1
fkp9utQtTaUVXWYYJ+Axa/xbkn+FUrObyFlFSpSRz4+Pyv5uxqs/3G+LLAk1orgrwWD0vtVBDr9D
iH0lGsHVgB+eSXG8iMF6YQs5D3NxGtfIxFHDYwVyD0zM9Q2k0cRQVruCiAvCJ7kb7wkItixHy26t
0MxOQm+vQEu1BV8p6EUZXHr5iBnF13ru9tuRzHuEuy6gcNfYn89yy/xehvYL15mk4PTgbTCrU7UQ
jonEB4hNIpZ2Q2dBh+2EmtJIu79B/3R0VcOAbxWB4dDhXTavZm8325TMMIy9BsnUT1CTY75P9xHT
XdyjVySJF5fqXpM1IFqpe123QCVufQ96sZ1wQKxiM86Wbf7/Lrzw/z8JiZyHGTPl40E+Y8mgLjSX
OAT8F/Eo97JQMN//ez4c+Pxz4J23wnK16LIg7vATxvItEhCJhfRThsYvxAKiv8M0qH627frQs0zE
vnFK6oTEGVzZ+/T7gu811rneFcgrHlJtvHB3Dk2gBPkNQ8BM5MbNqmIYdDRh5s+4L9kE7f2C2SWW
FAgR0zvCGZeoYimxrj9bcrAhqJDpie2vKC+J/wEgzbx1V938F7lQmlRT28LJM5u9XYmKf/25Ibzx
J3Kg0Cbkd9AdLS+Jc/sfiJ59cISr9IcaBrnPntKbDqtfWVsMn48c3qJLK7jfCizzzbKQQfFltJNb
w1AwGo6+DcYqV1rXv4FiEwPxTcmBt3p1A8hZMxY7/gsUwN+Ad/JD7NC+XZgk5OH/X5HQRXsOplOB
H4BP5/0PWRLVrr6SY+7RqubbGhLaSXD7oKWPGab8d6dosIhIN8xfpZpws9RVwI7dkMcqBLp5Bb7o
Ma5LXYRGu0wE/yhpKtyyhSdGb+uA6FNiWzof+5MCKWMIfUTC3Wh9iXRlHBUrOaVvzfK9LMfCumld
eSMIIgZYWJJPcCFZpcphmciY5NFgjHo3y/4nlIvREZhqc+eXQweVys3Sp2uW6OBhxYFVp4jtbo0c
rNZi+A2lUAsZeG5zvAXQosWTOpOe6pKTgEX37tPtbRw6h7aDt27lOjLA+44uahbCD3ZJJ1I0QbJb
qSZdSZeinh9X00tAs/lF0JwWt7kYeGWxxh0lr8dceSY0bl/CdPQsqkd22zt/O1o3jG6ReeB0vfJ7
QCfbIRozg86CSzVRiJuZ5P+TmPX7c2rk+FuvI1FtZoHnnd7f497qsI2T4cVw8QUmlEo6B1ndtHUt
HmYm3zlStlYXaRK91yg2+Tns9iLOdR6UUF54LMG7x4JHTGmY0rReFO4O2lDajJ/1XgoAWI+ihx/T
XDklK7ZzFhHrOm5Kw+QYX8uA4CHW3FEMTTFUqNhFpzLg8pyg8V/AIoha/lAB7Jiqk2FPEQuTqjwv
ja0yDhqA899bOduw0+p8B3G6u9e0B4JW0w0Uzngpdiff7VYmJLWhYWcfveKJUMom797YlNcLRVWA
dJgdgygGH0LAlmFD9k8EIO5Qpq1lt37zCGRewsEQBYlcPYt37TBuPQoCUEN6YCWBMjIOnnfDsI0q
sDGfD3PpKDJ9ZPAW9e/myUYvujSeAk1zk+AiePFJfXDMxTlnRux2+LNQ2gryiW8TjJO5DlKkX8Sp
HxAegBG0uFaSakMPQSfRfJa7Uw8nUhEcWx6gnkSuabRKPbH1dJj+6UnNdA7l9G6A4l0F+JO96HGa
rz1LcQrG0iTVuPkScYp7nKgDiHeSaMBXucxLl5gIFBJ496y8fsH/0/IcmpB9UzuUKhYNKY4CL+lm
nE802pNZ4DI3iUt+1HNJyduXY2v0gvykW8La8nOuA7v9LHp6XG7cZTsADzPc/A4Yd2ruFaVOM/I1
V6jMxfcvYHtBARQRAFJaNHpNM6dT8BCwNxB/LFQWgECmLSuuidjlkoKJzgEFeJknzFkf/w0OXbIb
G135iAYwhLx8Dh18unq0Qo/SR+vdQcVDRKND/MhhzBJIMqGkQIvPD3Ci8HpCv/etJbUHUNs1fo9C
OnTxdTvirvicPCKWQsfSs8Vjgn3PkEdypFLq3Rudg/8x0sDZcmltQ3uh2/qOW1Y0S7ids5xFHQn8
9wrGk/Hz8FlWHpcjRXqQ4LaD8gSfWveWNGWmB6IG+uwBiRkRpW92ANJQ+myGACNM8esZdzJpn9Wy
ymIS+5hQlaYYdIoPKu7AJylB1a6C2qdidlmJeFVvbuHqS7VZ3IaU31X4/iKsjteC1uKVBvtt2NWG
dFsB14KughsBNh/nFEp8A2KSs8R2J917AM0OCZTIHGN45TObeEP1krCG04RLc2ao8FIO9oD3xISq
bWaklmL/kDIWphqW2QCu1QKUSpg1rDfHk3z2v2eZhr2AlUqAjXs1aYkl/1pr6fjD9fa1dcpfCSq3
U8G3t2dLoYi7nVzCXbfz4+Cb/+JyZwtz63jdqC4KiI1Wj+Z8uZa8WMcxEL1RYFyOTeeR3KJebzxQ
wBdngTkrwEMNv1ZljIy7rSyoXKTagbX8oLjGC7FAtT951LyYPHIrg8vdVqfMmlw69cAz9EYp+E+R
72E0BDXWwa/3poxFtGb6CaL9jdy1Jpl+EqV2dMekcsU+FIMrV3dKoDFBEbV3jIKA20awgH4rOkjt
lks+KQSTRIOyBKHKeT5dGysxoEtNHBQNDsU/kodXocHqQsbDW3WT+C/H63+owaijEh1Gv5wzcFXu
ouN1oVNjAWt1Xrnw+S/PLrkMJpdn5bB+7BYqec3j2f91fQaKsdLpUW/MX2QayhQ6t/Tn9NedxsUI
0NAhwQMoI2OHRO8FXbiy0X8TssPC1UBTwAkIFZu+RtjGhP8SH8HP41535C/nzWYgrXSII5peNDG4
E4fIPhbKd/s3rnfMVwC5X3JXpRrkutzQYbY0DNljNrNrucaPAtkODmiQEkL4D9oofN/Rjds+ZYaQ
2ImVjT1Qutuc0IGgV79EdQpjm6GxV+KgqMo5lGWoHN0Okfo3W1NUjBMSO+gMRIdsotiGKaNYuNe3
U8HyrLqGZkBc3fMIH6iAywJBOJmX73xeKAdCEDknJT8WhmniL8mt7geY+i90LWBKlUklN2mEuj3x
IWG4xKwEoemp/0+IsDOfw/2SIdXBorUq3bYk73JHJ7TndObsLO25XvJXIOoF2xW6Jixn+wNtGTkz
RQJfVHXV9XCih61g8M+d2b0RDPnzGe80/qjE4Hjy6KBQd51Nv8qSPFGmELpmS6qcEmCIpx2W7ALy
s0QC8U+/K9YDmZW15CW3TH8JxQM20stF4tynGFQ1UwXjjRxZCNfRR20SWXJLpDvNPqp8G9vmOgl8
yiMZh5iKs4DQntZcjsuaesAte2om7Fd5JiyNqSRbFKavCVzCS/AjMbNbhiQo8NfA/Jn3jTmpIc0D
abY6bApdcmNGP+4QjSztZolqdnY1529RUfWZp/WOr1UrWxkfW101Zix8VKii0plmven9v9NKD3cJ
+sfjDVk9Vlbyh2V18m1T6Lakqa9EbLcpno6ZK8kWsv2trc4nnJS6admXIwF9w4DrmXwQhZNwQbhR
m/4lLIl3aDsxdQJudf+TBKd94ZAoNjGXcVByFpamjmZrI4NuukLIecegkfLNikodhHQXr6Uv59Sx
UhMDg8+vJpWXYg8437CCqX12zLSQAOttAYB1TOPyw2E0S+0U1ZJo78B3hpFznHPKj4vgF2jsTnbp
LmEwsOAurqpLj+YjUAniq4X26zgke+e6SZFBha0AFglxmQEDO0+o+AmyNSxP7NiiZjdTA/rPTzKu
xDCARhZXMWcTeGIHbgimUc/1THf4VPzBNKSAB30OwYuBRxWDusT8vw4ZGJ/gTiPPf2w3r4AdS7t3
RR1G96ZzV5bs5y1qik9eIuaFDnBxj0/A0q9o8tSJoDUMCrP+wcww/rA7tbYNuZD5ByztpTax+SWk
alg3Id/TLdQ/XDmFoYQ+oIekb7wLxJoevRp8EZp8TYp1oiBha5KHvzIxUVSoRABBfuHdo1RTKBhV
9dxt84IjiH0R9qdAVKj+JX+bliCsDP2YOQMbVjGLrVPlJMruKbVLeWg9txSOZgsp3HrCJZ/eKhcW
pJHk2T9+DeqoQyl7H0ZJ+S8l0Q1OTDiPgR+cRJ6eBQjDW5DvBVu9shOR0YCsAtrQDnLWIFNmIHvn
O7X5isDh9hNU7wU/B0bwYZn13kVq/WLitcU1dVZDKrBUBP1kX4rc/YXBzASNtuJAlsEHj3WpY665
CaS6FPfbPAtRhkX5LpmKb7zt4JJ++BZ1KWLlJoATgybD7WiEvrDkaaOCwHoH0cOtgedrKkWVtidv
rVXShKUPISqxwyE9DwjjD4em8zsYT2GjOMzKkVKETkHdJcCfA6Jd8Q8+RRLhCBwoQ0vUOr6qONPz
q3P053aOvGhlTsDrqZ2o91WV3j03kJATeMW2pe9T28szuUM5NR/gvrXjaOeDSg3ThKCyFkWRzGIh
0Hbe4wGPtjEAEWniRDEnj0e4bcwND8oPeBW2LwdyvGz+XVCcVNnvZf4hToTG5NCBaHYqmxqh+QRX
trPQpwYSltBBaXeJpzWu4Pl/wLVo+EjHscG3zZwiqMqWno2kDiqAUAwbHTHjigCJhgFXsLiVxks8
xttMyQyb0a7B/mnSxOgAxCUe86/CA3YNuGm2iSjLfyQShZ/8N7hIpcx8dOocjZutOx08bu/xRJZk
45iYfh9qC+3C80jqQ/PHNUyYv66wgF+Iagjv5laINk/Y46y6O1h27KpS/W3PzgPbzOhEP6qFRIhu
ut0RXnsy7P2rmOv5j+PUj94h6JLO91a178u/3bk3YwdnEFAHgxDknRQ47wzsOvjwNpsdVGeEqpl9
qChMB03UZH4kyj1oZO1kqYSPKPNuYlnlcin3Fb/eDfEti9ehgIIMtS0btFdrQCEcIMP0OsBvj9KG
cjj9PCAtHWjd2WMe8Ud3lhyKDWapH5JuZEmI51W3tNb4AR564YUivsFY37S6OIukleAisSXnagUo
wdBJ0FbGIKXMM70MNu8sR8qhRO8D17+RmgTGaReQ7cRZm1iutQvGKzXTXs81ypxQisj2Yh1LlPb0
i0/uBWCZABDzYbRK4KNh/zWCLYkWezZ7fLvreP3+1b/7TNt4StCSzVVd4fGYXnKKsj9FA7bXQyDD
Pp+7iyq6c2kX2ykxBczuEauc9PGd46IEfFDebMg7bxnp6QZQoaMNNhiv1J/a0+w0zWAumt4ttAnl
G1tloCSGVYs3T0vfnv8KDM5s3GyEpqQxh+y2jiutmAa31ymDQsSgIjxwR9GAdMVLRyRomWKRM9Mw
YMT+VFFyii/xdl58hNngNVAPdGEYoYILgP31U5DgUvN19qaU3mwYfq2VDx8w7Q/KfmKcGBZUor83
MhVB++9D7AcfZhuFVfYYj/dWZ0wh5TBXuEyxRUEzogI5SH/a92R+WiKXVL3ZT+DndAHEdwwFSZcO
n58rhPWZyTWHa//8yAEXe9wZV5Hl46Joi/7Vt0Yw/rTB9LsTRv4Q5ln1vN/FA0GYNDHdTMtqNCyW
RGfARM/hGzLh9ql97TUlVcwyYz5OvAi1Ul4FUneBcbfbXAhi63zWQyK6Db6L0XXmDzyW964FEQwu
AVVoJqS+CfATxCg3lJ3RGBuTuZ5vhTVclyJzkgGZQXoK6DIRqlsJ6ZPxp6zr4BGHA9UbOVOaPZ2Q
p5a4HzrRjnwLq5G+7Miw6+rnWep9TTkArnP2k58nRjxtGKG1AAyyCXrJJV8zqcSK3VzohxqHxPTY
53Um/9T4AiM1FMO5l7IgfSQng/yTXZQI6SE7dYAs2J8+afme+u0i45zR1X5aMvPdt4l7TnRvPEOa
WqYty9AsJYVXzceF8P2B+XU6Bfck8bJhATetMdg4qSLSDcG66IljXn7yiHj1v4TqCm547YU2faDF
/Qxd3MhHoPi9Ps+Fwlo94rAl+whrvw2Qx4YEWqWBgKCeW6YDMKOjxM+wUpBaOBpwkFhO7J37hOnM
m6e290fAa+aA3S82LdMOrAcy7o0exC0/EOP0uTKuzvugKHm9Xh0Ed8osxsNvS96lnhJATnPIq8du
Y5em4d3iV1JIHCyElUuz9PUUMvyRRU5U7uP922Nbg3ueY2BKSW1aepXO2tE8y4s79p349q3ZUUfp
AWXT57TA46jIOGc6LzYiZ7xAHRzlTv3iPl3VdlZa5PmBOu/t2eLdkB7eUPhT4OioQsnCXnDIHPp/
jseRV2FP1pBuzqBAKJUD1w2Us8xdaEtZTj4BPuG4Kf7nB4AaV3+4YUIaaSxPIw1Ks/CJDGjw4pTR
qOliSzahoj/VxQlKvGcP8STFA0I7AVkW4HvtjUlfCTYdcvyRNwMvzPO3rFzcMswF4oISgIN1tzhV
ybaeTjQXLBTZd5UIrcQkmyCNO7V40JymnsUFC5nHKNxtGkO4Y9/9lWFGx2NSnjizyOkdig2ZgY1X
HIwZCnOJofdsCjG/BW3gDStnIPIEdiA0G/LQZmpUzwVdbN3tySAONkrtLRCaWayosqE8VsMnYdTI
IM7IKb9JWR6vXnCVObvcc+am7imtNphHbsmvnGTCk9TlzC0g9yWBrBT5EcpAfgsUM60uZOsui8B5
tdkeWU9o6lVgL6/IupiZOveud3wjT6oW9kLVHq3eodmSZbooFxEucXBGGySWLM3cHZUmrn21Vwp1
hGiUT1xsfLDD6VSrzHsUayrnwVTVP0jJOOKwhCeUxg1Oxn/oPGywn7XGCH5YTJbyyQCAewhXl3ZP
zBkKbL85w+1Q8tT7GR6w4IAj26m4ptQY+ZydTlNBE2LhOiZSw8rquGzBCvXQW7V02aSNihiyxvfT
G9TzPLrWAtFoMj9Lf+k7ZDz01E2atfvjSHP/UuNGdNMtFSgqyLRl27bvwK8wK63duKjUJ+7yAWUN
4r96RJieC37A7vw6ViMLJRdzMEAyCMuO6t/quOCsYfe2wy6Gb7oIXs2V6u8bmRzmduWPUFieI3bD
XN6w/oGYq4c4ymDGM7EX4XXZkaV5HP69GVFlrrtPqqP0LzmoB9RR+E3cQQ1XbkQCND39vbLu27MJ
8vmkk9K/UY97iwGWdn3RkwpXKnDsiO5rgDfI1otNNG5WcpMb9XyYo/phMAOngch6TR+qsXOmB4o9
w8OEw7scM7JsCEjbnkxX6LTe/hTE2kPpKFO1ugxEgnaEsZshhgmb6SuK/Vj5k1Xuq8v7iikKsrKo
WgFZpLzy8AqhVKyj7qd51c1nMxqJHQJoNjYIyTQSvGIlqBBpuQ2yJv70YaOcSHp3sWE1xAUhp89N
pq+nBA+9C3SwhI3L+YO0O6/EWtvbhjMLVV45LcuFdNrWq+ibw6j4Ru8DRfrAx+kg3fkXpyvbp6kx
Szz+bnG0Cka2unQv2ZGsWHupPBZlyJ+iZW6Gzq98Y2MZETCusjYZHtN/EkrpY4SiR2tnpCm8jQ0M
G7jR83XLKa85ATBIvv8pP/UI0/PlJgUTrmwxGZTbccudyzPi5j7o3xpTSL+ANqUbIM6fCTPA67Fq
vEvXMgnloDmdudrtcfyNVD9R7EfEPfyY3ctfa31S/JVKrMNDSqAzAYe5P1w3MALCuE/Wjyg7VIuv
UeTYrF8j7LyPvZyUirKg6n3lJMDjTraEcLo=
`protect end_protected
