-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
bwvodibBOSlZVhwHp9f/jcmmYqTs0Tjoe69QFqj0dy7mAgigduDTutDTqpZ9QZSF
uqbz87pE6Pzoy4BB7gwNsRjDekjA2n7LANlCaotopu2ZGX6QnpwcPn8t8/bp8iet
WjI8JQCRoNUIVXHi7jVt8gg6j5pL1r7scDfC9eMRJJw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7957)

`protect DATA_BLOCK
TtADn9i8fx8Bi48uZ8RjHEKZNB3am3SZ1Qvt+3YxOMCMB+bNWi9ZEnOEfxN1s2eA
nnGEQtQ0oqp0rhBB4mW+7NimpHQwBmJnk9aJYw6C9hYMRKZSAlCJuocHsRvBWlVu
iVx1E9TjR+3aZshnGeiXL4PVzH5hWjZPIWf/0REUaW4Kxbu/mnJjyizly64zboFT
JKJgFNhNP3d/8VQONYus+5TlxTqUnCkFxp+39TegPt0SmXfrHhF8e93c8IKHHX0S
hWl0mM0ABdm4pK/nEribuLCfClOnm12KUTFhIPJnKIAgRz+sSqMob0eGIHjgszsp
NoxlaTX1s7l5gPCGQuew9DcY5b+7TKwrYvbpt7FleWM4JlBjBFVUzthxRzhd3Sn8
lXPZzC1idppqZf2tKac/CNsLVr9a4YECaeYYdD3T1BKIhNdMi5qDfh8rb2GzuvLg
aIXsXJoNIQ/jCMKGv76jVFx4EjotIErEItoGekR5ZP29VwF146Msuej3xToOfGR0
VwLPXuscPd/QgZK0ELmYlx9Pf4Dd9CkjgkL/y8TMVbTm+S6sEN5wZHlGh4QrGFsF
kl4BoInPH7kGn36I9pi9L7ixJ3cO9uHv0SeP29M6BKM6/IH/14rdwFpLrluayNg9
W3Qm/DC+IlFrPZNaHgK47Nifpk05rZHSo8l1WnuYbgx8MHBkpnjrlBfoDKTTLqr3
a0rTNoHuB5vam2LjSY5Ng/x2Hxz0CevEsM6mWAw0XdLn/tsbDYIEMoyELJ1CU3tj
Q38PR271zVCVncyfu4ei5ySlAHvogptVB4+xOrXqviWr/WED8xRoePZaEQMaWN4o
kXo6+WFjKNsMYfd4n/8JuMMaTGOyplWES5xOaicdYHLo1BU/lZ2eB7lpeb9hUjbY
T/qZzvuXrw5AXq4UmTsGe0BVMLi1JOKfwnCahpVgo31OyzoVDf02OagUzTBjKug/
wmy8FZkqX0AP8rkJ20rbVS8i9mkeHZlZZj2qkARx/2xlsYg8Zk1apJnKHKJhVwxW
6WltCTAfdscW5Olfhx4+iMfMLJeiKnlDE0IdBM+RNZVNnhCccm+jaaW2Smw3Fnxq
lkwc+JOi1mHQdQInf0JVIv3kTNSbKLTl63Ra3I9r/wW6HToIzX8Zw+iTzibmG+Fl
WfFNcfoOW4L69kT5dpoYs7TcYxn9Eua9ImGdPYDdNmt2dxKh3vrVUKUxaxOGP5/w
aCxPPKIfz9x4I805Qu+Vd9Hrw9L/LOwPP75sW+ZCJE8d1WEC9X3NeoQgMXtaw4+d
V12o58s2ACHgsCT3TnTPJsAMxSeustN6jWhEEyisB2g55ys4EUrrs+fZTvJMcXXm
WTfJiabDN9bFTfWKrgkSrC3aLwWGLRveMVbF5FdCiSN081HL8XW/18WBTPHo58fv
A0Js/dmJM68nbdFJ3M7SjT76XHSdQUj5z8bRhlEevHqrW1qWxUpMv6ATqoUfZm/L
EQg/Kvay7mT2N9cFEPVLlrkXnsk9X81M3UNsQxmtqlTAz2Sm2p/JQ1ShN82RManK
iJyt8sQEmLaEWBLL0RYryz1ooOPK70xWvdzl+AtZ/m13zs9SIqf9svXJZ9AcfbsP
p8JdMEOBaQCxJbbn/hUqXByUw5FB1P76p//qWcfktGai0koAi12fq57TNOXFIAvt
+Z4ZT3ycXGXFFUMMvz3eVuPSHJmpb6AgwUtN5yHgCFMWOMvC0u/UEYpbRvkXv0mP
hSH922cCxXjuMqXLqALYYN+lzDitouEmsnnxNgfUHW6JmJxnp3XWAKExzQs599vp
sboYgade4YPTMgHk3bXeaDgQR7dqK5cEni0GhdDKQwITINEeP+70ZU2pjheFF0f8
SwIs5JERT4BAULuPnaALHCpEM4553B3BwyE6v1wWIp02MRxUvEHhbQx7Eap+/qrG
xQIvvJxm2AOEZQ1ZI14pVSLEzTVdZnvox892gJc29/cvK8wz2QZF2illj8jMHHRd
/m4v7JKciUBv7alU5lYr+HLsbKi8KDMvJVg1GqyrbaBGPst6r3ajYKmvzI24P9ke
zQOCrlOKS761oOGI7Oxiz5ddvOBVOznTuY/PT45c++/0lL9qgqftgt0iOrz4rsTV
u6yhQsQhEEopp9Fqlz8nGW7Xlm71frCyk1oUG2wV9hDcNE03/wmehsBuuvV4VhKo
Dlm/Lig7zjK4ifw83pFv2JcY7PDzMOh2V5iuWubPvihgoOphnUCASqQRjWn+f2E/
9p6GtANA9b1euugkmcyua17ORwsfp3cr7WMKteuFcYM018cq5VjDcbkcqOQY6/OX
Gdic9NF043g2WZqh3dLYuuRodPyJK9MWd/s3thyw0IL1S4jPIUmJsd1e7aiXWcHX
GGglF1xI+jXS9H2GvvLZhFSBeDHtAYXknsmkYlb8DgsV0QbPR4YWIz/9TTcK2GJX
4sm4sszdYEKIuw1UmVc2hezPQLRCukMCpYlQLeUf/65CkpqDMbNez4PA7dHdAt9H
Eud55zUcVVNMwyKh0JonA2O5FPVV/DhP0NcupvHYRVKSV25k+ghdgNCdo9PKNU2m
Z0yYc1Cymv0sgGT70K44UsCNI6Wy+MO10H10AF7xNwfaOmaoljXVzREnfSx1iQjk
2livFABP/rm1K7zF7+QkmqoioyTiRYGNHLjvmcYmj2mJrwU7q9K9TUQzRSSGvyvD
YaXuR0sowPzWQQlD7ATxBHxdvXhnMCS0ll95v3ZFyqYGP267kF798iqYyk1tIHYi
YB3HOyoZLyJ7LcSUaexFuNeXeOpGopCrfzS/p3IPzqUaDjaL9cyEk/Eo/lweMj+d
g4kccSqTObiu7/dr5hTQE+V09rbPHgz0Vbiy3B5ue0vRKyWmbpyTSs/VLnQ965T6
5jj98Hk8CH6D5MLY1MotiDKBl4IDYsggoaX7tmuyWIZrEQPpYOtE9uvOleZzP7Cj
cJYZR96sVIQ4nbNd65pOvnuli2p9Y7M4OEcrEXQc2/duvO3FyMuNx/FhMEcGylr6
IASb4p2deXYJwJ9tiw3wDFCPO852AagNdJAKmjFNN6Sap4RdO7+E3Sgv75I5n9u2
u5seJt3ZQCa8IsE68Gtae8b4KrXRTq7zeEKsnapWmthCfc4jVZaOnlwTc0Lhpywq
lCAeLmStpmko6Bg6Y57u0GImmO5upVgWPuAPN8WadcPaNBdVHwKNVReHiwPMBqEO
CTicmjK0NoWjqUffcFAmVRJHuiGvfrQUfTJLXOUy6c/twP4VJW31kLOW5TAfbC31
14UJYCUBUeqqjxZBHl7p9WcIlCNTDXpKJ1dTyLne7GResZR4hs7G7BLFu7P8nEgX
aE7sBv/WZUV6tieiP3+DT87CsICm9LGC/H97Frsp7mHGPL7OvCbRJbgbPu7+QR4I
06YMs/66ayyhDU8c3N0C3xWIXMc2vaCxIzuRfXF1dfT56uM/IbXD1uqYV14uM6Zu
2sEM4uUqStKRINDzCNJecTaSVtDsEhitJQWdnn71s/fnqv+1TgoaICtDnzHSkGS0
2cSOEv9mcm0P08cowJ4lChtDFdO40enIGtwnXJTMjq5Mxn7HSa8UWPCA3bKdiySY
gXC7lUTbvWE+s4cXwUOy9HtR1zwxtUQzcWWLurAVYEzx5TGJJb0FaDZsTqB1biiG
1SVpzLF+Ooahk3ij1t9uEG1IERgkT94+pb6go4FcSbBp46iN9RFy27DXznlqT7i1
TajLOuaWURMMpzMoEqvpTSLU95ZLG9hVWhMIeuUZmVirDnHsapQwawDPVS6DiR/A
OtMzp2KfzpewdoTWOkdRNtJFEQDrE3vbI+08Lfr4I6FMuYOWuyVZY+YcIZFqzU5f
4ZW6F8kBO56uZGsMyMK+nvwHmTYXJtO4XeccxFg/pCx981GpbgC2ADyc2tHzTclN
SQq5z1L9tdQUZF5aQyGbzHYneZQHolOSZeClD5CbBFxLkwPzZSjzIB3LPcyyxFnM
H1O5EDCC2G7yU9mPHN/I0vzo5us/dNotIVKcsr/e/ChbkFC7DHR6ujTAuP4sk3vg
aXIQ3/FQ3fljgEIEzVV2kYre00ROeXxEf32vVDx4qlKbRX2EXlAZgnT9HBRv+ktA
FZ1B4gu2LL44/d8eR6NlT1ANOzx3STs/qLyQiA1CNtDUZUz+XoFklWEJN70WsTwo
ZPHgf+RXzntA+geTgnBMV8460Y0W3up8YkHe9Bz7Bq/wV0OqhhOcgmbWlnJqI2L+
Cm3GwGrP5XzlTSAO89v3Bf+MI6tTXBQjLa0NhiSav7BKusZZ/1YbcQJ1cMB0ES8m
wA5XVJ4yir0HX9A5iJDCpSBouAm5eAwIK9AS0zpsbIRXuZfu40G0276msvgEJHF/
9KuDH7knsRuYk3Y1K+wv9swvrUNSyJQ1Yj1rBvLYkXBw+Jgau6ZPfzTEE8RYPY7B
1E0Pw7cioV+D9tyFpfftqc6B7+218xsudJDO3oiiXnU6lTRFRaUHeRInSPAT6hCI
Qt+k9Pb89d5GUv45QTWTxGjmgoCEKh8THP265hlUFIHcWYEqiWkZTFBj1KNcRAUh
Msz8w88Z+LTBjL/fQN+ec+C6M0LDmkM1OdKYnNH8PrWnmKfISACvVPmWjkD41wrf
jNi7kckGWXBDW5e3/l9fYuC2jRS0PrgPEK47PM7LzoxjihXjnZpKJ0jo6+gZrYeP
ZtmaQrYSAsshn+gGKE86HdSnt4rm2G8plGlGeu4WIkce+dGbZ8uSVuYzeD9Sa/vZ
Ve975M79ihH3zVRbs/+x6W1kMLsxUI8NezWADeR2w/W7mX22wFBORgxg6LzZASsk
g7WNcFd53rS7r2/MLavQdMJV0mzOJnQ6LzTMPMy6Zi3XGXFRPMTMrPFtu49j/6yo
3Ji6/0v4pkeAWdJfwgW0JOYBF1DuiOZbErJToWP0BGtXWOxxWl5jpxXGNuOTXtxY
zeiOnPU1gDUaDWy4z1isctsGnaP1D4Y0Wahsh9BP4fpB1PH3NKYI8uSox1w/o3p9
ho/8euW0H/AjeH1eseMvS8f+bkDQTzcG02n8tWMO6Fu5tYYb+2yCLga76dO8luCH
SYpQE9U4lfmqQTJetwvU//MZCnjVHU2uvs51iXLGrJgpgPs7w9gUJUPptGMNE0es
mCSmexG7gIGweyVXdKjoEsihwPp9d2y6bHrMjxTEw2enBVa9V7OxaV2r7XumhoEV
nDkgO6VQmtOebXFKXPvXPV3XOThfzbpISsKUEuhhFJCBwMGJI6rjCNMKYFo2vArP
JvH64IHlt4BMXHgaGkhP+CyaSY0krCjwJsRUoH7NSo/WZD7u7E01fY5XlbMOzrmS
y5t9Dhz3H3UlY+9NdACrlwT5ago3izAGHTa+BjZ3xglSFO6CeXJOPj3DnsQSlwnm
jffEry7cKgia65Yj8J4fdk5sLlr+7dXcQzeu04TXEa3r4Xm2TKTrc3MfT4zvoeji
ue4uuHAiwXTQvWF6d/jParNA/6Fz0HpdyM0DhZv2Q/aIb8WOS+rk3n2U+xsxm/Uk
L1J+Sx6cDE+YcJMq9tpxSorTmWUFJX0Ytb0JIQtXrju7Q+ZEXmnLjPKaaNO50eUp
XrH6zIPSUlrR4Szb1CUL8yxMmssJPibKto6fOaEY+smwSLxheNYyztkb0WcYvn3s
YLkLfao2DgLMIKvdaBAqax4KwY0VZmuJV6YNqhxOOMQn2g43w1q77DeFMjhLshOf
3xJN+aLWkP9kmv1iA5PWJPH0g28D3y+PILOuwbweTCPZINZgBsDToLFWdxlE+fFd
AvBu3/tGwjBvz/Bc0U9zGO5h63uoqMenuFfmhBEX4ExUGa6cztV/rkaEzXgROpj9
lDQKtKZ4QaX3h2oULjllrkPR8T7unDqHAow5zFtwgVYHmEhvzq6vGV9nj5XAUAuy
XoY1zHbp2KIXsJ/mHzlpYXg5BBZctMK/Ikf8SEJz7yioRmwvkph7PlYz37jxuWw4
0Lf7s8eePzSgEj2pwn5cNg64BgDuOYd8+LsmmXno1alwMnLPtHtSOpddosK4pdFl
yI/cO2o9q/qfQw8Rj8dCn6XLGRA5NYROkEz8XxiXJsHVz1hIaRvyVAanlx0c97SG
LI4M5iQatIpLnp69ndUsPxK237D0Ibi2RbXDwjfHwv+yg8pg1/2q6fNdc5MBeTb0
PACeVNFrNyqZG/uAtoMnkON6AQJTJzSGVm9tYni6a+z9WkehLEEOK2yzu+D/Ues5
ouSJx/WOXpnT/7E2nAfULQVSuCZP1B6ORzL1A5DHkpb8k/c5MS67DND/ExpFSW/K
QW6QBTHPaMXJfEFGAXwqsDzV8WKDDZkqSBdtWYa2NgZmBktmXc+i3pqm79NNxvq8
dRtLUK+1NElwpLr5AuixTvpU6t/1299lEvUuDJO/WSRLo5HWiESgOcAzH9eCOOvw
kqbuh881wav2cpx/6KaPtLVvEdKTXNEKgINInmqra3Hc1RDCvsTqhoJ7sidfD6C0
+pacnryLGzCEEHdmqafPi4tHNgFs/OgwxwS3IcrAC61VLC7kfJuvzSY6NbSzcpmj
KoztpJAKgdtZf+S7cAFy90cy1/loicBbw5MmZisRGnzOT+gvUwR0JqGRv8M4it+Z
Q12zds//v1eG5JB3TRJzTJiR9dhz1CjUEVNLOncbK6zcWMed6JRMdvxaEycmeriT
vOIBoqXIztTSiJ6mXlv1hzXlAeMAV3QuoKhNVdoyKiNpOqSgFNRlHta7MjrLrakr
52+fk+O1QMUdCM7Jop2S23+oLclthioNqjZBTLyF7soTzj/lFeC+EENg5bd1+1OD
ZrLgzRNOBmwhQNffwTKY2+KrZegEMSMSDTPN/mnna3Qro3f/l+33XoS7JLfWjig6
Tso2I9XDwLHE8i56ynoBM904XfUD8XsbZkOcsxJTZrjE3bP3/mNa/iU1ruXtBvo+
03O7pGH4bMh5eZMiwLbB1iP7wC0ttnsLnvwRZXMOlpl96uNPugo13/zH5ocIu2TB
po3Q3V5IYBHUWazxDPPVxdud4OY0qub3GDDITr4f/TSiTRIxOK1DIJfK9ol5BEYY
VwEoyjc3TXSbp6hKu4AheyTPmU+UsmDczrSZmwyaJMMMiZlBS5gaMbHw5XN8b8Ms
R3KgQt9lDmEdR6ahOXfmQLVc8nuyEACIcBau6+gCIF2i6ShP+2T4jlt2RtXehXWy
wXOtEAViE1ETFKyL+cptrFCoYbY0YrliU3bFl0YhE6XiD/L7LBF6JUe4+JmYBDCM
3keltCHs3wd5SaXbh5XYEvibf27LKB9nd8z2aGxFy999I7PPJ6Wr0XY4kiqTTVQN
h01jeKSqxfnkhJTBHhp9N6pvQWs3KePd1iacUbVbqrnNJBQ++ZqOrVqFs18fwGLx
6gbQIsw+XNQdOHmNj31wkIbaZCNJSyeSPYvFPB5Qsm54ffzyswMxG4G0ev5L6zMZ
85N+roiavCf9IZqmoAr00Gx/bMUVV/cmflGR0jbumQoXqYqwlhupDR/HYC0CssRU
HYNRvMFDC3vFBmyNzXNxpuHhspFMvJXGiwxUbUmBNqrY37SfiACNTcC+o37Jt3lz
QvO5DTLTYyvGLUAu67iXuLGoYbnRq9QRcHmoC9NAoOUxXfhXJ9nF7/LjDtCMwKUx
7bfAfHy/xYcCQ+VPKuUXLrm72ua75GcGLp5vlM1qwGittMBsVduASO4vf6dRQ2lE
z1Vc0UUuQGSmr29ut8hlZu1+DzYuIeNGeDA3XkbvRIG2bALDjBp97crJYtEs04aC
rTkzkLNpaeBlOLplPjUSUMLL2weEAhvaaZJ59RKQh4s4B/iOZFmYA7NLjqsWWN/M
9M/0Hns98ER+Mbe7RIuxnjDX4bNXDN04Gz2I8Hta+OoeLswKwzDXUPdad9345Q++
8LGH7vyLfnEUGLSDP0lLUI3fsaca+ZtVxADMoxddb+IBLxKjj5RNwQ7IiTW+PHeF
P5E8VfKeNcGRW/ZXFJnpY6Ektmhk356iC8v+ebwZPVTYZ4a66qKuN5WNIqKcarqx
IHsE/kaeBdvUnY+qgTbqEPFQPQevBEoN/JcIGM9lXhVec0DI2xJNT6jOT2Xhzqr4
+is6WJNLIeo3T4h4mxaMj2LxhlO9uZnzwoB8yU8/IBmyIm5Qq58Coy3uMKWnWCr0
8BWomr31VZqPqnusCQT5YPEVZGYx81P7wCfuA5RW8VvB7+rRU1bq6coGBZxDh5WE
jVKwWnVmscwblQNDqjiMb8T9pSVxokH0yklAeuGBXnFgjP94uxomUZ853VYDBkzh
Vjj7HxoU0ugc19/L4+0woKBiMXkPfv9DAP5aDVvmgVntoP2+V6ad1jbZQs6Q4oLp
3RIVyYf65Ty/1MXJgqWz2C2i6+GS+q8vLqRSdVaFwtrRDBYu1mWlDwthEn9KIvFN
Oz81R55b27mJPANB+/cwKhHZM/3ty0eSYIe78cX2dDtP8f7xNSR4b3N5EthF9kLz
ZwHGa2VInVzUU0sSEtUDRUucAEKnmx9GK3qSWoIAD5m6X7mok8L2JK8Q17bgLsxU
q0D8+xGbr30YChKL0PnkjO1eimtxxDIoOP5zKbDmMyyBZX7j9g8akM1RakOCjpgs
mpCod3tGrsyJWo0n9VqlRe0jBTh7cDnO+aclOc/7egi2ainW9TeWhlK9fdSNmVp0
pzotwHodvjkxyAXpADuZXHlRyi68hs4ekTWWfrjhQXpM9zb+gNNl5nLzACQFnkmn
avu+sv50qyCleoU457ywTU+lr+NKybF7vDAv3D0wOL2iA7+hkEJPq6n7Vjtbcxjt
tE2cL0/m8uATGAKN+fmlLxAKaWnj9XQAUqUspap9OdzpZNQUzqNSqDjEEl428mTS
L5rQ3350s1WDtN2WqoIfextRQ3Io2YHLzZYQpBtMxjM1Xjmio7mBL2UNFszz7UHw
QADTG2epVLsx4YtYMurpnWr+BGnOsUXeKXo9mJSIMs1tQxm2HXs3yEoquD78n6hD
SDS6tZSqHE8DoIg8jC1N3V2QxjpSKuxbvLizQqzG0SmnemL6JxIy2zF4MlZwh8vk
25M68QYtGeElbdNmKqAf57kvLgRxl/T92+9Kn8T6/CRsmhec8xaXJWL0P9ACcPAy
+Vrw/+tf7AI/dYsggbDED9osics0DOokEzDCdmiPlzo82Td6X+AV/0QiDx4HuzkV
3nf1GTMvUuXhQMzNF3EcbUK6rv91kzxUvYxJLcfPSUaF/++WiUGAzOk00t42f0gp
E8ODY6sYGbMZ3vECKElfo6bSSu1GJmj0AXUDNpGtsT9z5HaYq7X3zHb0yLKvCiIk
z3a+7ewkRmodh4MJpZJ+rm5DK3wUpXEyeWuPJEYy8pB+uOzzioELmbGIP90U0as0
MWoVK5STMEAexqaN+cpKAMCdIsINh489mC8gvD5n08mP3xrijmC1kzM0aAoipx3w
ILfpiqSzjl/QV4iYfsWL7xsY6xpppDxEmZgqjVpgo7lt/L+318TXU4oFGm/xaqU0
Cszgrdn2BFmH/p+3lGN1P5vvolnd3p7M531p+oLm02WrQtARkREAkITGlOM9znOu
wAkMvGDjW+0dYxKSaJ7Qu9qv2u0Sbr+2b8lbg5r8KO6G6ZTgOWW/GWY/xzMU3K+j
KXXQ+0SX8Zx/9OnoGJ6KTIogqfU3nnM6VX0pBgQqzPIDNrfYvYCMvsNQ4kV2LC1M
yO7oMpEmEPXlIbsqJ7M/30/OM6EarTuVEKPal4UotRnMJeVKaYqhLuTW/TRRt0M7
zNw6HY/ARpw8BkuCsvctTofHT0DGvr+ngyqN1nvoM4E2W5B2Rgl0/0YlV2WnSiBD
MTjhW3fxE2U59J0+LhowCbBHsN6z8LdoljpKmAziyPDU1h999CFHNxZf7evrHdue
r4hwCxRVTTxKPILMUJs0Z0/sf4Z3g/SjP3hsJkBq9Z3J+sB/akD++HczleZNMODN
sFPt4RpMd1HR7ZW7kpFSNxf+aloS6F4mQ9ukcDA7RkPfaRYLuYGPIaZb6sBRN+rE
1QqoZpvIhZNPMsu7a1eqxFA2/GROITtXANZV6PUC0IvnbQuiNepCbKOCgjzKImvb
I2VXEboNed7lxOwd34fT9OB/WHzW8zhj7Qy2xOlZP6uMLcxMIsHbcyd3UaDxZtem
YZwoLl6he5FQL0d85zKn79J83A82SrtIzKe0yrX6dB2jaeai9fCSk+7BLTns3wsG
o4mUGIklkJRUjoLt3MvJPMyDPUJET/xgweLzlIYA03kFmCNOy+o9fZa8BJO6DQDV
7lyvTh41+rWwRMGZhQ/yLTagZ27DeYJZcooQfHg6/TLm7fraL6sctKObFDaDSnQ+
c3iKlEMaanI6TQRVKSd/8c9Cb22GeIDybPTHlzHaBITLPh8Kf9p6wLOLBVxAXANE
Zjtruv70RFZqUc911Lj37S3DRSOkJJmH4r5nDDf2QhP4PNqZ3sIWy3d+OS77h4IH
Us7rv62nRQ+4ErZCQRNWb1CYZ2d6+VJ/FpPEz9fxXrTsVvrc3tzvJl9xxfqQdcON
UamvHzn2iiNNzHp1Agecy8UrOV18S0nUm/JcNjf4bte6q1PmUVppPcQz3b95Usrg
vHAX8u1Utk16I87ERa1oyh6I/g58/K+XczUjx1bOSy6VsJFWxi40s+z6iJ78/Iyf
CkJzxOnWXrXWT7zrCOU8dw==
`protect END_PROTECTED