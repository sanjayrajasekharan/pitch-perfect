��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x���
����S�M�hkF��1~� Ά�``0Hɿ��b��i�<�1�SzFĐ�48��ch�iIQ���H����:4(c��_V����&��}�w9B
��T#�_qx35t���D��<��R*�E����nK�N���������19N3a7K�0~��!�@ըfG#�=V�[��&@0Xy8�U�N�
�y��I�S���j�kU�,���87��u�:]q�Ƒgh��8�i;�f��ܐWq�Re�R^Y�˒�
�1h��{�%z��1(Q�,1:k��S�pv�p�$�듮Z�����C;�y�A֚��Au��*��1�-�_��e�(� $��d8T4���z"�������0����W���j�Eզ�$f\��W�t�(;�g���u��A�j(���g.��=�kz�7݅cִ10m�OɅ��1YW��F�O�`�,�w#{�iR�{���X%>�w�?U4�re�C�E��C&�i��r0��vf�8�ԫ�ft�cY!h�����Ϸ����q�ׇ��/j�"(@��c������mI�kru��)��2��*��0�r4�������i:3a����-�������g=���\6A9l�6ιB������:p��Y�Y�[*i�29��w_�\�&�h+!�)�v<�}�!&��V� !/��y17�&�ţ�*�Ҕ} �2]�H�,�nV���˻u%x��[�n^j^���XԞ:��
v�9Q�����3.O?����Խ��@��5�RlCN=ۛR�J�%���oP���'�̐Ӓ�J�嫃C�EIg,�	кOY�y�f�����{I��xBE��e�[��a����-���;_4 �R�y�D7f3�ݛ���N�v��{,��ı�2°K�ui��:K���5rp�FJ�Z �ca�v����Ӟ�onHa_D�ޜ>��SD̈́E�8��>n�X��Y8|���"�UҚ�sq��x/?l��$z~և��NU
�[�I�I,? [���RN�zZ|mc���LM*JHOe	�WH</=<>m�hD98@@�b/ iD���z��$���o�o^��~po���;G����<�>���5ؤ�?)�ܲ^ʶ6�����P�9|����_�E�+�3P�F��0�w��XBȀ��>kH�%��C	)8� ���2�����Z�`�3�;$�sQR��_��]Z	Q͋ZY=�kNC��o���a���a��9*����� ��n�t-!��ǩ��*��qn�*��.�j�+�2�D!��!v@N����-k��b�T\?��{��w���,;a �b��1��'e,j�y+���9^��r`/P���*��ǒ�2l�c+��F`���v��!�����t�s�̺�0��@�������N٠��KN�͢I��}����/{��ܵ����2��	�E�y�� ���WDV>3e0/R��;H�U4*�´jf2�aJ�I�X���=16z�<MX����N�d�C�g��&��ӟ����l\��y��Ϫ(�Z�\6�'��8�ߋW+SV�+&Dw�)#"(�����Cg�m��Sm����w�����?L�n۶R�q˕�w����#��?������j�yB-�Z`�jү3�r\�B�;�A��L���څ<���%uCB���¤F�'��ֆ��K�I^+���P�v��-7M������z��@��5����mQ�aT��N�H@l�A/�?�B����Aa�+f�����𵂬ԩ�4�>�r�����(���M��M+���8
l�?^���`����P#����_�����X�v�N]��bI4��'��`,IA�K��?�3$�_̺��7�!/(��0��`J�\�H�/�XWeS�3\��q�0����;t�o�}����1i�`�f�H��M��b�'�d����8
i�0��&n$w��o�F���ތ m��D��x��!6�l�T�(;�H�.耶p��HK��$����q����X�r\�����S5gO/���q~[��B�º�X�.a��i�^4z�Kv8ã��M�a2�6�8*�(C�fע|�2N�C�k0?��y`��$?DgJ��8�4D���?�<:���aֹ�d�0'繦�M�q뀡�~�ZAZɑK4l��SNp����	~2�Md�|{��>�=���h;�E���%n'������� �-k��o��'ڍ�#�:�Y�&n\':>@�7.�N�	�Z���=B�5o,k[��]��Cx��psS)�PE�t��z���
���������7"w6I�����)"�ڹ]|"�� ��r��);e�T�`��@����Hh�3��E�N�{mn�q�-�⒧��<�.�Ip�oV�)b�ͣ��׆4]�!T�QM����Ji���j7!u��L�y��Bd��^jO"~+�a�.�]��8��yta���WsVt�R]��=�l�^0KW<�_#��O{nᶲ�Z�y�7a�8�IKI���������)��m?�Q踨�k%I�yF��ji�H^�t27�%�9'gx�:�pR7Y�:P���[� b(�%�[���>[�q^AyL"��S�9�_ Vܶ_y��,�s	C��r��6���!۽�~~�������7ˁy�(�>J81L;�n�\�؜w��M6���~��^��W* ։���k0�,b ��,܈��b�O<^��P�AP�я+�b�_JO]����]��Paxk�U��2�|	�x��_7+D�cg�g�ǒ�������.Տ���������N..?��ss4i��uT.�!|p�-�N���}`'���&�ep�hA3��s�]��ʽ��&e�����R��[�jR����tzRB�9���-N�wGɚ�?�ZF|�|Պ}H��/��W�>��=�aPBڿgs�>�d�T��zD�ېG���א���끵��auGm{�w�D��I��^9KpMQ]�l�<l�ؔC>4d��r�.Zˊ�n��+�(_!	�� �-���t�\y���-ݠC濒�
��������+O��/��2|�le�΃��e��iT�fl�%�Dx�C�p�d�v�홥�`�,�p8_h�_a=e���l�j�0� b��M^��צ�A���W������������:�.J#CP����J��+(�k�p�-�a#�Φ>�J:�8�M��&�9��:�|����ֶv¯y�}2i���={QA`ײB�q�vR�X+�3� z�J�}yٌ������[4���02�!p�k�F��҉kS��[����JA�$����&lT���^�:G	��a��C�\Z�[�Ny���o��N?�}|dN��ėZ�P��TJN�A*�Ɉ�²���H?����i��6��R1��q�Q_�P��. �/��l����X���+�=>�a:�� |�4�tAq��o"A�:�@���1���uZ2��5��P >���B�<3��"����]�;���W�������Vnq`���
�d6��b��
�B��v��$Z��P��S��t�B��1��Spy�fQŷh������1D�$i�>
�i�����P�ۃa����%-$�i{㊜����R��Xŝ<��&�AU�~��y@+l�cZ�0,�v��ĺ'��Ƣ�����Q1|y���3e����i%�S�~���Q�]�Iy	�����(k�q��g�c1��~��nU�	Q���ӋւH,T<�a��V�M�I��6�ҧc'�D���i>�*Y#��U�G����05�Ͷ׼ֵiK{I���0�NZ�cS���5־�8��S]yw��<��wp�=��aq�Τ���n��[� +� ���Ah\n��o�x�o.��Y�|
ʑ7�J�����ڇT����%��
���l.���p"5�wq�i6�/�YԎ��6HҬkl��?!+C��n��G؀ˣ�U�&\�}v2�n@��hX�j⢻����0��W	��)O�p�J��ւۺ��\�����8�[�^�H�Q�ܲ�����}����������(�7h(a��k�Ju�&�7�!�SÄӢ���[���t�93�������_,!-]��nf3�<&�c��6��k�ێ��\Akf�AZP����=��9Z*'r.E4{qV͟�@܆�f_.mh����L	��>���}w�$�
V1�l�3���[E�h��Z�%TV�Ӳp��ݗ�\�jf4ڜqf,B���R���
�ǍJy�]E��R*�-n.6�%�$r���I��Ár��f��opɭ�sC�0ޡ^�пIO�������K=c�e�Rd����jB�(�-S�%�AR$wx�����-�U�(�ߞ���� ��O>��61zI0D�U�v�M�0LM��+>g_o|_&&J̙ $�5��fR1��5������>����q���*�g\�p�PJI3�@��&������v٧]1��20�u��k���Xr=����V5��i���$��S�&m����:t|� ��=)J�z���\���"��Ccz��ߒ#0�ƶw5��`df�t�Gk'���b��@����jV�����\�H3�����R�	R�W�ݒw=�/"�S�9����L�9Wiy�h�h�G#0�4��Q�S��y���^��/A��3��p�o��hM<�\���{>\w�|DJU����ُ�4H7�'�bu�*�[�5��� dS��;��ކ�Y,�������U�o���$T^x�VPU�-��%#��>g��������\��B��p�!=�/�X�gWH�]c	��3r�>BNH�yK҂��nHs�.~-Ŷ�YE�i�S�~���ݞ4����/v�;���%�-Z6��p��!v���	4��Y,��f�@��B��T��~@5�J`towlD�)g�����}���w�Rp�� `w�;uw�T7ޔ 7�D����)�r`��*l�J���� �6���kK�&)���C���pO��&t��ae0�LȀ�ctI=@��.�Q�I�@�"0�O`�-6\���K"j�x	�T4�[Nv�����VG�8N�,;�{w����
�k��9�kd6�e���/۟ka�G���3˳g��GR��'���8C<`��Z�$I܅��ۉ�-nU��6� ��PN��cJiP�>�^`w(E^��-2Ŋ?b�ib��V㤱v�w��B��?�\�������/8s`H�y�.S;YB�U�.M��A�>G���)L-a�&�qj��d��S<Y�4�E�	�mך���?j;A#�/dD�qIv
'�H|n�5�������&�b-ȿ��	4��8��zRX3�3���d+,t���&>c�MN
�-�?w(<��")P��s\����4p�c��Z�\e;3y0���#��F�/&�?#�T(�aS��lߙG�:|mwء���&3fug���T#�*/;����HS�����*�����h�9kMO�ar�#��L#�`��o���S�f����f�ms��1�ݶ�CqH�,:jȝ[�Z1I���#O�b������,ٌ����_�2e�P\�1��.	 �N�cz?���
�V���B0���OH��!A�#��ku3�2"#L6:�E(�ۑ1�{���ÝLDj��7fB5j�b�D��5K���9R���`c�q���<�Zod�B"U�p��{��a�~�������K�ʙ�)xʄ2Ϭ��E��aܵ���������k��Gѵ��u{�#���m � ��PU�C�S�ΐxd�� b}�ְ�D��Hm����1X����u�6[ ���� �}�@=���%k���7��y���awC/�.�	�3.Y@��ND���jL<�La�e���I��T � �'�
��$�Z���jFj���]�7�ޠ�=��깵�'���99��]W�����eU��s�xϮ�j�𹴷D%�S�O
'�ʣJ�^%�ؑ9���v�R�b��g'>M�`��6)�ڨ��}4�����a_��^�ج�&�d��ݚO-����i\@u(#�;$�ł��.��j�H�Q�/��^���eI���Ϲ��}�ē��4��V����I������Q�Ȥ�&߼��(pD�&:uN]Y����S&�:s� ʄ�CwR��xku0��A���(*xգC�iމ��QƁ�D�g�COK�v�W�"|2I�����ٸK��_F�����D�hE��-L,$b?5H�4b����1zm�����b{�/7g�Qs��������W��ծ��
�-�]�c���/}��"�?s�E1�w�����؛2�U�� �Z�?��y��@2��%r���#u�'Lה7X��m]�u��h*���ZvO3��Xy�x� �Ǡ��|g�
gǳ�kv���qeB�����a�����rpF[�M���x����e(%��¨N�%ٺ/�P�kèn9� �x�����T0�Nt�H��1�.�BJ=�0U�(?�T�o},S24�����a�N{��ڈ):R�,o�� i�c��r�}��-�^:�P~6�i�x�)����6T�T���q2��l��m�R����mh�t�;h�[v�A���8�L���7#\����u�Қ$ѱ"�PJ�:��ꥋ�Z[���^�v/�m��<�X��W��Y�B��J� %i0�,�>x_�H�R]��l8|}�~{v9"l`��;W����A�
��5�i V-9��?��_�~?�Rsr00Yf�Ľ�EO��  ed<��8�k�`�Al�{�Ž�'��A�[�vA��㭩;<����]Fo��O��F����5¢L��TX�In�9\�K�Rf1��fr��b��G�S��~�O�;�8K�}t���f������fut�(*ް+_8��s��䟮T��"w�����L�?4�e��$�6�by�D�6{]�c�����>ߧ�)�����|�kCScۼ�DKdi�$��$�p��B-�do1���*�/΄��$�,�Ni�	R`i�z��%A��������ĽJo52;���8e�-�3�Es��Z�\:�.dH�ci�(���R�۶�ap�'}'
2au;�R}�O�P⛚�f9$�:a&gb1=�׮���iWd�:P+x��; ɺ5�Q�}���\O��l��/��(L��,�mW�"��0c#SE��B}��Dtu�@��!�\U��&�=M��N%@2rOA)n�ե�v�S��,���f�Ū��!d8?��O��M�*�jK���_e�=Eȴ@�	�~57IM��a$Ҕk�L��<���VLo�^���l�_q'A�?w�K��HƯ����-i	y�ִ���
�Né�#]��<G��HD�'����X�	��i�� �jk�Y��r�r�λ��L�]u��w����������9��eg�%���Fhґ�4�����N�0g��q��Q���.�+$�p�����,
bj��P9�%.��	 ����|�w,I�Y_���� .�F0�*%����&�߽���<�V�<�g�xb@%�z�4�� >2�Xh;���d{��~^bi�]��t	j���/ ��0��a'd.Ν�K������d�m?�4�5X�W��pyT��:��ǦS��:��%U���������R�yۡK'8����։���݊MbZk�nqj]���H*[t#�f�}��.u(G�i����x�M��3| g�30�^ɗ�s�X�J�t
��Ud�*��Q�V[;"�/�#�dF �
��i���E�>Oߢ����sv�Ӡ�;E�B����f(���ܤ[hTo.R7�j���*M*��c#������E�jHUC��6�	#��t����	�P�<C��U�,w,[!9�-ݮ'�)� uu�5;@�g��`�
���ǛҊ���;i�F���;��$Zw~�ǲ暽��[z�z��։�	�Ϊ��Q)���v�SU�����B j���zߟL�5�3�����1�]�����؂����K�U���;2"�nh�5{�*��Ì�����ے:�6mg���U��&/�+��8��qD#"�Q u���N�؊��wXs���f��}ó������w�?�qd�||��D_��]���PQ8�^��*�1Ũ�!5�����Ʊh���.�z�Ī#_jsPKY�����g� #+w�k�O�Sª�CmX�J���
fI��z0�o�|�
.G�	t�r�"n����L��lDd& ~	58��X����-�D�n���qI�k<��P$�XQ�«�q���7k����$�ŕ�ܶD �ʺc���bֳ�0���4�[�9
bݡ�����t�g�㘃���|��W@M�3��*M��x�K�m�����[� ���x�.�b�
�\����c��[}������Fɩ��V�Q���$�H�i�?�����NTG�pkAt� ����L��/��Ŭ��O�&�
�0�ލ.�D��;z�-�����vn�y�>�m)a��������ޞ�$^�f/r��P	���VA"���A���߮s�DcIU���6�L�^� [` #�E�m� L�8BkW���vV�L��~Y/`R
%�x��<���ge_Gn�U�<g�!�R��Ƥ8�'ۻ�5�N�v�?jwb2�ȝ�����(Ұ%�Id1Q��0y2�%���'�}�x�[��,��}}6ˑ��K�ʣ��!��T4<��|Ts�L��zQ��G�thr�!]��~Ѓ��P�lLoW��X(w"=�BsQs��N��0��a4��\���雞P�XE�1����b?����7�m��;���/d ��ݮ�#�dG��6_e��7Ua0FM���YR��Z�#��z8�Ӕ��~����ˑȡh
�Ь�lƯ�@�+�0yE� c:ny��i-��
+�cA��-aɹAY��E0�@'�����G~�=���t��:��Tv�p�z.׊`}K��~�p�,�����$���d�����$U��Ky�"�[����]bC��5�WB��0 ������1D�|�ם�Q�Lf�T9��!��WclEE<�u�r��1!�Z��S�XۯM�0��&���J��,d��cu^�Q��ʈ��ia�����3�u]��<����rW/�HC�U��˓^��|��<�F�����ӑ�/��������O��-��0	-��OR���h��!�� �R;����8c5����k��W�M�uOGcwq�5���4��|�gW&����K���\�f��D�v���v�x:�3*[��~�K�+&y�C��R^4��[;����揂�ZV?�{�O\q0=^��l���M�����5R�J���3�����U޿�e�)�<��[.2�zO��A��k5)q��t@��u�A/�m���	C&]Z�.gz�s�)*���� WU�2i'�}C_�پ,..�h�o?c+��I�
�r1�Z?Z͆�#�z�T4��3��Gڔ܇�M����#���E#�°Bq-k4�T��|�[8KT�[�Pa�2���Ԓ=�s)����!��:P�,�[^�a@gu�=�J��<�r{�^6ݵ�?��8I�ƹN5��k=#u܅�A�p_� �TA$�E<���\�v�MM�7�$�\�x-��Ú1V&�z~̹�X9��o���צH� ��Eq#��&�����?J�z�W�g
����%��H��X�����y#?�:*Ky�B=��Uo����w�P�9���7�U��W�D��瀨���l6��:�"~��
2ݓ���s�N��q�R�*�3�#{a���t�@Xa�]�O�o��Nf2�Q׉̪�(-���������=G��D{[�Ì�}���X8Q`��m�����G'~����JLCK�8a{���O;�3� Y>��BD�I����`y^�}8�q\������s��m%>����Y�ӊ�53�?v�j�]�!�I�aӫ#u���e9؉V�����V`��߮��r�K�e?s�HK	J+j�VN�s0#׵.ׯ���Q�|[åMkI%��_?�簧�
�)��T�g�e�O��u����4�΅W��`M����If<�&e}�ȇ)�8h�e�αL���`��/]����d�iQ5J�������ӗ�t�)���12�G$o��:�3�f��T��C�Dfd���q�G����w�
E�q#�ڛv�G(��3���'<���_E6Un/RG}$����7�Mܾ�<���e��Ҳ���"t/#�Mu��$�4_d�$�?�|őR^8x��uX��ٱ��G7�?�@@�j���W.cf��j���v�ۄY��<������+���[�M.I�F>�=�l��:R�-�m���y��>�eҏZ��q'��}�P]�Y+�R �`��a�q����z=��C�P����G�����ޥ�9����^H�]Q@BȰK��"�GH���&�`�D���t}���9P�e`>T���۝6�.�+R� �i�%�{0v�&dC�WKYZ��u��y$�3�[#�<�qUÉ"28 � �obת���'K.��γt�����qOA�N ��ɸ��m蘘p�D��%���oa��\e�q=4�ȷ���@q!�����|¸N���F۹��S�Gm}%����,-ǁ�[qҘ�:�0�pd�t4<Bת���H{��kT��f7S�Si^��	A��+�@h!��|�&�M~O.˖�ǝr��DaiiݐG�����'1;նD�M�-�����1�*����T�>Nc!��i�m.��4dJ���i������C*D�R��a�A��.SEث)Mވ���Xub���RQ%̆
K9ܤ�:6�U�6����3� a0��X*Rc<�=�Z=��:G]��.Ζz�C\��p���2���D�c�@w�z�@M�^�-g/�&O�������>�������@`jϪ�^3��{�5��?�m0�12�5���[���ul�?z�Q=��RJ�ź�Ն�1�28����+PKS� ��o�>�i�췼A�'��H+� k�,���l8AJ��s�X(�o��:p<ӱl˛��Ѳ#t�+d"/���Y�F[��Wd��P9D�fVa�r�g~��Ҥ	*9��F)a��ț�N ����P�LF)
U@��o��3B��w����'4�ܑ��}~�f�J ���&`�mQ�^F5&y��`��$�d_.����87��TX��9 ���Sm�)�g�����3�H�\��7J5WtIP�PF��hMN(�5���)�J��E�Ç59��~[k�Ie?_�m�L�@d�3�=�:��d���\��\�Դ��ɘ��j�O��#/`}{�۵�9�R�B���xtc��X�&����q�{.ړ�[��׹��^_X����֢�J��@����H���t��Vi�6{��ak�(�6=���Tď�8!C�ˀ�a=R�0p�JfQ���jMg�a�6�+R��ճ�1�S��I�Zũ��FP� Y�"��ˍ�u��mG{\���������z��RS�V��o�-]��1�p�0eB�)_��3*�$�b�;~u���g%\,>cߣm��ط?������!*�S�Q�aR�A،���&��Dـp�F�@5�����JX��6��Ux��p�=Ŋ���"�Wk���2U��$�$�ݴ,��Ȧ�,(�&�h�y*Is
L������=w��s+���S2u�6������b;���IE�G�r��T7�v*M,q��	
!�a�����M�f�?��r�T�(s7�D	J�����m��zh[�CJE\����l��y˶�`����R����Bҏj$�;���a|���W3�AX��7��7 Yh����?$|p�-?��#6���	�Z��OH����ܥ�%X������#J������-�	<i	�(BW^^�ɿpU�Rş�M��hojWߥ��	��F�}��r�?���ǐ��0�	�U�z�=,�V�>�DR�S�\�����c.D�k&y�;���i�+�'/��x'����5��̷�!T�*�
o9.MD�G�!¾�1�t��G&�E X�+���~b�i}M|u�}ռZ�͂B۹�1�Ҋ�E�"{�#H����Ӂ�(~��A%o�z	8o��<su�4==cĒ"�����m�\x��M��9��T��wZ���Y�c�ׅZ�s:�ڔr����#��n�Y����l�{�$ءKCiQ�"�j�:+���wo����A���D�$����N���m��{�Hf��6I�ґ_槝�,���YP�랿�UFlr��Q�J 1=�صb�U�XPN�V{C��k��9e᳖*j���-)�����B��xU�DXl�E\���iEh��0Cܚ@\q^�Z�GRA�'¨kY��u'����~���5��!�J��˝�
�Yկ/"��1���H�r��)�թg��b0�`�\�D�;R�2<�ռ��%u�����)�N��[����Ӌ�o������m�E�	Uuذy�>{�v�g��l���d�ӿ٦A4�t�#�T��bǇ�2�a۳��aM#>��[t	�Vb�;�9����C`�W܈��AQ�#V�BcF�t�2�$5�
�5k��pV��j���-o��yп�p���׵�>�����\�����^�c{tM:.�S2�|a�X�įxhQJ|�R���f
~F�D�����a���`FN	�

��Ƥ�15���k:d��	�g�.׾�K�����9"��� ��z^���pl��C�
���W�Z����#����T��K@*�0�mD�0d�>Hd��|o4G90a`� ��ٔ�k6��{�����m�0�C��=�X�+oᘱ��֌u�+]g�) ɸ���2m�'�1�o1!ַk���Z�,��xz�{�G�F&Gt��IHR	}��Ք�e�����Tb��.{�IV�b=L ��ݝ�J����J���X��o!��E:f`5�:��I�.��	�gc�&9 � ы���o�P�e����oF���F~�CY�~�9'"�8��6�@��7�{&���ު��A���Q��Mq�ċ��F4>/=Q�������G)�#��f�^:G��?�'���#��s^q��-��=����e�tb5GUT������	?��|�]��`^�����?� �Ls����C(E:,���MZ�wP��+���Jm��k�(:��.��̾	��t!��r���Y�בz𛝂>Q	 ���5��˅���7m����TԆ�T��@e�R_[�q>�o�
?�%I�QX��*S��s��#�P8nFjh.զ���L��%�BqEЫ���^��I��qY�z�����.��[�	N����_u�(���������A�}b�?S^~r«������vjw#!���b��D��d�#HN�b���i��GnV6�'��9�|�E��Q��L�Ql{�E�!,�_7�q�l��y} S��8����/����/��~r�;�Oq�q��DI�l(}Cmx�N�"z��!�Z�mM$ۓ���T]�s$�Ǩ�0�n�P�;�Ns�W��LL��v�r�̹�Ru�a;_����ˠ�X	*U�
�u���4^7{e����훵^���\��OˡͱH/��\ʢ�ѧ ���5��%x��LS��s��d �H�z��,{ʜ�Qm�Ef�φ�:�+�}�@����B ܅LX�W*����l-c��OX�J4�K^��]>�������)*�{!uҍ���	{��*RVX��D4�[���/���N��Q�&y�l��ޱ�$�a9D�<��*���a���.*��6��Y�&�<��6�?�nu��J�+BU�� �׵�2܃�P�߻m�X�}��u���f7��q�n	8D˚��p�
���G/���������XK�߂�,E���T��V})�H�QQ|:�s�s��W�@�O�~�X���; �S];��6����ꚉ��KCn*Wt���4]���}�f�nPh���v[�HoKC3�?%2	)�M���*�QH�h�Bt�j0�@?uk�D�2���;�>�%9���jMT#%� ���2����1;�����-
η��?���R�7uy���$���F�vй<�Gx�N�_U)�H�ی)6��E~����3�.x���0�6t�jr�Bv������+���v��D���3���+�0���d^���|/���p#.��p�&���礨.��f�`�؍B/5�n��
\�nk#>�(C�8�_�����:a�@�
���E�V#�C�M��04ۖ��
��:�GdLг�x�4�ۺ,'��]'{*��E	q�N�#-�<���M����������F}�߭T-�Ol�`��S(�p�l�Q�h{Y��&�E]�;� P���S����L}cRl��T�� RWM9��~`Ϭ�F:�]�Z���0|�e���/���GQ\{N�a,�@�C���:�]z:�t��@rD�3� ��b��=��Iՠ�^��c�f`v�`m��s��T)Nޏ5�Fc{3]�%��\��N�%�.�&)�u؅���_N_�?��$��y�)pS��+� F;˕w.R�2�!tO���M"�����\��?���͉�*�� %*�,Ɛ�#�@�4��;��u%��#LR��<&`�4��t�ݖm�����4���.�-�@I`Ȑ�}�%B�8�~K��g��BXuvDoa�֖�k$�v�n
FQ�s����J�MeE�L\��c�6QL*�����wY�Kr���7�ee�@�r%"Ķ[~ �Ko��ٝg�d��I{t�V�fD�:B��U!��4="mA�n
<�ĕ ����*�G�[&ldnԭ�G�Q$-�$D*�� ���b��X��6؞z�><n���p���j�;����̟�_��(G�e	��7��Oo T��3A��ş�NP�9��=��RP�w���j���8I��լrK��v�{�<0 z ��Y9��-)��ȡ�Y��������Ab!ܡ�R{�(��)�݀SFS�����0����tp�ݖn�"��SﱞI09؃ӹ�Ԑ��oY�EM?��zv���~��U�UTXa�y�4��G+I��[�s�إQ�x��R(~����4�v_����!$Ҁ�KlL�r�Q��뾯��������닽s���ʆ+Y��X/�B�z�;`�r?�x*�͖r���SYI��/fzzu��x��_�T��M���*�x���}V�ȯ��1���(ʍV?���yP�6^��(G��e�����H�?��|{a������(�;�+��m�Lw�q�c�WڏdĐ랟���>�}�_|k����Ҳ��3�6�Jx��j�&U)ܤBK�\���sI�$pi~�#���By.�2�yh�C��j5l���5y Ń#\5jN[�lf�= i����p��¨l�?����)�l�I��/$4���_5(8[f��sC܉�-3I������BʴOV�w�.��4$�H���6�$G���7S)�z��#����#�f�x-�<��:�
D��I�]�
n����\�b0�v�k]<�-w�s��}���sP���s�9��7���i���Y�?�X�n"(�F��|��S�y�=����OF����?�
�f{���Q�8`d��dgh�}hW�g���+�D��9Z'��F�����v���l��m/2w�X�%˯���VX��5w�f��; �*�6[Y��E$�^Er�NzIN*��t��q5��f�����~ͥʁ}Wo-r.q�_��~#Ms�k�%�I,V�؜l���}#�_��c�g&���C�����9�_�i"K�:_Ksމ�8]���w59�����{�f��M�´;V6yE��|!��.�+���_soо�*C���35�KX�nf���2&{r���H&�k/x��+x�\�͎M T������}e�O^�h���=���T�m�v<`jvK2�W�y���g���{F/'W����3Ȅ簔-%���ֈ���*4�R<-���}A�������5�y�\5�Rh�Wl�f�k��m#f(r�y��8�c=f�j��+m�E��q��
����cX����M9U��]8h��F+ʶ�Ա�t~��g�}�I�@�o@z*;D� ���X��+��J� �U�J((����nc㟉|�#r��a|˻H}N�yuW�\�~������ >�̢����p���������{.̏��H�r��b���pC?
����Ni�7��=TFC,Wع+�(f?#F�o�0C����~)��^���'Y{�CԸ���@,��֭�ܾ4�g)ꑝuG#q�Rq��r_{
1T�->m�$�f����o�=�c2�&,F��jx3�:b1�Et�� �9w3�PZ�m���?lW�� 󒼜�b��LW��;�l	�=���F���
�#ƔD�T)����Ɵ��뚒�|�Z��}9�):I�1?�Az��^�N-ז����G�_��K�e���jX�E�.9���b���ӽA��:�4؝�z��8W�/�pi�O��nx�(b��㟿	I����_�wC�t@*��6���}%ç�:�V&a�b��K��!�Ik�iL8�./q�W$_�$9C_�������_�ƻ�1��������_��	���n8t�ǩ�1��W	��*�ЙҦ��N��W��,�b�6l�����3���j����/%�x��� �L�23�������u}#��ӺwCk�?���e�W���2��!�Jlv���_w��Sv#�̽c�Q�+�I �k�yq\5�IW�f�]^R��й����kZ��
��0]�(@���&-n�YM3�f��MSa��]H$aT�r�X��_�!BKv����#ե�9��9'��PW����䠽�vj5a"��wSyM�����|3� P��E���hG��$a��m���ͥ������k�L3��xLM�[�t����Kl���W���?�w+ȫgQ�TL����R���>�u��.Jifȧ����^?��	�*����m���f&kE�mn���B�%��|��L�#�f�kz�<aӭ��=��ݎA)sO��62����u0�iZGyAݼ�Z�(�%80{}��#�ժ�|S��%�O8���*�J#wLb�6ʴ�hZő��#�&./���JُT����z��m��ۣ_�A�l��PWZ��-�j��H��T��U�)�����V��+wv'����4
�΋נa���kK�5��09d37�/,:��bV��A���>|��acF����ڳB�o�}��jr�bXp��m̑��o���!�����]��&(��bss *I�� ��N�?�c݉�!��e���N�|����I=[����{� yms��$d�d��+��Q����l�����B$��Ac�������!]�&~8�&K���	����t����#�9ͅ�b,p�͋!��`"8�K��!���c�8Y��
'6�Mq�j��F��wv9c�6߄N�N�{���.[!!���}q:��6�,n��Ll��ʎm�q����ST:S��9�u4Jʞ�Fw "�ߵH���M&H"�R4P����-?����C����F�z�gNDp^9�%.��_�A�a�|�5I�)�v}�l-A�=R��3�I=�z�S��m�`����&���/OY�q���s6�C��go���0���*=2�g��y�����Dv.�uYZ��G�� ]Sڒ�x���Ϯ�o�lES��9^�@9�#��r{��G.��L�z����J��C��&UVz����~����$�����Q:���H̀�)�Oԃ��K�t��q�)|������G�����d��Iud".�X���Y�-GdOt��;�5Iy�;d��(��R�1����:w���=��}�$����c��Ҫ�6�O<e���C\�p�R�QX2W�P5�����^wwV��Φ����;����t������)���.'��7f kp�u,+�!�
�X"@�}����}&���y9��9�x'�S�?���N��P	k�3���;R��T�B��C��R�^�o�U�,���\ݦ�6R^;�-f��Q|�0Z�βy�soVSBO��{��n�G)l)���,/�����A����g��pehSw@~�u�&I���>��g�H�ֻBDH�pz1�nă(�.3�L�v��˫Lu(��T��Q�ul��Jʷ�6Y��%�?�*�15�3�Q+W�{/����E�₥���=3!1"��*���Z��N�k��Uݰ��$F��pȤ�e��s��|�b{3T� �Sѱ=8y��89����o��}"p��,�4��c����𥪽N�642e�#��+�`����K�\����b,������V���P_����K�&�ڭ{���v"cC&*�Zܠ �]��!d��]����Z9���>E_�l��B�D���P�rs���|�B�D��D{hh� G��`q��}а�{6��6����E���3����tKqW��@��Zf�����6u%j�Yr���b�Τ��r!`�Se"f�׋B3Y$�O�R�ӪʻP}����)n�2z��:�Z�Aآ-���)���ͭL�3�q㰯ۇ�b���*�oJV�ZG�	�w"�ߨ>oʃ����	�P�7/�?�7�@�o9�4����׽��qk(�~����o.�p����J���[�\���?��_������{,��A�v9��`̡��޳Z䘇6�t9jd�{8�($B|S^/��NU}��/Z���ڃ!/��&�ʖqf䵂��F-|	�u�u�R�7.�E]E
�:l��0����7Ug�;1L/%(�-mȵ��`�2E�
eD���U��͊����Oz�oSM�+��~*�J�%�߸m�Jqf�}_�"CRR �L%�,�6=)H=7�a�1���︵f5�k����˺"�4�*��`�e8�|�|Àk�_�aY�֠�>s���_�\��E٠�����"�C�3�|��C~w
��^�SK[ôP	־�ƺ͈lɌ�w]�����"z:C`7�Q�h����Go��7L΃u�s߄
���x����N��mp�5��>��|�=�9�UE�H�޲���=�eX���%<ܓ?���n�*��.�.���_mLf{7�\S���K�}��W� ��3뒰gw�[��^�l���G��TT\8����2ǖݨ �a�d
�c�GJ�Lؙf�i��U��)�DhP�F��-���OOE<�a�1�&[�]�!-��:���A��Z� ����`�B�
U^~�-EW�2��7V���'�M�Ѵ��z�=U�1f�0~�N��$ z���QR�i%kC�Q�x����gS�ͩC|ً���= Z֣�Y��!ăj�m�+�� ���? y���}4`�8�B�}��4��I/ �����<���40i~C��U�&��P�0�$PX(�C�M�v�� @dJ�>�aQ�+n��ʿJk��3��VI�VZc�M<��V~|���f�鹶T�|�-��K��WOI�бW�;��Ŭ��|u4h��cX�_0��F{´B�Fu���MrF\�����pǀ��KZ�}�]rfC	�twQ�s�C��0�;������5���J~��0qV&�:��m�w�;�?H���i�����u摺?No=�����\͘=�;,�����<�X�uGz�e���*�&M�˶�+��PG�t��
���a1��Y�'v�X������+qM�
Ui�G�)���0�3������:�n(�i���� >R&nl�*Sj�����6�����УY�7
߅�����	�{���5J�;�p9�ƶR,��[&ѕA�h1���������ɭ�&���g~�}��]R���<��|s�4/AÇP�/E,��VA��#\5��\����{6>Af-�O��J(��Hb�6c!�2ѳ�^�Z\�{���-�������!&95yw���Aꭁ��!j��#1ԑ^`o����YJQ.{�S'(��}�e���"���?��C�����EOp���%�_~X�����.r�[Nšdd�@��Ot���ߕ9��\0(}���'˽�,��.��Z����x�_;�S9i��tt\�e�!2�m5��%v�_��<���?��Z#���ڲG��$ƪ1t��뽧:�80��2����(Y�|����
 A"{.��e"��H���d�޽F@�i���9#��J�Ҟw?��Vh�<�5n��ӠL	��샢����h}s�ۤ�@+;��G$teDS�sAe�#ak%�*�17�>H$����"����G�>:Z�"�	Ǭ�� �-�M�O&��������AÔz����J�0RC[U���=�ݴ�(�I��\������t1��r��冾?�}�(�S�Y�t
�cY		���̶ϑA�Y ��>n�k6�Z;p�����s�/��χ�B��*�:؞M]��Q�ް�) �4������������?7�����݅�R0:��E�f�&�ۍ(��ܱ4a<�cy�?�rx�̢=O��Hā��b��_�ǣ��(�2�IXO%${�K���G�ҧ&%��FhKIbuv@G+�I�4�1z�TRPE���Gފ�l���ݮT���o3�����8ӌ�u.Ojh2Jr�	���5.���	rH���`��z�?���z8�����oV�BO��@G������v�n��j���Rgl]{�4��H��?�w�Q�Q��k���?�t���Mb������x48.:DX�����>��9n�4���J��l.� G}q�Jt�Y�������Xya�u�W��,�j|<���&cMk�$!*�����%ˇV#Ԇ�OB\�_�Gex�������@�᝺`���>���ňn�5�}~ɱ���y�E�⇗ݭ�WƜ��c�!֬[k�݇"7�y�`?�l��U����piT�xp� �Uw�
���Ϗ��A�O�c���6﮺�4��;�;�b��v�o���Pv��'r��M��CcItv���B��_Rx,��q���t�fn�)��n>}���.�ʾͅX ��=�L���] ]��!�"�6AqT|����eb)۾n��������0S[5�xa�0���sf4T�`[}Ş�1����$r�{�E�5��?�_��^� 圹���S{膼Xj���	RڭP�ڶ���x>ApN
۸L*�<���Yq�͚�@nBE���*R1�����1&zDI*?�n��Xm������92A@�O^	�>G�Ԣ�6��E<11<�Z�M��O�5�v6w�4����MΚ�9�y�R]�Eo��*4�X*��� ���k�]/��X���G���M�VN�W�x*��u�>���9^��eF ����C��"gsV�@��IV�罢��Bלh�E�����@ȿ!� �5�F�YSÏz~7�%�s,&өx�!��Na
��6X�7@RIۈ�1V~Kaf�>ha&������w��3*�2�e���0�0��S��yỲ�Q{�gCꔹu1��q$\^��U�]#	<v�^E�X��ӵ�e�5���4h�dS_`y�&�{��`삡��a*f�m��Tw���˷a��Q*,���S��#�:��h�F����1���`ݵ.�o�H�lmU/s�R懜[BC�H|�E��E�b".�zb��wL҂o���d:�'Y � ��r��McimaA��]`r�v�!�=G_LΔ�4*���9Yp��J��"�۴�6;,{���<�� 
�'!����F�V�ZLs�����~ca�v�o�!p�D����*N���?hհ+�K'�L�����Bn8C� ����ii��%��og�M��8r��zݦ���O�m�R-P9Y��{'��U�P2�Ε��i�ҡ����2��vU�G���,_P�H�O����� �ߤ��[�=B�i`�v*� ѿ_u��dK�(�a^\2�I��?��l��ʅ�jix��>\���S�Ip&='���ЪΠ���ǵ&8p���y�'IC���@ �r#�`ݎΓ���́�wEJ�c��M�R�x@�^�V?Ϻ�k�BH��ÉlY�#w`>G��A��*g?�<�N1�yW.��̡4P4�!+�歎�K �o�����Xti��7s{P�x8��o�v�" <+���QZ��Δ�|��$x�3_[E]l?�O�yR*���U��7��W"�2|܌)�ҭu�����s��L~��.P��	��>��I�A��8��E�6�\��b���~�a7��bYFz>�oٞ�Ƹ?����=��P�!L���.u>S�}9���~.VD�/��MP����yB�W_���0��o8� X�o[� $���'�����b�,�'�!P-����׉T��:_]&���?AG@#��k�7�/6�q|O=D^�`��ya��%�����/�Gh2
Ir�(d���h1i{�E,�8g#��;�r��M�༖��4]�$F&iO��F�ԟ<�G�_[Dw���J9O�L��i��-�n�ƞ�ArsE���ߨo��q,�ò�rZ����p$ p���E�d&�d��ȣ�O������!"pb`��8xٙė�)�Z��8s���&�7�M^����t�+RB�f��K���"���x��ԩ�b���뤹X�����E�������[�>��!5�� c��Ȉ�j�V��Fc�V..�a�P���ض��(�8U���e�Dо�Xbr���X��
�U�?E��{o��8�b����G�v��]�[�/<��78�����>�#��b����\�a}��#��~���Q����a�%�>E,�>D����ذ���rt�P�1�� MWh�1c����u_C���r�$s�t��8����$cC_�>Yr�i�KA�uO�B�}���)��IL��Z�U8��[��c"�)����ao!�jI+���+����С�����y���z�J���˼m9Z��i���n{Du��9�hNT��0q