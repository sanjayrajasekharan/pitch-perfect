-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1rXJF0bwo8jkDzkLQvOhCvmNgpue8SZ3FNQzKXwlLqHbfRjK02xl66FtCo8zcZhh
ACVyLCJXkUKGV7KnKBqVL/dxpWufuhhHPe+3ISUBy0nMDFR4F3URSeo4/UQ189iz
p8z9TlWvgN1tmBvfO+P3mdIw+mGoteCjhtnD4GT5f/4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24704)
`protect data_block
A6kIfvmpkkYPytcsoXf2KVDlWOBl4uBPLTSji6xNvZcKrHH7juvjxeP2hlT9BISL
h/LTMphbHeJV7ehARhJlfhICIoHmFYpXM+5gdnreSMAqNDdH3i6TQNjE2OrpYlNN
gpslRcIZl7V34lQ5LvO3zN5yzqJeaM1FhIgyCJmJkA9oTMEYDHxp8IYNsIiJxxDQ
peu3TGAbbMZsq+eeAfUcEwyaoSd8KPjA7vgQ5q6r063I3UsGHl64z25JDb0T3DZY
TifJFuE2HqzpldYstJNEC9ZVdB1/Qj/51IB+GLCxGZFxzC6d+yKv5k+QPlcCkn47
s+mz63kui9+5R8T7cRiMOxRb9SAvlKoVX4MO6tUntb1sRe5CYOUjKTzfzSKfeioL
6A9yhhJO5JTTgwPEz18HxRPNsoK1YzZFSLHGZcXEh59DOnz/8D1yv0FJvTs8dW7c
FCkhfTWCZBJVqMxEjLiUFgqEQIPAedUVU7fljp/IYOQNtW87j/7Tg5t41cqx0u6f
HdDVMfe4aCJBvqLkMHzXpvZfXknp2jf8AZqHO4WBRdSvB1e48m9ENv3+QNFk37Em
mHE2mwHzMp9saTDrtf5xsuL8C5B3r1ke/BMHSnnlYaRNqQZzZ925Ua9vY3XmALZR
vocWiSZRdoflbz56t/a7X/TQJFM0w8lafbSUeVZ09oiCUXhzOsBTh68+PueUYjV4
/sAtIci11ycR8P0P+xFdd35j+i2/FRI8Q2N6SFAh/dXl5ZafKpsXdKxhtbTXye82
WhwzpEHLEr93BWgk2HiKBbO9JPwoPkaeAQt2y9uJju3QkKCrAuGXaIoubVewhvQu
sU6DQN5wPH45C/LOzmpm/8SwOB/nN/FsQSQDvRKgKLJN7jzP/1ShKoCnmt71OCo8
tpQr3sZWnI5rfs2rOmMyHPLddo2Swk6TSA/D7DUcxhFwgzoEZ4v9hSmtnpMM5bIM
XsOaWyxbt7k0eCSk2lyqMeNfznJGNsvQlG9g3AXYe/ip/do8lWvA7YRZkGkI9vJN
69hsWd+7ZHT5X4Yp5UhLb3fyPQxzAjB2IiaLMYCK8qvj8a/tJb8V4v2g3e1I/J/H
N20DZlR88ZSbUSgO3seX/9lIhTnaH8Kx7FF2sglpk3AUk8ejm61YOOxIbEcSUEbY
rnrJxVXsGCSJNS+P7/3xl40UJpAa8nqye/xtA0PHC3eXIT880q6xvsO6J+4mAHxL
ghCMot3LDHrhIy+rvplpMOesntgeCAmoUFURBhNIam6rVfE1KZ7y4aIlk+e+KBxy
+2TOmLLTL2SEpfKt/0er26uFyZ22IxCm4gMcpgNKk9rJB/RyMNw0++ZHyLxsBGCG
VCTEx55+obmHgHL+jyeNpAZpcUWMRf1urEa8bGkC3uPj29FHbwwIkdR9VEhqPBjt
ZO1lETkWRnycBf2fU9XgDGXrgbQo3JNUDjwmDuMrKoMZ48NXWF0pgiA532xq5hV3
2fHYKHLjKJ1+2DuFvTk6cxEB0hlEqx+n2U/+p5DnFMRwBXdJBZ9ORYZo3bA0npnD
PEOTXPItgLnJrfRPC3JIhMyxUTcBlp/r+hj4cRHw+6UXVVq06Wdrjy4xXstC+XED
Xs09VW+5t2RiSVBmImP7cRi3OxDROE0ILSGrg/OZl9nsmPmGnavLJLQe5m3b470M
MG56FmCzx5/4Ag6JXxniwkCYEK/9OyX/Gm43QkSH6Twl4VJd5ha7Q/7JWDhjEEBe
yhcv/a7MEFQSxX/RM9+zHEpKfjmEfpQ2nbFWJBOMoDqhntdrKe75PgfzGriMCZHQ
Y3hDYWrfMRiPsPFUePZ4suINAtbPRm2wXjyjvNta2GUkqkl3I9DS6R1I+j0RK+MX
0tExk4OD+4NGi3M8wNtKnW8ywqyOw9jWpxfuxcDkONHaB3mfS+fZcT+YHJnQxUk1
LtIdlEwPI47Oqv03ayp2ceA1kXixXCCnwaxzCtyh4mPpFK26K22o0aKs97JOcIZE
HQGORz2N/eKkaePhIzHwGoKGiwdq9z5uvwey8Js8zAgRbyb3/hML+hmQphbTE1m9
WQObOV3RLQFOBnl8YphwWi46z7FxB+lXSGVAoz2ncgnReTCtdtpQTS8mw+JTAIL3
91sN/JvXVgdlEet1f98fpiw9W8G32Iu0VStByyoX3Efb6Qgdem9tpi9fnAUYNOu1
R2WNEE3PyGhg3qKs8ulwVyAD2ucAzyZ9h2ECedT4YWiFJkWAZo1TvSF0FjFO3/FJ
RjIZCUzNsNBQ7N9Z9b72GxOLqy7GIjEroYlFhCKXJ05maigYG6iP7ytUH2gMZDL9
msS2gSB2rIDWvOsUFoP4bOizElBEOs8sWcUDPgrCArRim989+SdB2Ps0mZ4XfICE
DutSZlm1ba8tsjpyr5NEP0fJzbNBcA8zkKDVgOkjhHKDjohocgn8NB3VLrJqDTF2
HosGRAtGMTXaBppiQVHWgtaxDUoShWw/247WAqPlOZ+KTd+bAkfP4Ea4rpMS5vu/
YOR0RNZTgFcM6asxKIlgOc4ETp7hTaie2qi85l45hm0fz14n/XmoE3l1MIvvYWGR
WfRt35s5k/njnp3sDIvLdtRj4jPWbmDwOYppjTdS4jDIrXnCOb0dVq3Fn+3tyyQD
FIYuMBwWTPQOWRtqckfDm0vO3zVQ8P653TPEYofu//AQJvgGgFGzNM9mU99jTzBD
IysGgdhT7/MmKvzxa66FeGKixcbnUvrdLcE2Z1K5HTYz0lGkCPbYR8B0L3fr0WXm
5mdl/Cdpe9LA6cmppswD/zccqc726hTc5JUI8SQJGVDnl4305Hq6gd9Ck6qTXaYZ
qPZqusmphmy9PCcRZMMi6bC8QqiBE7OgmsoVWBPQZttse6NgN0ea60EezEna+7zI
4VfADLY9vb1/m64VnIod1cikIBXYWj50fiz1bcVucagP2N9o4Wy6FtoPfckEgv/y
WX0NAXyGDMEq2/dy8x2+9cKNhX6GKoi/hH5DkRbEc3qim/FaK0piad15GBdXYf/e
3cXyW+s3Ngtr6obL1fIOnUyUD7MHWPaJDyApwsBdo1+8QX0XREqviZQHLuHhN66Z
G7k3rNYkkW1kxCroPCa5ieMvwM18ejxDKbBL9PEu4JHze3Ud3B6oycSargyPJRcX
kAd45ykuPqGMsEKQD1YDrfJvB7+0OtzPbF7LVsKv5zr7nIBfvcsnkA/YjKmXON9F
0RSJg90ng/RcJBph6nlFwVDd/Oebrsfp6ZPiIXm2nRsFxMVJSCICdHMN67psQuYT
kN0d9ZZ9uhAUM9diPwvHmPsgQIZiPhORi4sXf+tOkogb+dDLbkJJF3KqsJQGLo3M
C3B0sv+KBiuAnYFZHvbXWdkghu+fQHgEPnXuklFTZVXDQiRkgTGMTImFACegoOQt
M97rZ45LLddx/LLnQpkijWMnwuXU+hl05XEIzwkAhB0NiJLoajcLGZr20hDmNAiv
vCqBE5okDXT2yRyXgaruld4llYG8Sb60JUviI4Jgh0Cz6PIkLjl9zIusk/eEDYbD
aoFoBuHWAPV66a1RhcPz/kpnou/fzbhu1YXs6fDwnVdBXyufPk4u37LXH1Qeloh5
FncD34g6tu3Mvf+XwckndaggHMLhyxQ0nS0+Bg0uTV5uKtiDVSlctCXPtQMZp2AH
2SgJ93iIqiMS8eWtYylQ08gVC2ipdQ1geIolQVTiKtVEwz77zWfMvm3vLSirX+dJ
0uPckd0E4I5Woun82SatKzk8rVaw11anFbveRz1Xu4FBFyxL98kU5y0qVnoPd3F4
YyVut0w+jGQ2LjZLHi+uM0V/bQDIVFKg1mGrUHoSjA0QWs2GTUAs4UhKHJFlTxoj
GaCXKKa9pSePLV8lvyj7zOVxRtc0UNhtkuaj5C9W6iJOkFvNfoP8e68AerM7iRiy
9VBimN0fYF40Y/x63HgZwnqe1eSXg/oxy03OwI/d34XZxt7WaCdo3IZwRnK5Lh90
XBX/1JgkL+yBzH1ab31yEbNnQAw6iBv/t8jI19X4JmYQsh/IWRrrY7PQkmUjdQ6x
v5+PucDh6kSeVnoHm5ikfNRvZL83eOTpNp10k27YhPTwuCOACL2sRt9YwSUcNhnz
s5yA3xpkeW656S1+BRSELTM7otNt562zUh7bE5lEr7ITO6EiWANzAp/wH8UW/jAY
SLRezM+9exhkJw5qJ1ctlumj9g6DK6rEns4+kcvkdm8hJCINlgpjr3qdE6XG4VUC
wFnJHRTMaOEFkTN4a5axmcSFMD9wdDSwUFZUqe+TVIbFsWaBZFyrkyWm04hKGOrd
5tya0b6rpgpyGbsA5WDJV/hpk4sIl7/yRSXwoPcOis/vOQHoUni7Q99DyP9Vbl8k
ui6pPaUHWSgdEcB0seAFb6i+XF/ufKm6v65UKC9YyjJgxIvJKdzd49DKilkpLobu
MGR2PKbAlN72EBYPaOHZQOZANrVf3nb6tqW58Q6SA66i/UfMhRFmKAOf1zZDUQci
rgMw9gqBGf2DVsPcvKcbLUJ+Guc6Aeo1lc2FNl1aD5a09AEK6Od+Pcu5mAs3jqZB
m38ns4NjWb6U6GirmF0i8izUbHaDkDIIrWMsRrPmmK/Q/Fc4oxZQiaWn/i2Xo7H3
KS6F35VzUhZZb4QAB9Vd30gNzQGqvWkuEovKv1CLT0m20AiAkIb1jPPVUYKsGX2+
mk5P0jw8FAOFAnnx+c4pIU4y3A1hTWdIURbZT6vSNUP26hnGJrTteyfUx9eiYBZz
mcrsFWCMcgSuFhAL59/mSCxP9iS/mCOFwpuS3UZwinG2GdFOHwmi+I/Wfshwe/oz
CMPV/XiXHaiFxnUuYZVg37Yw+x4kwd+LS6SnYwh4cdytQoAqrQVx4alGd3bRvSnG
twdGEJzIrW6rPPk+qb9Yn/SBsPNBPGgQSAQW0pS/PGvnRGZwXt/gWYndNGhu4Itq
6JpTeuTsbL+Re3hdX2doLD2XhDoTkQvN8z1KNOMTlK+N53fbvP3rHHC3yfVRNiuf
jxf+O1USZDZhpJ5hfq+nvnFiMZZKHNfmqPaCEWNto+e7VQl4KwQLiKGUR/mZszAp
tC5mQRX3JPHBWM2kXZK0fqiwguJcKeJlx90jfGtNluJzu2KgiFUuzkmSGoWqy4Px
YSfNXVnsOEBbQHdNQP6GIdxGxKAikh4vZ4/gbQe/pAyRVqE6BodtcivQKQ2Kg/oU
eQjmgTtP79EtRa5PxR2qsXLhS9eLaHg1XFrAHDVSUJ/EbWwqNEAQrrbwkiSsBSar
n/6OIgxcqfKscMjRXj1vyBIcGG8XOZC5inaADmLqOtp4eyK1wVJkOse2i0dSwonh
e+36ehqFNNi5Cel4OJPldewHgoJ8tEkEiVj/MebU8uDPBrmJe2xiZvfV4Yyg0U+K
TNnmQj0wCv4ITMWPEwtGEGn/BXtiX/sIsDvT1mj+cuxyYpzmRM/Fbf0IFl46wg+s
riUYGlBQDwTmVS921vBUIt/vaR8AhUQvPccIhEcbin64C0oQXyaZgtF9qntVs4i+
roXOlMQVLU8fktWMeSXtZNiyPInFelZ8cGciqkAzLBEwOVusEMFIwrsKOGXFSskr
h+3ykJO4rfUja5gtvH51HFRqJGAzJfRq+6g/7WfjEb89R/DrEOwtmGQDsshtpFuz
v6fzPWcCukJjwOuGA9NDTKEyj2n/Lzno67QxeUKRuKTG8Yt7qB5Dk1N46om7EvsD
emr4PwXauro0fASIczOJDKqX2jF6QUgwCgLb5MO+Do9wHHy6rDFM58tfEkYq4VZZ
5NZBK4ynpzlJ08UOn5QCKimdizy+bEtJZa0mU/+VNOjczut1xKW5CEksUq0N8Pv6
g6l0tHsPdFQ3ypswHo9PqJ8nvoraJ6KnKm3nYMNyCwcvTzfL7vRzX7FQkrRlswSg
rKShuadOpPXCUVPMgxqtKtEK94OrYwDOkgy3ZRYw1en6V48oWLOuzGZlKYgi1jaV
wLldwddT9OqgH/KhkJX28FGsok0lICBI+hMpz2oKJunKsvFshZD3Kj5lvSos2Yq4
kH10GGlw2TThf+4eTRN/SBc+E1mdB4qnSJ0dQVZSTzQGUoqb94YGGx4v0nQho0zI
rusw5gQ9de2wc668LNTvG9aPJfcjZEd3RDi5iuFLxFXRbf1PKhhN+gZUCv4MTbsT
YM9vLEh6ilUBm21n9HkfIaaUYhQNrgs9+N/NLq/una1d2V6Nt2VSb2lddse6LKNV
jHwKxWNn3w5mACe19Bxi50Ueg09IhDcUqQKRbXxp11I3k5vYP6Z7kmB0BEXKAAaQ
ZGgZdY4QMXDiU7508eG/bEeZXo2Yh6ZRB62E5y6Ynk7I+rLYARBwYKZJQvbxufOS
MVTW4tFjCDJ/dOMc5SuJbMGGkGnsHWhewoTL1onTfEQ+WsiyMPHV4lDspv2Hgk8I
BpRDMlckd6DMi6vH1tEZPqqhngzbZAE4YRpGPBW9Wd+uGXwqeZVVD4EmKchSGA2S
ul2L9SYhEVxrWSyV83Hsm4vR5Ol2IBJYJuXWOdZNjEAkEoUniLwBHzdmqyNwIHaU
Ey9NlGbyD7rm6qvDADoZfVujI5pl8O1ZPOqeGcap8cL/+u9kyreJteMNDxWXXhjh
jxGbQoDaT8iGaeGM5Pdm+KN9Np/Ti7fbQnCJdXWWxXThIyWd+7tlEl2MAN1mmM1Z
IloKD9MdoNvSY2rAccZGUtoakN0sLShciWcXUCwLAvj2hlZi1nrSn0lKGxCJQeLY
P2pS+MvcPSsBUMkuBjg9nf4vm+gjtQrbIuuBSIm+Qgu1CLUDNMD/BbGOsf1o2Q3F
CyFn2PvKBmYO/lc4b6SuV/LN0+FUe49UJ0dIGgAJ9jl7nP6Bm2HwvTIx7KfHOYUS
vuecy46qbO3yxSCQd84Fm9qdFLRcdJhdQ0kGAE7TQP8tXeT7au1LXLGsjQE3SSNZ
1hg1bXyHjWyNMdTNLzwLnFm51A6REdN3/u33r5BOiEyISkSnMElIa53fxAMP2ERy
kVxBPx3Oii1UWsQXC/1GfktS2X+P8OKTSq+S5KxvsttxAHKC3tlB9FfZlrePhtxS
lEnukMrbiymB57pn3zDxw/QuCt6Och8kWiYbcXJiEF3u2JpmBtS2G7kS02WTakLk
g2BA4Sp6w6DGzixOgVFn5GiURV71hXItu1UbRzttbtkTCyemUC1YTPUIBB3LKDnn
O+R0d229TBwv98N/kZVA1/nW7bWssfLW8BAViW7kBRK9wfNAG6nDJThki8EoAnVY
xHsXvRIAwRQMpSin5n+kf+ZvgUR9VvoW6GmBBF9LBhSAUJmPPpXbzTxsrUeBQx8t
wKEUvXoul/iWtM4eikdMN7GxviRC8w+/2VeBD01/UM2jvWMZyhcPogTx231QZSht
evhR0C6eXgdcdE9JiHpJ39vvAvgHqy2MxiOGbLh9pogexf5wLK9NterE/5uJny0T
WH1lEO+slOpWBYg82szDn4HutbNdncOR06APP0I2zYCqa/a7u55+VetEoHKCr+Na
mWmqrub+3bC+LBK2YgtiJ61dyq9e8uZMx8Jpe8r0l/3zgMO3nWy6bI/l3mxMIMEG
GOVVCDeSH+DIDZxUHFu5auEMYeDhvEJdjJa3S15dwgeYn3jeH60gm1PKNjLgpPu9
gS4FcVIqqnOv5F9R+wy3aE2GMmuNvCKx8caEpjgjGJSjjEXYxR8nb8bjAgMSJ540
tkSfo1Z15y/gDbQA12xjXh1ko8uRBaGTbBxS/ESL3ai2sb07A6foOG9qAnYvdfTM
dt8HEtsNiqZZzf/nm2vv06niPhqAC9WFcaMsrUTXG985R2BMxgDnIRJkqqtJNUQt
iGqAIP6KGXVH8d0tz6eU9LgYq064JyZJqT6EpEKM2RFwk28shbn3aDFfU0n7B38k
AVvpo/XCHWRPZiCcgzbN3RgyF11lEEkkNsq09Lx58AUfwX+09q/jRJTl30BCbTL3
vc00vbOGfOOt6F7njwjq4LmXpWhX7CJY0WE3KpmEWzb8ya4dKbvtwb/QCGqjw+BK
0oBkQNuWFOiUvMYlwly3JOdxnu0P6+XPjVkHP8W1RFGnEmXByOEMOHegZGxTI4KK
IF9+9cFBuzso8Xpz/6Lm2hFZbi1/QKc2Cgj1v8a3IecsxDlw2Sx8kKPO7Ea7Q1Ti
WQRp7nGxiOy5zWRp+12TrbJYQgeNvNen3lg04g2VtU/Q0uLGMM7W4nOmaVfF3pqR
47R04b/aaNDufrA1wgeipcc77E3yPEmr9UlaeHTlQJfKMCdeHjuVx25ljJTBUkYW
CJWdLR85RWs7Ng8IgyGE+Zmq60oi1Bt6oDH++pG1IwCSOnK8CTj7+gGswySX9mcI
TEZErrOrlLd8bA2afIC6g9V8JrNmdnkhr5BtASvbAzo4QfXyoPLVbijsdObYPccn
I8BXYPuk/geY3tLCCsE+PR19qxlZMPcIukF8jDYNrVc/2C+1lK2lC5vnxK31ZJ8v
3/pb9ADbM244HWdaOWVkMXRBkU8hNRwHacONDMU4o41qr+qZKG2GvKzzqY1dM8dz
lAZY8zJQcLdN/VGUcZVbpH+s7rLP5g66qYgRIbUjjoYVG50aporoVCWHFVLTmSOe
eYEyfbTSEP7P3G9i2bf3m9WOFkA4BIpjMfpLdHaq8XDHRP2Jq3okgCjikmDdfx94
JmUnmNGy9zxg3q7ZS6Lv1hZGCpXM/93+9at/YQO/8fKU9PAyx3bNArJSo2pboZys
bBYxBCYHTSdhUxSaxVbyLnpvUmPF8//hRZuVOGHcUQrI8cKtgwpesRD64ojoiKkp
gaUagojQVVGYU1O5imBG78rh9rVT6QmCDKj33Xyp4UUDn2VF1axCibiBRH4iklLz
b78NNgsUoMTGGXS2tZwhcbYJtfLRzBHs4/tUveUZzDvMDvCvENUrY8XL9MMYvADt
3iegXqa+u67dYwCiLtIsP3+huzf6oL53TSh2YdWdJFy5BCK91bTCGohXjt4nCgoc
kWQevRauRUj8tYT8l+Rh90G7HP8FZbpyR2gFNUC9Pmr9jLe9o0rEoNgCAaiYDTi7
NNu7P87p86awBSFXLVNvl+c2k4cn7sSIIoZD2PZws2AofoWWByavN0f0s9+ItAkO
c3q5Y7dfuPL7NjkkFbppO9FAXxWRW7hOR2/NKS8NBuR/UZZ4FvsRBLqwse3sww47
Nk+997QHU+WW+URptnf28aW0aobpAS/iVOKfqfPRjc6H+gP9NClaVRfEauvs0sXY
pI8NslflLhOk/tiyGsIcyOmpMLJkJsneXFp25xWczAwtQB4n7mTpqPfYcOnyhSwQ
v7WBi72+Fe2jABmrYpLX/E+nZ6mqJ2UCG/hLdQzja7k0kmrF7vQogjOgtm2aY9ik
Gc/aOsz54iJNpFa3mPlZOvgyOEsQCM0fUzX2jtlkxgvpVtJe4unhDtWlBY+/8JJZ
a/KQY01teqTYewLo73NQ6TZEWauOP5vgFY/IWhzgnX2gs5fnynDOKudeaEWW1GVn
hfV2NXhMXDnt8sSMS12U+Z18L2xiicEXHOXJLian+Sa+5+gBosYZHg7ElU/UrlcM
Oktw1Hho5Gatsr0F+KcBnybD8MiVtNXPA2l9KSEDn1EZm00ixhxuFl/Juf8CBPoa
sv4rs+57XJBgPvrNI49OkAjc/MZYLq8c6cdt2MmG9urBrpbym7qKBlgwrvjDtmEZ
7APGOwbFC3OY96PjIF1pjZlH4gcCZrtb5+0rC6wXHNLFqvb4sbapj2r+T3ipSRbN
s8F9WkiZ5t4PSbMOFaZXjK4vfSk4CGbfU6wP8YWHR4oHKbkqpLptjRq+OAOQmT4i
2hE2MIunaNXLLTyWr/lsxmKSrbkk5lj6wMzbxBE8b/SeYhYXogunsZARFBeRghDk
uVf4PHN83bNrf+kx1HoiDGDOS/DZuBkW5Deiw6BjsS2w4ugfFmC+AfELn8WQV+2l
M2FgchTrEb+H5/xawPm/KrpjRG/7FTe9ZD1zm+Hg21GVj7m1l/VGamlNncdJ/6/m
IX8x+UkwE2ivQFYmXhJqTSw5DpTzNiQR6SRRpnpZfuT2Ov1Ww+DnEY6Ca0cMFuYj
Y46phs6iyGbqn9EiNshsb13k9ATqREFlmiI+0NkSQZ09bvf+bl0B7VlzLPeGt0ST
xdUHM0rUuqvX1xLTVVvN7JubUcVNHhFvLpX2cQOnljHD1zfF4Khlj5jSMmwAzlgV
aQME3U7sRBteJUgIFz5BI/VvzfM1tDyEWkBFij2fyYN1ayG14pMWrdTmCSarDM52
Ayihk9jIaPlBMkfETuYryPD5JQWkJcEeYSwr9zev62ZXNkmxcb3ZON9+zK4uRlwQ
L4heR32U45aolobb1kDFU9cVbsB5swo0Kt23njW4pJpfVe1Ibcn6GPXUAxSdhwHt
y0Gh7BeShPujGnkEuCVhnPAF1sFqUbXKOKYKwmJMIQa+vhrMvafxHnCUVFAt3g37
XsGvdz5jlCi8SDm74vSCQQgWBol874c7hcUIky1Kc62VIUVdg1JwZ6yda68sZtS3
aq9SzpSbK6Wf2M2irFUzfALe7QB01ajqS+jqBsmt2RrxMMG05uQznWx6z/VZO6/S
JntCfgYX3NCpHsXfybMRHW21ZMfk9LFkNxsU9YJfoIUSim/AcS2BBXMg3RJQudZs
Yi0/yQMqHwYJ8loW2M74ZdYvZ0IuHBd4FPbHvqkuAvRGmNB7blVmf82+O4HFYQs2
nuzk1FL+9ve37rHpCKulLo8hbiiuTUBL0ES6wjYT+lyGu20y9p+xfYZLWhxyudgN
JBul11g5A80AAPKuUnGepmbaKx0eEUyINOfCXnVaMbaUQlqD4wWhZhV+cdyp/qzb
uNRCMPd/V0Ro68yodhGRmAguurnEEhi4lq+8TSz+qhKhAJtz29cmMR/8Ld5SI9nf
0rXx9X18DBwgmlSOEtZVMAFgo6O2WkDth3rAbduItdwQJ7qs2wBnfudeNFR+fmk0
RrPlsyDsjlFBRcCABbQyk222Fcow5Is7SdMZHeMdlU5vlPDS8WybYXjusrbl1Emg
N8Gxl8LjBIHvtPJKF30RhZ/JBiH4k9YJ5QvC7DnZf4RrKmLZdLfUhYz/MtynJb4E
XFa4CRyrlogrKwHTUu46lxMG6T5r6u5us1VS4aIGNcuoBenPz7SANml2YTdkWZRm
lYBo5nUsXTIu2KNeyOJaOaRw/jnC5yFIrMylz+M2zMz9EOzTz5iEN30WGE8P9jkU
M++klql5SNHFwp1VFW0Wxy13qJ4/9eWGH0tYMhqBWzl7WJBLjeadi8bAwBH+efEk
GGAp6y7w/Eky8wnW8RZys3p6GTHZB5Fff6+2f/JLal7YuaL/yPDNhdf51AGBnvfH
tPJFNJL+rOK0hbVEJgbOc6lt9VRiqWwxcBH9g7om5UsN/Udf2UOD9z/iBpSZRlDE
IWS1id4PRYxzp9UMzob+8Q7d5VFZbND3+sWdmBFPMjhx13NBAj+hjNl233ZA85EA
lYlrnrijBU02PLMjWftBL+JkVsFyCYzL8tgvQZU/nrdYZCa/vQPgIJQCmJNdcwVk
ZTJl1XE92DLw4gpknM/GsEBymZbWpTUDLXAPQSGhC+3Xm7SAtp6Ah4sBP5+hn1WO
A9fo9tmuQ3YfQGTYcJXiF+n5gKsF7pGTOlLC5mx5edegWOBokTgQ2EZBWHmoIwfC
v0xKIP+GCqUEGn51twYpkUzMloe8Q574qwsu1AZV7PQSWWXmN/46pSDjsLBxJgNG
8A/aYo8cDP88SmtdqnQhmq7lNoCawZPUoSoYV3v0zeTdYsecKjwXDZgDPTwgLGJd
eOERyl9qHhLT54tn/Ax3ZfJohHg1y+khykrmD7jTu3008MCbTFllFt16vgN/Wmak
sOFgfcKNkYlpFtXtAbnvNVsMrwUJaM2YtL2c3xoHOt9QNPw5L4vfxQltbXbX6zfu
EzRf/xhwc04kp2tH10O43khlfELkO/iQ8wDKavbLq6QIyQGo76VUDEmaWZDnc3fg
BnRZxPZ2ty3QAnHWfzSd6DRUvDCp3qRi5jKpra0iYut5WfBwAYM8fvarMFKl5ob4
CJnsSQ+OE1KdylsjLdRDyeHFhIeJnN8E292TjBt3gu7LiGPtMtDqgM+WMTzGOOP3
p/YeYqr2kOWI6j+xPKLNjwvynM17in/yL6HryeKBDJGT8QSFrgB3VuCHK0zgxnTc
OESseltlS/pQvy8+v+OdNcLkLXITqGkVRTuaQumdPYphqM0GEJzoW7CHxOGe7NTx
8g6VYjrs9jTPvdiczc03yAguz1ceYiyfPdPjrqkSC2ntWyUaqyxmajX6tkHqNL8B
MalbeZLAA9pwvTHvZWaTISf5JmvyWLNki4p155N88CW4xc1O+9xoKW8xEyBJEZif
PbuYv/ue6fgrjBNEHWp5Kt70+fhH9F/Slgwypihqm3iohQGUR/meZHFUVpqtb5Fi
/fUZpnCtGZe9mS/CF4Ougjocv1gBKsyR4rQFHfne9jr1zh17pejgkWPq22DuEFsw
ItQp1pTCZUpN+ApCgl/Dec6iEwYEZdEWPHDxM+9aH1y16EvgKxOCx0xjFb84SJP5
NJTACawnVbOEGpJ8gie0EFto/O2zhzL5ATIu2da+H8QKBqJJEw2SSE732nTOQSNM
qe3GT3LJBAnzd0zYLBOlLQIGE4tZPk7bd6VMvUyPUSQTEUaNOIGUW0dDsxU3vna1
uVQO2yHRLutreXFUhWQe9ooR8nPPSt3l7xicnlLAqd45HXs3EjFxYaT4Anu77Ns8
h8wVy8B5jQIokXEoWiFSiS8YGoras9zU692VRcAcTKXQKwvqNSrE6aDPyBV8D2cr
0MOgu3pnvf3JLGAX+Ndafd+UmJ3Szuxxfp/g9rIHK/WMqQ3ApN00yezGJtlFphgi
vov4iX7rpWaXDm0GUixVOihgLaIc3j4FmG5wlMP/2QFdVGU3EaaaDurpefnwdnUh
cnjh1C1Ufe/Bta11nZ8RSGTUrfvwHo1aHW+kCFFMoO8VnE+OwYbg65zDLC8sZQOl
+mJQdXDCzzrhNZfjPTcSDBmr0/fQfeLntAE8enANQiNZS2vMkpZzjPm0SVVtpe9n
XhFI6SPp5S3a8Rlpk4wR/vSnq9m58x4fm9tIi3yInEzICkesZwketRV3lMr6Knp5
HGfr0qnrPF5TDgNCW4HCpK+53tQ2v6PjCMX1l9w2N78CRG4hwXDdu9QjPhzvFnsf
i6BhlnnzR6nJkBP+3uePDRsYZRGql50sdJpEgolps0nUqIlvVnzj6jcsXmMTd6Oi
ryLj+Pi/DL/BiRLKAdz96diTifbEdBJocTvFx1B4L5NduL2uQJ1gKLiALqJGUvB7
p13/qTrxnYX34VfMYOHE4+Mz2M813VgQzHGeVXPvDN7rCqhJE9i4y8nykj7sF1d5
bqRrsdvnw9gWdgWZ9op1V9Ll1txfb6fvvSOzAu/VV/IvrRburqdC0yY6C2Nm1PxR
iy74QDbHGI9IsqaY9/ZnLMn0gdRJSjQ/MlWFtjX4LkWdf5z7ajY3eb5a/q+r+JHi
pWtXkDl6VDsXJhVTks8MxmOA92aySL07prFjgr4Qx2kIRiL8X7jONFk7FYk0tTXK
v+Ygc9C97UxtoTWH09XacOp2gFlPBbsAjBLpyahm22T9YRxvWZ8cwk2Jkid0s1Qr
cxky5RplxCpwpsTxs0jPYVkbQLvItaAIzHT2XV8MYqria5aWBaDDVbm6y3cQYxUp
HtRJKTlbwjKbMDshtqZmzG50auF6GkVDYmEQUsScAs9KUs18iaEZ4YhQeb4QwGLo
QaYq0Am17zmEH9dLiQibBoqHEEqeOXTzvg8OcYgDYflwEpfTcnoTcoBz77oH1Wdg
zuBok/z7HcHEg+gsvFvUoHYlxJDh4FTRAsoYAQXyQiHS22+W6+9G7DSRQUM1iw0P
9f+JeHQvOLCqeAwW3XmjIQypCbh1v+mWWp9NgxIiXIiQntMexbfPmkHhMOut/3sk
1dtyQSYkR+gsEVx7XtONNaNTomh47J9lLSeoRhy/l3wMh7PSVNLNBM9xxomlvMbf
EoDHSsM7T0PjMxEqlznJEfuBB00+mna+O0+fXQ1pA/ncEVX0osA7r5xbRKeN4xVt
nXPrF5z4YbpHU1rd8ZRegucCFi9dHDBxzRjK8/K37Hwmy+Ss7YRrmMjLOhvJY1kL
2k/BUAPlj3f5FTfXm6gfNOk83a1sPNpSOyHABkaB0bb8F5o06FhUwy1FNZILmXOi
0nXG1wnASerfBwhiYK5Rrxqccdyjj3CP/mh5N1VCCfDSUxS0nzHJZLdM3SPzmmiG
D/P+ES8TNpR98CDG6+JXaQDTXBn9d0dFRA/u9sOc/+GlsBJ3P+32dyFS/qrdt/Ce
iPR4wrHNKz9j3SlnCL2S9sZdcST58eVMWLDHVdsKwUANzvrqS9J6j9NVcyn/A6TC
p/Lznhwydxz/aPxAPaefTBl5WH/3VGcxMzlU69P3EhxdQyMNdjomUyNqFOPjjSVy
9WMQqKAmd2B5YcLg2BAjKqk3a56d2yFKuXTzU59Lzykpqj3Cazl1qpDT6EQivhrP
wBBwKpRh3VbTdjWZAZcBmPTZFvUvvEE2kNRtN0jOShhaQ4BHdJmo25A80ILuUUVr
d36y16N0mf2Wj7Yo4AKGoiRnNfyfQGK/NcNInN6G1+wfZWMOV0w3uzE9GbBoHrPc
nMAEfwcwEKn059f8Vh3X02DrGidGJUiPA6IAuxs41PrpvyBwD3UEZgzfvT60JTrB
1CU+qQZO4Gt11fXSYZ/SLuwfWh2sjhhhJoLX1xwBpm3wMJ5dYfA6UkEHFekFqRD4
jnCoY+ait/eJxrYNCsd0ttDDKJElz0nEntQTKxeP2l4M87no0jHun732/T8KdCnT
EFcTJb+9y2ZO+VowC0UeZq4D6OJUKySelZDajGeQoAoKvdyqWnZ/eoqKIKxQP/WG
0Mh8eeuiK6T2kwGuHJD16KAuN8EjTfULL6VmHt2zpX+7aghenj16QfyVTRdbqgDX
oASU7ywOi4JdCXVJGIJyxDfnDC3Qz1gz2tXK7YnX99sFVduKTGUS5i712IsBBZ0l
NyMJofMPR18d3RknnkxeYTeB0d5hv7/z/JM1PXfrUxl5D6T89deCDHAhzg3GMqtV
IDKCG/tgrqY3ySHvRX8wh5BQMbbH/rtuUy5gfImkj0MKfie5KxlET3sjtjMrdxkc
PcWwOg/lFGFpg/2F7nWn6cg6h3SMSKTG33ydlRtLm97NXlAAtCA3xg9EgB1J4rg5
Fjcd68Bo18/42n3hyRcw2aVR89G8TpohJbwLq3JtcOBhHIThKYhPYM31RD3ywxJt
F237ThYYA3tIMPlMzHkN2bpKuRBHEM5qAE+ff23716612XyhaqYbR6JaxdrTdSRG
GS+xmCEL3FcgmblJrogI2zZxRgG/5fP6/OfbhXdCLK/1TEoQnNXLiQXVQh7p7XsM
PHUGPfP5Wr4kV41FdKHC/UoYuIdPbqNfLb9vuuDUuXyEhd9/Kdw7F6ie1xzN/ebi
1pMopGeNV/dlm7xvxBIDpD48baIPGl3rBBTcSjpAVCDP9H3q3NWi+7JzSbQ0bqG6
VA3cVYgYHcljxy8sDQYfDxTiuv4sLa+VVaHMeHz+UmrzYMkoE/1yN30Ba+WcV5Ad
Lum0j0pGoOT8DqCwPU3l1N/vrdUJKq1aoLfSTnZf2KIrEQypyWPinCbeWFIXhjev
yjAUCQ7+cRzL9x+RiJAaQ0GCGNx940dyQ2QK6h4iO2fiJoleDFMwmidjyYXn12TQ
IouiIAQgGz1ksUKpHmaD2GOmFp/y0LPbWweNyxK72mpCf8Uf//0g0xq6D6BlrnlF
rHrO5UHLKxW0wbgCT/5aCMHyGvFhsl7FfGtjyOhQQLNS5CieewH/VYxzI8pp/xvn
v/UzBntGNjoYDI+QpFY5yaHfEb8JRFQCIruhWouNjRV9hA2E6GRpSYL7ClKasnrj
vdF+72K4M2IBwzUDOnvf7KV8vS9Hexo0eZNQ2cJytNyTBBMEyTaJDJHlxlgBTq0a
CbQQCIRBHhHKbgBtiAEG0wg4u8DrNZGsITJf3VEPzVl/AOH1TYI7QbbCbnahePx/
x0ciqG7F9W+60YumSZgUxpk0V1bqciVoPo7Ul06nGSqhrQnTNIeXmN4NaAiJyJBr
+qHfWtHOOWVDd6HQiJcEz+hmRSTM8lsT+AIoDAximmuwPHipqofzrjG3ngQVJ0j9
jK1N4uFj7hOocucUoQPRlJ/r2J4s30Jsyo/z89ymp1pcB19eE4sAxJ4aL5/p4BLS
ZYThmmVml9udc0SmwtNekQ98uH02LAmhq+iu9OHeiOO0vu8AAQy/QPYpA29oEaf1
+si789BgK9fcHjFh4YprLuE+CMNQ+e5lb3E0CjHzDs8vnAvqHwG0zFUgrwyeVNNh
VPyL19rGva45aOLeKDZCstEqaanVqSG9zyWeL0QYY49zgDoBh26gxp9/tOOdggZk
mS7DZYJiOfhfFexzhD9ZSdMzzjFP4wShytdvotXDhd9iNDiUD6pHxi8j6rXjvn5f
4uDrruzPeTf2jsctf1tBN/gJC5ow7ZJpoDutkpwOwe51W8VSqa6M2XsGZ9fmkpEr
C3Iq213Y8Pzq4d7DY4dTU8f3QNF5JXttvK6f0GR16RjvQvNB7slmoFl/REBxwFRv
X9IvyR3DOerrPB+48jBQLQeF6Tza5H2tlALz0bq0fjL88Q/QTELnsA2FMwZKkYIT
O99XdZqPOAcazhyH3b+QXr+qALOdmy3vXaNgOyzYwnpPxi8Xrj+vw3eDoBIusq34
j50BlqkvtE3Lnhs1i8+vDW6GnXPzUIHUeHZ5Owzx7gfW11hXPoKV/RKYOtLQAEGB
f5vyxPzbRr3np2lyFKB5FVWsGN7/6Ju4kEbljbwXCbLSZp4dhMGONoWQFKDMD4Gm
Uv3+3m2JE92+/znfVyS6ZRTfLemKPxaVqQOM+HMTFE2iGb+SSb8+WtU3iPp54l5a
Ti2f739ULetVi7c+Ly8b+h2eGrtWJPVBsPmHeSLo5pBM0MGmqROb1rx/YrGSw6HG
Rh+/v8qZsMMGdn53GP8ZboQIbRkpffb1JBnm9GxJ+1Swv8LAt9vwzwWzZUHcRtL9
NkkdKB9P+x6vnRosPxpPzS0rh32as2+EPGSh+JBh4cvx58I5wzpFz93D2uje4FFh
c6Hr7XJUD1MRKiZjIR6fIwQHd8ktx+XIej0nPhH177rKe1vVfia56AlwOcZBqsre
GAAsaiDPses8P9HdcUO+S938Xja3ZAtdBNP665Yha19zPUzNTz3L1/AuoA74ckhC
8dBbW9d26YR1Izw7kNAvG1PAHZtBFoSxjGjm33mbgnLTmgK9gdZP7aid8wVbInwJ
zK8TL+2cc1YVjPQ619Km6rx/zYk4HIlS35nIed66BOVMniVGqQN1/O7Pi8z4J0nZ
ZQhclMcDJ7aG7C0qY7KuHWpS+rmVKtyybiCWvRCnKXtYOv150gmBm2X+gBN60dp7
RkJQj/vD28Vs1zuOecgrh5kq9kl3RfQqxd1BwtziLohmRLxA+/jFou9QMHuR/OoK
shxB9VYsg2h2pZ4fjbTNZRxV0U3AgxJ4uR31JZwcILCk1bSeszTRPyZJJh1BBwjn
I3pqNwuOb/AmGRSHmJjgB5cylWK6Ym0euNUJ4gUy0jiGi49ZqaXBk5OrQPE9gB5y
mkveNO4DvNjrFkPSl6b2OFb2JdiRwqC5PsgKM3IzssEOww5NLov7WW8kRnrrvkdv
Jz5a56zM7DNmzFjR3iXbS51qI3e11BsN10SrGTTucT7borU85X2erJYfJYDm+svG
JzrWnam1ImGM0yS6JO5y572TDdLtKq8jIoZiI5FHl9oKNs1oU5qlLSkchd2F+Lv4
h3voGF5vuBXVLG3ZDE8+ff4e9IoTPihok4Wl8TyebNmArbFOXN/XJSvIkPCUx0hp
Iov3630Ufh2ghThl1S1fmJ/NHYN2guNtgZYNoYvgtZBe2+SUB3r4o0+48Y3CJ32b
RNcYXYBO5Y6TICsW8gs3YtxLLGe7XVEtse0AZw1ZAQyqo5qNCNs5LCDtSoopMRfl
yiHTlWsyahiYVAq8bdzzwporwVsd+Jiwwj8DJ+TJ9nXVAuy9VDLe7LkKlQ/NiOaC
yXjkjgqs79BOPbpVp2tolU/LXixzNttV+hiLri/9Pxwnyy9ODrXvNVCBzNowt3xt
n0XLHVsaGJMrL57TsEgDWXVoKWw6UCH4XNPma9J9buXmw2mtb9G0qW+GLbl7tED7
R/ByNWZB0RH0586jx6sT6t/AmtzL70UI+CGXQtMDnnJmhgnSGz16JQGwYOZJpozi
mPNM6eAWoVAjomI25NCU/DgzdoRWiG3gWyLt9/eNFntH9jduFFL2lfhFJ5Muqg5Q
L4YCp5zQRKyJnwV4TsfLc21BOyzyanb8ew7+oE19O7nk4h9SoaR26ZqqpQBNVWr7
lrHUxBW9viAJcrdPXpEH2kOuPgmKbyvjYJYbKaQXRu9flUyUudPlM29XBhk9sg0c
ABksqRhWOW3jBe61n2z0uPQ2iuE7vdgbspbty2BZH1ekdKQHwFk0zb9KX6zZxSkn
GvnQ07faAixpj3v1RpVV+ON56VnZlGb09h5rKeOqR5MwubSOCUkQZYXv7TIsVZ4k
K63hCZES9HcwtkLT3J1frGRW3FPOyYflPW9g+MSjrfsPrX+ep4oDOlCqg7i26x5r
tmdbXmjB92ketejUBrwWB51HNAs4OF6eK/t6b0hkP1kMcR7Q9Zjvsftbky72p1Bn
yFCEOrry5yoUAqaBs4Kwlci2+eVFEZWZ+foZrrpHEntwOe1SPqZcLsiVFTIyUX36
O9Vhjwb1zVKkyAlz/z0QhP85769eSKiakFR6UKG89LPZRNP3hLJZU7pAEFeBbYfA
sueCXipPKmoeHa2sB1Iv0vw/cS/PD5/BdILRd1euDOdaGUOVXwsRxanUAlPQhfNt
iFxceDP5NAoe2kZXYuoQC2KE9F0RbBgfmiMDB6ZN4lJOF1IilKyqYrEkAkvm6uQg
Q0O7EVEDSbsFasvOP/XcVp/1NMacV4bbhhbuyIe7vUowPj8sxax/j4qs51r252DZ
4dKTlGqeTb+Mv0AMZTXEwrI0RspJVIW25MRJQVWWWnUx6yNjnpDqf2URtXRrJcp/
e7sXKaqkS0f2oF0VwfYlDc+Avv7J6Res77GzM6awZGVFKtADYGtcc3qb4eOa42wX
HISHgzcIdqyUJucHyoueRg5TVtO85SGcUAwlfRxiIT6pu4SyeKNyWUrJHycor+Ek
frydb8sQRVVgHSSm386GJRGXF3JbcaG/EBlvnCruXyULVT9qeIzftQ+xZ62HzR9s
myrQxJBvIXcMvbb2t9rkkXcBJpfc0duCR7452pt3EKWUFax+OOYyZ748UX/ca5wt
4Cvfy8lf6NSj3V/SqikTyNhPXA9L45FuXJtKBJPekBx4ElZ2PhfICBjojWIsRa5D
7rWD4RxqkNZ59IWd1sTZGramAbMF1OBQMpd0e9DjaCprp8/wSFlwdOgP6rvOPq/A
kehA7bgbkCtjpgsaVf0a3tMVJrYwo+hPWNwiqPyRqY+EEJoJY3qxb6GIb4ahsnHB
vejQVMq8JBlB+ve66gLQedI0ewF6C6x4FqM2p86yjjYh9NZF5S24UCPh1HmZJbKf
2VuoYSZ5sWgKfNGiGKNGiS5DCUamBLy4eTZTuo5UGK8THjlaeQ+r4ADpa84dTPy4
GbyLIAOcL8ZJ3yYBcCYcJIXeDVG3ZoYIvsmM/QE8C0T/f5djgAbQfdqVfP1p7LTC
SOdkZ0yhM7BVmKnriUZ8s7LR6ha7beT7C/0Rmk/5qXEAuu0vjiB1Be/cZKxyMtVa
d2GMdED6BMBSqK9cUjRls6Y7C3X5J3DVQsK2dufD4vAgD72858Hc7u/B76Sk+GTR
Fu4J62x7O6JefoNcfLXN17/ycK6wZI6kM+sMN0kOtIzowj0374qPtPL4gfZZjqjf
mL0nDbQ87bMSNDtC+r0uSyF33xOQpP+bw2BCi+e0PZ/g6uvkMnhYpZVwGczqz+ck
VtuYUWeZII2Z0qg5ztKVteGwjXfoWqkJnXaNKS0AfHRgCHsnme/vBCF3AXV1RGLT
tUnN0UWoOOwgFrYrPIv/pHNuKpvFTrUESamu16U7zhe92vobE3C9BQeC07QULdLp
bXgp5e8iorP7hzG1yfqZjNwMlajO9z5kGJGduCJfLg/vFXKSHAFKlpLhWvMX/Hq7
c7xN8YP6GGD+hy9xx2bZWOmzQfbwU5YKRwx5YQ5qXgK3+QpGO7twWJwbdaIKUWhQ
r0MCtl9QoewSSDSZBTUOVwb1ujB53dK1NmB/iUqS9iffzFq+FQGEHtuj1uHDaQS6
CzhCeIMAx7yfmMfe8PmgOlmk/tj9zjwNxKNLlfwyXsUaijkZjoujR20W1pB1L0Fi
m35k1okRds2bme/OdKAewjrOSXpbijMS9dVKcBlsJhrNscHPAs6mLs1YyXZe/o6h
WayhmKtjwR9y5ekXtB6JMCXxzXAVl1BVrxqCLgjJ/R/nzqYGaPEPlhruxYCX5PGe
aNbPK2EuC9PhR+Zko/1d0JeO5hh0Gjzl9tLBE1eLBM6b7EntAA6C1sY762eVlYxM
9+d9oXjEUfoX1hCjIlZDOy3pyaK5bMlei/8bXp18oLIWGjMOnCOms0FVYmKmhTIK
Fb3UMiMGj6bVG3oB/AHxSkGUt7nzbAuYMQaGWDQeUwABindpt7Q1iBwiNDIA7eIS
jphRVE88pODvdfm9kvfDvCfmo6kHsPlgQ5z2ggtITeCXl6nV4L2JBzqfp4RrAQIM
77eQBN/bs3w8nleEyXaQ1NypkaLjc9S2IZzj+8IdwM7nrmGZacMqUbH1rL3dJJpj
PcEcxFKvkkIyOwF2FssNhk4GjAyLkmjZZdOjVQgw5GE6EQCnfLTFRvosypNplMwU
J2qPYXpSaWNUFpAAtiPc0r7bOo/Iefm6LCDartxtFdozVTqA3q68d4dHLaSLJqwZ
ZHBSK6XWcfSBFAKS2aIwnN9sN37tp05mJF7uqbhBxtYtHwiwi1V66/aZmegSSxB8
RriDIzhCNj18gHxmZIlVsTgDFaVZtti65Fb84NEI6TkedV8jYbs6MCf/9M8O0K56
6+6e+iKJctCx2dnt3UtPjAsY2zODdVpKjZKekGnIP2g3nUAvromVtdmqIQLloiVq
rgVXuMlJmzK5IpvrEF+JeE6GDJgJ89jfVXCqXIP5bhfPT8r31XgYOtae5XayUQd7
w6myeM82WMeLDoGk8LabuASmCue5yfLb7ninFLueirsOEl2wSrNtkBLXWyU0i7M/
OfXuJnfTDOrILrGF4DNzdG2vfcGTnqXycJXrVOsG29ki4/uIV1B1r3pTHNR0mkAq
CuIv4DmZlBsP/sfjQsr7y22yYNn3kdR4Uh63qko2R/C8Ggjr9adewzjoD+EIjBHC
6q9C4CKDyZNfKR3D71GQDs7lnIlS25STA/fobiSnx+22pIvdzrFKgMy3PB2nXIFG
4h+xpebBfNUNButhhhD0sHdJW23NdcxHu7CKmyRrsi9xfADEcMPhu+31MylNnlX2
nsq+U3Q9C3Z1A/60emoPFVfEfAvWvpOVO1fjyvbfmEwTzEbcWpAYPDCVAPansjg2
1EAAjBDmvHfS5oWsQuCC3J5iB5t9L5VC1O7qInhmjkNRGgOCrY9qceLML9u0mgMt
pYjAOU8a5PTirEUMtHd90PZ+fpEznMDN6YllIYxFd/gmzkwSz48XUBYXMloDxrsw
ZOLZU6xs7L1/KkgpWGW52ho8Dxyk0mlvxRP1W9FZ1EgFpLpYYO0CPB458feILFMb
hs38XEzSJxIwOZoTx1g53HYYzn01h806CQxegk3G7G3KLc7KVs7yAW+4D2nmIaBv
mGfXQZH2TG1GSKPTkI8ls1hwvQ+WYudlyROAKHwlpLrZG7bhvWXmOu6f11rB2yPz
QKdIghTkx+Xg3EY3cNC3FIcXokjPHSTdfCJtQAgn+mkiqWQR6kuIVIFLvW4IttXk
behyV5Og7Xhv0a5vuwiMwOTPqPO8s+lUPVO3DSnmzlPUUTzZsAFWqAM5locRrXcg
MNaj+QAIeqvLaz35dImFzvxDedyO8/Ymj2NTB8gsP7MXGoEKsOPpVxbiIpT19iM4
iS3zx8aRKUiA9euYrA9F0t8YAGU1Fely2BZ079mcmWGaKOYE3rt7ow7N31MG5Lf8
I5Y/vhfDgr5ifR04ch9b0vdIjl77mXEx3dE+oeh+viuE69YbyHKh5hFN68zq7LiO
bcZ+H/md621d6XenzLpfDrPNJOGmetnzQgcYdyvpHFIvLkRcEKs1BU6yRbNB+tvE
ATNVQgishCZe51Kn+RDG3WoFK+5RcJdPhM9W2Z+XXGCGCL+QbXZL2skQHZ+Ei2uo
4iCXwx4c5IwTdtp34PJUNkJw6qIMFM5iyE6mFmBJSCdjJslvcLrLG86A7R/fqxbW
tpTD/ryklWwIseHHFLFG8vFgwJljRJFnMRBDO89g7L13pYwuZpf4wBZVBys6taEJ
eH13BKwM8ULMYF2b01AQVJx5EtnXcGWeWTnBDkzoE/70uQl7skWbl+UoIhT4N16o
J5Ta5yYQN6hnR7wEVh6RrrVDBq48nFK8T9SuBcagijeunadis6982KwFtR8z+7TM
8IiWyHp8BrwLwMGkC81wNwXjarP9Z3GwJbJfsnwQPldQl7glwaacylxcRV1eXh47
w00roYg8U/8Avxvj2OLOD22ENwnt4iuOZNVIwKePoEt2qFSN8OXliR4F48F3+Ws7
/4BXWuSTWlbu6QjpJdsPBzj3acqH1y6ZSHUD5nmM/1HZPx9IgLM1RmDMA1+zzNp4
EvlZCRjhDKiD9nCmCzUwOfIqcCfZq58LHG6Q6N/Q79sLOSXLTgCWDkipvGLY81ns
AuMpJkSqpO2fGyOfbhvobCsGxFtvo8lt5K99pQ+8PDOIj1lyw7Zv+Etz4ozZ8KfY
JfhPb97dZTteEVky75i6XcDjb54Xn32k64FkFBCp+AtFU7iza5VzeF1oH2Mgz/0Y
QFLW2z6kiF/M5ryJM6cIwf2tNC5XEqVg2YdTfM/+TgMPEuR0qZtEl9tQX2j7IKk5
+7FEP3XwaiR/hzMieGwsFv60Pc8irH4EJA5j2KegDTr9nLD/JQxT0/EcvcLDU4YU
EBqGjoLofmLXFQmuvPASCoGEa1bSjEsUNf00IMMuqJXIMt0sbh69BTE+GYuUmwAj
UYVZJUSq2hy9xCyV0MXfgn+9XqKXg61MP1EbkeEG8sVvClFG2O3jIGeZcgreHfTZ
PEsDbfwtCKPyO+kZABz8P8YjjUhx3QjSv4LpyrzIYmsP6GBu//mLP4z1DQzL6bf8
V8mlxDePAhjVU8/f0yE/LCHkQX6wSheC0WETdy2VA+1EZiDfSuXBGeLMC7GyAbZz
KEzYUlgrpMGFDoDK5zCVN/rPttvpZRMavRbsYnRoT6hFz5mYCn4bcdA02m1U0Zrt
IsfHHALc/jyrt8+gCbiU+NQ69FS+v4DjMmEpq809KV23pRdgTgk20e9q5CQEH0XL
GrSlBtNfVcQo5amuFCbBgnIbpN8Wa4rcehaLJny5ZXUGeMma6nw0t39YtwxIbKDD
qmkkSbUTaHuR/3OfLSi225cAopQLNY+dC4j0LHINZKyebztSrewjxM3LkdIPuUgx
K5u9yMQrKcJg+13OiBo9qOr8YGjg1x2BxRGRN5jzGJxRNnzxVvfVjwJF4tDjHJqp
ewzp3lhp/U4IXUhJ9F+q89iF1frzr+YZKeQ6Ciotpz7gKN1+536tVQRfQ7XTLdTU
Y9/yxmybwTNRECueEPAOvyMGRk2ERlP/68bP1sA0HASAdZwRWxgGPGEV+NOb4hl7
iEcVqVfdF/AFLgLgUqp3IkuioYAkAdOPhssAFJvL74Tk1wrkdRB4dKPDw+wq5F/R
fT+BaMofHLTssgbuz7NyXBdobDpgBsNYAlkF0GoW4N3XztAG2232rrLtO0FrXVFC
q9185pUcyHkFTLdR5vufhjj05yu+JSmzaTU6fzT1Cl78tD36ZHJEcJWsd+6QoIUh
f7OVo1yrO9kUXJKtigZWbn4NMBvYKa/d93jcTgW+aFru1LLKz+jV2wnIFILg7KDN
GdpySL85YHXuWfvtAEBwJgMKGbJWT1LD7MjRQCcVQ9V96Gfs9IFkHAfbeavUELYf
CVkqV3P9oc5QAkMBmuzYejxoQliQY+Aj3/Tcgi5hVxH3wDC9kC/IwXTOn+l2NMTE
t4Btb7f2O1RcwrznQf/I6Jw/GPMMykh57wpmJ0MnCR4j4Cb4emKMwTG4AjRSQeDD
+DCCIaK65aYYxNoORGqtXdCao4YyruB+tdOxT8nVGI5Wz05XNcixZCNkAg4/XThR
d/lAud5d4YQPRdFx8vFpjQf+wTJ7t74H/L30BRJ815BxbMFyzU2ejgyb+fb/0oHi
LVjL6T0wq2v8ol2BbIosRuF/QRF2T8yBfBSRqFG3SkU5KX6U2LTywcltgKp9k/eq
aF/+IsSQOZssokyiyoRdFaT3HEtPe6qqD8+uu/2H0/m41xYU/K1l6UevxfqBNpEG
HbXgZTitjmwP6t8Fum8RNF9FpdaUQ0LnPCHm+2jG80D0OqZ0P834LTjhaLwZl8Cp
NiFFwGRSHglXd9L+XIPfr+qRM90UIC/OKcmS4EYa064SqqXSwLk55D09+AqFlBCm
z9Lz61jrjLm33VBD0MWadG7qMc4cyeouSJaTyclFtjAP3J1oEyvvNy93zCNbproc
BNnmVrHwT6hUYjC8RAgsZ29HxCJ8MJ9lIVyPu9zMHnsJGIGUXacx9M7r8PTJYDkH
svJp1JiLZmXGS4svMMRPCofgjIp2iP54H3QhBTGUBCgnNYH+ecRBvUlGS0MfzSM8
Q2zZev7pYmVuSQa+X87xa+YJPN/XoK14h7x/HfJjgJYItdz1iFd760SeQcAbz1Ay
l+c7Sa2uigskIyAMAK3SjbldpBkI4Ld/1H0UzTQrivjlpkmst714gxNTsPJFj8mW
wisj/3TaW2w8xXMXysTUbBb95L6nFD3N563npNMy0Yol6lL1HGicOShvUf3dEpm0
v1R1tsHxdS3OzmLQbsZnrFPbKAxGJEmvBjLkrCTiV1as8ioaoM3hcUJsSiw+jliA
DgprCFJJ0A6rYsYq8UoyAAZrsmw0KJbIw+enjNWmpqvJU3bSTFfw8eqTjz5kfDaB
8giuhrxFMTeFP8tbBrt6+3r1iTJu14KTbxdrvGRsSmQ90W4wMz0BQt5OrqrmBB/y
GXc3PbncLKN2P55mkj3kns0E550tzwDpsnhst/qJLIExbC60mgQdsXNt4HNnRWWc
zKtKEvI23+amLSL4RYqNsSQYbQBosCK8Pvl8+HscarvFghIvbdvT4MLRMJm+sZE3
JVKhsEFBq3EtymWqYIjT/EGts7ADfaxmgYoeAIzgFEK4yUm2dJZ635Hq5x6nn/ga
aR3ew7aVA+htkHFkmnQ7gWakJcDCXgUzdrOqTq30T3Wg4Wdd6FxrdTNX0KVXpRjJ
bltaY/0N5sQJbE5bmo2JBufOMRAX/s44tUPjlwEOTRjzAU/g6neE2K5U4kiZ29qw
C9m6ccz30fO/NRExm/ttJqpviwdUddrLVz4Nq8h9iM0BS4/KoJpMi7TJYglds1Sz
QwA8Y3ggHpHRo+UINErtg6GPvPjLZ+1ftkAM34GEjMiIvC5Zz8nD/AsU/zNSmL6w
7z25cAal1828aesmMQuhCELIXc9a7PyHsKUGSA+WEbAJToWUb1kAQg+Y3VncuUsU
pyrNJCEHDPs9CvT8mBg7Bb6Pgj1G4nyfNKps+ThICHg4FjN+hv5D1988hdOgj8tr
z05OoYAqP3kB5oTdadLcopUzaMZHSih8SPHB28coxZb6wV3i23JO3VvJabHAqLHg
eUykU4uGXu86pGt7k2dHIPdYdsa50F4LEvxqRzU7n3cQrnNDrXJMFV7/leUIrs9X
G0D0HOoEpkDD0G3m3B3Bvz3+Gr6AxQh8fNZ9/LvWez6SgzcMd6GX8E5UpHnwoqEV
TtB/udpihwo/x6mXRli8q25Ure2hDZcinzxI/EP9SXDKVdHLf953LZSndNENPFqD
P0WenXgrCpoPeZHc27yh+WM6clJEhc/moLHy40cr+Xp+kyaAwxbOViCKgJnQwtMa
B3IQC4+9vNWKA+OP0xAvmzLaHZVKUdah2vpNjwc4x7pce1Z6Do+sbP2utLH/hHjl
lHkIDozQd98F8D2AlfSMrsVHtG537UWttq2+g/5jlm1aBicR9dUa9q6OIKJQZQWb
MpVVn7Uh6xNYAay+HztpKKU3VnK6viwEcRaaeCg6PmNZNFi5Bmg2ONrsLiC06VNM
8suvLzB/Nckd3Pce6dnBAVdK+gx0DHFzPnoRs4O1GL+r3bevTqDCtdM0hwn2PYIG
HIgtY1xpdgmM67CPNKewZVmzUe7Jni2Ib5h1r0DBxjTI0zHGQgf+IBVUzcslcDm4
nsXECAKZtRl85MAIyPBd4OQRUEu32I8mxmV5BWtmC+TMJRLjzYs0pyz4Kiq2H3NL
Gc1TEzxePEuOBddlaOoyAB2vGn/ILFD0NLcKuyW+PhQNYckx8fThRBS6VCTHzmoG
e1eXWfqJ45/3uOUo36GGkdyK/WK2RWc7ZfxbS9uLVhQkHWgsMNk6fNdy2M+31bnI
binrhqV8KadqiipFq4SLtkM8jLKwF7p5hY0v3txYF8XIMx98v98lj7vWEWXc1u88
bbH+go236C8rAVzyhEPZYwajpC2hZFNqSKsLfWB4V76byRv+M2eXhJuL4l2emp5+
8znyLdXcN9M/0OXxqeoe6d8Yjxgp3x6SOTgZSc2BFRQU8qA0ppTge4e8Hwjiht9G
cInIuPlY99UL0SsDgqWNmI+EO7aBBf2db4mYWZLiNUEyRWc4+jXs9FQl1fu1jGCT
UWsH84bjHhs+z6nlKjjLLOI/JnGb3hpyAGaDZtbam5jc+E5bLwhmK2vcTMwrlfUu
/h53TPCgjiZfPLnuwOvb5Rjf4d7ntXfjX7HXsQg926spf5BhBNm0qq/BZgHtZe11
hzoelzK6gRXlAO4JhFMYy11MaMTogH1ubaeu9aL4I44Qtibxai9Ll83qXkUvosad
b6fG7wNeD9bcTUNLoFJ/wHKowGdL51QAVQZMLQLnu/iLuc0r+6OTmekmN7j3LIQ/
kv4s41zD0ENEskPN8/jWKDTCkzmwb9FsPrNw+F7LayAIf7d1tcxQusBdY9qNuFTe
LjjknKa+BXqAjbhcleAYFeMaa567WJGh0zn71/0XtPiK+Ume7TS96N3uSudJN4XK
ySpxJG21uWeUTCbS3ntZVdJ3wXewaToTrbFlJBuzrGmbKMSMb+0ZjdSj3pvm5T7S
zxCkgO8sjzdWL2EWedFAjkPFyjvaGa/+VN7xNuvslfeFQ7Nwu9R6v9/5MxLJoaYw
IaN9/ygcsmLFG7mSh/otfrhnXsJOto+8ofO2hX7X8YB6+tT0DbHnEnsp9JIKfrxL
LzACtiISBTCY8UQaQqQkAzSL8IQJCMLQfAHs1QaHaiVOJEYRvj41JE+Nk37qkiia
j4hGpr1Xl+1k7JFBV+iUOCNpOSIgNe9N8fLyMOE5MUusI9sSr4cHU4VyRLs9HXVL
GMAiGRM28p/yoxMlHVMKf5onpEuveiWPU9lru25IQ78knGuwU+++gnUcH9OU4K1j
lGt444sGYXtxD/4fmFi8H+t6H6IFm79w6McuQg8ZLZOp/t6l9Ubcuv9anwlcaKkn
YYJyxxy3bSsaMuLkV6qy7IlxqTBl44RkTOI/nVTGijXKjoIMmY+6wUbeBM3jpP5i
1wnoHQsUcyG4SBoKBFkz9MNJ4UVJXZ9kQiHf7G5Q78A4t6Db61mjcNul5u/1Knrj
BrddVxLuke0YHgz7XPkDG+pb9KBRCPy9oBxqLfdw3lDYodR/VHdX8vPK/NZ4iutN
mirovvxC1UbQX5408h3f7fKMtBQ8tJ5pD2rDPxDawdzHjXzAtxhDlZM6i9C6blXO
ii3PqdVddyvzvma7pgG97H8QzWgnNZ80oIn2m5rmmkInGKmDpSvkXzOHjLmFsv+P
GRd/IQEQwoKMqTaQvM7UNslrnBnhf1YsqO7+59CrWj49QMeREndLsd+Sg6Q606/p
yKpaqc80ZL3xBrrM2151MM04LM6i5YAJ5EsLF4k5MFhJdmuAX/xF4EvDQfmSSg3n
d/4ngjBj62Q5pQHm1HgQ/wSQ9AHZ9XPWq6y4n4wm+F7aCpxigDK4yb267njtT7jU
Bg9OP2kvee7Di0fYOAIRjtE1cjM1C2bdIMJB0xnY8+h+SlkAJ7fQsTiPQhza/vax
+/EolLeus88VFSBjukSlhg0K2JfHR4RQHq0zx3KCc10xVEG3IodKExp0n/r6x3PQ
430TU1Mm+MJqI2cSvVJTQp5yrq7jFEq/hjrjdaTUrCG0adFaqb2poxmS2QqcRjy9
RpZOyupzRnEjfCf2usWxTjz3vdHC8NJHzrWaqnKUtCtSU2K2n+jVESRYtYj7fEX9
1XdtdrysYklx3oUA3xrVbEMmkG7e92ryey4KvIkHaVwcOeW3oOeW1+J6yKvU7SLI
f5MLTXAsbmM9Bf1X84kYkwzFM4Nm0fWxa9M1Atlqs+IOaUxYKNeMlzrl5Z3gw/KR
j429JpvJ819O4KTqjWSSf7A7Fz6nwySTYVaEgV90If602cIS1CHMBXUEfI3VCSdM
RUxRvGRG4kT6Eg8vj5x3Oimz/h1zfBtKRy186sJSNfMghGv9A4U/yWLndVLLNZlC
y7j5QrJpt1qW1c6gWdo/CmEoEtQa9A/UW0MrNKP/OGtW4EUFVENkeF7OnkkVQtNq
UB/YRqBrOjgqaI95paMQ0cZvlekYPYeuXkLhth6jmXb0HMPdqFAIrUH0xOQBl9m/
/sQe63BVo1OVX5l+23c5o2Rqozhy7iBHI1s8KccjrhN2U29QtycgBW1lPTuMAgVJ
jtGGAcwMlCLfuOONjc4f26fRcoDTFPCvzj7fsUm1AdEMXV938Hwnn9HATHcuJ9kv
WOFg/LX1+Sm0Hqev1upxNVqydnRSZSVZNanc5dLwYbexj+MddcDhYeAzIxAqvNws
F2W7r4thAp8mjX7OwDQi2aqW2u0xQ1QGA2qha6lJeo2ZNd250vk+83HgfwL54MT0
G1a2SzncjcAEEKMDoiHNDRZtp36Kq9omnBtmgHLUVAVfLb+VgjzJGkavwbrIC+OU
t3Xx0J/X6vYq7rbT4QZ5ZDxrfM0hhSsi6R3BfRmGuiHxYQWyeKm33HqZPG5NzjRO
o4GSpZ2US2bzBAaDirH7hRahyt3joB2AeTRJnuSjrJz/LhLNC0y+nqf/czFd0Gl0
iMP7L0cZ9NWMIpOFe+5+zY1q8lQ6N2K3HHoSS4yyc1VStW7U8xxlTadxM3kyzKSz
d/9iuBtIiXyFWhkkhQytQI+KbsGwRIKFu05P0PeWSgCyAQTTJolpfLtA1vCTNSjY
szvHSBOHMKABO+NNDXfDvgXrBcFxlyxeV81tRfKFa7ZVExRXUB4pIt8c/N8+PR7/
VcjveYRoTBKm5Ne1v9RanTmbhbAJJUFgdNQoyj7kkj4LQkFKMm17CvEJez2d9Ddi
FkPKkaqFAwJ1K+kJSlKCQyC0tgRYxDS2dzKXp7P+lvfL/von/BuWGIkAJ2AG9WWk
uy6M2/mJ1Kbwt37ngFlwgpv6O4fRSEFdLmsk+VM2eys3xnn02/HZTEJwhGW6HRNY
y+SU7rAH0a8ebzfRE2W9GgLnzFmPKLzdmFeV+7Qq5IkCQDO0XlsnqD+K4332oSqg
bKkeSvxYFsvhV2S7rYJUJM9VM4isPHlyANRZ+tlO8QvtGAq/cByo2fUrhKxfug5Y
5mz6r1+/oVP3QFpA78FwTJarJ/pTF4R8E6ZBmLN/r2k5/LFcSdIlbTG8ZtmrAwh4
FJFB2qPiDGPq9ztTxeC7ws+sIvNilG6fAyilO3saF4ZaFQjFjnPhNKsFVVoNMu80
3TCd3UI+d6RmSwCfCrmTvBNR8JSCxnLSi15+8rNHoJKMfWR0h3kk9nR/7COtTa3U
lOkvrvcAFZ3eSaNwSZPgDK6fcsatdeuXhrVWRC4y4zqlpZXkKbpURh/1bB48FgyC
C11MbjrZ1YH799C4joXTyTE4m4CnC5I8rfzWJE1z3dMU9pJ6DB1EjqczGs37c+hj
VUSgczqMy3v8lTaZLtTHG66qibR6/GlAhVPyqY9XcoEaNmcNrxe0JG2Vhv1+pAjw
LZYz7uMINDHL34Dl3ZkFbLEVDSFl/mzMsIjNcqpWAZc1Qc1ECAOAZlAIUElAoiLB
terTH7xBiIpS8gewPvE0rvpNABqLvRnnmQ/UnOR1NSg34YjWv3ovOZCRoPSxhI6+
FZW0IsPB4Ng6bRe0Pi2JYRmM2vgoJr0YpRFCV5SukvPsJUpFVqH/OWgNRO/9Ihpg
xWh2MNBt+fazHSZxROItNeXi4HSNKx5YVYJpo3mVN2WQ0U5YhxRrsBzTwsld3hBb
NzvBHo23SjNT6b+WX5LWdbtxNCnRMoxBdAU5piTXcsFYmgwqAwTxKkI50qQP4Swu
eXd5+u1kMto8IW2KsZZ9yznWcLVbeLbJx19/WnHZIcI9ofPE4KsLW6xgnxb9MB5D
r4is4ct6dVvw7qQxRKbZGxecYaB3U6R7sc/z4jsMMqqccXa3XETzN9AVqCGtaEDa
4n3O0KrlxXHwgCrl9xXjtBXs9bCxRwtsDu1+o5/2xFMvnrS4PXcaePeC216NXeTf
NAkErkcdH+N40UXwTJCZ1xDXXEzjSmzHyUZlIa+A+Cr0diW2SylWcW/Bwcrg0Z3Z
0Vo0LVE28CnnhbTjLuJMSFIvms3ydBXLtDhOh8zMWr1MuJ2fRdqI8SGLRfZZHQSe
n27Tt2nrlqfzTVkjb89KzuVxSIO4Wvby0iP9ggGZ7tSwExgAUhIg3UfTmt85epD/
b3m1kdeuWLuG+xS+9xgSGErvurDPs1Xn4VTF16wMHOrsQ1f97MeO1d4rQW2QtrIv
FikXpkCUfGsdGEZWyoUYgkEfxL/ktpIARD1EBKQf0qBp9+RPUlz488EdDtGjHcjd
mhuUwnK4YdO1WwJZYxza9BsesUUO2DjqMT3mUdXMRHi62RHpbXOTO3ol7uP8MJ2w
+Of4mhpdU9VtY/EjuQFL7ny/V6dz8bn0yawgurFdKmyQseqk+lvZm+ZxnymrDNpl
0VYBcWDGendtLTwoeKxbGzVCLVphowVy1P5OT1lAnkZA9Mga9x+fAIeg3OT6EGuz
+WrId4++Gxn0eWV7kObWPtJL617Wr7pIzsxC2+YlLSqDkSDuaeN5gyxlTOTxxKqo
JMpxgu8XklPLrq/s1TOuuAC67f3IW7CLEbOE5AUFMpJdDQzBwfFV1Gf+9m3abN0c
FRlvZ+sq6xjhjgcwhT62/w5Zwd2s4x25f6xsRPWomqJ93tiX7l1O4/yHkJdGmtqC
KyyZMDBz4/2kiqB+kVQS8IzaYzWH2GCWNsgVSr4e5CCiyIRwwka24g3QqD/V/1ri
TaP3F0RSflenLtUolbGXeWX0kdfsR/tF8mMF+KFP3VqprICubLyqiGohEqjoZcJZ
iPo+aAo1tIFGlyuS4nq7NMRlXMxu/fP4tRoKjsuk/i8+f/MOh0ZbLY7mq6AIF17P
UNmDRvgjproE0B1tyObRD8bn+HI/bzL3CLf20BWuFZoPEwtGEbkvkYvoJ7isyPJ/
Z+LwJM/MsqBFdsNmZ5a1INlu4ZMVP96royz7liPsW3j6lAvg7BaRS0rV7iztdiby
8iNyobwKG99Fq+JuLsqLBJ7+heX3ldujrUi/71zImt682xfFXMFLjiSByojyjLfY
N+nVFGT4YzIDVagEkL90K7OBcA3HjmHSMcS4eT71NI8Pu6qJFUSfNomdPQjbGxJE
tmSbAiGprag/8b/qJpULhYv0FV5UTgcTSP2rvW/+tmyyd03mJJvTDwpqIT/Mcdbc
0uaPqGUXdPz7zROPMB/1L5xTOZ99SmYCi5w8EoKWTMzhPZqd1BBqZ/7eBVwTG5Rh
aFYAMtLmeAPim9qw6kN1dmixhz1voSydNiUXmYSDEJ9LUpnSr804IjMdZKBM301q
ZI5oTuLBT0CaldGQiFZVWgjiaBwX3Uzr/Dcp+L4DcGW/p+mOLFL9ewfrMbtyUb2P
w+7WdJV+XQHso+F3VLVb8ACLGRTWU1ROsPjKvfUNom4ewRriXair53g7D+W6mv3u
Aq+mZ07khcHr0SlEnTwDdMhPD5XI/5IiP8OG63ZPWT3Tof5R1Zlxyq6GsSfHg3j7
7jLZjTnOBjFyxOzKDUKkSSeh14Vw3e8Oeyokick7j4Ty8Xh0znv5bF+MBDromlBe
7M6uJmjAs8KurKYKabxKH0q8XSNk1FgfzbGwPvK3JAvfz7RWbYuQHSGa1oqS4kbz
CXjDcT81RgoFFVDNcdJjw1h4glZY8Gj/nkBREpkBMp3yuGLRr7gS2ts6um3S4p/i
e+VLKYsbhJT5MEiU/N2FjDlff5sbAIQ7cJYSNIS13rxrmWISatnpiFaZ7/S3ONVo
Y0CnFuIjQlVZQyn2rnMABEv2vX/ZVySh81XyaweqYcrLZT8xDIzxRZ7yGbvs7gCr
06QfEp6KAO3Bz2gTXOnOY5dg8OZ85HkwVgMsg78JQ6M72akSfa5tSWtJWPxTcqxN
8BL8sEjePblkbOMS/o5KNtpynCffjNKgBa/GNICBzCAZn2dyK5dQpb9PRzbchgrO
NsDUat87MLwf3DA2OsqeHOZ2gboALSkKlQfKuzz4uX7fXi0RTmd1eCg17LSXZlv0
MGIBDmilOW8QvYWeTKl8of780uwSzXEpm0QtIpiXHLUwm5/vyNBGsKl+MbsMUSOU
GUtP1kAmLL2jg9PhHUjuT3+J+1M83p2Yl3oN78YDLHM=
`protect end_protected
